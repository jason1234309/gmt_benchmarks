module top(
  input LIOB33_SING_X0Y50_IOB_X0Y50_IPAD,
  input LIOB33_X0Y51_IOB_X0Y51_IPAD,
  input LIOB33_X0Y51_IOB_X0Y52_IPAD,
  input LIOB33_X0Y53_IOB_X0Y53_IPAD,
  input LIOB33_X0Y53_IOB_X0Y54_IPAD,
  input LIOB33_X0Y55_IOB_X0Y55_IPAD,
  input LIOB33_X0Y55_IOB_X0Y56_IPAD,
  input LIOB33_X0Y57_IOB_X0Y57_IPAD,
  input LIOB33_X0Y57_IOB_X0Y58_IPAD,
  input LIOB33_X0Y59_IOB_X0Y59_IPAD,
  input LIOB33_X0Y59_IOB_X0Y60_IPAD,
  input LIOB33_X0Y61_IOB_X0Y61_IPAD,
  input LIOB33_X0Y61_IOB_X0Y62_IPAD,
  input LIOB33_X0Y63_IOB_X0Y63_IPAD,
  input LIOB33_X0Y63_IOB_X0Y64_IPAD,
  input LIOB33_X0Y65_IOB_X0Y65_IPAD,
  input LIOB33_X0Y65_IOB_X0Y66_IPAD,
  input LIOB33_X0Y67_IOB_X0Y67_IPAD,
  input LIOB33_X0Y67_IOB_X0Y68_IPAD,
  input LIOB33_X0Y69_IOB_X0Y69_IPAD,
  input LIOB33_X0Y69_IOB_X0Y70_IPAD,
  input LIOB33_X0Y71_IOB_X0Y71_IPAD,
  input LIOB33_X0Y71_IOB_X0Y72_IPAD,
  input LIOB33_X0Y73_IOB_X0Y73_IPAD,
  input LIOB33_X0Y73_IOB_X0Y74_IPAD,
  input LIOB33_X0Y75_IOB_X0Y75_IPAD,
  input LIOB33_X0Y75_IOB_X0Y76_IPAD,
  input LIOB33_X0Y77_IOB_X0Y77_IPAD,
  input LIOB33_X0Y77_IOB_X0Y78_IPAD,
  input LIOB33_X0Y79_IOB_X0Y79_IPAD,
  input RIOB33_SING_X105Y100_IOB_X1Y100_IPAD,
  input RIOB33_SING_X105Y149_IOB_X1Y149_IPAD,
  input RIOB33_X105Y101_IOB_X1Y101_IPAD,
  input RIOB33_X105Y101_IOB_X1Y102_IPAD,
  input RIOB33_X105Y103_IOB_X1Y103_IPAD,
  input RIOB33_X105Y103_IOB_X1Y104_IPAD,
  input RIOB33_X105Y105_IOB_X1Y105_IPAD,
  input RIOB33_X105Y105_IOB_X1Y106_IPAD,
  input RIOB33_X105Y107_IOB_X1Y107_IPAD,
  input RIOB33_X105Y107_IOB_X1Y108_IPAD,
  input RIOB33_X105Y109_IOB_X1Y109_IPAD,
  input RIOB33_X105Y109_IOB_X1Y110_IPAD,
  input RIOB33_X105Y111_IOB_X1Y111_IPAD,
  input RIOB33_X105Y111_IOB_X1Y112_IPAD,
  input RIOB33_X105Y113_IOB_X1Y113_IPAD,
  input RIOB33_X105Y113_IOB_X1Y114_IPAD,
  input RIOB33_X105Y115_IOB_X1Y115_IPAD,
  input RIOB33_X105Y115_IOB_X1Y116_IPAD,
  input RIOB33_X105Y117_IOB_X1Y117_IPAD,
  input RIOB33_X105Y117_IOB_X1Y118_IPAD,
  input RIOB33_X105Y119_IOB_X1Y119_IPAD,
  input RIOB33_X105Y119_IOB_X1Y120_IPAD,
  input RIOB33_X105Y121_IOB_X1Y121_IPAD,
  input RIOB33_X105Y121_IOB_X1Y122_IPAD,
  input RIOB33_X105Y123_IOB_X1Y123_IPAD,
  input RIOB33_X105Y123_IOB_X1Y124_IPAD,
  input RIOB33_X105Y125_IOB_X1Y125_IPAD,
  input RIOB33_X105Y125_IOB_X1Y126_IPAD,
  input RIOB33_X105Y127_IOB_X1Y127_IPAD,
  input RIOB33_X105Y127_IOB_X1Y128_IPAD,
  input RIOB33_X105Y129_IOB_X1Y129_IPAD,
  input RIOB33_X105Y129_IOB_X1Y130_IPAD,
  input RIOB33_X105Y131_IOB_X1Y131_IPAD,
  input RIOB33_X105Y131_IOB_X1Y132_IPAD,
  input RIOB33_X105Y133_IOB_X1Y133_IPAD,
  input RIOB33_X105Y133_IOB_X1Y134_IPAD,
  input RIOB33_X105Y135_IOB_X1Y135_IPAD,
  input RIOB33_X105Y135_IOB_X1Y136_IPAD,
  input RIOB33_X105Y137_IOB_X1Y137_IPAD,
  input RIOB33_X105Y137_IOB_X1Y138_IPAD,
  input RIOB33_X105Y139_IOB_X1Y139_IPAD,
  input RIOB33_X105Y139_IOB_X1Y140_IPAD,
  input RIOB33_X105Y141_IOB_X1Y141_IPAD,
  input RIOB33_X105Y141_IOB_X1Y142_IPAD,
  input RIOB33_X105Y143_IOB_X1Y143_IPAD,
  input RIOB33_X105Y143_IOB_X1Y144_IPAD,
  input RIOB33_X105Y145_IOB_X1Y145_IPAD,
  input RIOB33_X105Y145_IOB_X1Y146_IPAD,
  input RIOB33_X105Y147_IOB_X1Y147_IPAD,
  input RIOB33_X105Y147_IOB_X1Y148_IPAD,
  output LIOB33_SING_X0Y100_IOB_X0Y100_OPAD,
  output LIOB33_SING_X0Y149_IOB_X0Y149_OPAD,
  output LIOB33_SING_X0Y150_IOB_X0Y150_OPAD,
  output LIOB33_SING_X0Y199_IOB_X0Y199_OPAD,
  output LIOB33_X0Y101_IOB_X0Y101_OPAD,
  output LIOB33_X0Y101_IOB_X0Y102_OPAD,
  output LIOB33_X0Y103_IOB_X0Y103_OPAD,
  output LIOB33_X0Y103_IOB_X0Y104_OPAD,
  output LIOB33_X0Y105_IOB_X0Y105_OPAD,
  output LIOB33_X0Y105_IOB_X0Y106_OPAD,
  output LIOB33_X0Y107_IOB_X0Y107_OPAD,
  output LIOB33_X0Y107_IOB_X0Y108_OPAD,
  output LIOB33_X0Y109_IOB_X0Y109_OPAD,
  output LIOB33_X0Y109_IOB_X0Y110_OPAD,
  output LIOB33_X0Y111_IOB_X0Y111_OPAD,
  output LIOB33_X0Y111_IOB_X0Y112_OPAD,
  output LIOB33_X0Y113_IOB_X0Y113_OPAD,
  output LIOB33_X0Y113_IOB_X0Y114_OPAD,
  output LIOB33_X0Y115_IOB_X0Y115_OPAD,
  output LIOB33_X0Y115_IOB_X0Y116_OPAD,
  output LIOB33_X0Y117_IOB_X0Y117_OPAD,
  output LIOB33_X0Y117_IOB_X0Y118_OPAD,
  output LIOB33_X0Y119_IOB_X0Y119_OPAD,
  output LIOB33_X0Y119_IOB_X0Y120_OPAD,
  output LIOB33_X0Y121_IOB_X0Y121_OPAD,
  output LIOB33_X0Y121_IOB_X0Y122_OPAD,
  output LIOB33_X0Y123_IOB_X0Y123_OPAD,
  output LIOB33_X0Y123_IOB_X0Y124_OPAD,
  output LIOB33_X0Y125_IOB_X0Y125_OPAD,
  output LIOB33_X0Y125_IOB_X0Y126_OPAD,
  output LIOB33_X0Y127_IOB_X0Y127_OPAD,
  output LIOB33_X0Y127_IOB_X0Y128_OPAD,
  output LIOB33_X0Y129_IOB_X0Y129_OPAD,
  output LIOB33_X0Y129_IOB_X0Y130_OPAD,
  output LIOB33_X0Y131_IOB_X0Y131_OPAD,
  output LIOB33_X0Y131_IOB_X0Y132_OPAD,
  output LIOB33_X0Y133_IOB_X0Y133_OPAD,
  output LIOB33_X0Y133_IOB_X0Y134_OPAD,
  output LIOB33_X0Y135_IOB_X0Y135_OPAD,
  output LIOB33_X0Y135_IOB_X0Y136_OPAD,
  output LIOB33_X0Y137_IOB_X0Y137_OPAD,
  output LIOB33_X0Y137_IOB_X0Y138_OPAD,
  output LIOB33_X0Y139_IOB_X0Y139_OPAD,
  output LIOB33_X0Y139_IOB_X0Y140_OPAD,
  output LIOB33_X0Y141_IOB_X0Y141_OPAD,
  output LIOB33_X0Y141_IOB_X0Y142_OPAD,
  output LIOB33_X0Y143_IOB_X0Y143_OPAD,
  output LIOB33_X0Y145_IOB_X0Y145_OPAD,
  output LIOB33_X0Y145_IOB_X0Y146_OPAD,
  output LIOB33_X0Y147_IOB_X0Y147_OPAD,
  output LIOB33_X0Y147_IOB_X0Y148_OPAD,
  output LIOB33_X0Y151_IOB_X0Y151_OPAD,
  output LIOB33_X0Y151_IOB_X0Y152_OPAD,
  output LIOB33_X0Y153_IOB_X0Y153_OPAD,
  output LIOB33_X0Y153_IOB_X0Y154_OPAD,
  output LIOB33_X0Y155_IOB_X0Y155_OPAD,
  output LIOB33_X0Y155_IOB_X0Y156_OPAD,
  output LIOB33_X0Y157_IOB_X0Y157_OPAD,
  output LIOB33_X0Y157_IOB_X0Y158_OPAD,
  output LIOB33_X0Y159_IOB_X0Y159_OPAD,
  output LIOB33_X0Y159_IOB_X0Y160_OPAD,
  output LIOB33_X0Y161_IOB_X0Y161_OPAD,
  output LIOB33_X0Y161_IOB_X0Y162_OPAD,
  output LIOB33_X0Y163_IOB_X0Y163_OPAD,
  output LIOB33_X0Y163_IOB_X0Y164_OPAD,
  output LIOB33_X0Y165_IOB_X0Y165_OPAD,
  output LIOB33_X0Y165_IOB_X0Y166_OPAD,
  output LIOB33_X0Y167_IOB_X0Y167_OPAD,
  output LIOB33_X0Y167_IOB_X0Y168_OPAD,
  output LIOB33_X0Y169_IOB_X0Y169_OPAD,
  output LIOB33_X0Y169_IOB_X0Y170_OPAD,
  output LIOB33_X0Y171_IOB_X0Y171_OPAD,
  output LIOB33_X0Y171_IOB_X0Y172_OPAD,
  output LIOB33_X0Y173_IOB_X0Y173_OPAD,
  output LIOB33_X0Y173_IOB_X0Y174_OPAD,
  output LIOB33_X0Y175_IOB_X0Y175_OPAD,
  output LIOB33_X0Y175_IOB_X0Y176_OPAD,
  output LIOB33_X0Y177_IOB_X0Y177_OPAD,
  output LIOB33_X0Y177_IOB_X0Y178_OPAD,
  output LIOB33_X0Y179_IOB_X0Y179_OPAD,
  output LIOB33_X0Y179_IOB_X0Y180_OPAD,
  output LIOB33_X0Y181_IOB_X0Y181_OPAD,
  output LIOB33_X0Y181_IOB_X0Y182_OPAD,
  output LIOB33_X0Y183_IOB_X0Y183_OPAD,
  output LIOB33_X0Y183_IOB_X0Y184_OPAD,
  output LIOB33_X0Y185_IOB_X0Y185_OPAD,
  output LIOB33_X0Y185_IOB_X0Y186_OPAD,
  output LIOB33_X0Y187_IOB_X0Y187_OPAD,
  output LIOB33_X0Y187_IOB_X0Y188_OPAD,
  output LIOB33_X0Y189_IOB_X0Y189_OPAD,
  output LIOB33_X0Y189_IOB_X0Y190_OPAD,
  output LIOB33_X0Y191_IOB_X0Y191_OPAD,
  output LIOB33_X0Y191_IOB_X0Y192_OPAD,
  output LIOB33_X0Y193_IOB_X0Y193_OPAD,
  output LIOB33_X0Y193_IOB_X0Y194_OPAD,
  output LIOB33_X0Y195_IOB_X0Y195_OPAD,
  output LIOB33_X0Y195_IOB_X0Y196_OPAD,
  output LIOB33_X0Y197_IOB_X0Y197_OPAD,
  output LIOB33_X0Y197_IOB_X0Y198_OPAD,
  output LIOB33_X0Y79_IOB_X0Y80_OPAD,
  output RIOB33_SING_X105Y150_IOB_X1Y150_OPAD,
  output RIOB33_SING_X105Y199_IOB_X1Y199_OPAD,
  output RIOB33_X105Y151_IOB_X1Y151_OPAD,
  output RIOB33_X105Y151_IOB_X1Y152_OPAD,
  output RIOB33_X105Y153_IOB_X1Y153_OPAD,
  output RIOB33_X105Y153_IOB_X1Y154_OPAD,
  output RIOB33_X105Y155_IOB_X1Y155_OPAD,
  output RIOB33_X105Y155_IOB_X1Y156_OPAD,
  output RIOB33_X105Y157_IOB_X1Y157_OPAD,
  output RIOB33_X105Y157_IOB_X1Y158_OPAD,
  output RIOB33_X105Y159_IOB_X1Y159_OPAD,
  output RIOB33_X105Y159_IOB_X1Y160_OPAD,
  output RIOB33_X105Y161_IOB_X1Y161_OPAD,
  output RIOB33_X105Y161_IOB_X1Y162_OPAD,
  output RIOB33_X105Y163_IOB_X1Y163_OPAD,
  output RIOB33_X105Y163_IOB_X1Y164_OPAD,
  output RIOB33_X105Y165_IOB_X1Y165_OPAD,
  output RIOB33_X105Y165_IOB_X1Y166_OPAD,
  output RIOB33_X105Y167_IOB_X1Y167_OPAD,
  output RIOB33_X105Y167_IOB_X1Y168_OPAD,
  output RIOB33_X105Y169_IOB_X1Y169_OPAD,
  output RIOB33_X105Y169_IOB_X1Y170_OPAD,
  output RIOB33_X105Y171_IOB_X1Y171_OPAD,
  output RIOB33_X105Y171_IOB_X1Y172_OPAD,
  output RIOB33_X105Y173_IOB_X1Y173_OPAD,
  output RIOB33_X105Y173_IOB_X1Y174_OPAD,
  output RIOB33_X105Y175_IOB_X1Y175_OPAD,
  output RIOB33_X105Y175_IOB_X1Y176_OPAD,
  output RIOB33_X105Y177_IOB_X1Y177_OPAD,
  output RIOB33_X105Y177_IOB_X1Y178_OPAD,
  output RIOB33_X105Y179_IOB_X1Y179_OPAD,
  output RIOB33_X105Y179_IOB_X1Y180_OPAD,
  output RIOB33_X105Y181_IOB_X1Y181_OPAD,
  output RIOB33_X105Y181_IOB_X1Y182_OPAD,
  output RIOB33_X105Y183_IOB_X1Y183_OPAD,
  output RIOB33_X105Y183_IOB_X1Y184_OPAD,
  output RIOB33_X105Y185_IOB_X1Y185_OPAD,
  output RIOB33_X105Y185_IOB_X1Y186_OPAD,
  output RIOB33_X105Y187_IOB_X1Y187_OPAD,
  output RIOB33_X105Y187_IOB_X1Y188_OPAD,
  output RIOB33_X105Y189_IOB_X1Y189_OPAD,
  output RIOB33_X105Y189_IOB_X1Y190_OPAD,
  output RIOB33_X105Y191_IOB_X1Y191_OPAD,
  output RIOB33_X105Y191_IOB_X1Y192_OPAD,
  output RIOB33_X105Y193_IOB_X1Y193_OPAD,
  output RIOB33_X105Y193_IOB_X1Y194_OPAD,
  output RIOB33_X105Y195_IOB_X1Y195_OPAD,
  output RIOB33_X105Y195_IOB_X1Y196_OPAD,
  output RIOB33_X105Y197_IOB_X1Y197_OPAD,
  output RIOB33_X105Y197_IOB_X1Y198_OPAD
  );
  wire [0:0] CLBLL_L_X2Y109_SLICE_X0Y109_A;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X0Y109_A1;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X0Y109_A2;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X0Y109_A3;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X0Y109_A4;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X0Y109_A5;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X0Y109_A6;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X0Y109_AO5;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X0Y109_AO6;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X0Y109_A_CY;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X0Y109_A_XOR;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X0Y109_B;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X0Y109_B1;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X0Y109_B2;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X0Y109_B3;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X0Y109_B4;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X0Y109_B5;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X0Y109_B6;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X0Y109_BO5;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X0Y109_BO6;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X0Y109_B_CY;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X0Y109_B_XOR;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X0Y109_C;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X0Y109_C1;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X0Y109_C2;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X0Y109_C3;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X0Y109_C4;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X0Y109_C5;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X0Y109_C6;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X0Y109_CO5;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X0Y109_CO6;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X0Y109_C_CY;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X0Y109_C_XOR;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X0Y109_D;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X0Y109_D1;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X0Y109_D2;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X0Y109_D3;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X0Y109_D4;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X0Y109_D5;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X0Y109_D6;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X0Y109_DO5;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X0Y109_DO6;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X0Y109_D_CY;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X0Y109_D_XOR;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X1Y109_A;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X1Y109_A1;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X1Y109_A2;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X1Y109_A3;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X1Y109_A4;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X1Y109_A5;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X1Y109_A6;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X1Y109_AO5;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X1Y109_AO6;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X1Y109_A_CY;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X1Y109_A_XOR;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X1Y109_B;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X1Y109_B1;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X1Y109_B2;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X1Y109_B3;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X1Y109_B4;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X1Y109_B5;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X1Y109_B6;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X1Y109_BO5;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X1Y109_BO6;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X1Y109_B_CY;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X1Y109_B_XOR;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X1Y109_C;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X1Y109_C1;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X1Y109_C2;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X1Y109_C3;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X1Y109_C4;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X1Y109_C5;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X1Y109_C6;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X1Y109_CO5;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X1Y109_CO6;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X1Y109_C_CY;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X1Y109_C_XOR;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X1Y109_D;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X1Y109_D1;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X1Y109_D2;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X1Y109_D3;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X1Y109_D4;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X1Y109_D5;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X1Y109_D6;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X1Y109_DO5;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X1Y109_DO6;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X1Y109_D_CY;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X1Y109_D_XOR;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X0Y110_A;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X0Y110_A1;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X0Y110_A2;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X0Y110_A3;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X0Y110_A4;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X0Y110_A5;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X0Y110_A6;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X0Y110_AMUX;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X0Y110_AO5;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X0Y110_AO6;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X0Y110_A_CY;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X0Y110_A_XOR;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X0Y110_B;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X0Y110_B1;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X0Y110_B2;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X0Y110_B3;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X0Y110_B4;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X0Y110_B5;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X0Y110_B6;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X0Y110_BO5;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X0Y110_BO6;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X0Y110_B_CY;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X0Y110_B_XOR;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X0Y110_C;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X0Y110_C1;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X0Y110_C2;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X0Y110_C3;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X0Y110_C4;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X0Y110_C5;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X0Y110_C6;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X0Y110_CO5;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X0Y110_CO6;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X0Y110_C_CY;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X0Y110_C_XOR;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X0Y110_D;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X0Y110_D1;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X0Y110_D2;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X0Y110_D3;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X0Y110_D4;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X0Y110_D5;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X0Y110_D6;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X0Y110_DO5;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X0Y110_DO6;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X0Y110_D_CY;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X0Y110_D_XOR;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X1Y110_A;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X1Y110_A1;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X1Y110_A2;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X1Y110_A3;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X1Y110_A4;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X1Y110_A5;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X1Y110_A6;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X1Y110_AO5;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X1Y110_AO6;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X1Y110_A_CY;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X1Y110_A_XOR;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X1Y110_B;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X1Y110_B1;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X1Y110_B2;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X1Y110_B3;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X1Y110_B4;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X1Y110_B5;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X1Y110_B6;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X1Y110_BO5;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X1Y110_BO6;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X1Y110_B_CY;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X1Y110_B_XOR;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X1Y110_C;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X1Y110_C1;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X1Y110_C2;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X1Y110_C3;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X1Y110_C4;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X1Y110_C5;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X1Y110_C6;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X1Y110_CO5;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X1Y110_CO6;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X1Y110_C_CY;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X1Y110_C_XOR;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X1Y110_D;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X1Y110_D1;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X1Y110_D2;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X1Y110_D3;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X1Y110_D4;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X1Y110_D5;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X1Y110_D6;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X1Y110_DO5;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X1Y110_DO6;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X1Y110_D_CY;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X1Y110_D_XOR;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X0Y111_A;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X0Y111_A1;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X0Y111_A2;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X0Y111_A3;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X0Y111_A4;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X0Y111_A5;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X0Y111_A6;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X0Y111_AMUX;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X0Y111_AO5;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X0Y111_AO6;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X0Y111_A_CY;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X0Y111_A_XOR;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X0Y111_B;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X0Y111_B1;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X0Y111_B2;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X0Y111_B3;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X0Y111_B4;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X0Y111_B5;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X0Y111_B6;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X0Y111_BMUX;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X0Y111_BO5;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X0Y111_BO6;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X0Y111_B_CY;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X0Y111_B_XOR;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X0Y111_C;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X0Y111_C1;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X0Y111_C2;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X0Y111_C3;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X0Y111_C4;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X0Y111_C5;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X0Y111_C6;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X0Y111_CMUX;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X0Y111_CO5;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X0Y111_CO6;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X0Y111_C_CY;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X0Y111_C_XOR;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X0Y111_D;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X0Y111_D1;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X0Y111_D2;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X0Y111_D3;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X0Y111_D4;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X0Y111_D5;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X0Y111_D6;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X0Y111_DMUX;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X0Y111_DO5;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X0Y111_DO6;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X0Y111_D_CY;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X0Y111_D_XOR;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X1Y111_A;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X1Y111_A1;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X1Y111_A2;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X1Y111_A3;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X1Y111_A4;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X1Y111_A5;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X1Y111_A6;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X1Y111_AO5;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X1Y111_AO6;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X1Y111_A_CY;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X1Y111_A_XOR;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X1Y111_B;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X1Y111_B1;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X1Y111_B2;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X1Y111_B3;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X1Y111_B4;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X1Y111_B5;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X1Y111_B6;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X1Y111_BO5;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X1Y111_BO6;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X1Y111_B_CY;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X1Y111_B_XOR;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X1Y111_C;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X1Y111_C1;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X1Y111_C2;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X1Y111_C3;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X1Y111_C4;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X1Y111_C5;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X1Y111_C6;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X1Y111_CO5;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X1Y111_CO6;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X1Y111_C_CY;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X1Y111_C_XOR;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X1Y111_D;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X1Y111_D1;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X1Y111_D2;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X1Y111_D3;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X1Y111_D4;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X1Y111_D5;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X1Y111_D6;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X1Y111_DO5;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X1Y111_DO6;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X1Y111_D_CY;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X1Y111_D_XOR;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X0Y112_A;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X0Y112_A1;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X0Y112_A2;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X0Y112_A3;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X0Y112_A4;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X0Y112_A5;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X0Y112_A6;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X0Y112_AO5;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X0Y112_AO6;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X0Y112_A_CY;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X0Y112_A_XOR;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X0Y112_B;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X0Y112_B1;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X0Y112_B2;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X0Y112_B3;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X0Y112_B4;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X0Y112_B5;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X0Y112_B6;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X0Y112_BO5;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X0Y112_BO6;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X0Y112_B_CY;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X0Y112_B_XOR;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X0Y112_C;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X0Y112_C1;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X0Y112_C2;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X0Y112_C3;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X0Y112_C4;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X0Y112_C5;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X0Y112_C6;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X0Y112_CO5;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X0Y112_CO6;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X0Y112_C_CY;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X0Y112_C_XOR;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X0Y112_D;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X0Y112_D1;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X0Y112_D2;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X0Y112_D3;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X0Y112_D4;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X0Y112_D5;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X0Y112_D6;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X0Y112_DO5;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X0Y112_DO6;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X0Y112_D_CY;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X0Y112_D_XOR;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X1Y112_A;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X1Y112_A1;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X1Y112_A2;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X1Y112_A3;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X1Y112_A4;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X1Y112_A5;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X1Y112_A5Q;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X1Y112_A6;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X1Y112_AMUX;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X1Y112_AO5;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X1Y112_AO6;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X1Y112_AQ;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X1Y112_AX;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X1Y112_A_CY;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X1Y112_A_XOR;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X1Y112_B;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X1Y112_B1;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X1Y112_B2;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X1Y112_B3;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X1Y112_B4;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X1Y112_B5;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X1Y112_B6;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X1Y112_BO5;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X1Y112_BO6;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X1Y112_BQ;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X1Y112_B_CY;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X1Y112_B_XOR;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X1Y112_C;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X1Y112_C1;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X1Y112_C2;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X1Y112_C3;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X1Y112_C4;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X1Y112_C5;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X1Y112_C6;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X1Y112_CLK;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X1Y112_CMUX;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X1Y112_CO5;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X1Y112_CO6;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X1Y112_C_CY;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X1Y112_C_XOR;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X1Y112_D;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X1Y112_D1;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X1Y112_D2;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X1Y112_D3;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X1Y112_D4;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X1Y112_D5;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X1Y112_D6;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X1Y112_DO5;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X1Y112_DO6;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X1Y112_D_CY;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X1Y112_D_XOR;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X0Y113_A;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X0Y113_A1;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X0Y113_A2;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X0Y113_A3;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X0Y113_A4;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X0Y113_A5;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X0Y113_A6;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X0Y113_AMUX;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X0Y113_AO5;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X0Y113_AO6;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X0Y113_A_CY;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X0Y113_A_XOR;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X0Y113_B;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X0Y113_B1;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X0Y113_B2;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X0Y113_B3;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X0Y113_B4;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X0Y113_B5;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X0Y113_B6;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X0Y113_BO5;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X0Y113_BO6;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X0Y113_B_CY;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X0Y113_B_XOR;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X0Y113_C;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X0Y113_C1;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X0Y113_C2;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X0Y113_C3;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X0Y113_C4;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X0Y113_C5;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X0Y113_C6;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X0Y113_CO5;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X0Y113_CO6;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X0Y113_C_CY;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X0Y113_C_XOR;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X0Y113_D;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X0Y113_D1;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X0Y113_D2;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X0Y113_D3;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X0Y113_D4;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X0Y113_D5;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X0Y113_D6;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X0Y113_DO5;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X0Y113_DO6;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X0Y113_D_CY;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X0Y113_D_XOR;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X1Y113_A;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X1Y113_A1;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X1Y113_A2;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X1Y113_A3;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X1Y113_A4;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X1Y113_A5;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X1Y113_A6;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X1Y113_AO5;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X1Y113_AO6;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X1Y113_AQ;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X1Y113_A_CY;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X1Y113_A_XOR;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X1Y113_B;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X1Y113_B1;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X1Y113_B2;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X1Y113_B3;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X1Y113_B4;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X1Y113_B5;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X1Y113_B6;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X1Y113_BO5;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X1Y113_BO6;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X1Y113_BQ;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X1Y113_B_CY;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X1Y113_B_XOR;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X1Y113_C;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X1Y113_C1;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X1Y113_C2;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X1Y113_C3;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X1Y113_C4;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X1Y113_C5;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X1Y113_C5Q;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X1Y113_C6;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X1Y113_CLK;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X1Y113_CMUX;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X1Y113_CO5;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X1Y113_CO6;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X1Y113_CQ;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X1Y113_C_CY;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X1Y113_C_XOR;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X1Y113_D;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X1Y113_D1;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X1Y113_D2;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X1Y113_D3;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X1Y113_D4;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X1Y113_D5;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X1Y113_D6;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X1Y113_DO5;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X1Y113_DO6;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X1Y113_D_CY;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X1Y113_D_XOR;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X0Y114_A;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X0Y114_A1;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X0Y114_A2;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X0Y114_A3;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X0Y114_A4;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X0Y114_A5;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X0Y114_A6;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X0Y114_AO5;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X0Y114_AO6;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X0Y114_A_CY;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X0Y114_A_XOR;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X0Y114_B;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X0Y114_B1;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X0Y114_B2;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X0Y114_B3;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X0Y114_B4;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X0Y114_B5;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X0Y114_B6;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X0Y114_BO5;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X0Y114_BO6;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X0Y114_B_CY;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X0Y114_B_XOR;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X0Y114_C;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X0Y114_C1;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X0Y114_C2;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X0Y114_C3;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X0Y114_C4;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X0Y114_C5;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X0Y114_C6;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X0Y114_CO5;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X0Y114_CO6;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X0Y114_C_CY;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X0Y114_C_XOR;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X0Y114_D;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X0Y114_D1;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X0Y114_D2;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X0Y114_D3;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X0Y114_D4;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X0Y114_D5;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X0Y114_D6;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X0Y114_DO5;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X0Y114_DO6;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X0Y114_D_CY;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X0Y114_D_XOR;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X1Y114_A;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X1Y114_A1;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X1Y114_A2;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X1Y114_A3;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X1Y114_A4;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X1Y114_A5;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X1Y114_A6;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X1Y114_AO5;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X1Y114_AO6;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X1Y114_AQ;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X1Y114_A_CY;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X1Y114_A_XOR;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X1Y114_B;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X1Y114_B1;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X1Y114_B2;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X1Y114_B3;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X1Y114_B4;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X1Y114_B5;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X1Y114_B6;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X1Y114_BMUX;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X1Y114_BO5;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X1Y114_BO6;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X1Y114_B_CY;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X1Y114_B_XOR;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X1Y114_C;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X1Y114_C1;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X1Y114_C2;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X1Y114_C3;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X1Y114_C4;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X1Y114_C5;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X1Y114_C6;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X1Y114_CLK;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X1Y114_CMUX;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X1Y114_CO5;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X1Y114_CO6;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X1Y114_C_CY;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X1Y114_C_XOR;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X1Y114_D;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X1Y114_D1;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X1Y114_D2;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X1Y114_D3;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X1Y114_D4;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X1Y114_D5;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X1Y114_D6;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X1Y114_DO5;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X1Y114_DO6;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X1Y114_D_CY;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X1Y114_D_XOR;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X0Y115_A;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X0Y115_A1;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X0Y115_A2;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X0Y115_A3;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X0Y115_A4;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X0Y115_A5;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X0Y115_A6;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X0Y115_AO5;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X0Y115_AO6;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X0Y115_A_CY;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X0Y115_A_XOR;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X0Y115_B;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X0Y115_B1;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X0Y115_B2;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X0Y115_B3;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X0Y115_B4;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X0Y115_B5;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X0Y115_B6;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X0Y115_BO5;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X0Y115_BO6;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X0Y115_B_CY;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X0Y115_B_XOR;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X0Y115_C;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X0Y115_C1;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X0Y115_C2;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X0Y115_C3;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X0Y115_C4;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X0Y115_C5;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X0Y115_C6;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X0Y115_CO5;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X0Y115_CO6;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X0Y115_C_CY;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X0Y115_C_XOR;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X0Y115_D;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X0Y115_D1;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X0Y115_D2;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X0Y115_D3;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X0Y115_D4;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X0Y115_D5;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X0Y115_D6;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X0Y115_DO5;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X0Y115_DO6;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X0Y115_D_CY;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X0Y115_D_XOR;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X1Y115_A;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X1Y115_A1;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X1Y115_A2;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X1Y115_A3;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X1Y115_A4;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X1Y115_A5;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X1Y115_A6;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X1Y115_AO5;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X1Y115_AO6;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X1Y115_AQ;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X1Y115_A_CY;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X1Y115_A_XOR;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X1Y115_B;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X1Y115_B1;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X1Y115_B2;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X1Y115_B3;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X1Y115_B4;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X1Y115_B5;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X1Y115_B6;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X1Y115_BO5;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X1Y115_BO6;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X1Y115_BQ;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X1Y115_B_CY;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X1Y115_B_XOR;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X1Y115_C;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X1Y115_C1;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X1Y115_C2;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X1Y115_C3;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X1Y115_C4;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X1Y115_C5;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X1Y115_C6;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X1Y115_CLK;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X1Y115_CO5;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X1Y115_CO6;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X1Y115_C_CY;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X1Y115_C_XOR;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X1Y115_D;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X1Y115_D1;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X1Y115_D2;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X1Y115_D3;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X1Y115_D4;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X1Y115_D5;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X1Y115_D6;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X1Y115_DO5;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X1Y115_DO6;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X1Y115_D_CY;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X1Y115_D_XOR;
  wire [0:0] CLBLL_L_X2Y116_SLICE_X0Y116_A;
  wire [0:0] CLBLL_L_X2Y116_SLICE_X0Y116_A1;
  wire [0:0] CLBLL_L_X2Y116_SLICE_X0Y116_A2;
  wire [0:0] CLBLL_L_X2Y116_SLICE_X0Y116_A3;
  wire [0:0] CLBLL_L_X2Y116_SLICE_X0Y116_A4;
  wire [0:0] CLBLL_L_X2Y116_SLICE_X0Y116_A5;
  wire [0:0] CLBLL_L_X2Y116_SLICE_X0Y116_A6;
  wire [0:0] CLBLL_L_X2Y116_SLICE_X0Y116_AO5;
  wire [0:0] CLBLL_L_X2Y116_SLICE_X0Y116_AO6;
  wire [0:0] CLBLL_L_X2Y116_SLICE_X0Y116_A_CY;
  wire [0:0] CLBLL_L_X2Y116_SLICE_X0Y116_A_XOR;
  wire [0:0] CLBLL_L_X2Y116_SLICE_X0Y116_B;
  wire [0:0] CLBLL_L_X2Y116_SLICE_X0Y116_B1;
  wire [0:0] CLBLL_L_X2Y116_SLICE_X0Y116_B2;
  wire [0:0] CLBLL_L_X2Y116_SLICE_X0Y116_B3;
  wire [0:0] CLBLL_L_X2Y116_SLICE_X0Y116_B4;
  wire [0:0] CLBLL_L_X2Y116_SLICE_X0Y116_B5;
  wire [0:0] CLBLL_L_X2Y116_SLICE_X0Y116_B6;
  wire [0:0] CLBLL_L_X2Y116_SLICE_X0Y116_BO5;
  wire [0:0] CLBLL_L_X2Y116_SLICE_X0Y116_BO6;
  wire [0:0] CLBLL_L_X2Y116_SLICE_X0Y116_B_CY;
  wire [0:0] CLBLL_L_X2Y116_SLICE_X0Y116_B_XOR;
  wire [0:0] CLBLL_L_X2Y116_SLICE_X0Y116_C;
  wire [0:0] CLBLL_L_X2Y116_SLICE_X0Y116_C1;
  wire [0:0] CLBLL_L_X2Y116_SLICE_X0Y116_C2;
  wire [0:0] CLBLL_L_X2Y116_SLICE_X0Y116_C3;
  wire [0:0] CLBLL_L_X2Y116_SLICE_X0Y116_C4;
  wire [0:0] CLBLL_L_X2Y116_SLICE_X0Y116_C5;
  wire [0:0] CLBLL_L_X2Y116_SLICE_X0Y116_C6;
  wire [0:0] CLBLL_L_X2Y116_SLICE_X0Y116_CO5;
  wire [0:0] CLBLL_L_X2Y116_SLICE_X0Y116_CO6;
  wire [0:0] CLBLL_L_X2Y116_SLICE_X0Y116_C_CY;
  wire [0:0] CLBLL_L_X2Y116_SLICE_X0Y116_C_XOR;
  wire [0:0] CLBLL_L_X2Y116_SLICE_X0Y116_D;
  wire [0:0] CLBLL_L_X2Y116_SLICE_X0Y116_D1;
  wire [0:0] CLBLL_L_X2Y116_SLICE_X0Y116_D2;
  wire [0:0] CLBLL_L_X2Y116_SLICE_X0Y116_D3;
  wire [0:0] CLBLL_L_X2Y116_SLICE_X0Y116_D4;
  wire [0:0] CLBLL_L_X2Y116_SLICE_X0Y116_D5;
  wire [0:0] CLBLL_L_X2Y116_SLICE_X0Y116_D6;
  wire [0:0] CLBLL_L_X2Y116_SLICE_X0Y116_DO5;
  wire [0:0] CLBLL_L_X2Y116_SLICE_X0Y116_DO6;
  wire [0:0] CLBLL_L_X2Y116_SLICE_X0Y116_D_CY;
  wire [0:0] CLBLL_L_X2Y116_SLICE_X0Y116_D_XOR;
  wire [0:0] CLBLL_L_X2Y116_SLICE_X1Y116_A;
  wire [0:0] CLBLL_L_X2Y116_SLICE_X1Y116_A1;
  wire [0:0] CLBLL_L_X2Y116_SLICE_X1Y116_A2;
  wire [0:0] CLBLL_L_X2Y116_SLICE_X1Y116_A3;
  wire [0:0] CLBLL_L_X2Y116_SLICE_X1Y116_A4;
  wire [0:0] CLBLL_L_X2Y116_SLICE_X1Y116_A5;
  wire [0:0] CLBLL_L_X2Y116_SLICE_X1Y116_A6;
  wire [0:0] CLBLL_L_X2Y116_SLICE_X1Y116_AO5;
  wire [0:0] CLBLL_L_X2Y116_SLICE_X1Y116_AO6;
  wire [0:0] CLBLL_L_X2Y116_SLICE_X1Y116_AQ;
  wire [0:0] CLBLL_L_X2Y116_SLICE_X1Y116_A_CY;
  wire [0:0] CLBLL_L_X2Y116_SLICE_X1Y116_A_XOR;
  wire [0:0] CLBLL_L_X2Y116_SLICE_X1Y116_B;
  wire [0:0] CLBLL_L_X2Y116_SLICE_X1Y116_B1;
  wire [0:0] CLBLL_L_X2Y116_SLICE_X1Y116_B2;
  wire [0:0] CLBLL_L_X2Y116_SLICE_X1Y116_B3;
  wire [0:0] CLBLL_L_X2Y116_SLICE_X1Y116_B4;
  wire [0:0] CLBLL_L_X2Y116_SLICE_X1Y116_B5;
  wire [0:0] CLBLL_L_X2Y116_SLICE_X1Y116_B6;
  wire [0:0] CLBLL_L_X2Y116_SLICE_X1Y116_BO5;
  wire [0:0] CLBLL_L_X2Y116_SLICE_X1Y116_BO6;
  wire [0:0] CLBLL_L_X2Y116_SLICE_X1Y116_B_CY;
  wire [0:0] CLBLL_L_X2Y116_SLICE_X1Y116_B_XOR;
  wire [0:0] CLBLL_L_X2Y116_SLICE_X1Y116_C;
  wire [0:0] CLBLL_L_X2Y116_SLICE_X1Y116_C1;
  wire [0:0] CLBLL_L_X2Y116_SLICE_X1Y116_C2;
  wire [0:0] CLBLL_L_X2Y116_SLICE_X1Y116_C3;
  wire [0:0] CLBLL_L_X2Y116_SLICE_X1Y116_C4;
  wire [0:0] CLBLL_L_X2Y116_SLICE_X1Y116_C5;
  wire [0:0] CLBLL_L_X2Y116_SLICE_X1Y116_C6;
  wire [0:0] CLBLL_L_X2Y116_SLICE_X1Y116_CLK;
  wire [0:0] CLBLL_L_X2Y116_SLICE_X1Y116_CO5;
  wire [0:0] CLBLL_L_X2Y116_SLICE_X1Y116_CO6;
  wire [0:0] CLBLL_L_X2Y116_SLICE_X1Y116_C_CY;
  wire [0:0] CLBLL_L_X2Y116_SLICE_X1Y116_C_XOR;
  wire [0:0] CLBLL_L_X2Y116_SLICE_X1Y116_D;
  wire [0:0] CLBLL_L_X2Y116_SLICE_X1Y116_D1;
  wire [0:0] CLBLL_L_X2Y116_SLICE_X1Y116_D2;
  wire [0:0] CLBLL_L_X2Y116_SLICE_X1Y116_D3;
  wire [0:0] CLBLL_L_X2Y116_SLICE_X1Y116_D4;
  wire [0:0] CLBLL_L_X2Y116_SLICE_X1Y116_D5;
  wire [0:0] CLBLL_L_X2Y116_SLICE_X1Y116_D6;
  wire [0:0] CLBLL_L_X2Y116_SLICE_X1Y116_DO5;
  wire [0:0] CLBLL_L_X2Y116_SLICE_X1Y116_DO6;
  wire [0:0] CLBLL_L_X2Y116_SLICE_X1Y116_D_CY;
  wire [0:0] CLBLL_L_X2Y116_SLICE_X1Y116_D_XOR;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X0Y117_A;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X0Y117_A1;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X0Y117_A2;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X0Y117_A3;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X0Y117_A4;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X0Y117_A5;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X0Y117_A5Q;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X0Y117_A6;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X0Y117_AMUX;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X0Y117_AO5;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X0Y117_AO6;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X0Y117_AQ;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X0Y117_AX;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X0Y117_A_CY;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X0Y117_A_XOR;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X0Y117_B;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X0Y117_B1;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X0Y117_B2;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X0Y117_B3;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X0Y117_B4;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X0Y117_B5;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X0Y117_B6;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X0Y117_BO5;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X0Y117_BO6;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X0Y117_BQ;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X0Y117_B_CY;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X0Y117_B_XOR;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X0Y117_C;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X0Y117_C1;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X0Y117_C2;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X0Y117_C3;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X0Y117_C4;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X0Y117_C5;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X0Y117_C6;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X0Y117_CLK;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X0Y117_CO5;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X0Y117_CO6;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X0Y117_CQ;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X0Y117_C_CY;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X0Y117_C_XOR;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X0Y117_D;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X0Y117_D1;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X0Y117_D2;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X0Y117_D3;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X0Y117_D4;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X0Y117_D5;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X0Y117_D6;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X0Y117_DMUX;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X0Y117_DO5;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X0Y117_DO6;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X0Y117_D_CY;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X0Y117_D_XOR;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X1Y117_A;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X1Y117_A1;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X1Y117_A2;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X1Y117_A3;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X1Y117_A4;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X1Y117_A5;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X1Y117_A6;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X1Y117_AO5;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X1Y117_AO6;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X1Y117_AQ;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X1Y117_A_CY;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X1Y117_A_XOR;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X1Y117_B;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X1Y117_B1;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X1Y117_B2;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X1Y117_B3;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X1Y117_B4;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X1Y117_B5;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X1Y117_B6;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X1Y117_BO5;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X1Y117_BO6;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X1Y117_BQ;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X1Y117_B_CY;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X1Y117_B_XOR;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X1Y117_C;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X1Y117_C1;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X1Y117_C2;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X1Y117_C3;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X1Y117_C4;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X1Y117_C5;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X1Y117_C6;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X1Y117_CLK;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X1Y117_CMUX;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X1Y117_CO5;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X1Y117_CO6;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X1Y117_C_CY;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X1Y117_C_XOR;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X1Y117_D;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X1Y117_D1;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X1Y117_D2;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X1Y117_D3;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X1Y117_D4;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X1Y117_D5;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X1Y117_D6;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X1Y117_DO5;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X1Y117_DO6;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X1Y117_D_CY;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X1Y117_D_XOR;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X0Y118_A;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X0Y118_A1;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X0Y118_A2;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X0Y118_A3;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X0Y118_A4;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X0Y118_A5;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X0Y118_A6;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X0Y118_AO5;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X0Y118_AO6;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X0Y118_A_CY;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X0Y118_A_XOR;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X0Y118_B;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X0Y118_B1;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X0Y118_B2;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X0Y118_B3;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X0Y118_B4;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X0Y118_B5;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X0Y118_B6;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X0Y118_BO5;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X0Y118_BO6;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X0Y118_B_CY;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X0Y118_B_XOR;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X0Y118_C;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X0Y118_C1;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X0Y118_C2;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X0Y118_C3;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X0Y118_C4;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X0Y118_C5;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X0Y118_C6;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X0Y118_CO5;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X0Y118_CO6;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X0Y118_C_CY;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X0Y118_C_XOR;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X0Y118_D;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X0Y118_D1;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X0Y118_D2;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X0Y118_D3;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X0Y118_D4;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X0Y118_D5;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X0Y118_D6;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X0Y118_DO5;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X0Y118_DO6;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X0Y118_D_CY;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X0Y118_D_XOR;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X1Y118_A;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X1Y118_A1;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X1Y118_A2;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X1Y118_A3;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X1Y118_A4;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X1Y118_A5;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X1Y118_A6;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X1Y118_AO5;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X1Y118_AO6;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X1Y118_A_CY;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X1Y118_A_XOR;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X1Y118_B;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X1Y118_B1;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X1Y118_B2;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X1Y118_B3;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X1Y118_B4;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X1Y118_B5;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X1Y118_B6;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X1Y118_BO5;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X1Y118_BO6;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X1Y118_B_CY;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X1Y118_B_XOR;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X1Y118_C;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X1Y118_C1;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X1Y118_C2;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X1Y118_C3;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X1Y118_C4;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X1Y118_C5;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X1Y118_C6;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X1Y118_CO5;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X1Y118_CO6;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X1Y118_C_CY;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X1Y118_C_XOR;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X1Y118_D;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X1Y118_D1;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X1Y118_D2;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X1Y118_D3;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X1Y118_D4;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X1Y118_D5;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X1Y118_D6;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X1Y118_DO5;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X1Y118_DO6;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X1Y118_D_CY;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X1Y118_D_XOR;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X0Y119_A;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X0Y119_A1;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X0Y119_A2;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X0Y119_A3;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X0Y119_A4;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X0Y119_A5;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X0Y119_A6;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X0Y119_AO5;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X0Y119_AO6;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X0Y119_A_CY;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X0Y119_A_XOR;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X0Y119_B;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X0Y119_B1;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X0Y119_B2;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X0Y119_B3;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X0Y119_B4;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X0Y119_B5;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X0Y119_B6;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X0Y119_BO5;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X0Y119_BO6;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X0Y119_B_CY;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X0Y119_B_XOR;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X0Y119_C;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X0Y119_C1;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X0Y119_C2;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X0Y119_C3;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X0Y119_C4;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X0Y119_C5;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X0Y119_C6;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X0Y119_CO5;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X0Y119_CO6;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X0Y119_C_CY;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X0Y119_C_XOR;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X0Y119_D;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X0Y119_D1;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X0Y119_D2;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X0Y119_D3;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X0Y119_D4;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X0Y119_D5;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X0Y119_D6;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X0Y119_DO5;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X0Y119_DO6;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X0Y119_D_CY;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X0Y119_D_XOR;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X1Y119_A;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X1Y119_A1;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X1Y119_A2;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X1Y119_A3;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X1Y119_A4;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X1Y119_A5;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X1Y119_A6;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X1Y119_AMUX;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X1Y119_AO5;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X1Y119_AO6;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X1Y119_A_CY;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X1Y119_A_XOR;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X1Y119_B;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X1Y119_B1;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X1Y119_B2;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X1Y119_B3;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X1Y119_B4;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X1Y119_B5;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X1Y119_B6;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X1Y119_BO5;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X1Y119_BO6;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X1Y119_B_CY;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X1Y119_B_XOR;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X1Y119_C;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X1Y119_C1;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X1Y119_C2;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X1Y119_C3;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X1Y119_C4;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X1Y119_C5;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X1Y119_C6;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X1Y119_CO5;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X1Y119_CO6;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X1Y119_C_CY;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X1Y119_C_XOR;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X1Y119_D;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X1Y119_D1;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X1Y119_D2;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X1Y119_D3;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X1Y119_D4;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X1Y119_D5;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X1Y119_D6;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X1Y119_DO5;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X1Y119_DO6;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X1Y119_D_CY;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X1Y119_D_XOR;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X0Y120_A;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X0Y120_A1;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X0Y120_A2;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X0Y120_A3;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X0Y120_A4;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X0Y120_A5;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X0Y120_A6;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X0Y120_AMUX;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X0Y120_AO5;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X0Y120_AO6;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X0Y120_A_CY;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X0Y120_A_XOR;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X0Y120_B;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X0Y120_B1;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X0Y120_B2;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X0Y120_B3;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X0Y120_B4;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X0Y120_B5;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X0Y120_B6;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X0Y120_BO5;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X0Y120_BO6;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X0Y120_B_CY;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X0Y120_B_XOR;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X0Y120_C;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X0Y120_C1;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X0Y120_C2;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X0Y120_C3;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X0Y120_C4;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X0Y120_C5;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X0Y120_C6;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X0Y120_CO5;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X0Y120_CO6;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X0Y120_C_CY;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X0Y120_C_XOR;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X0Y120_D;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X0Y120_D1;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X0Y120_D2;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X0Y120_D3;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X0Y120_D4;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X0Y120_D5;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X0Y120_D6;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X0Y120_DO5;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X0Y120_DO6;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X0Y120_D_CY;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X0Y120_D_XOR;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X1Y120_A;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X1Y120_A1;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X1Y120_A2;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X1Y120_A3;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X1Y120_A4;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X1Y120_A5;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X1Y120_A6;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X1Y120_AMUX;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X1Y120_AO5;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X1Y120_AO6;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X1Y120_A_CY;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X1Y120_A_XOR;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X1Y120_B;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X1Y120_B1;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X1Y120_B2;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X1Y120_B3;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X1Y120_B4;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X1Y120_B5;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X1Y120_B6;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X1Y120_BO5;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X1Y120_BO6;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X1Y120_B_CY;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X1Y120_B_XOR;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X1Y120_C;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X1Y120_C1;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X1Y120_C2;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X1Y120_C3;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X1Y120_C4;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X1Y120_C5;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X1Y120_C6;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X1Y120_CMUX;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X1Y120_CO5;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X1Y120_CO6;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X1Y120_C_CY;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X1Y120_C_XOR;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X1Y120_D;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X1Y120_D1;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X1Y120_D2;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X1Y120_D3;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X1Y120_D4;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X1Y120_D5;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X1Y120_D6;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X1Y120_DO5;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X1Y120_DO6;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X1Y120_D_CY;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X1Y120_D_XOR;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X0Y121_A;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X0Y121_A1;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X0Y121_A2;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X0Y121_A3;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X0Y121_A4;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X0Y121_A5;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X0Y121_A6;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X0Y121_AMUX;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X0Y121_AO5;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X0Y121_AO6;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X0Y121_A_CY;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X0Y121_A_XOR;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X0Y121_B;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X0Y121_B1;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X0Y121_B2;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X0Y121_B3;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X0Y121_B4;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X0Y121_B5;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X0Y121_B6;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X0Y121_BMUX;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X0Y121_BO5;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X0Y121_BO6;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X0Y121_B_CY;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X0Y121_B_XOR;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X0Y121_C;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X0Y121_C1;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X0Y121_C2;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X0Y121_C3;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X0Y121_C4;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X0Y121_C5;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X0Y121_C6;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X0Y121_CO5;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X0Y121_CO6;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X0Y121_C_CY;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X0Y121_C_XOR;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X0Y121_D;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X0Y121_D1;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X0Y121_D2;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X0Y121_D3;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X0Y121_D4;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X0Y121_D5;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X0Y121_D6;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X0Y121_DO5;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X0Y121_DO6;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X0Y121_D_CY;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X0Y121_D_XOR;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X1Y121_A;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X1Y121_A1;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X1Y121_A2;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X1Y121_A3;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X1Y121_A4;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X1Y121_A5;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X1Y121_A6;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X1Y121_AMUX;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X1Y121_AO5;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X1Y121_AO6;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X1Y121_A_CY;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X1Y121_A_XOR;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X1Y121_B;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X1Y121_B1;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X1Y121_B2;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X1Y121_B3;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X1Y121_B4;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X1Y121_B5;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X1Y121_B6;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X1Y121_BMUX;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X1Y121_BO5;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X1Y121_BO6;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X1Y121_B_CY;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X1Y121_B_XOR;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X1Y121_C;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X1Y121_C1;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X1Y121_C2;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X1Y121_C3;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X1Y121_C4;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X1Y121_C5;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X1Y121_C6;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X1Y121_CO5;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X1Y121_CO6;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X1Y121_C_CY;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X1Y121_C_XOR;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X1Y121_D;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X1Y121_D1;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X1Y121_D2;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X1Y121_D3;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X1Y121_D4;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X1Y121_D5;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X1Y121_D6;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X1Y121_DO5;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X1Y121_DO6;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X1Y121_D_CY;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X1Y121_D_XOR;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X0Y122_A;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X0Y122_A1;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X0Y122_A2;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X0Y122_A3;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X0Y122_A4;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X0Y122_A5;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X0Y122_A6;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X0Y122_AMUX;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X0Y122_AO5;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X0Y122_AO6;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X0Y122_A_CY;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X0Y122_A_XOR;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X0Y122_B;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X0Y122_B1;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X0Y122_B2;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X0Y122_B3;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X0Y122_B4;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X0Y122_B5;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X0Y122_B6;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X0Y122_BO5;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X0Y122_BO6;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X0Y122_B_CY;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X0Y122_B_XOR;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X0Y122_C;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X0Y122_C1;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X0Y122_C2;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X0Y122_C3;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X0Y122_C4;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X0Y122_C5;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X0Y122_C6;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X0Y122_CO5;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X0Y122_CO6;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X0Y122_C_CY;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X0Y122_C_XOR;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X0Y122_D;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X0Y122_D1;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X0Y122_D2;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X0Y122_D3;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X0Y122_D4;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X0Y122_D5;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X0Y122_D6;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X0Y122_DO5;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X0Y122_DO6;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X0Y122_D_CY;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X0Y122_D_XOR;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X1Y122_A;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X1Y122_A1;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X1Y122_A2;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X1Y122_A3;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X1Y122_A4;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X1Y122_A5;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X1Y122_A6;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X1Y122_AO5;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X1Y122_AO6;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X1Y122_A_CY;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X1Y122_A_XOR;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X1Y122_B;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X1Y122_B1;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X1Y122_B2;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X1Y122_B3;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X1Y122_B4;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X1Y122_B5;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X1Y122_B6;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X1Y122_BMUX;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X1Y122_BO5;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X1Y122_BO6;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X1Y122_B_CY;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X1Y122_B_XOR;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X1Y122_C;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X1Y122_C1;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X1Y122_C2;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X1Y122_C3;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X1Y122_C4;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X1Y122_C5;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X1Y122_C6;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X1Y122_CO5;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X1Y122_CO6;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X1Y122_C_CY;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X1Y122_C_XOR;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X1Y122_D;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X1Y122_D1;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X1Y122_D2;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X1Y122_D3;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X1Y122_D4;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X1Y122_D5;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X1Y122_D6;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X1Y122_DO5;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X1Y122_DO6;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X1Y122_D_CY;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X1Y122_D_XOR;
  wire [0:0] CLBLL_L_X2Y123_SLICE_X0Y123_A;
  wire [0:0] CLBLL_L_X2Y123_SLICE_X0Y123_A1;
  wire [0:0] CLBLL_L_X2Y123_SLICE_X0Y123_A2;
  wire [0:0] CLBLL_L_X2Y123_SLICE_X0Y123_A3;
  wire [0:0] CLBLL_L_X2Y123_SLICE_X0Y123_A4;
  wire [0:0] CLBLL_L_X2Y123_SLICE_X0Y123_A5;
  wire [0:0] CLBLL_L_X2Y123_SLICE_X0Y123_A6;
  wire [0:0] CLBLL_L_X2Y123_SLICE_X0Y123_AO5;
  wire [0:0] CLBLL_L_X2Y123_SLICE_X0Y123_AO6;
  wire [0:0] CLBLL_L_X2Y123_SLICE_X0Y123_A_CY;
  wire [0:0] CLBLL_L_X2Y123_SLICE_X0Y123_A_XOR;
  wire [0:0] CLBLL_L_X2Y123_SLICE_X0Y123_B;
  wire [0:0] CLBLL_L_X2Y123_SLICE_X0Y123_B1;
  wire [0:0] CLBLL_L_X2Y123_SLICE_X0Y123_B2;
  wire [0:0] CLBLL_L_X2Y123_SLICE_X0Y123_B3;
  wire [0:0] CLBLL_L_X2Y123_SLICE_X0Y123_B4;
  wire [0:0] CLBLL_L_X2Y123_SLICE_X0Y123_B5;
  wire [0:0] CLBLL_L_X2Y123_SLICE_X0Y123_B6;
  wire [0:0] CLBLL_L_X2Y123_SLICE_X0Y123_BO5;
  wire [0:0] CLBLL_L_X2Y123_SLICE_X0Y123_BO6;
  wire [0:0] CLBLL_L_X2Y123_SLICE_X0Y123_B_CY;
  wire [0:0] CLBLL_L_X2Y123_SLICE_X0Y123_B_XOR;
  wire [0:0] CLBLL_L_X2Y123_SLICE_X0Y123_C;
  wire [0:0] CLBLL_L_X2Y123_SLICE_X0Y123_C1;
  wire [0:0] CLBLL_L_X2Y123_SLICE_X0Y123_C2;
  wire [0:0] CLBLL_L_X2Y123_SLICE_X0Y123_C3;
  wire [0:0] CLBLL_L_X2Y123_SLICE_X0Y123_C4;
  wire [0:0] CLBLL_L_X2Y123_SLICE_X0Y123_C5;
  wire [0:0] CLBLL_L_X2Y123_SLICE_X0Y123_C6;
  wire [0:0] CLBLL_L_X2Y123_SLICE_X0Y123_CO5;
  wire [0:0] CLBLL_L_X2Y123_SLICE_X0Y123_CO6;
  wire [0:0] CLBLL_L_X2Y123_SLICE_X0Y123_C_CY;
  wire [0:0] CLBLL_L_X2Y123_SLICE_X0Y123_C_XOR;
  wire [0:0] CLBLL_L_X2Y123_SLICE_X0Y123_D;
  wire [0:0] CLBLL_L_X2Y123_SLICE_X0Y123_D1;
  wire [0:0] CLBLL_L_X2Y123_SLICE_X0Y123_D2;
  wire [0:0] CLBLL_L_X2Y123_SLICE_X0Y123_D3;
  wire [0:0] CLBLL_L_X2Y123_SLICE_X0Y123_D4;
  wire [0:0] CLBLL_L_X2Y123_SLICE_X0Y123_D5;
  wire [0:0] CLBLL_L_X2Y123_SLICE_X0Y123_D6;
  wire [0:0] CLBLL_L_X2Y123_SLICE_X0Y123_DO5;
  wire [0:0] CLBLL_L_X2Y123_SLICE_X0Y123_DO6;
  wire [0:0] CLBLL_L_X2Y123_SLICE_X0Y123_D_CY;
  wire [0:0] CLBLL_L_X2Y123_SLICE_X0Y123_D_XOR;
  wire [0:0] CLBLL_L_X2Y123_SLICE_X1Y123_A;
  wire [0:0] CLBLL_L_X2Y123_SLICE_X1Y123_A1;
  wire [0:0] CLBLL_L_X2Y123_SLICE_X1Y123_A2;
  wire [0:0] CLBLL_L_X2Y123_SLICE_X1Y123_A3;
  wire [0:0] CLBLL_L_X2Y123_SLICE_X1Y123_A4;
  wire [0:0] CLBLL_L_X2Y123_SLICE_X1Y123_A5;
  wire [0:0] CLBLL_L_X2Y123_SLICE_X1Y123_A6;
  wire [0:0] CLBLL_L_X2Y123_SLICE_X1Y123_AO5;
  wire [0:0] CLBLL_L_X2Y123_SLICE_X1Y123_AO6;
  wire [0:0] CLBLL_L_X2Y123_SLICE_X1Y123_A_CY;
  wire [0:0] CLBLL_L_X2Y123_SLICE_X1Y123_A_XOR;
  wire [0:0] CLBLL_L_X2Y123_SLICE_X1Y123_B;
  wire [0:0] CLBLL_L_X2Y123_SLICE_X1Y123_B1;
  wire [0:0] CLBLL_L_X2Y123_SLICE_X1Y123_B2;
  wire [0:0] CLBLL_L_X2Y123_SLICE_X1Y123_B3;
  wire [0:0] CLBLL_L_X2Y123_SLICE_X1Y123_B4;
  wire [0:0] CLBLL_L_X2Y123_SLICE_X1Y123_B5;
  wire [0:0] CLBLL_L_X2Y123_SLICE_X1Y123_B6;
  wire [0:0] CLBLL_L_X2Y123_SLICE_X1Y123_BO5;
  wire [0:0] CLBLL_L_X2Y123_SLICE_X1Y123_BO6;
  wire [0:0] CLBLL_L_X2Y123_SLICE_X1Y123_B_CY;
  wire [0:0] CLBLL_L_X2Y123_SLICE_X1Y123_B_XOR;
  wire [0:0] CLBLL_L_X2Y123_SLICE_X1Y123_C;
  wire [0:0] CLBLL_L_X2Y123_SLICE_X1Y123_C1;
  wire [0:0] CLBLL_L_X2Y123_SLICE_X1Y123_C2;
  wire [0:0] CLBLL_L_X2Y123_SLICE_X1Y123_C3;
  wire [0:0] CLBLL_L_X2Y123_SLICE_X1Y123_C4;
  wire [0:0] CLBLL_L_X2Y123_SLICE_X1Y123_C5;
  wire [0:0] CLBLL_L_X2Y123_SLICE_X1Y123_C6;
  wire [0:0] CLBLL_L_X2Y123_SLICE_X1Y123_CO5;
  wire [0:0] CLBLL_L_X2Y123_SLICE_X1Y123_CO6;
  wire [0:0] CLBLL_L_X2Y123_SLICE_X1Y123_C_CY;
  wire [0:0] CLBLL_L_X2Y123_SLICE_X1Y123_C_XOR;
  wire [0:0] CLBLL_L_X2Y123_SLICE_X1Y123_D;
  wire [0:0] CLBLL_L_X2Y123_SLICE_X1Y123_D1;
  wire [0:0] CLBLL_L_X2Y123_SLICE_X1Y123_D2;
  wire [0:0] CLBLL_L_X2Y123_SLICE_X1Y123_D3;
  wire [0:0] CLBLL_L_X2Y123_SLICE_X1Y123_D4;
  wire [0:0] CLBLL_L_X2Y123_SLICE_X1Y123_D5;
  wire [0:0] CLBLL_L_X2Y123_SLICE_X1Y123_D6;
  wire [0:0] CLBLL_L_X2Y123_SLICE_X1Y123_DO5;
  wire [0:0] CLBLL_L_X2Y123_SLICE_X1Y123_DO6;
  wire [0:0] CLBLL_L_X2Y123_SLICE_X1Y123_D_CY;
  wire [0:0] CLBLL_L_X2Y123_SLICE_X1Y123_D_XOR;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X4Y110_A;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X4Y110_A1;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X4Y110_A2;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X4Y110_A3;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X4Y110_A4;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X4Y110_A5;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X4Y110_A5Q;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X4Y110_A6;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X4Y110_AMUX;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X4Y110_AO5;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X4Y110_AO6;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X4Y110_AQ;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X4Y110_AX;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X4Y110_A_CY;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X4Y110_A_XOR;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X4Y110_B;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X4Y110_B1;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X4Y110_B2;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X4Y110_B3;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X4Y110_B4;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X4Y110_B5;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X4Y110_B6;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X4Y110_BMUX;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X4Y110_BO5;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X4Y110_BO6;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X4Y110_B_CY;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X4Y110_B_XOR;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X4Y110_C;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X4Y110_C1;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X4Y110_C2;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X4Y110_C3;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X4Y110_C4;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X4Y110_C5;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X4Y110_C6;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X4Y110_CLK;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X4Y110_CO5;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X4Y110_CO6;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X4Y110_CQ;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X4Y110_C_CY;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X4Y110_C_XOR;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X4Y110_D;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X4Y110_D1;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X4Y110_D2;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X4Y110_D3;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X4Y110_D4;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X4Y110_D5;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X4Y110_D6;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X4Y110_DO5;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X4Y110_DO6;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X4Y110_DQ;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X4Y110_D_CY;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X4Y110_D_XOR;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X5Y110_A;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X5Y110_A1;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X5Y110_A2;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X5Y110_A3;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X5Y110_A4;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X5Y110_A5;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X5Y110_A6;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X5Y110_AO5;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X5Y110_AO6;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X5Y110_AQ;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X5Y110_A_CY;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X5Y110_A_XOR;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X5Y110_B;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X5Y110_B1;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X5Y110_B2;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X5Y110_B3;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X5Y110_B4;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X5Y110_B5;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X5Y110_B6;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X5Y110_BO5;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X5Y110_BO6;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X5Y110_BQ;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X5Y110_B_CY;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X5Y110_B_XOR;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X5Y110_C;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X5Y110_C1;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X5Y110_C2;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X5Y110_C3;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X5Y110_C4;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X5Y110_C5;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X5Y110_C6;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X5Y110_CLK;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X5Y110_CMUX;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X5Y110_CO5;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X5Y110_CO6;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X5Y110_C_CY;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X5Y110_C_XOR;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X5Y110_D;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X5Y110_D1;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X5Y110_D2;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X5Y110_D3;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X5Y110_D4;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X5Y110_D5;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X5Y110_D6;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X5Y110_DO5;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X5Y110_DO6;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X5Y110_D_CY;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X5Y110_D_XOR;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X4Y111_A;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X4Y111_A1;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X4Y111_A2;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X4Y111_A3;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X4Y111_A4;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X4Y111_A5;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X4Y111_A6;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X4Y111_AMUX;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X4Y111_AO5;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X4Y111_AO6;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X4Y111_AQ;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X4Y111_A_CY;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X4Y111_A_XOR;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X4Y111_B;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X4Y111_B1;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X4Y111_B2;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X4Y111_B3;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X4Y111_B4;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X4Y111_B5;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X4Y111_B6;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X4Y111_BO5;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X4Y111_BO6;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X4Y111_BQ;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X4Y111_B_CY;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X4Y111_B_XOR;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X4Y111_C;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X4Y111_C1;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X4Y111_C2;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X4Y111_C3;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X4Y111_C4;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X4Y111_C5;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X4Y111_C6;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X4Y111_CLK;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X4Y111_CO5;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X4Y111_CO6;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X4Y111_CQ;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X4Y111_C_CY;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X4Y111_C_XOR;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X4Y111_D;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X4Y111_D1;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X4Y111_D2;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X4Y111_D3;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X4Y111_D4;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X4Y111_D5;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X4Y111_D6;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X4Y111_DO5;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X4Y111_DO6;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X4Y111_DQ;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X4Y111_D_CY;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X4Y111_D_XOR;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X5Y111_A;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X5Y111_A1;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X5Y111_A2;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X5Y111_A3;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X5Y111_A4;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X5Y111_A5;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X5Y111_A5Q;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X5Y111_A6;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X5Y111_AMUX;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X5Y111_AO5;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X5Y111_AO6;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X5Y111_AQ;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X5Y111_AX;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X5Y111_A_CY;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X5Y111_A_XOR;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X5Y111_B;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X5Y111_B1;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X5Y111_B2;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X5Y111_B3;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X5Y111_B4;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X5Y111_B5;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X5Y111_B6;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X5Y111_BO5;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X5Y111_BO6;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X5Y111_BQ;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X5Y111_B_CY;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X5Y111_B_XOR;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X5Y111_C;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X5Y111_C1;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X5Y111_C2;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X5Y111_C3;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X5Y111_C4;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X5Y111_C5;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X5Y111_C6;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X5Y111_CLK;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X5Y111_CO5;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X5Y111_CO6;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X5Y111_C_CY;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X5Y111_C_XOR;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X5Y111_D;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X5Y111_D1;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X5Y111_D2;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X5Y111_D3;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X5Y111_D4;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X5Y111_D5;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X5Y111_D6;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X5Y111_DMUX;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X5Y111_DO5;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X5Y111_DO6;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X5Y111_D_CY;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X5Y111_D_XOR;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X4Y112_A;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X4Y112_A1;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X4Y112_A2;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X4Y112_A3;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X4Y112_A4;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X4Y112_A5;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X4Y112_A6;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X4Y112_AO5;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X4Y112_AO6;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X4Y112_AQ;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X4Y112_A_CY;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X4Y112_A_XOR;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X4Y112_B;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X4Y112_B1;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X4Y112_B2;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X4Y112_B3;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X4Y112_B4;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X4Y112_B5;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X4Y112_B6;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X4Y112_BO5;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X4Y112_BO6;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X4Y112_BQ;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X4Y112_B_CY;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X4Y112_B_XOR;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X4Y112_C;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X4Y112_C1;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X4Y112_C2;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X4Y112_C3;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X4Y112_C4;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X4Y112_C5;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X4Y112_C6;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X4Y112_CLK;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X4Y112_CO5;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X4Y112_CO6;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X4Y112_C_CY;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X4Y112_C_XOR;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X4Y112_D;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X4Y112_D1;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X4Y112_D2;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X4Y112_D3;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X4Y112_D4;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X4Y112_D5;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X4Y112_D6;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X4Y112_DO5;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X4Y112_DO6;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X4Y112_D_CY;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X4Y112_D_XOR;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X5Y112_A;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X5Y112_A1;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X5Y112_A2;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X5Y112_A3;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X5Y112_A4;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X5Y112_A5;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X5Y112_A6;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X5Y112_AO5;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X5Y112_AO6;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X5Y112_AQ;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X5Y112_A_CY;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X5Y112_A_XOR;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X5Y112_B;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X5Y112_B1;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X5Y112_B2;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X5Y112_B3;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X5Y112_B4;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X5Y112_B5;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X5Y112_B6;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X5Y112_BO5;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X5Y112_BO6;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X5Y112_B_CY;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X5Y112_B_XOR;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X5Y112_C;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X5Y112_C1;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X5Y112_C2;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X5Y112_C3;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X5Y112_C4;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X5Y112_C5;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X5Y112_C6;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X5Y112_CLK;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X5Y112_CO5;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X5Y112_CO6;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X5Y112_C_CY;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X5Y112_C_XOR;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X5Y112_D;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X5Y112_D1;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X5Y112_D2;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X5Y112_D3;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X5Y112_D4;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X5Y112_D5;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X5Y112_D6;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X5Y112_DMUX;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X5Y112_DO5;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X5Y112_DO6;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X5Y112_D_CY;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X5Y112_D_XOR;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_A;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_A1;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_A2;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_A3;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_A4;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_A5;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_A6;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_AO5;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_AO6;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_AQ;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_A_CY;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_A_XOR;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_B;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_B1;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_B2;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_B3;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_B4;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_B5;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_B6;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_BO5;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_BO6;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_BQ;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_B_CY;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_B_XOR;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_C;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_C1;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_C2;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_C3;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_C4;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_C5;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_C6;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_CLK;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_CO5;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_CO6;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_C_CY;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_C_XOR;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_D;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_D1;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_D2;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_D3;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_D4;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_D5;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_D6;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_DO5;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_DO6;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_D_CY;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_D_XOR;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_A;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_A1;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_A2;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_A3;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_A4;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_A5;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_A6;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_AO5;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_AO6;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_AQ;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_A_CY;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_A_XOR;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_B;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_B1;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_B2;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_B3;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_B4;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_B5;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_B6;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_BO5;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_BO6;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_BQ;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_B_CY;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_B_XOR;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_C;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_C1;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_C2;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_C3;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_C4;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_C5;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_C6;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_CLK;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_CO5;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_CO6;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_CQ;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_C_CY;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_C_XOR;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_D;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_D1;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_D2;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_D3;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_D4;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_D5;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_D6;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_DMUX;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_DO5;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_DO6;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_D_CY;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_D_XOR;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X4Y114_A;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X4Y114_A1;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X4Y114_A2;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X4Y114_A3;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X4Y114_A4;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X4Y114_A5;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X4Y114_A6;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X4Y114_AO5;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X4Y114_AO6;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X4Y114_AQ;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X4Y114_A_CY;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X4Y114_A_XOR;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X4Y114_B;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X4Y114_B1;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X4Y114_B2;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X4Y114_B3;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X4Y114_B4;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X4Y114_B5;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X4Y114_B6;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X4Y114_BO5;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X4Y114_BO6;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X4Y114_BQ;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X4Y114_B_CY;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X4Y114_B_XOR;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X4Y114_C;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X4Y114_C1;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X4Y114_C2;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X4Y114_C3;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X4Y114_C4;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X4Y114_C5;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X4Y114_C6;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X4Y114_CLK;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X4Y114_CO5;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X4Y114_CO6;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X4Y114_CQ;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X4Y114_C_CY;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X4Y114_C_XOR;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X4Y114_D;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X4Y114_D1;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X4Y114_D2;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X4Y114_D3;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X4Y114_D4;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X4Y114_D5;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X4Y114_D6;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X4Y114_DO5;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X4Y114_DO6;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X4Y114_D_CY;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X4Y114_D_XOR;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X5Y114_A;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X5Y114_A1;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X5Y114_A2;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X5Y114_A3;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X5Y114_A4;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X5Y114_A5;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X5Y114_A6;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X5Y114_AO5;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X5Y114_AO6;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X5Y114_AQ;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X5Y114_A_CY;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X5Y114_A_XOR;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X5Y114_B;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X5Y114_B1;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X5Y114_B2;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X5Y114_B3;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X5Y114_B4;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X5Y114_B5;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X5Y114_B6;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X5Y114_BMUX;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X5Y114_BO5;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X5Y114_BO6;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X5Y114_B_CY;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X5Y114_B_XOR;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X5Y114_C;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X5Y114_C1;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X5Y114_C2;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X5Y114_C3;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X5Y114_C4;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X5Y114_C5;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X5Y114_C6;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X5Y114_CLK;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X5Y114_CMUX;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X5Y114_CO5;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X5Y114_CO6;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X5Y114_C_CY;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X5Y114_C_XOR;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X5Y114_D;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X5Y114_D1;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X5Y114_D2;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X5Y114_D3;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X5Y114_D4;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X5Y114_D5;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X5Y114_D6;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X5Y114_DO5;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X5Y114_DO6;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X5Y114_D_CY;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X5Y114_D_XOR;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X4Y115_A;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X4Y115_A1;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X4Y115_A2;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X4Y115_A3;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X4Y115_A4;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X4Y115_A5;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X4Y115_A6;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X4Y115_AO5;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X4Y115_AO6;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X4Y115_AQ;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X4Y115_A_CY;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X4Y115_A_XOR;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X4Y115_B;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X4Y115_B1;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X4Y115_B2;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X4Y115_B3;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X4Y115_B4;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X4Y115_B5;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X4Y115_B6;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X4Y115_BO5;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X4Y115_BO6;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X4Y115_BQ;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X4Y115_B_CY;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X4Y115_B_XOR;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X4Y115_C;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X4Y115_C1;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X4Y115_C2;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X4Y115_C3;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X4Y115_C4;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X4Y115_C5;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X4Y115_C5Q;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X4Y115_C6;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X4Y115_CLK;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X4Y115_CMUX;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X4Y115_CO5;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X4Y115_CO6;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X4Y115_CQ;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X4Y115_C_CY;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X4Y115_C_XOR;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X4Y115_D;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X4Y115_D1;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X4Y115_D2;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X4Y115_D3;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X4Y115_D4;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X4Y115_D5;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X4Y115_D6;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X4Y115_DO5;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X4Y115_DO6;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X4Y115_DQ;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X4Y115_D_CY;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X4Y115_D_XOR;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X5Y115_A;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X5Y115_A1;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X5Y115_A2;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X5Y115_A3;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X5Y115_A4;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X5Y115_A5;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X5Y115_A6;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X5Y115_AO5;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X5Y115_AO6;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X5Y115_AQ;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X5Y115_A_CY;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X5Y115_A_XOR;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X5Y115_B;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X5Y115_B1;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X5Y115_B2;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X5Y115_B3;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X5Y115_B4;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X5Y115_B5;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X5Y115_B6;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X5Y115_BO5;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X5Y115_BO6;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X5Y115_BQ;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X5Y115_B_CY;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X5Y115_B_XOR;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X5Y115_C;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X5Y115_C1;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X5Y115_C2;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X5Y115_C3;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X5Y115_C4;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X5Y115_C5;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X5Y115_C6;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X5Y115_CLK;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X5Y115_CO5;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X5Y115_CO6;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X5Y115_CQ;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X5Y115_C_CY;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X5Y115_C_XOR;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X5Y115_D;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X5Y115_D1;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X5Y115_D2;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X5Y115_D3;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X5Y115_D4;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X5Y115_D5;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X5Y115_D6;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X5Y115_DO5;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X5Y115_DO6;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X5Y115_DQ;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X5Y115_D_CY;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X5Y115_D_XOR;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X4Y116_A;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X4Y116_A1;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X4Y116_A2;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X4Y116_A3;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X4Y116_A4;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X4Y116_A5;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X4Y116_A6;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X4Y116_AO5;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X4Y116_AO6;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X4Y116_AQ;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X4Y116_A_CY;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X4Y116_A_XOR;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X4Y116_B;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X4Y116_B1;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X4Y116_B2;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X4Y116_B3;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X4Y116_B4;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X4Y116_B5;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X4Y116_B6;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X4Y116_BO5;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X4Y116_BO6;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X4Y116_BQ;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X4Y116_B_CY;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X4Y116_B_XOR;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X4Y116_C;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X4Y116_C1;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X4Y116_C2;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X4Y116_C3;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X4Y116_C4;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X4Y116_C5;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X4Y116_C5Q;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X4Y116_C6;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X4Y116_CLK;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X4Y116_CMUX;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X4Y116_CO5;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X4Y116_CO6;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X4Y116_CQ;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X4Y116_C_CY;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X4Y116_C_XOR;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X4Y116_D;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X4Y116_D1;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X4Y116_D2;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X4Y116_D3;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X4Y116_D4;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X4Y116_D5;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X4Y116_D6;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X4Y116_DO5;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X4Y116_DO6;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X4Y116_DQ;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X4Y116_D_CY;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X4Y116_D_XOR;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X5Y116_A;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X5Y116_A1;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X5Y116_A2;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X5Y116_A3;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X5Y116_A4;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X5Y116_A5;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X5Y116_A5Q;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X5Y116_A6;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X5Y116_AMUX;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X5Y116_AO5;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X5Y116_AO6;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X5Y116_AQ;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X5Y116_AX;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X5Y116_A_CY;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X5Y116_A_XOR;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X5Y116_B;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X5Y116_B1;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X5Y116_B2;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X5Y116_B3;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X5Y116_B4;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X5Y116_B5;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X5Y116_B6;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X5Y116_BO5;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X5Y116_BO6;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X5Y116_BQ;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X5Y116_B_CY;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X5Y116_B_XOR;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X5Y116_C;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X5Y116_C1;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X5Y116_C2;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X5Y116_C3;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X5Y116_C4;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X5Y116_C5;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X5Y116_C6;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X5Y116_CLK;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X5Y116_CMUX;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X5Y116_CO5;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X5Y116_CO6;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X5Y116_C_CY;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X5Y116_C_XOR;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X5Y116_D;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X5Y116_D1;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X5Y116_D2;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X5Y116_D3;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X5Y116_D4;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X5Y116_D5;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X5Y116_D6;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X5Y116_DO5;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X5Y116_DO6;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X5Y116_DQ;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X5Y116_D_CY;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X5Y116_D_XOR;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X4Y117_A;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X4Y117_A1;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X4Y117_A2;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X4Y117_A3;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X4Y117_A4;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X4Y117_A5;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X4Y117_A6;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X4Y117_AO5;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X4Y117_AO6;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X4Y117_AQ;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X4Y117_A_CY;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X4Y117_A_XOR;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X4Y117_B;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X4Y117_B1;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X4Y117_B2;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X4Y117_B3;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X4Y117_B4;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X4Y117_B5;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X4Y117_B6;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X4Y117_BO5;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X4Y117_BO6;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X4Y117_BQ;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X4Y117_B_CY;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X4Y117_B_XOR;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X4Y117_C;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X4Y117_C1;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X4Y117_C2;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X4Y117_C3;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X4Y117_C4;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X4Y117_C5;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X4Y117_C6;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X4Y117_CLK;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X4Y117_CO5;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X4Y117_CO6;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X4Y117_C_CY;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X4Y117_C_XOR;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X4Y117_D;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X4Y117_D1;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X4Y117_D2;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X4Y117_D3;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X4Y117_D4;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X4Y117_D5;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X4Y117_D6;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X4Y117_DO5;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X4Y117_DO6;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X4Y117_D_CY;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X4Y117_D_XOR;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X5Y117_A;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X5Y117_A1;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X5Y117_A2;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X5Y117_A3;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X5Y117_A4;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X5Y117_A5;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X5Y117_A6;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X5Y117_AO5;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X5Y117_AO6;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X5Y117_AQ;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X5Y117_A_CY;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X5Y117_A_XOR;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X5Y117_B;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X5Y117_B1;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X5Y117_B2;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X5Y117_B3;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X5Y117_B4;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X5Y117_B5;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X5Y117_B6;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X5Y117_BO5;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X5Y117_BO6;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X5Y117_BQ;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X5Y117_B_CY;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X5Y117_B_XOR;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X5Y117_C;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X5Y117_C1;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X5Y117_C2;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X5Y117_C3;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X5Y117_C4;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X5Y117_C5;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X5Y117_C6;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X5Y117_CLK;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X5Y117_CO5;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X5Y117_CO6;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X5Y117_CQ;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X5Y117_C_CY;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X5Y117_C_XOR;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X5Y117_D;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X5Y117_D1;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X5Y117_D2;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X5Y117_D3;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X5Y117_D4;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X5Y117_D5;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X5Y117_D6;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X5Y117_DO5;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X5Y117_DO6;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X5Y117_DQ;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X5Y117_D_CY;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X5Y117_D_XOR;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X4Y118_A;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X4Y118_A1;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X4Y118_A2;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X4Y118_A3;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X4Y118_A4;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X4Y118_A5;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X4Y118_A6;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X4Y118_AO5;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X4Y118_AO6;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X4Y118_AQ;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X4Y118_A_CY;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X4Y118_A_XOR;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X4Y118_B;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X4Y118_B1;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X4Y118_B2;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X4Y118_B3;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X4Y118_B4;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X4Y118_B5;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X4Y118_B6;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X4Y118_BO5;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X4Y118_BO6;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X4Y118_B_CY;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X4Y118_B_XOR;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X4Y118_C;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X4Y118_C1;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X4Y118_C2;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X4Y118_C3;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X4Y118_C4;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X4Y118_C5;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X4Y118_C6;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X4Y118_CLK;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X4Y118_CO5;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X4Y118_CO6;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X4Y118_C_CY;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X4Y118_C_XOR;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X4Y118_D;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X4Y118_D1;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X4Y118_D2;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X4Y118_D3;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X4Y118_D4;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X4Y118_D5;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X4Y118_D6;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X4Y118_DO5;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X4Y118_DO6;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X4Y118_D_CY;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X4Y118_D_XOR;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X5Y118_A;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X5Y118_A1;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X5Y118_A2;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X5Y118_A3;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X5Y118_A4;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X5Y118_A5;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X5Y118_A6;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X5Y118_AO5;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X5Y118_AO6;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X5Y118_AQ;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X5Y118_A_CY;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X5Y118_A_XOR;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X5Y118_B;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X5Y118_B1;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X5Y118_B2;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X5Y118_B3;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X5Y118_B4;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X5Y118_B5;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X5Y118_B6;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X5Y118_BO5;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X5Y118_BO6;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X5Y118_BQ;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X5Y118_B_CY;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X5Y118_B_XOR;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X5Y118_C;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X5Y118_C1;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X5Y118_C2;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X5Y118_C3;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X5Y118_C4;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X5Y118_C5;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X5Y118_C6;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X5Y118_CLK;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X5Y118_CO5;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X5Y118_CO6;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X5Y118_CQ;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X5Y118_C_CY;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X5Y118_C_XOR;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X5Y118_D;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X5Y118_D1;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X5Y118_D2;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X5Y118_D3;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X5Y118_D4;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X5Y118_D5;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X5Y118_D6;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X5Y118_DO5;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X5Y118_DO6;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X5Y118_D_CY;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X5Y118_D_XOR;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X4Y119_A;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X4Y119_A1;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X4Y119_A2;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X4Y119_A3;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X4Y119_A4;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X4Y119_A5;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X4Y119_A6;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X4Y119_AO5;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X4Y119_AO6;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X4Y119_AQ;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X4Y119_A_CY;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X4Y119_A_XOR;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X4Y119_B;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X4Y119_B1;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X4Y119_B2;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X4Y119_B3;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X4Y119_B4;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X4Y119_B5;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X4Y119_B5Q;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X4Y119_B6;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X4Y119_BMUX;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X4Y119_BO5;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X4Y119_BO6;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X4Y119_BQ;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X4Y119_B_CY;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X4Y119_B_XOR;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X4Y119_C;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X4Y119_C1;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X4Y119_C2;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X4Y119_C3;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X4Y119_C4;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X4Y119_C5;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X4Y119_C5Q;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X4Y119_C6;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X4Y119_CLK;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X4Y119_CMUX;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X4Y119_CO5;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X4Y119_CO6;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X4Y119_CQ;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X4Y119_C_CY;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X4Y119_C_XOR;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X4Y119_D;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X4Y119_D1;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X4Y119_D2;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X4Y119_D3;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X4Y119_D4;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X4Y119_D5;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X4Y119_D6;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X4Y119_DO5;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X4Y119_DO6;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X4Y119_DQ;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X4Y119_D_CY;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X4Y119_D_XOR;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X5Y119_A;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X5Y119_A1;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X5Y119_A2;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X5Y119_A3;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X5Y119_A4;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X5Y119_A5;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X5Y119_A6;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X5Y119_AO5;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X5Y119_AO6;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X5Y119_AQ;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X5Y119_A_CY;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X5Y119_A_XOR;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X5Y119_B;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X5Y119_B1;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X5Y119_B2;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X5Y119_B3;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X5Y119_B4;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X5Y119_B5;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X5Y119_B6;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X5Y119_BO5;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X5Y119_BO6;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X5Y119_B_CY;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X5Y119_B_XOR;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X5Y119_C;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X5Y119_C1;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X5Y119_C2;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X5Y119_C3;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X5Y119_C4;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X5Y119_C5;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X5Y119_C6;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X5Y119_CLK;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X5Y119_CO5;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X5Y119_CO6;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X5Y119_C_CY;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X5Y119_C_XOR;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X5Y119_D;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X5Y119_D1;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X5Y119_D2;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X5Y119_D3;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X5Y119_D4;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X5Y119_D5;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X5Y119_D6;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X5Y119_DO5;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X5Y119_DO6;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X5Y119_D_CY;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X5Y119_D_XOR;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X4Y120_A;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X4Y120_A1;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X4Y120_A2;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X4Y120_A3;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X4Y120_A4;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X4Y120_A5;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X4Y120_A6;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X4Y120_AO5;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X4Y120_AO6;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X4Y120_A_CY;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X4Y120_A_XOR;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X4Y120_B;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X4Y120_B1;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X4Y120_B2;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X4Y120_B3;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X4Y120_B4;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X4Y120_B5;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X4Y120_B6;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X4Y120_BO5;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X4Y120_BO6;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X4Y120_B_CY;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X4Y120_B_XOR;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X4Y120_C;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X4Y120_C1;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X4Y120_C2;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X4Y120_C3;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X4Y120_C4;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X4Y120_C5;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X4Y120_C6;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X4Y120_CO5;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X4Y120_CO6;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X4Y120_C_CY;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X4Y120_C_XOR;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X4Y120_D;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X4Y120_D1;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X4Y120_D2;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X4Y120_D3;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X4Y120_D4;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X4Y120_D5;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X4Y120_D6;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X4Y120_DMUX;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X4Y120_DO5;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X4Y120_DO6;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X4Y120_D_CY;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X4Y120_D_XOR;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X5Y120_A;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X5Y120_A1;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X5Y120_A2;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X5Y120_A3;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X5Y120_A4;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X5Y120_A5;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X5Y120_A6;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X5Y120_AMUX;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X5Y120_AO5;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X5Y120_AO6;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X5Y120_A_CY;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X5Y120_A_XOR;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X5Y120_B;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X5Y120_B1;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X5Y120_B2;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X5Y120_B3;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X5Y120_B4;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X5Y120_B5;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X5Y120_B6;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X5Y120_BMUX;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X5Y120_BO5;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X5Y120_BO6;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X5Y120_B_CY;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X5Y120_B_XOR;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X5Y120_C;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X5Y120_C1;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X5Y120_C2;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X5Y120_C3;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X5Y120_C4;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X5Y120_C5;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X5Y120_C6;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X5Y120_CO5;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X5Y120_CO6;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X5Y120_C_CY;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X5Y120_C_XOR;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X5Y120_D;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X5Y120_D1;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X5Y120_D2;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X5Y120_D3;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X5Y120_D4;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X5Y120_D5;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X5Y120_D6;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X5Y120_DO5;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X5Y120_DO6;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X5Y120_D_CY;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X5Y120_D_XOR;
  wire [0:0] CLBLL_L_X4Y121_SLICE_X4Y121_A;
  wire [0:0] CLBLL_L_X4Y121_SLICE_X4Y121_A1;
  wire [0:0] CLBLL_L_X4Y121_SLICE_X4Y121_A2;
  wire [0:0] CLBLL_L_X4Y121_SLICE_X4Y121_A3;
  wire [0:0] CLBLL_L_X4Y121_SLICE_X4Y121_A4;
  wire [0:0] CLBLL_L_X4Y121_SLICE_X4Y121_A5;
  wire [0:0] CLBLL_L_X4Y121_SLICE_X4Y121_A6;
  wire [0:0] CLBLL_L_X4Y121_SLICE_X4Y121_AO5;
  wire [0:0] CLBLL_L_X4Y121_SLICE_X4Y121_AO6;
  wire [0:0] CLBLL_L_X4Y121_SLICE_X4Y121_AQ;
  wire [0:0] CLBLL_L_X4Y121_SLICE_X4Y121_A_CY;
  wire [0:0] CLBLL_L_X4Y121_SLICE_X4Y121_A_XOR;
  wire [0:0] CLBLL_L_X4Y121_SLICE_X4Y121_B;
  wire [0:0] CLBLL_L_X4Y121_SLICE_X4Y121_B1;
  wire [0:0] CLBLL_L_X4Y121_SLICE_X4Y121_B2;
  wire [0:0] CLBLL_L_X4Y121_SLICE_X4Y121_B3;
  wire [0:0] CLBLL_L_X4Y121_SLICE_X4Y121_B4;
  wire [0:0] CLBLL_L_X4Y121_SLICE_X4Y121_B5;
  wire [0:0] CLBLL_L_X4Y121_SLICE_X4Y121_B6;
  wire [0:0] CLBLL_L_X4Y121_SLICE_X4Y121_BO5;
  wire [0:0] CLBLL_L_X4Y121_SLICE_X4Y121_BO6;
  wire [0:0] CLBLL_L_X4Y121_SLICE_X4Y121_BQ;
  wire [0:0] CLBLL_L_X4Y121_SLICE_X4Y121_B_CY;
  wire [0:0] CLBLL_L_X4Y121_SLICE_X4Y121_B_XOR;
  wire [0:0] CLBLL_L_X4Y121_SLICE_X4Y121_C;
  wire [0:0] CLBLL_L_X4Y121_SLICE_X4Y121_C1;
  wire [0:0] CLBLL_L_X4Y121_SLICE_X4Y121_C2;
  wire [0:0] CLBLL_L_X4Y121_SLICE_X4Y121_C3;
  wire [0:0] CLBLL_L_X4Y121_SLICE_X4Y121_C4;
  wire [0:0] CLBLL_L_X4Y121_SLICE_X4Y121_C5;
  wire [0:0] CLBLL_L_X4Y121_SLICE_X4Y121_C6;
  wire [0:0] CLBLL_L_X4Y121_SLICE_X4Y121_CLK;
  wire [0:0] CLBLL_L_X4Y121_SLICE_X4Y121_CMUX;
  wire [0:0] CLBLL_L_X4Y121_SLICE_X4Y121_CO5;
  wire [0:0] CLBLL_L_X4Y121_SLICE_X4Y121_CO6;
  wire [0:0] CLBLL_L_X4Y121_SLICE_X4Y121_C_CY;
  wire [0:0] CLBLL_L_X4Y121_SLICE_X4Y121_C_XOR;
  wire [0:0] CLBLL_L_X4Y121_SLICE_X4Y121_D;
  wire [0:0] CLBLL_L_X4Y121_SLICE_X4Y121_D1;
  wire [0:0] CLBLL_L_X4Y121_SLICE_X4Y121_D2;
  wire [0:0] CLBLL_L_X4Y121_SLICE_X4Y121_D3;
  wire [0:0] CLBLL_L_X4Y121_SLICE_X4Y121_D4;
  wire [0:0] CLBLL_L_X4Y121_SLICE_X4Y121_D5;
  wire [0:0] CLBLL_L_X4Y121_SLICE_X4Y121_D6;
  wire [0:0] CLBLL_L_X4Y121_SLICE_X4Y121_DMUX;
  wire [0:0] CLBLL_L_X4Y121_SLICE_X4Y121_DO5;
  wire [0:0] CLBLL_L_X4Y121_SLICE_X4Y121_DO6;
  wire [0:0] CLBLL_L_X4Y121_SLICE_X4Y121_D_CY;
  wire [0:0] CLBLL_L_X4Y121_SLICE_X4Y121_D_XOR;
  wire [0:0] CLBLL_L_X4Y121_SLICE_X5Y121_A;
  wire [0:0] CLBLL_L_X4Y121_SLICE_X5Y121_A1;
  wire [0:0] CLBLL_L_X4Y121_SLICE_X5Y121_A2;
  wire [0:0] CLBLL_L_X4Y121_SLICE_X5Y121_A3;
  wire [0:0] CLBLL_L_X4Y121_SLICE_X5Y121_A4;
  wire [0:0] CLBLL_L_X4Y121_SLICE_X5Y121_A5;
  wire [0:0] CLBLL_L_X4Y121_SLICE_X5Y121_A6;
  wire [0:0] CLBLL_L_X4Y121_SLICE_X5Y121_AO5;
  wire [0:0] CLBLL_L_X4Y121_SLICE_X5Y121_AO6;
  wire [0:0] CLBLL_L_X4Y121_SLICE_X5Y121_AQ;
  wire [0:0] CLBLL_L_X4Y121_SLICE_X5Y121_A_CY;
  wire [0:0] CLBLL_L_X4Y121_SLICE_X5Y121_A_XOR;
  wire [0:0] CLBLL_L_X4Y121_SLICE_X5Y121_B;
  wire [0:0] CLBLL_L_X4Y121_SLICE_X5Y121_B1;
  wire [0:0] CLBLL_L_X4Y121_SLICE_X5Y121_B2;
  wire [0:0] CLBLL_L_X4Y121_SLICE_X5Y121_B3;
  wire [0:0] CLBLL_L_X4Y121_SLICE_X5Y121_B4;
  wire [0:0] CLBLL_L_X4Y121_SLICE_X5Y121_B5;
  wire [0:0] CLBLL_L_X4Y121_SLICE_X5Y121_B6;
  wire [0:0] CLBLL_L_X4Y121_SLICE_X5Y121_BMUX;
  wire [0:0] CLBLL_L_X4Y121_SLICE_X5Y121_BO5;
  wire [0:0] CLBLL_L_X4Y121_SLICE_X5Y121_BO6;
  wire [0:0] CLBLL_L_X4Y121_SLICE_X5Y121_B_CY;
  wire [0:0] CLBLL_L_X4Y121_SLICE_X5Y121_B_XOR;
  wire [0:0] CLBLL_L_X4Y121_SLICE_X5Y121_C;
  wire [0:0] CLBLL_L_X4Y121_SLICE_X5Y121_C1;
  wire [0:0] CLBLL_L_X4Y121_SLICE_X5Y121_C2;
  wire [0:0] CLBLL_L_X4Y121_SLICE_X5Y121_C3;
  wire [0:0] CLBLL_L_X4Y121_SLICE_X5Y121_C4;
  wire [0:0] CLBLL_L_X4Y121_SLICE_X5Y121_C5;
  wire [0:0] CLBLL_L_X4Y121_SLICE_X5Y121_C6;
  wire [0:0] CLBLL_L_X4Y121_SLICE_X5Y121_CLK;
  wire [0:0] CLBLL_L_X4Y121_SLICE_X5Y121_CMUX;
  wire [0:0] CLBLL_L_X4Y121_SLICE_X5Y121_CO5;
  wire [0:0] CLBLL_L_X4Y121_SLICE_X5Y121_CO6;
  wire [0:0] CLBLL_L_X4Y121_SLICE_X5Y121_C_CY;
  wire [0:0] CLBLL_L_X4Y121_SLICE_X5Y121_C_XOR;
  wire [0:0] CLBLL_L_X4Y121_SLICE_X5Y121_D;
  wire [0:0] CLBLL_L_X4Y121_SLICE_X5Y121_D1;
  wire [0:0] CLBLL_L_X4Y121_SLICE_X5Y121_D2;
  wire [0:0] CLBLL_L_X4Y121_SLICE_X5Y121_D3;
  wire [0:0] CLBLL_L_X4Y121_SLICE_X5Y121_D4;
  wire [0:0] CLBLL_L_X4Y121_SLICE_X5Y121_D5;
  wire [0:0] CLBLL_L_X4Y121_SLICE_X5Y121_D6;
  wire [0:0] CLBLL_L_X4Y121_SLICE_X5Y121_DO5;
  wire [0:0] CLBLL_L_X4Y121_SLICE_X5Y121_DO6;
  wire [0:0] CLBLL_L_X4Y121_SLICE_X5Y121_D_CY;
  wire [0:0] CLBLL_L_X4Y121_SLICE_X5Y121_D_XOR;
  wire [0:0] CLBLL_L_X4Y122_SLICE_X4Y122_A;
  wire [0:0] CLBLL_L_X4Y122_SLICE_X4Y122_A1;
  wire [0:0] CLBLL_L_X4Y122_SLICE_X4Y122_A2;
  wire [0:0] CLBLL_L_X4Y122_SLICE_X4Y122_A3;
  wire [0:0] CLBLL_L_X4Y122_SLICE_X4Y122_A4;
  wire [0:0] CLBLL_L_X4Y122_SLICE_X4Y122_A5;
  wire [0:0] CLBLL_L_X4Y122_SLICE_X4Y122_A6;
  wire [0:0] CLBLL_L_X4Y122_SLICE_X4Y122_AMUX;
  wire [0:0] CLBLL_L_X4Y122_SLICE_X4Y122_AO5;
  wire [0:0] CLBLL_L_X4Y122_SLICE_X4Y122_AO6;
  wire [0:0] CLBLL_L_X4Y122_SLICE_X4Y122_A_CY;
  wire [0:0] CLBLL_L_X4Y122_SLICE_X4Y122_A_XOR;
  wire [0:0] CLBLL_L_X4Y122_SLICE_X4Y122_B;
  wire [0:0] CLBLL_L_X4Y122_SLICE_X4Y122_B1;
  wire [0:0] CLBLL_L_X4Y122_SLICE_X4Y122_B2;
  wire [0:0] CLBLL_L_X4Y122_SLICE_X4Y122_B3;
  wire [0:0] CLBLL_L_X4Y122_SLICE_X4Y122_B4;
  wire [0:0] CLBLL_L_X4Y122_SLICE_X4Y122_B5;
  wire [0:0] CLBLL_L_X4Y122_SLICE_X4Y122_B6;
  wire [0:0] CLBLL_L_X4Y122_SLICE_X4Y122_BO5;
  wire [0:0] CLBLL_L_X4Y122_SLICE_X4Y122_BO6;
  wire [0:0] CLBLL_L_X4Y122_SLICE_X4Y122_B_CY;
  wire [0:0] CLBLL_L_X4Y122_SLICE_X4Y122_B_XOR;
  wire [0:0] CLBLL_L_X4Y122_SLICE_X4Y122_C;
  wire [0:0] CLBLL_L_X4Y122_SLICE_X4Y122_C1;
  wire [0:0] CLBLL_L_X4Y122_SLICE_X4Y122_C2;
  wire [0:0] CLBLL_L_X4Y122_SLICE_X4Y122_C3;
  wire [0:0] CLBLL_L_X4Y122_SLICE_X4Y122_C4;
  wire [0:0] CLBLL_L_X4Y122_SLICE_X4Y122_C5;
  wire [0:0] CLBLL_L_X4Y122_SLICE_X4Y122_C6;
  wire [0:0] CLBLL_L_X4Y122_SLICE_X4Y122_CO5;
  wire [0:0] CLBLL_L_X4Y122_SLICE_X4Y122_CO6;
  wire [0:0] CLBLL_L_X4Y122_SLICE_X4Y122_C_CY;
  wire [0:0] CLBLL_L_X4Y122_SLICE_X4Y122_C_XOR;
  wire [0:0] CLBLL_L_X4Y122_SLICE_X4Y122_D;
  wire [0:0] CLBLL_L_X4Y122_SLICE_X4Y122_D1;
  wire [0:0] CLBLL_L_X4Y122_SLICE_X4Y122_D2;
  wire [0:0] CLBLL_L_X4Y122_SLICE_X4Y122_D3;
  wire [0:0] CLBLL_L_X4Y122_SLICE_X4Y122_D4;
  wire [0:0] CLBLL_L_X4Y122_SLICE_X4Y122_D5;
  wire [0:0] CLBLL_L_X4Y122_SLICE_X4Y122_D6;
  wire [0:0] CLBLL_L_X4Y122_SLICE_X4Y122_DO5;
  wire [0:0] CLBLL_L_X4Y122_SLICE_X4Y122_DO6;
  wire [0:0] CLBLL_L_X4Y122_SLICE_X4Y122_D_CY;
  wire [0:0] CLBLL_L_X4Y122_SLICE_X4Y122_D_XOR;
  wire [0:0] CLBLL_L_X4Y122_SLICE_X5Y122_A;
  wire [0:0] CLBLL_L_X4Y122_SLICE_X5Y122_A1;
  wire [0:0] CLBLL_L_X4Y122_SLICE_X5Y122_A2;
  wire [0:0] CLBLL_L_X4Y122_SLICE_X5Y122_A3;
  wire [0:0] CLBLL_L_X4Y122_SLICE_X5Y122_A4;
  wire [0:0] CLBLL_L_X4Y122_SLICE_X5Y122_A5;
  wire [0:0] CLBLL_L_X4Y122_SLICE_X5Y122_A6;
  wire [0:0] CLBLL_L_X4Y122_SLICE_X5Y122_AO5;
  wire [0:0] CLBLL_L_X4Y122_SLICE_X5Y122_AO6;
  wire [0:0] CLBLL_L_X4Y122_SLICE_X5Y122_A_CY;
  wire [0:0] CLBLL_L_X4Y122_SLICE_X5Y122_A_XOR;
  wire [0:0] CLBLL_L_X4Y122_SLICE_X5Y122_B;
  wire [0:0] CLBLL_L_X4Y122_SLICE_X5Y122_B1;
  wire [0:0] CLBLL_L_X4Y122_SLICE_X5Y122_B2;
  wire [0:0] CLBLL_L_X4Y122_SLICE_X5Y122_B3;
  wire [0:0] CLBLL_L_X4Y122_SLICE_X5Y122_B4;
  wire [0:0] CLBLL_L_X4Y122_SLICE_X5Y122_B5;
  wire [0:0] CLBLL_L_X4Y122_SLICE_X5Y122_B6;
  wire [0:0] CLBLL_L_X4Y122_SLICE_X5Y122_BO5;
  wire [0:0] CLBLL_L_X4Y122_SLICE_X5Y122_BO6;
  wire [0:0] CLBLL_L_X4Y122_SLICE_X5Y122_B_CY;
  wire [0:0] CLBLL_L_X4Y122_SLICE_X5Y122_B_XOR;
  wire [0:0] CLBLL_L_X4Y122_SLICE_X5Y122_C;
  wire [0:0] CLBLL_L_X4Y122_SLICE_X5Y122_C1;
  wire [0:0] CLBLL_L_X4Y122_SLICE_X5Y122_C2;
  wire [0:0] CLBLL_L_X4Y122_SLICE_X5Y122_C3;
  wire [0:0] CLBLL_L_X4Y122_SLICE_X5Y122_C4;
  wire [0:0] CLBLL_L_X4Y122_SLICE_X5Y122_C5;
  wire [0:0] CLBLL_L_X4Y122_SLICE_X5Y122_C6;
  wire [0:0] CLBLL_L_X4Y122_SLICE_X5Y122_CO5;
  wire [0:0] CLBLL_L_X4Y122_SLICE_X5Y122_CO6;
  wire [0:0] CLBLL_L_X4Y122_SLICE_X5Y122_C_CY;
  wire [0:0] CLBLL_L_X4Y122_SLICE_X5Y122_C_XOR;
  wire [0:0] CLBLL_L_X4Y122_SLICE_X5Y122_D;
  wire [0:0] CLBLL_L_X4Y122_SLICE_X5Y122_D1;
  wire [0:0] CLBLL_L_X4Y122_SLICE_X5Y122_D2;
  wire [0:0] CLBLL_L_X4Y122_SLICE_X5Y122_D3;
  wire [0:0] CLBLL_L_X4Y122_SLICE_X5Y122_D4;
  wire [0:0] CLBLL_L_X4Y122_SLICE_X5Y122_D5;
  wire [0:0] CLBLL_L_X4Y122_SLICE_X5Y122_D6;
  wire [0:0] CLBLL_L_X4Y122_SLICE_X5Y122_DO5;
  wire [0:0] CLBLL_L_X4Y122_SLICE_X5Y122_DO6;
  wire [0:0] CLBLL_L_X4Y122_SLICE_X5Y122_D_CY;
  wire [0:0] CLBLL_L_X4Y122_SLICE_X5Y122_D_XOR;
  wire [0:0] CLBLL_L_X4Y123_SLICE_X4Y123_A;
  wire [0:0] CLBLL_L_X4Y123_SLICE_X4Y123_A1;
  wire [0:0] CLBLL_L_X4Y123_SLICE_X4Y123_A2;
  wire [0:0] CLBLL_L_X4Y123_SLICE_X4Y123_A3;
  wire [0:0] CLBLL_L_X4Y123_SLICE_X4Y123_A4;
  wire [0:0] CLBLL_L_X4Y123_SLICE_X4Y123_A5;
  wire [0:0] CLBLL_L_X4Y123_SLICE_X4Y123_A6;
  wire [0:0] CLBLL_L_X4Y123_SLICE_X4Y123_AO5;
  wire [0:0] CLBLL_L_X4Y123_SLICE_X4Y123_AO6;
  wire [0:0] CLBLL_L_X4Y123_SLICE_X4Y123_AQ;
  wire [0:0] CLBLL_L_X4Y123_SLICE_X4Y123_A_CY;
  wire [0:0] CLBLL_L_X4Y123_SLICE_X4Y123_A_XOR;
  wire [0:0] CLBLL_L_X4Y123_SLICE_X4Y123_B;
  wire [0:0] CLBLL_L_X4Y123_SLICE_X4Y123_B1;
  wire [0:0] CLBLL_L_X4Y123_SLICE_X4Y123_B2;
  wire [0:0] CLBLL_L_X4Y123_SLICE_X4Y123_B3;
  wire [0:0] CLBLL_L_X4Y123_SLICE_X4Y123_B4;
  wire [0:0] CLBLL_L_X4Y123_SLICE_X4Y123_B5;
  wire [0:0] CLBLL_L_X4Y123_SLICE_X4Y123_B6;
  wire [0:0] CLBLL_L_X4Y123_SLICE_X4Y123_BO5;
  wire [0:0] CLBLL_L_X4Y123_SLICE_X4Y123_BO6;
  wire [0:0] CLBLL_L_X4Y123_SLICE_X4Y123_BQ;
  wire [0:0] CLBLL_L_X4Y123_SLICE_X4Y123_B_CY;
  wire [0:0] CLBLL_L_X4Y123_SLICE_X4Y123_B_XOR;
  wire [0:0] CLBLL_L_X4Y123_SLICE_X4Y123_C;
  wire [0:0] CLBLL_L_X4Y123_SLICE_X4Y123_C1;
  wire [0:0] CLBLL_L_X4Y123_SLICE_X4Y123_C2;
  wire [0:0] CLBLL_L_X4Y123_SLICE_X4Y123_C3;
  wire [0:0] CLBLL_L_X4Y123_SLICE_X4Y123_C4;
  wire [0:0] CLBLL_L_X4Y123_SLICE_X4Y123_C5;
  wire [0:0] CLBLL_L_X4Y123_SLICE_X4Y123_C6;
  wire [0:0] CLBLL_L_X4Y123_SLICE_X4Y123_CLK;
  wire [0:0] CLBLL_L_X4Y123_SLICE_X4Y123_CO5;
  wire [0:0] CLBLL_L_X4Y123_SLICE_X4Y123_CO6;
  wire [0:0] CLBLL_L_X4Y123_SLICE_X4Y123_CQ;
  wire [0:0] CLBLL_L_X4Y123_SLICE_X4Y123_C_CY;
  wire [0:0] CLBLL_L_X4Y123_SLICE_X4Y123_C_XOR;
  wire [0:0] CLBLL_L_X4Y123_SLICE_X4Y123_D;
  wire [0:0] CLBLL_L_X4Y123_SLICE_X4Y123_D1;
  wire [0:0] CLBLL_L_X4Y123_SLICE_X4Y123_D2;
  wire [0:0] CLBLL_L_X4Y123_SLICE_X4Y123_D3;
  wire [0:0] CLBLL_L_X4Y123_SLICE_X4Y123_D4;
  wire [0:0] CLBLL_L_X4Y123_SLICE_X4Y123_D5;
  wire [0:0] CLBLL_L_X4Y123_SLICE_X4Y123_D6;
  wire [0:0] CLBLL_L_X4Y123_SLICE_X4Y123_DO5;
  wire [0:0] CLBLL_L_X4Y123_SLICE_X4Y123_DO6;
  wire [0:0] CLBLL_L_X4Y123_SLICE_X4Y123_D_CY;
  wire [0:0] CLBLL_L_X4Y123_SLICE_X4Y123_D_XOR;
  wire [0:0] CLBLL_L_X4Y123_SLICE_X5Y123_A;
  wire [0:0] CLBLL_L_X4Y123_SLICE_X5Y123_A1;
  wire [0:0] CLBLL_L_X4Y123_SLICE_X5Y123_A2;
  wire [0:0] CLBLL_L_X4Y123_SLICE_X5Y123_A3;
  wire [0:0] CLBLL_L_X4Y123_SLICE_X5Y123_A4;
  wire [0:0] CLBLL_L_X4Y123_SLICE_X5Y123_A5;
  wire [0:0] CLBLL_L_X4Y123_SLICE_X5Y123_A6;
  wire [0:0] CLBLL_L_X4Y123_SLICE_X5Y123_AMUX;
  wire [0:0] CLBLL_L_X4Y123_SLICE_X5Y123_AO5;
  wire [0:0] CLBLL_L_X4Y123_SLICE_X5Y123_AO6;
  wire [0:0] CLBLL_L_X4Y123_SLICE_X5Y123_A_CY;
  wire [0:0] CLBLL_L_X4Y123_SLICE_X5Y123_A_XOR;
  wire [0:0] CLBLL_L_X4Y123_SLICE_X5Y123_B;
  wire [0:0] CLBLL_L_X4Y123_SLICE_X5Y123_B1;
  wire [0:0] CLBLL_L_X4Y123_SLICE_X5Y123_B2;
  wire [0:0] CLBLL_L_X4Y123_SLICE_X5Y123_B3;
  wire [0:0] CLBLL_L_X4Y123_SLICE_X5Y123_B4;
  wire [0:0] CLBLL_L_X4Y123_SLICE_X5Y123_B5;
  wire [0:0] CLBLL_L_X4Y123_SLICE_X5Y123_B6;
  wire [0:0] CLBLL_L_X4Y123_SLICE_X5Y123_BO5;
  wire [0:0] CLBLL_L_X4Y123_SLICE_X5Y123_BO6;
  wire [0:0] CLBLL_L_X4Y123_SLICE_X5Y123_B_CY;
  wire [0:0] CLBLL_L_X4Y123_SLICE_X5Y123_B_XOR;
  wire [0:0] CLBLL_L_X4Y123_SLICE_X5Y123_C;
  wire [0:0] CLBLL_L_X4Y123_SLICE_X5Y123_C1;
  wire [0:0] CLBLL_L_X4Y123_SLICE_X5Y123_C2;
  wire [0:0] CLBLL_L_X4Y123_SLICE_X5Y123_C3;
  wire [0:0] CLBLL_L_X4Y123_SLICE_X5Y123_C4;
  wire [0:0] CLBLL_L_X4Y123_SLICE_X5Y123_C5;
  wire [0:0] CLBLL_L_X4Y123_SLICE_X5Y123_C6;
  wire [0:0] CLBLL_L_X4Y123_SLICE_X5Y123_CO5;
  wire [0:0] CLBLL_L_X4Y123_SLICE_X5Y123_CO6;
  wire [0:0] CLBLL_L_X4Y123_SLICE_X5Y123_C_CY;
  wire [0:0] CLBLL_L_X4Y123_SLICE_X5Y123_C_XOR;
  wire [0:0] CLBLL_L_X4Y123_SLICE_X5Y123_D;
  wire [0:0] CLBLL_L_X4Y123_SLICE_X5Y123_D1;
  wire [0:0] CLBLL_L_X4Y123_SLICE_X5Y123_D2;
  wire [0:0] CLBLL_L_X4Y123_SLICE_X5Y123_D3;
  wire [0:0] CLBLL_L_X4Y123_SLICE_X5Y123_D4;
  wire [0:0] CLBLL_L_X4Y123_SLICE_X5Y123_D5;
  wire [0:0] CLBLL_L_X4Y123_SLICE_X5Y123_D6;
  wire [0:0] CLBLL_L_X4Y123_SLICE_X5Y123_DO5;
  wire [0:0] CLBLL_L_X4Y123_SLICE_X5Y123_DO6;
  wire [0:0] CLBLL_L_X4Y123_SLICE_X5Y123_D_CY;
  wire [0:0] CLBLL_L_X4Y123_SLICE_X5Y123_D_XOR;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X78Y126_A;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X78Y126_A1;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X78Y126_A2;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X78Y126_A3;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X78Y126_A4;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X78Y126_A5;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X78Y126_A6;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X78Y126_AO5;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X78Y126_AO6;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X78Y126_A_CY;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X78Y126_A_XOR;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X78Y126_B;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X78Y126_B1;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X78Y126_B2;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X78Y126_B3;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X78Y126_B4;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X78Y126_B5;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X78Y126_B6;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X78Y126_BO5;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X78Y126_BO6;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X78Y126_B_CY;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X78Y126_B_XOR;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X78Y126_C;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X78Y126_C1;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X78Y126_C2;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X78Y126_C3;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X78Y126_C4;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X78Y126_C5;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X78Y126_C6;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X78Y126_CO5;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X78Y126_CO6;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X78Y126_C_CY;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X78Y126_C_XOR;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X78Y126_D;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X78Y126_D1;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X78Y126_D2;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X78Y126_D3;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X78Y126_D4;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X78Y126_D5;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X78Y126_D6;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X78Y126_DO5;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X78Y126_DO6;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X78Y126_D_CY;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X78Y126_D_XOR;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X79Y126_A;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X79Y126_A1;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X79Y126_A2;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X79Y126_A3;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X79Y126_A4;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X79Y126_A5;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X79Y126_A6;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X79Y126_AO5;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X79Y126_AO6;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X79Y126_A_CY;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X79Y126_A_XOR;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X79Y126_B;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X79Y126_B1;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X79Y126_B2;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X79Y126_B3;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X79Y126_B4;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X79Y126_B5;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X79Y126_B6;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X79Y126_BO5;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X79Y126_BO6;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X79Y126_B_CY;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X79Y126_B_XOR;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X79Y126_C;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X79Y126_C1;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X79Y126_C2;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X79Y126_C3;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X79Y126_C4;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X79Y126_C5;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X79Y126_C6;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X79Y126_CO5;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X79Y126_CO6;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X79Y126_C_CY;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X79Y126_C_XOR;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X79Y126_D;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X79Y126_D1;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X79Y126_D2;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X79Y126_D3;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X79Y126_D4;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X79Y126_D5;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X79Y126_D6;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X79Y126_DO5;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X79Y126_DO6;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X79Y126_D_CY;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X79Y126_D_XOR;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X12Y110_A;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X12Y110_A1;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X12Y110_A2;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X12Y110_A3;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X12Y110_A4;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X12Y110_A5;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X12Y110_A6;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X12Y110_AO5;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X12Y110_AO6;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X12Y110_AQ;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X12Y110_A_CY;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X12Y110_A_XOR;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X12Y110_B;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X12Y110_B1;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X12Y110_B2;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X12Y110_B3;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X12Y110_B4;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X12Y110_B5;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X12Y110_B6;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X12Y110_BO5;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X12Y110_BO6;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X12Y110_BQ;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X12Y110_B_CY;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X12Y110_B_XOR;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X12Y110_C;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X12Y110_C1;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X12Y110_C2;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X12Y110_C3;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X12Y110_C4;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X12Y110_C5;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X12Y110_C6;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X12Y110_CLK;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X12Y110_CO5;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X12Y110_CO6;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X12Y110_C_CY;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X12Y110_C_XOR;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X12Y110_D;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X12Y110_D1;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X12Y110_D2;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X12Y110_D3;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X12Y110_D4;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X12Y110_D5;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X12Y110_D6;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X12Y110_DO5;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X12Y110_DO6;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X12Y110_D_CY;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X12Y110_D_XOR;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X13Y110_A;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X13Y110_A1;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X13Y110_A2;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X13Y110_A3;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X13Y110_A4;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X13Y110_A5;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X13Y110_A6;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X13Y110_AO5;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X13Y110_AO6;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X13Y110_AQ;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X13Y110_A_CY;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X13Y110_A_XOR;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X13Y110_B;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X13Y110_B1;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X13Y110_B2;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X13Y110_B3;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X13Y110_B4;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X13Y110_B5;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X13Y110_B6;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X13Y110_BO5;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X13Y110_BO6;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X13Y110_BQ;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X13Y110_B_CY;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X13Y110_B_XOR;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X13Y110_C;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X13Y110_C1;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X13Y110_C2;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X13Y110_C3;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X13Y110_C4;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X13Y110_C5;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X13Y110_C6;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X13Y110_CLK;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X13Y110_CMUX;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X13Y110_CO5;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X13Y110_CO6;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X13Y110_C_CY;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X13Y110_C_XOR;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X13Y110_D;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X13Y110_D1;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X13Y110_D2;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X13Y110_D3;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X13Y110_D4;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X13Y110_D5;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X13Y110_D6;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X13Y110_DMUX;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X13Y110_DO5;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X13Y110_DO6;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X13Y110_D_CY;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X13Y110_D_XOR;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X12Y111_A;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X12Y111_A1;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X12Y111_A2;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X12Y111_A3;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X12Y111_A4;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X12Y111_A5;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X12Y111_A6;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X12Y111_AMUX;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X12Y111_AO5;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X12Y111_AO6;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X12Y111_A_CY;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X12Y111_A_XOR;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X12Y111_B;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X12Y111_B1;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X12Y111_B2;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X12Y111_B3;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X12Y111_B4;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X12Y111_B5;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X12Y111_B6;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X12Y111_BMUX;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X12Y111_BO5;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X12Y111_BO6;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X12Y111_B_CY;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X12Y111_B_XOR;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X12Y111_C;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X12Y111_C1;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X12Y111_C2;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X12Y111_C3;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X12Y111_C4;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X12Y111_C5;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X12Y111_C6;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X12Y111_CO5;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X12Y111_CO6;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X12Y111_C_CY;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X12Y111_C_XOR;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X12Y111_D;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X12Y111_D1;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X12Y111_D2;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X12Y111_D3;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X12Y111_D4;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X12Y111_D5;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X12Y111_D6;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X12Y111_DO5;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X12Y111_DO6;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X12Y111_D_CY;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X12Y111_D_XOR;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X13Y111_A;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X13Y111_A1;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X13Y111_A2;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X13Y111_A3;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X13Y111_A4;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X13Y111_A5;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X13Y111_A6;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X13Y111_AO5;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X13Y111_AO6;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X13Y111_AQ;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X13Y111_A_CY;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X13Y111_A_XOR;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X13Y111_B;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X13Y111_B1;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X13Y111_B2;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X13Y111_B3;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X13Y111_B4;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X13Y111_B5;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X13Y111_B6;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X13Y111_BMUX;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X13Y111_BO5;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X13Y111_BO6;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X13Y111_B_CY;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X13Y111_B_XOR;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X13Y111_C;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X13Y111_C1;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X13Y111_C2;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X13Y111_C3;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X13Y111_C4;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X13Y111_C5;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X13Y111_C6;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X13Y111_CLK;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X13Y111_CMUX;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X13Y111_CO5;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X13Y111_CO6;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X13Y111_C_CY;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X13Y111_C_XOR;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X13Y111_D;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X13Y111_D1;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X13Y111_D2;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X13Y111_D3;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X13Y111_D4;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X13Y111_D5;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X13Y111_D6;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X13Y111_DO5;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X13Y111_DO6;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X13Y111_D_CY;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X13Y111_D_XOR;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X12Y112_A;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X12Y112_A1;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X12Y112_A2;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X12Y112_A3;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X12Y112_A4;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X12Y112_A5;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X12Y112_A6;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X12Y112_AMUX;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X12Y112_AO5;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X12Y112_AO6;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X12Y112_A_CY;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X12Y112_A_XOR;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X12Y112_B;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X12Y112_B1;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X12Y112_B2;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X12Y112_B3;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X12Y112_B4;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X12Y112_B5;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X12Y112_B6;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X12Y112_BO5;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X12Y112_BO6;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X12Y112_BQ;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X12Y112_B_CY;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X12Y112_B_XOR;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X12Y112_C;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X12Y112_C1;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X12Y112_C2;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X12Y112_C3;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X12Y112_C4;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X12Y112_C5;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X12Y112_C6;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X12Y112_CLK;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X12Y112_CO5;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X12Y112_CO6;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X12Y112_CQ;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X12Y112_C_CY;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X12Y112_C_XOR;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X12Y112_D;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X12Y112_D1;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X12Y112_D2;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X12Y112_D3;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X12Y112_D4;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X12Y112_D5;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X12Y112_D6;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X12Y112_DO5;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X12Y112_DO6;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X12Y112_DQ;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X12Y112_D_CY;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X12Y112_D_XOR;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X13Y112_A;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X13Y112_A1;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X13Y112_A2;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X13Y112_A3;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X13Y112_A4;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X13Y112_A5;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X13Y112_A6;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X13Y112_AO5;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X13Y112_AO6;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X13Y112_AQ;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X13Y112_A_CY;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X13Y112_A_XOR;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X13Y112_B;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X13Y112_B1;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X13Y112_B2;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X13Y112_B3;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X13Y112_B4;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X13Y112_B5;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X13Y112_B6;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X13Y112_BO5;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X13Y112_BO6;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X13Y112_BQ;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X13Y112_B_CY;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X13Y112_B_XOR;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X13Y112_C;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X13Y112_C1;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X13Y112_C2;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X13Y112_C3;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X13Y112_C4;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X13Y112_C5;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X13Y112_C6;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X13Y112_CLK;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X13Y112_CO5;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X13Y112_CO6;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X13Y112_CQ;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X13Y112_C_CY;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X13Y112_C_XOR;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X13Y112_D;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X13Y112_D1;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X13Y112_D2;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X13Y112_D3;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X13Y112_D4;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X13Y112_D5;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X13Y112_D6;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X13Y112_DO5;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X13Y112_DO6;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X13Y112_D_CY;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X13Y112_D_XOR;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X12Y113_A;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X12Y113_A1;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X12Y113_A2;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X12Y113_A3;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X12Y113_A4;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X12Y113_A5;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X12Y113_A6;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X12Y113_AMUX;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X12Y113_AO5;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X12Y113_AO6;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X12Y113_A_CY;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X12Y113_A_XOR;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X12Y113_B;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X12Y113_B1;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X12Y113_B2;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X12Y113_B3;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X12Y113_B4;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X12Y113_B5;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X12Y113_B6;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X12Y113_BO5;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X12Y113_BO6;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X12Y113_BQ;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X12Y113_B_CY;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X12Y113_B_XOR;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X12Y113_C;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X12Y113_C1;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X12Y113_C2;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X12Y113_C3;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X12Y113_C4;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X12Y113_C5;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X12Y113_C6;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X12Y113_CLK;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X12Y113_CO5;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X12Y113_CO6;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X12Y113_C_CY;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X12Y113_C_XOR;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X12Y113_D;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X12Y113_D1;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X12Y113_D2;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X12Y113_D3;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X12Y113_D4;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X12Y113_D5;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X12Y113_D6;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X12Y113_DO5;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X12Y113_DO6;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X12Y113_D_CY;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X12Y113_D_XOR;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X13Y113_A;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X13Y113_A1;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X13Y113_A2;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X13Y113_A3;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X13Y113_A4;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X13Y113_A5;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X13Y113_A6;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X13Y113_AMUX;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X13Y113_AO5;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X13Y113_AO6;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X13Y113_A_CY;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X13Y113_A_XOR;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X13Y113_B;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X13Y113_B1;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X13Y113_B2;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X13Y113_B3;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X13Y113_B4;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X13Y113_B5;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X13Y113_B6;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X13Y113_BO5;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X13Y113_BO6;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X13Y113_B_CY;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X13Y113_B_XOR;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X13Y113_C;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X13Y113_C1;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X13Y113_C2;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X13Y113_C3;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X13Y113_C4;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X13Y113_C5;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X13Y113_C6;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X13Y113_CMUX;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X13Y113_CO5;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X13Y113_CO6;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X13Y113_C_CY;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X13Y113_C_XOR;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X13Y113_D;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X13Y113_D1;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X13Y113_D2;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X13Y113_D3;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X13Y113_D4;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X13Y113_D5;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X13Y113_D6;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X13Y113_DO5;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X13Y113_DO6;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X13Y113_D_CY;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X13Y113_D_XOR;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X12Y114_A;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X12Y114_A1;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X12Y114_A2;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X12Y114_A3;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X12Y114_A4;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X12Y114_A5;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X12Y114_A6;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X12Y114_AMUX;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X12Y114_AO5;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X12Y114_AO6;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X12Y114_AQ;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X12Y114_AX;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X12Y114_A_CY;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X12Y114_A_XOR;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X12Y114_B;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X12Y114_B1;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X12Y114_B2;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X12Y114_B3;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X12Y114_B4;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X12Y114_B5;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X12Y114_B6;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X12Y114_BMUX;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X12Y114_BO5;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X12Y114_BO6;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X12Y114_B_CY;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X12Y114_B_XOR;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X12Y114_C;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X12Y114_C1;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X12Y114_C2;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X12Y114_C3;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X12Y114_C4;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X12Y114_C5;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X12Y114_C6;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X12Y114_CE;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X12Y114_CLK;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X12Y114_CO5;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X12Y114_CO6;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X12Y114_C_CY;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X12Y114_C_XOR;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X12Y114_D;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X12Y114_D1;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X12Y114_D2;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X12Y114_D3;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X12Y114_D4;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X12Y114_D5;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X12Y114_D6;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X12Y114_DO5;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X12Y114_DO6;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X12Y114_D_CY;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X12Y114_D_XOR;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X12Y114_SR;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X13Y114_A;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X13Y114_A1;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X13Y114_A2;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X13Y114_A3;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X13Y114_A4;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X13Y114_A5;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X13Y114_A5Q;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X13Y114_A6;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X13Y114_AMUX;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X13Y114_AO5;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X13Y114_AO6;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X13Y114_AQ;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X13Y114_AX;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X13Y114_A_CY;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X13Y114_A_XOR;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X13Y114_B;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X13Y114_B1;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X13Y114_B2;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X13Y114_B3;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X13Y114_B4;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X13Y114_B5;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X13Y114_B6;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X13Y114_BMUX;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X13Y114_BO5;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X13Y114_BO6;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X13Y114_B_CY;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X13Y114_B_XOR;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X13Y114_C;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X13Y114_C1;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X13Y114_C2;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X13Y114_C3;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X13Y114_C4;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X13Y114_C5;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X13Y114_C6;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X13Y114_CLK;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X13Y114_CO5;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X13Y114_CO6;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X13Y114_CQ;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X13Y114_C_CY;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X13Y114_C_XOR;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X13Y114_D;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X13Y114_D1;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X13Y114_D2;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X13Y114_D3;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X13Y114_D4;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X13Y114_D5;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X13Y114_D5Q;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X13Y114_D6;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X13Y114_DMUX;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X13Y114_DO5;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X13Y114_DO6;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X13Y114_DQ;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X13Y114_D_CY;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X13Y114_D_XOR;
  wire [0:0] CLBLM_L_X10Y115_SLICE_X12Y115_A;
  wire [0:0] CLBLM_L_X10Y115_SLICE_X12Y115_A1;
  wire [0:0] CLBLM_L_X10Y115_SLICE_X12Y115_A2;
  wire [0:0] CLBLM_L_X10Y115_SLICE_X12Y115_A3;
  wire [0:0] CLBLM_L_X10Y115_SLICE_X12Y115_A4;
  wire [0:0] CLBLM_L_X10Y115_SLICE_X12Y115_A5;
  wire [0:0] CLBLM_L_X10Y115_SLICE_X12Y115_A6;
  wire [0:0] CLBLM_L_X10Y115_SLICE_X12Y115_AO5;
  wire [0:0] CLBLM_L_X10Y115_SLICE_X12Y115_AO6;
  wire [0:0] CLBLM_L_X10Y115_SLICE_X12Y115_AQ;
  wire [0:0] CLBLM_L_X10Y115_SLICE_X12Y115_A_CY;
  wire [0:0] CLBLM_L_X10Y115_SLICE_X12Y115_A_XOR;
  wire [0:0] CLBLM_L_X10Y115_SLICE_X12Y115_B;
  wire [0:0] CLBLM_L_X10Y115_SLICE_X12Y115_B1;
  wire [0:0] CLBLM_L_X10Y115_SLICE_X12Y115_B2;
  wire [0:0] CLBLM_L_X10Y115_SLICE_X12Y115_B3;
  wire [0:0] CLBLM_L_X10Y115_SLICE_X12Y115_B4;
  wire [0:0] CLBLM_L_X10Y115_SLICE_X12Y115_B5;
  wire [0:0] CLBLM_L_X10Y115_SLICE_X12Y115_B6;
  wire [0:0] CLBLM_L_X10Y115_SLICE_X12Y115_BO5;
  wire [0:0] CLBLM_L_X10Y115_SLICE_X12Y115_BO6;
  wire [0:0] CLBLM_L_X10Y115_SLICE_X12Y115_BQ;
  wire [0:0] CLBLM_L_X10Y115_SLICE_X12Y115_B_CY;
  wire [0:0] CLBLM_L_X10Y115_SLICE_X12Y115_B_XOR;
  wire [0:0] CLBLM_L_X10Y115_SLICE_X12Y115_C;
  wire [0:0] CLBLM_L_X10Y115_SLICE_X12Y115_C1;
  wire [0:0] CLBLM_L_X10Y115_SLICE_X12Y115_C2;
  wire [0:0] CLBLM_L_X10Y115_SLICE_X12Y115_C3;
  wire [0:0] CLBLM_L_X10Y115_SLICE_X12Y115_C4;
  wire [0:0] CLBLM_L_X10Y115_SLICE_X12Y115_C5;
  wire [0:0] CLBLM_L_X10Y115_SLICE_X12Y115_C6;
  wire [0:0] CLBLM_L_X10Y115_SLICE_X12Y115_CLK;
  wire [0:0] CLBLM_L_X10Y115_SLICE_X12Y115_CO5;
  wire [0:0] CLBLM_L_X10Y115_SLICE_X12Y115_CO6;
  wire [0:0] CLBLM_L_X10Y115_SLICE_X12Y115_CQ;
  wire [0:0] CLBLM_L_X10Y115_SLICE_X12Y115_C_CY;
  wire [0:0] CLBLM_L_X10Y115_SLICE_X12Y115_C_XOR;
  wire [0:0] CLBLM_L_X10Y115_SLICE_X12Y115_D;
  wire [0:0] CLBLM_L_X10Y115_SLICE_X12Y115_D1;
  wire [0:0] CLBLM_L_X10Y115_SLICE_X12Y115_D2;
  wire [0:0] CLBLM_L_X10Y115_SLICE_X12Y115_D3;
  wire [0:0] CLBLM_L_X10Y115_SLICE_X12Y115_D4;
  wire [0:0] CLBLM_L_X10Y115_SLICE_X12Y115_D5;
  wire [0:0] CLBLM_L_X10Y115_SLICE_X12Y115_D6;
  wire [0:0] CLBLM_L_X10Y115_SLICE_X12Y115_DO5;
  wire [0:0] CLBLM_L_X10Y115_SLICE_X12Y115_DO6;
  wire [0:0] CLBLM_L_X10Y115_SLICE_X12Y115_DQ;
  wire [0:0] CLBLM_L_X10Y115_SLICE_X12Y115_D_CY;
  wire [0:0] CLBLM_L_X10Y115_SLICE_X12Y115_D_XOR;
  wire [0:0] CLBLM_L_X10Y115_SLICE_X13Y115_A;
  wire [0:0] CLBLM_L_X10Y115_SLICE_X13Y115_A1;
  wire [0:0] CLBLM_L_X10Y115_SLICE_X13Y115_A2;
  wire [0:0] CLBLM_L_X10Y115_SLICE_X13Y115_A3;
  wire [0:0] CLBLM_L_X10Y115_SLICE_X13Y115_A4;
  wire [0:0] CLBLM_L_X10Y115_SLICE_X13Y115_A5;
  wire [0:0] CLBLM_L_X10Y115_SLICE_X13Y115_A6;
  wire [0:0] CLBLM_L_X10Y115_SLICE_X13Y115_AMUX;
  wire [0:0] CLBLM_L_X10Y115_SLICE_X13Y115_AO5;
  wire [0:0] CLBLM_L_X10Y115_SLICE_X13Y115_AO6;
  wire [0:0] CLBLM_L_X10Y115_SLICE_X13Y115_A_CY;
  wire [0:0] CLBLM_L_X10Y115_SLICE_X13Y115_A_XOR;
  wire [0:0] CLBLM_L_X10Y115_SLICE_X13Y115_B;
  wire [0:0] CLBLM_L_X10Y115_SLICE_X13Y115_B1;
  wire [0:0] CLBLM_L_X10Y115_SLICE_X13Y115_B2;
  wire [0:0] CLBLM_L_X10Y115_SLICE_X13Y115_B3;
  wire [0:0] CLBLM_L_X10Y115_SLICE_X13Y115_B4;
  wire [0:0] CLBLM_L_X10Y115_SLICE_X13Y115_B5;
  wire [0:0] CLBLM_L_X10Y115_SLICE_X13Y115_B6;
  wire [0:0] CLBLM_L_X10Y115_SLICE_X13Y115_BO5;
  wire [0:0] CLBLM_L_X10Y115_SLICE_X13Y115_BO6;
  wire [0:0] CLBLM_L_X10Y115_SLICE_X13Y115_B_CY;
  wire [0:0] CLBLM_L_X10Y115_SLICE_X13Y115_B_XOR;
  wire [0:0] CLBLM_L_X10Y115_SLICE_X13Y115_C;
  wire [0:0] CLBLM_L_X10Y115_SLICE_X13Y115_C1;
  wire [0:0] CLBLM_L_X10Y115_SLICE_X13Y115_C2;
  wire [0:0] CLBLM_L_X10Y115_SLICE_X13Y115_C3;
  wire [0:0] CLBLM_L_X10Y115_SLICE_X13Y115_C4;
  wire [0:0] CLBLM_L_X10Y115_SLICE_X13Y115_C5;
  wire [0:0] CLBLM_L_X10Y115_SLICE_X13Y115_C6;
  wire [0:0] CLBLM_L_X10Y115_SLICE_X13Y115_CO5;
  wire [0:0] CLBLM_L_X10Y115_SLICE_X13Y115_CO6;
  wire [0:0] CLBLM_L_X10Y115_SLICE_X13Y115_C_CY;
  wire [0:0] CLBLM_L_X10Y115_SLICE_X13Y115_C_XOR;
  wire [0:0] CLBLM_L_X10Y115_SLICE_X13Y115_D;
  wire [0:0] CLBLM_L_X10Y115_SLICE_X13Y115_D1;
  wire [0:0] CLBLM_L_X10Y115_SLICE_X13Y115_D2;
  wire [0:0] CLBLM_L_X10Y115_SLICE_X13Y115_D3;
  wire [0:0] CLBLM_L_X10Y115_SLICE_X13Y115_D4;
  wire [0:0] CLBLM_L_X10Y115_SLICE_X13Y115_D5;
  wire [0:0] CLBLM_L_X10Y115_SLICE_X13Y115_D6;
  wire [0:0] CLBLM_L_X10Y115_SLICE_X13Y115_DO5;
  wire [0:0] CLBLM_L_X10Y115_SLICE_X13Y115_DO6;
  wire [0:0] CLBLM_L_X10Y115_SLICE_X13Y115_D_CY;
  wire [0:0] CLBLM_L_X10Y115_SLICE_X13Y115_D_XOR;
  wire [0:0] CLBLM_L_X10Y116_SLICE_X12Y116_A;
  wire [0:0] CLBLM_L_X10Y116_SLICE_X12Y116_A1;
  wire [0:0] CLBLM_L_X10Y116_SLICE_X12Y116_A2;
  wire [0:0] CLBLM_L_X10Y116_SLICE_X12Y116_A3;
  wire [0:0] CLBLM_L_X10Y116_SLICE_X12Y116_A4;
  wire [0:0] CLBLM_L_X10Y116_SLICE_X12Y116_A5;
  wire [0:0] CLBLM_L_X10Y116_SLICE_X12Y116_A5Q;
  wire [0:0] CLBLM_L_X10Y116_SLICE_X12Y116_A6;
  wire [0:0] CLBLM_L_X10Y116_SLICE_X12Y116_AMUX;
  wire [0:0] CLBLM_L_X10Y116_SLICE_X12Y116_AO5;
  wire [0:0] CLBLM_L_X10Y116_SLICE_X12Y116_AO6;
  wire [0:0] CLBLM_L_X10Y116_SLICE_X12Y116_AQ;
  wire [0:0] CLBLM_L_X10Y116_SLICE_X12Y116_AX;
  wire [0:0] CLBLM_L_X10Y116_SLICE_X12Y116_A_CY;
  wire [0:0] CLBLM_L_X10Y116_SLICE_X12Y116_A_XOR;
  wire [0:0] CLBLM_L_X10Y116_SLICE_X12Y116_B;
  wire [0:0] CLBLM_L_X10Y116_SLICE_X12Y116_B1;
  wire [0:0] CLBLM_L_X10Y116_SLICE_X12Y116_B2;
  wire [0:0] CLBLM_L_X10Y116_SLICE_X12Y116_B3;
  wire [0:0] CLBLM_L_X10Y116_SLICE_X12Y116_B4;
  wire [0:0] CLBLM_L_X10Y116_SLICE_X12Y116_B5;
  wire [0:0] CLBLM_L_X10Y116_SLICE_X12Y116_B6;
  wire [0:0] CLBLM_L_X10Y116_SLICE_X12Y116_BO5;
  wire [0:0] CLBLM_L_X10Y116_SLICE_X12Y116_BO6;
  wire [0:0] CLBLM_L_X10Y116_SLICE_X12Y116_BQ;
  wire [0:0] CLBLM_L_X10Y116_SLICE_X12Y116_B_CY;
  wire [0:0] CLBLM_L_X10Y116_SLICE_X12Y116_B_XOR;
  wire [0:0] CLBLM_L_X10Y116_SLICE_X12Y116_C;
  wire [0:0] CLBLM_L_X10Y116_SLICE_X12Y116_C1;
  wire [0:0] CLBLM_L_X10Y116_SLICE_X12Y116_C2;
  wire [0:0] CLBLM_L_X10Y116_SLICE_X12Y116_C3;
  wire [0:0] CLBLM_L_X10Y116_SLICE_X12Y116_C4;
  wire [0:0] CLBLM_L_X10Y116_SLICE_X12Y116_C5;
  wire [0:0] CLBLM_L_X10Y116_SLICE_X12Y116_C6;
  wire [0:0] CLBLM_L_X10Y116_SLICE_X12Y116_CLK;
  wire [0:0] CLBLM_L_X10Y116_SLICE_X12Y116_CO5;
  wire [0:0] CLBLM_L_X10Y116_SLICE_X12Y116_CO6;
  wire [0:0] CLBLM_L_X10Y116_SLICE_X12Y116_CQ;
  wire [0:0] CLBLM_L_X10Y116_SLICE_X12Y116_C_CY;
  wire [0:0] CLBLM_L_X10Y116_SLICE_X12Y116_C_XOR;
  wire [0:0] CLBLM_L_X10Y116_SLICE_X12Y116_D;
  wire [0:0] CLBLM_L_X10Y116_SLICE_X12Y116_D1;
  wire [0:0] CLBLM_L_X10Y116_SLICE_X12Y116_D2;
  wire [0:0] CLBLM_L_X10Y116_SLICE_X12Y116_D3;
  wire [0:0] CLBLM_L_X10Y116_SLICE_X12Y116_D4;
  wire [0:0] CLBLM_L_X10Y116_SLICE_X12Y116_D5;
  wire [0:0] CLBLM_L_X10Y116_SLICE_X12Y116_D6;
  wire [0:0] CLBLM_L_X10Y116_SLICE_X12Y116_DMUX;
  wire [0:0] CLBLM_L_X10Y116_SLICE_X12Y116_DO5;
  wire [0:0] CLBLM_L_X10Y116_SLICE_X12Y116_DO6;
  wire [0:0] CLBLM_L_X10Y116_SLICE_X12Y116_D_CY;
  wire [0:0] CLBLM_L_X10Y116_SLICE_X12Y116_D_XOR;
  wire [0:0] CLBLM_L_X10Y116_SLICE_X13Y116_A;
  wire [0:0] CLBLM_L_X10Y116_SLICE_X13Y116_A1;
  wire [0:0] CLBLM_L_X10Y116_SLICE_X13Y116_A2;
  wire [0:0] CLBLM_L_X10Y116_SLICE_X13Y116_A3;
  wire [0:0] CLBLM_L_X10Y116_SLICE_X13Y116_A4;
  wire [0:0] CLBLM_L_X10Y116_SLICE_X13Y116_A5;
  wire [0:0] CLBLM_L_X10Y116_SLICE_X13Y116_A6;
  wire [0:0] CLBLM_L_X10Y116_SLICE_X13Y116_AMUX;
  wire [0:0] CLBLM_L_X10Y116_SLICE_X13Y116_AO5;
  wire [0:0] CLBLM_L_X10Y116_SLICE_X13Y116_AO6;
  wire [0:0] CLBLM_L_X10Y116_SLICE_X13Y116_AQ;
  wire [0:0] CLBLM_L_X10Y116_SLICE_X13Y116_AX;
  wire [0:0] CLBLM_L_X10Y116_SLICE_X13Y116_A_CY;
  wire [0:0] CLBLM_L_X10Y116_SLICE_X13Y116_A_XOR;
  wire [0:0] CLBLM_L_X10Y116_SLICE_X13Y116_B;
  wire [0:0] CLBLM_L_X10Y116_SLICE_X13Y116_B1;
  wire [0:0] CLBLM_L_X10Y116_SLICE_X13Y116_B2;
  wire [0:0] CLBLM_L_X10Y116_SLICE_X13Y116_B3;
  wire [0:0] CLBLM_L_X10Y116_SLICE_X13Y116_B4;
  wire [0:0] CLBLM_L_X10Y116_SLICE_X13Y116_B5;
  wire [0:0] CLBLM_L_X10Y116_SLICE_X13Y116_B6;
  wire [0:0] CLBLM_L_X10Y116_SLICE_X13Y116_BMUX;
  wire [0:0] CLBLM_L_X10Y116_SLICE_X13Y116_BO5;
  wire [0:0] CLBLM_L_X10Y116_SLICE_X13Y116_BO6;
  wire [0:0] CLBLM_L_X10Y116_SLICE_X13Y116_BQ;
  wire [0:0] CLBLM_L_X10Y116_SLICE_X13Y116_B_CY;
  wire [0:0] CLBLM_L_X10Y116_SLICE_X13Y116_B_XOR;
  wire [0:0] CLBLM_L_X10Y116_SLICE_X13Y116_C;
  wire [0:0] CLBLM_L_X10Y116_SLICE_X13Y116_C1;
  wire [0:0] CLBLM_L_X10Y116_SLICE_X13Y116_C2;
  wire [0:0] CLBLM_L_X10Y116_SLICE_X13Y116_C3;
  wire [0:0] CLBLM_L_X10Y116_SLICE_X13Y116_C4;
  wire [0:0] CLBLM_L_X10Y116_SLICE_X13Y116_C5;
  wire [0:0] CLBLM_L_X10Y116_SLICE_X13Y116_C6;
  wire [0:0] CLBLM_L_X10Y116_SLICE_X13Y116_CLK;
  wire [0:0] CLBLM_L_X10Y116_SLICE_X13Y116_CMUX;
  wire [0:0] CLBLM_L_X10Y116_SLICE_X13Y116_CO5;
  wire [0:0] CLBLM_L_X10Y116_SLICE_X13Y116_CO6;
  wire [0:0] CLBLM_L_X10Y116_SLICE_X13Y116_CQ;
  wire [0:0] CLBLM_L_X10Y116_SLICE_X13Y116_C_CY;
  wire [0:0] CLBLM_L_X10Y116_SLICE_X13Y116_C_XOR;
  wire [0:0] CLBLM_L_X10Y116_SLICE_X13Y116_D;
  wire [0:0] CLBLM_L_X10Y116_SLICE_X13Y116_D1;
  wire [0:0] CLBLM_L_X10Y116_SLICE_X13Y116_D2;
  wire [0:0] CLBLM_L_X10Y116_SLICE_X13Y116_D3;
  wire [0:0] CLBLM_L_X10Y116_SLICE_X13Y116_D4;
  wire [0:0] CLBLM_L_X10Y116_SLICE_X13Y116_D5;
  wire [0:0] CLBLM_L_X10Y116_SLICE_X13Y116_D6;
  wire [0:0] CLBLM_L_X10Y116_SLICE_X13Y116_DO5;
  wire [0:0] CLBLM_L_X10Y116_SLICE_X13Y116_DO6;
  wire [0:0] CLBLM_L_X10Y116_SLICE_X13Y116_DQ;
  wire [0:0] CLBLM_L_X10Y116_SLICE_X13Y116_D_CY;
  wire [0:0] CLBLM_L_X10Y116_SLICE_X13Y116_D_XOR;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X12Y117_A;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X12Y117_A1;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X12Y117_A2;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X12Y117_A3;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X12Y117_A4;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X12Y117_A5;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X12Y117_A6;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X12Y117_AO5;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X12Y117_AO6;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X12Y117_AQ;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X12Y117_A_CY;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X12Y117_A_XOR;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X12Y117_B;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X12Y117_B1;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X12Y117_B2;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X12Y117_B3;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X12Y117_B4;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X12Y117_B5;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X12Y117_B6;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X12Y117_BO5;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X12Y117_BO6;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X12Y117_BQ;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X12Y117_B_CY;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X12Y117_B_XOR;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X12Y117_C;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X12Y117_C1;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X12Y117_C2;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X12Y117_C3;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X12Y117_C4;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X12Y117_C5;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X12Y117_C6;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X12Y117_CLK;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X12Y117_CO5;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X12Y117_CO6;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X12Y117_C_CY;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X12Y117_C_XOR;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X12Y117_D;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X12Y117_D1;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X12Y117_D2;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X12Y117_D3;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X12Y117_D4;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X12Y117_D5;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X12Y117_D6;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X12Y117_DO5;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X12Y117_DO6;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X12Y117_D_CY;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X12Y117_D_XOR;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X13Y117_A;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X13Y117_A1;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X13Y117_A2;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X13Y117_A3;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X13Y117_A4;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X13Y117_A5;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X13Y117_A6;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X13Y117_AO5;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X13Y117_AO6;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X13Y117_AQ;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X13Y117_A_CY;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X13Y117_A_XOR;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X13Y117_B;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X13Y117_B1;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X13Y117_B2;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X13Y117_B3;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X13Y117_B4;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X13Y117_B5;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X13Y117_B6;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X13Y117_BO5;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X13Y117_BO6;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X13Y117_BQ;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X13Y117_B_CY;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X13Y117_B_XOR;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X13Y117_C;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X13Y117_C1;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X13Y117_C2;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X13Y117_C3;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X13Y117_C4;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X13Y117_C5;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X13Y117_C6;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X13Y117_CLK;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X13Y117_CO5;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X13Y117_CO6;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X13Y117_CQ;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X13Y117_C_CY;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X13Y117_C_XOR;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X13Y117_D;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X13Y117_D1;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X13Y117_D2;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X13Y117_D3;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X13Y117_D4;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X13Y117_D5;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X13Y117_D6;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X13Y117_DO5;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X13Y117_DO6;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X13Y117_DQ;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X13Y117_D_CY;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X13Y117_D_XOR;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X12Y118_A;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X12Y118_A1;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X12Y118_A2;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X12Y118_A3;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X12Y118_A4;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X12Y118_A5;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X12Y118_A6;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X12Y118_AO5;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X12Y118_AO6;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X12Y118_AQ;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X12Y118_A_CY;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X12Y118_A_XOR;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X12Y118_B;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X12Y118_B1;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X12Y118_B2;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X12Y118_B3;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X12Y118_B4;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X12Y118_B5;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X12Y118_B5Q;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X12Y118_B6;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X12Y118_BMUX;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X12Y118_BO5;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X12Y118_BO6;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X12Y118_BQ;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X12Y118_B_CY;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X12Y118_B_XOR;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X12Y118_C;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X12Y118_C1;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X12Y118_C2;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X12Y118_C3;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X12Y118_C4;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X12Y118_C5;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X12Y118_C6;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X12Y118_CLK;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X12Y118_CO5;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X12Y118_CO6;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X12Y118_C_CY;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X12Y118_C_XOR;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X12Y118_D;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X12Y118_D1;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X12Y118_D2;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X12Y118_D3;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X12Y118_D4;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X12Y118_D5;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X12Y118_D6;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X12Y118_DO5;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X12Y118_DO6;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X12Y118_D_CY;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X12Y118_D_XOR;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X13Y118_A;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X13Y118_A1;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X13Y118_A2;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X13Y118_A3;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X13Y118_A4;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X13Y118_A5;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X13Y118_A6;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X13Y118_AO5;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X13Y118_AO6;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X13Y118_AQ;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X13Y118_A_CY;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X13Y118_A_XOR;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X13Y118_B;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X13Y118_B1;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X13Y118_B2;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X13Y118_B3;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X13Y118_B4;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X13Y118_B5;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X13Y118_B6;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X13Y118_BO5;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X13Y118_BO6;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X13Y118_BQ;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X13Y118_B_CY;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X13Y118_B_XOR;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X13Y118_C;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X13Y118_C1;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X13Y118_C2;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X13Y118_C3;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X13Y118_C4;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X13Y118_C5;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X13Y118_C6;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X13Y118_CLK;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X13Y118_CO5;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X13Y118_CO6;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X13Y118_CQ;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X13Y118_C_CY;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X13Y118_C_XOR;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X13Y118_D;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X13Y118_D1;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X13Y118_D2;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X13Y118_D3;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X13Y118_D4;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X13Y118_D5;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X13Y118_D6;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X13Y118_DO5;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X13Y118_DO6;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X13Y118_D_CY;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X13Y118_D_XOR;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X12Y119_A;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X12Y119_A1;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X12Y119_A2;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X12Y119_A3;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X12Y119_A4;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X12Y119_A5;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X12Y119_A6;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X12Y119_AO5;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X12Y119_AO6;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X12Y119_AQ;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X12Y119_A_CY;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X12Y119_A_XOR;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X12Y119_B;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X12Y119_B1;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X12Y119_B2;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X12Y119_B3;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X12Y119_B4;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X12Y119_B5;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X12Y119_B6;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X12Y119_BO5;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X12Y119_BO6;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X12Y119_BQ;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X12Y119_B_CY;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X12Y119_B_XOR;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X12Y119_C;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X12Y119_C1;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X12Y119_C2;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X12Y119_C3;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X12Y119_C4;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X12Y119_C5;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X12Y119_C6;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X12Y119_CLK;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X12Y119_CO5;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X12Y119_CO6;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X12Y119_CQ;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X12Y119_C_CY;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X12Y119_C_XOR;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X12Y119_D;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X12Y119_D1;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X12Y119_D2;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X12Y119_D3;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X12Y119_D4;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X12Y119_D5;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X12Y119_D6;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X12Y119_DO5;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X12Y119_DO6;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X12Y119_D_CY;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X12Y119_D_XOR;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X13Y119_A;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X13Y119_A1;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X13Y119_A2;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X13Y119_A3;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X13Y119_A4;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X13Y119_A5;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X13Y119_A6;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X13Y119_AO5;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X13Y119_AO6;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X13Y119_AQ;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X13Y119_A_CY;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X13Y119_A_XOR;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X13Y119_B;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X13Y119_B1;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X13Y119_B2;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X13Y119_B3;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X13Y119_B4;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X13Y119_B5;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X13Y119_B6;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X13Y119_BO5;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X13Y119_BO6;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X13Y119_BQ;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X13Y119_B_CY;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X13Y119_B_XOR;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X13Y119_C;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X13Y119_C1;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X13Y119_C2;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X13Y119_C3;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X13Y119_C4;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X13Y119_C5;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X13Y119_C6;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X13Y119_CLK;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X13Y119_CO5;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X13Y119_CO6;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X13Y119_CQ;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X13Y119_C_CY;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X13Y119_C_XOR;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X13Y119_D;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X13Y119_D1;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X13Y119_D2;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X13Y119_D3;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X13Y119_D4;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X13Y119_D5;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X13Y119_D6;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X13Y119_DO5;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X13Y119_DO6;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X13Y119_DQ;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X13Y119_D_CY;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X13Y119_D_XOR;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X12Y120_A;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X12Y120_A1;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X12Y120_A2;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X12Y120_A3;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X12Y120_A4;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X12Y120_A5;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X12Y120_A6;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X12Y120_AO5;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X12Y120_AO6;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X12Y120_AQ;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X12Y120_A_CY;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X12Y120_A_XOR;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X12Y120_B;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X12Y120_B1;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X12Y120_B2;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X12Y120_B3;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X12Y120_B4;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X12Y120_B5;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X12Y120_B6;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X12Y120_BO5;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X12Y120_BO6;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X12Y120_BQ;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X12Y120_B_CY;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X12Y120_B_XOR;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X12Y120_C;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X12Y120_C1;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X12Y120_C2;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X12Y120_C3;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X12Y120_C4;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X12Y120_C5;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X12Y120_C6;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X12Y120_CLK;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X12Y120_CO5;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X12Y120_CO6;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X12Y120_CQ;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X12Y120_C_CY;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X12Y120_C_XOR;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X12Y120_D;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X12Y120_D1;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X12Y120_D2;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X12Y120_D3;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X12Y120_D4;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X12Y120_D5;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X12Y120_D6;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X12Y120_DO5;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X12Y120_DO6;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X12Y120_DQ;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X12Y120_D_CY;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X12Y120_D_XOR;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X13Y120_A;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X13Y120_A1;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X13Y120_A2;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X13Y120_A3;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X13Y120_A4;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X13Y120_A5;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X13Y120_A5Q;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X13Y120_A6;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X13Y120_AMUX;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X13Y120_AO5;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X13Y120_AO6;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X13Y120_AQ;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X13Y120_AX;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X13Y120_A_CY;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X13Y120_A_XOR;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X13Y120_B;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X13Y120_B1;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X13Y120_B2;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X13Y120_B3;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X13Y120_B4;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X13Y120_B5;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X13Y120_B6;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X13Y120_BO5;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X13Y120_BO6;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X13Y120_BQ;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X13Y120_B_CY;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X13Y120_B_XOR;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X13Y120_C;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X13Y120_C1;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X13Y120_C2;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X13Y120_C3;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X13Y120_C4;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X13Y120_C5;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X13Y120_C6;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X13Y120_CLK;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X13Y120_CO5;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X13Y120_CO6;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X13Y120_C_CY;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X13Y120_C_XOR;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X13Y120_D;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X13Y120_D1;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X13Y120_D2;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X13Y120_D3;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X13Y120_D4;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X13Y120_D5;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X13Y120_D6;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X13Y120_DO5;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X13Y120_DO6;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X13Y120_D_CY;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X13Y120_D_XOR;
  wire [0:0] CLBLM_L_X10Y121_SLICE_X12Y121_A;
  wire [0:0] CLBLM_L_X10Y121_SLICE_X12Y121_A1;
  wire [0:0] CLBLM_L_X10Y121_SLICE_X12Y121_A2;
  wire [0:0] CLBLM_L_X10Y121_SLICE_X12Y121_A3;
  wire [0:0] CLBLM_L_X10Y121_SLICE_X12Y121_A4;
  wire [0:0] CLBLM_L_X10Y121_SLICE_X12Y121_A5;
  wire [0:0] CLBLM_L_X10Y121_SLICE_X12Y121_A6;
  wire [0:0] CLBLM_L_X10Y121_SLICE_X12Y121_AO5;
  wire [0:0] CLBLM_L_X10Y121_SLICE_X12Y121_AO6;
  wire [0:0] CLBLM_L_X10Y121_SLICE_X12Y121_AQ;
  wire [0:0] CLBLM_L_X10Y121_SLICE_X12Y121_A_CY;
  wire [0:0] CLBLM_L_X10Y121_SLICE_X12Y121_A_XOR;
  wire [0:0] CLBLM_L_X10Y121_SLICE_X12Y121_B;
  wire [0:0] CLBLM_L_X10Y121_SLICE_X12Y121_B1;
  wire [0:0] CLBLM_L_X10Y121_SLICE_X12Y121_B2;
  wire [0:0] CLBLM_L_X10Y121_SLICE_X12Y121_B3;
  wire [0:0] CLBLM_L_X10Y121_SLICE_X12Y121_B4;
  wire [0:0] CLBLM_L_X10Y121_SLICE_X12Y121_B5;
  wire [0:0] CLBLM_L_X10Y121_SLICE_X12Y121_B6;
  wire [0:0] CLBLM_L_X10Y121_SLICE_X12Y121_BO5;
  wire [0:0] CLBLM_L_X10Y121_SLICE_X12Y121_BO6;
  wire [0:0] CLBLM_L_X10Y121_SLICE_X12Y121_BQ;
  wire [0:0] CLBLM_L_X10Y121_SLICE_X12Y121_B_CY;
  wire [0:0] CLBLM_L_X10Y121_SLICE_X12Y121_B_XOR;
  wire [0:0] CLBLM_L_X10Y121_SLICE_X12Y121_C;
  wire [0:0] CLBLM_L_X10Y121_SLICE_X12Y121_C1;
  wire [0:0] CLBLM_L_X10Y121_SLICE_X12Y121_C2;
  wire [0:0] CLBLM_L_X10Y121_SLICE_X12Y121_C3;
  wire [0:0] CLBLM_L_X10Y121_SLICE_X12Y121_C4;
  wire [0:0] CLBLM_L_X10Y121_SLICE_X12Y121_C5;
  wire [0:0] CLBLM_L_X10Y121_SLICE_X12Y121_C6;
  wire [0:0] CLBLM_L_X10Y121_SLICE_X12Y121_CLK;
  wire [0:0] CLBLM_L_X10Y121_SLICE_X12Y121_CO5;
  wire [0:0] CLBLM_L_X10Y121_SLICE_X12Y121_CO6;
  wire [0:0] CLBLM_L_X10Y121_SLICE_X12Y121_C_CY;
  wire [0:0] CLBLM_L_X10Y121_SLICE_X12Y121_C_XOR;
  wire [0:0] CLBLM_L_X10Y121_SLICE_X12Y121_D;
  wire [0:0] CLBLM_L_X10Y121_SLICE_X12Y121_D1;
  wire [0:0] CLBLM_L_X10Y121_SLICE_X12Y121_D2;
  wire [0:0] CLBLM_L_X10Y121_SLICE_X12Y121_D3;
  wire [0:0] CLBLM_L_X10Y121_SLICE_X12Y121_D4;
  wire [0:0] CLBLM_L_X10Y121_SLICE_X12Y121_D5;
  wire [0:0] CLBLM_L_X10Y121_SLICE_X12Y121_D6;
  wire [0:0] CLBLM_L_X10Y121_SLICE_X12Y121_DO5;
  wire [0:0] CLBLM_L_X10Y121_SLICE_X12Y121_DO6;
  wire [0:0] CLBLM_L_X10Y121_SLICE_X12Y121_D_CY;
  wire [0:0] CLBLM_L_X10Y121_SLICE_X12Y121_D_XOR;
  wire [0:0] CLBLM_L_X10Y121_SLICE_X13Y121_A;
  wire [0:0] CLBLM_L_X10Y121_SLICE_X13Y121_A1;
  wire [0:0] CLBLM_L_X10Y121_SLICE_X13Y121_A2;
  wire [0:0] CLBLM_L_X10Y121_SLICE_X13Y121_A3;
  wire [0:0] CLBLM_L_X10Y121_SLICE_X13Y121_A4;
  wire [0:0] CLBLM_L_X10Y121_SLICE_X13Y121_A5;
  wire [0:0] CLBLM_L_X10Y121_SLICE_X13Y121_A6;
  wire [0:0] CLBLM_L_X10Y121_SLICE_X13Y121_AO5;
  wire [0:0] CLBLM_L_X10Y121_SLICE_X13Y121_AO6;
  wire [0:0] CLBLM_L_X10Y121_SLICE_X13Y121_AQ;
  wire [0:0] CLBLM_L_X10Y121_SLICE_X13Y121_A_CY;
  wire [0:0] CLBLM_L_X10Y121_SLICE_X13Y121_A_XOR;
  wire [0:0] CLBLM_L_X10Y121_SLICE_X13Y121_B;
  wire [0:0] CLBLM_L_X10Y121_SLICE_X13Y121_B1;
  wire [0:0] CLBLM_L_X10Y121_SLICE_X13Y121_B2;
  wire [0:0] CLBLM_L_X10Y121_SLICE_X13Y121_B3;
  wire [0:0] CLBLM_L_X10Y121_SLICE_X13Y121_B4;
  wire [0:0] CLBLM_L_X10Y121_SLICE_X13Y121_B5;
  wire [0:0] CLBLM_L_X10Y121_SLICE_X13Y121_B6;
  wire [0:0] CLBLM_L_X10Y121_SLICE_X13Y121_BO5;
  wire [0:0] CLBLM_L_X10Y121_SLICE_X13Y121_BO6;
  wire [0:0] CLBLM_L_X10Y121_SLICE_X13Y121_BQ;
  wire [0:0] CLBLM_L_X10Y121_SLICE_X13Y121_B_CY;
  wire [0:0] CLBLM_L_X10Y121_SLICE_X13Y121_B_XOR;
  wire [0:0] CLBLM_L_X10Y121_SLICE_X13Y121_C;
  wire [0:0] CLBLM_L_X10Y121_SLICE_X13Y121_C1;
  wire [0:0] CLBLM_L_X10Y121_SLICE_X13Y121_C2;
  wire [0:0] CLBLM_L_X10Y121_SLICE_X13Y121_C3;
  wire [0:0] CLBLM_L_X10Y121_SLICE_X13Y121_C4;
  wire [0:0] CLBLM_L_X10Y121_SLICE_X13Y121_C5;
  wire [0:0] CLBLM_L_X10Y121_SLICE_X13Y121_C6;
  wire [0:0] CLBLM_L_X10Y121_SLICE_X13Y121_CLK;
  wire [0:0] CLBLM_L_X10Y121_SLICE_X13Y121_CO5;
  wire [0:0] CLBLM_L_X10Y121_SLICE_X13Y121_CO6;
  wire [0:0] CLBLM_L_X10Y121_SLICE_X13Y121_CQ;
  wire [0:0] CLBLM_L_X10Y121_SLICE_X13Y121_C_CY;
  wire [0:0] CLBLM_L_X10Y121_SLICE_X13Y121_C_XOR;
  wire [0:0] CLBLM_L_X10Y121_SLICE_X13Y121_D;
  wire [0:0] CLBLM_L_X10Y121_SLICE_X13Y121_D1;
  wire [0:0] CLBLM_L_X10Y121_SLICE_X13Y121_D2;
  wire [0:0] CLBLM_L_X10Y121_SLICE_X13Y121_D3;
  wire [0:0] CLBLM_L_X10Y121_SLICE_X13Y121_D4;
  wire [0:0] CLBLM_L_X10Y121_SLICE_X13Y121_D5;
  wire [0:0] CLBLM_L_X10Y121_SLICE_X13Y121_D6;
  wire [0:0] CLBLM_L_X10Y121_SLICE_X13Y121_DO5;
  wire [0:0] CLBLM_L_X10Y121_SLICE_X13Y121_DO6;
  wire [0:0] CLBLM_L_X10Y121_SLICE_X13Y121_D_CY;
  wire [0:0] CLBLM_L_X10Y121_SLICE_X13Y121_D_XOR;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X12Y122_A;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X12Y122_A1;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X12Y122_A2;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X12Y122_A3;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X12Y122_A4;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X12Y122_A5;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X12Y122_A6;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X12Y122_AO5;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X12Y122_AO6;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X12Y122_AQ;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X12Y122_A_CY;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X12Y122_A_XOR;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X12Y122_B;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X12Y122_B1;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X12Y122_B2;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X12Y122_B3;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X12Y122_B4;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X12Y122_B5;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X12Y122_B6;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X12Y122_BO5;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X12Y122_BO6;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X12Y122_BQ;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X12Y122_B_CY;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X12Y122_B_XOR;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X12Y122_C;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X12Y122_C1;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X12Y122_C2;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X12Y122_C3;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X12Y122_C4;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X12Y122_C5;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X12Y122_C6;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X12Y122_CLK;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X12Y122_CMUX;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X12Y122_CO5;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X12Y122_CO6;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X12Y122_C_CY;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X12Y122_C_XOR;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X12Y122_D;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X12Y122_D1;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X12Y122_D2;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X12Y122_D3;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X12Y122_D4;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X12Y122_D5;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X12Y122_D6;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X12Y122_DO5;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X12Y122_DO6;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X12Y122_D_CY;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X12Y122_D_XOR;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X13Y122_A;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X13Y122_A1;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X13Y122_A2;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X13Y122_A3;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X13Y122_A4;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X13Y122_A5;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X13Y122_A5Q;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X13Y122_A6;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X13Y122_AMUX;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X13Y122_AO5;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X13Y122_AO6;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X13Y122_AQ;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X13Y122_AX;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X13Y122_A_CY;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X13Y122_A_XOR;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X13Y122_B;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X13Y122_B1;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X13Y122_B2;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X13Y122_B3;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X13Y122_B4;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X13Y122_B5;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X13Y122_B6;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X13Y122_BO5;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X13Y122_BO6;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X13Y122_BQ;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X13Y122_B_CY;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X13Y122_B_XOR;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X13Y122_C;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X13Y122_C1;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X13Y122_C2;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X13Y122_C3;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X13Y122_C4;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X13Y122_C5;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X13Y122_C6;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X13Y122_CLK;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X13Y122_CO5;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X13Y122_CO6;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X13Y122_CQ;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X13Y122_C_CY;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X13Y122_C_XOR;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X13Y122_D;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X13Y122_D1;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X13Y122_D2;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X13Y122_D3;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X13Y122_D4;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X13Y122_D5;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X13Y122_D6;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X13Y122_DMUX;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X13Y122_DO5;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X13Y122_DO6;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X13Y122_D_CY;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X13Y122_D_XOR;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X12Y123_A;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X12Y123_A1;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X12Y123_A2;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X12Y123_A3;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X12Y123_A4;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X12Y123_A5;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X12Y123_A6;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X12Y123_AMUX;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X12Y123_AO5;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X12Y123_AO6;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X12Y123_A_CY;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X12Y123_A_XOR;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X12Y123_B;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X12Y123_B1;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X12Y123_B2;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X12Y123_B3;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X12Y123_B4;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X12Y123_B5;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X12Y123_B6;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X12Y123_BO5;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X12Y123_BO6;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X12Y123_B_CY;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X12Y123_B_XOR;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X12Y123_C;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X12Y123_C1;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X12Y123_C2;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X12Y123_C3;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X12Y123_C4;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X12Y123_C5;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X12Y123_C6;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X12Y123_CMUX;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X12Y123_CO5;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X12Y123_CO6;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X12Y123_C_CY;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X12Y123_C_XOR;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X12Y123_D;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X12Y123_D1;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X12Y123_D2;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X12Y123_D3;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X12Y123_D4;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X12Y123_D5;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X12Y123_D6;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X12Y123_DO5;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X12Y123_DO6;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X12Y123_D_CY;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X12Y123_D_XOR;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X13Y123_A;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X13Y123_A1;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X13Y123_A2;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X13Y123_A3;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X13Y123_A4;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X13Y123_A5;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X13Y123_A6;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X13Y123_AO5;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X13Y123_AO6;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X13Y123_AQ;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X13Y123_A_CY;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X13Y123_A_XOR;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X13Y123_B;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X13Y123_B1;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X13Y123_B2;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X13Y123_B3;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X13Y123_B4;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X13Y123_B5;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X13Y123_B6;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X13Y123_BO5;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X13Y123_BO6;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X13Y123_B_CY;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X13Y123_B_XOR;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X13Y123_C;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X13Y123_C1;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X13Y123_C2;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X13Y123_C3;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X13Y123_C4;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X13Y123_C5;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X13Y123_C6;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X13Y123_CLK;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X13Y123_CO5;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X13Y123_CO6;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X13Y123_C_CY;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X13Y123_C_XOR;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X13Y123_D;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X13Y123_D1;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X13Y123_D2;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X13Y123_D3;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X13Y123_D4;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X13Y123_D5;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X13Y123_D6;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X13Y123_DO5;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X13Y123_DO6;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X13Y123_D_CY;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X13Y123_D_XOR;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X12Y124_A;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X12Y124_A1;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X12Y124_A2;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X12Y124_A3;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X12Y124_A4;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X12Y124_A5;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X12Y124_A6;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X12Y124_AO5;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X12Y124_AO6;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X12Y124_AQ;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X12Y124_A_CY;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X12Y124_A_XOR;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X12Y124_B;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X12Y124_B1;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X12Y124_B2;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X12Y124_B3;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X12Y124_B4;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X12Y124_B5;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X12Y124_B6;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X12Y124_BO5;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X12Y124_BO6;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X12Y124_B_CY;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X12Y124_B_XOR;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X12Y124_C;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X12Y124_C1;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X12Y124_C2;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X12Y124_C3;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X12Y124_C4;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X12Y124_C5;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X12Y124_C6;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X12Y124_CLK;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X12Y124_CO5;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X12Y124_CO6;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X12Y124_C_CY;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X12Y124_C_XOR;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X12Y124_D;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X12Y124_D1;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X12Y124_D2;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X12Y124_D3;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X12Y124_D4;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X12Y124_D5;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X12Y124_D6;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X12Y124_DO5;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X12Y124_DO6;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X12Y124_D_CY;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X12Y124_D_XOR;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X13Y124_A;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X13Y124_A1;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X13Y124_A2;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X13Y124_A3;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X13Y124_A4;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X13Y124_A5;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X13Y124_A6;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X13Y124_AMUX;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X13Y124_AO5;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X13Y124_AO6;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X13Y124_AQ;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X13Y124_AX;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X13Y124_A_CY;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X13Y124_A_XOR;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X13Y124_B;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X13Y124_B1;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X13Y124_B2;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X13Y124_B3;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X13Y124_B4;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X13Y124_B5;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X13Y124_B6;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X13Y124_BMUX;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X13Y124_BO5;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X13Y124_BO6;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X13Y124_B_CY;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X13Y124_B_XOR;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X13Y124_C;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X13Y124_C1;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X13Y124_C2;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X13Y124_C3;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X13Y124_C4;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X13Y124_C5;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X13Y124_C6;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X13Y124_CE;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X13Y124_CLK;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X13Y124_CMUX;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X13Y124_CO5;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X13Y124_CO6;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X13Y124_C_CY;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X13Y124_C_XOR;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X13Y124_D;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X13Y124_D1;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X13Y124_D2;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X13Y124_D3;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X13Y124_D4;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X13Y124_D5;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X13Y124_D6;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X13Y124_DO5;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X13Y124_DO6;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X13Y124_D_CY;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X13Y124_D_XOR;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X13Y124_SR;
  wire [0:0] CLBLM_L_X10Y126_SLICE_X12Y126_A;
  wire [0:0] CLBLM_L_X10Y126_SLICE_X12Y126_A1;
  wire [0:0] CLBLM_L_X10Y126_SLICE_X12Y126_A2;
  wire [0:0] CLBLM_L_X10Y126_SLICE_X12Y126_A3;
  wire [0:0] CLBLM_L_X10Y126_SLICE_X12Y126_A4;
  wire [0:0] CLBLM_L_X10Y126_SLICE_X12Y126_A5;
  wire [0:0] CLBLM_L_X10Y126_SLICE_X12Y126_A6;
  wire [0:0] CLBLM_L_X10Y126_SLICE_X12Y126_AO5;
  wire [0:0] CLBLM_L_X10Y126_SLICE_X12Y126_AO6;
  wire [0:0] CLBLM_L_X10Y126_SLICE_X12Y126_AQ;
  wire [0:0] CLBLM_L_X10Y126_SLICE_X12Y126_AX;
  wire [0:0] CLBLM_L_X10Y126_SLICE_X12Y126_A_CY;
  wire [0:0] CLBLM_L_X10Y126_SLICE_X12Y126_A_XOR;
  wire [0:0] CLBLM_L_X10Y126_SLICE_X12Y126_B;
  wire [0:0] CLBLM_L_X10Y126_SLICE_X12Y126_B1;
  wire [0:0] CLBLM_L_X10Y126_SLICE_X12Y126_B2;
  wire [0:0] CLBLM_L_X10Y126_SLICE_X12Y126_B3;
  wire [0:0] CLBLM_L_X10Y126_SLICE_X12Y126_B4;
  wire [0:0] CLBLM_L_X10Y126_SLICE_X12Y126_B5;
  wire [0:0] CLBLM_L_X10Y126_SLICE_X12Y126_B6;
  wire [0:0] CLBLM_L_X10Y126_SLICE_X12Y126_BO5;
  wire [0:0] CLBLM_L_X10Y126_SLICE_X12Y126_BO6;
  wire [0:0] CLBLM_L_X10Y126_SLICE_X12Y126_B_CY;
  wire [0:0] CLBLM_L_X10Y126_SLICE_X12Y126_B_XOR;
  wire [0:0] CLBLM_L_X10Y126_SLICE_X12Y126_C;
  wire [0:0] CLBLM_L_X10Y126_SLICE_X12Y126_C1;
  wire [0:0] CLBLM_L_X10Y126_SLICE_X12Y126_C2;
  wire [0:0] CLBLM_L_X10Y126_SLICE_X12Y126_C3;
  wire [0:0] CLBLM_L_X10Y126_SLICE_X12Y126_C4;
  wire [0:0] CLBLM_L_X10Y126_SLICE_X12Y126_C5;
  wire [0:0] CLBLM_L_X10Y126_SLICE_X12Y126_C6;
  wire [0:0] CLBLM_L_X10Y126_SLICE_X12Y126_CLK;
  wire [0:0] CLBLM_L_X10Y126_SLICE_X12Y126_CO5;
  wire [0:0] CLBLM_L_X10Y126_SLICE_X12Y126_CO6;
  wire [0:0] CLBLM_L_X10Y126_SLICE_X12Y126_C_CY;
  wire [0:0] CLBLM_L_X10Y126_SLICE_X12Y126_C_XOR;
  wire [0:0] CLBLM_L_X10Y126_SLICE_X12Y126_D;
  wire [0:0] CLBLM_L_X10Y126_SLICE_X12Y126_D1;
  wire [0:0] CLBLM_L_X10Y126_SLICE_X12Y126_D2;
  wire [0:0] CLBLM_L_X10Y126_SLICE_X12Y126_D3;
  wire [0:0] CLBLM_L_X10Y126_SLICE_X12Y126_D4;
  wire [0:0] CLBLM_L_X10Y126_SLICE_X12Y126_D5;
  wire [0:0] CLBLM_L_X10Y126_SLICE_X12Y126_D6;
  wire [0:0] CLBLM_L_X10Y126_SLICE_X12Y126_DO5;
  wire [0:0] CLBLM_L_X10Y126_SLICE_X12Y126_DO6;
  wire [0:0] CLBLM_L_X10Y126_SLICE_X12Y126_D_CY;
  wire [0:0] CLBLM_L_X10Y126_SLICE_X12Y126_D_XOR;
  wire [0:0] CLBLM_L_X10Y126_SLICE_X13Y126_A;
  wire [0:0] CLBLM_L_X10Y126_SLICE_X13Y126_A1;
  wire [0:0] CLBLM_L_X10Y126_SLICE_X13Y126_A2;
  wire [0:0] CLBLM_L_X10Y126_SLICE_X13Y126_A3;
  wire [0:0] CLBLM_L_X10Y126_SLICE_X13Y126_A4;
  wire [0:0] CLBLM_L_X10Y126_SLICE_X13Y126_A5;
  wire [0:0] CLBLM_L_X10Y126_SLICE_X13Y126_A6;
  wire [0:0] CLBLM_L_X10Y126_SLICE_X13Y126_AO5;
  wire [0:0] CLBLM_L_X10Y126_SLICE_X13Y126_AO6;
  wire [0:0] CLBLM_L_X10Y126_SLICE_X13Y126_A_CY;
  wire [0:0] CLBLM_L_X10Y126_SLICE_X13Y126_A_XOR;
  wire [0:0] CLBLM_L_X10Y126_SLICE_X13Y126_B;
  wire [0:0] CLBLM_L_X10Y126_SLICE_X13Y126_B1;
  wire [0:0] CLBLM_L_X10Y126_SLICE_X13Y126_B2;
  wire [0:0] CLBLM_L_X10Y126_SLICE_X13Y126_B3;
  wire [0:0] CLBLM_L_X10Y126_SLICE_X13Y126_B4;
  wire [0:0] CLBLM_L_X10Y126_SLICE_X13Y126_B5;
  wire [0:0] CLBLM_L_X10Y126_SLICE_X13Y126_B6;
  wire [0:0] CLBLM_L_X10Y126_SLICE_X13Y126_BO5;
  wire [0:0] CLBLM_L_X10Y126_SLICE_X13Y126_BO6;
  wire [0:0] CLBLM_L_X10Y126_SLICE_X13Y126_B_CY;
  wire [0:0] CLBLM_L_X10Y126_SLICE_X13Y126_B_XOR;
  wire [0:0] CLBLM_L_X10Y126_SLICE_X13Y126_C;
  wire [0:0] CLBLM_L_X10Y126_SLICE_X13Y126_C1;
  wire [0:0] CLBLM_L_X10Y126_SLICE_X13Y126_C2;
  wire [0:0] CLBLM_L_X10Y126_SLICE_X13Y126_C3;
  wire [0:0] CLBLM_L_X10Y126_SLICE_X13Y126_C4;
  wire [0:0] CLBLM_L_X10Y126_SLICE_X13Y126_C5;
  wire [0:0] CLBLM_L_X10Y126_SLICE_X13Y126_C6;
  wire [0:0] CLBLM_L_X10Y126_SLICE_X13Y126_CO5;
  wire [0:0] CLBLM_L_X10Y126_SLICE_X13Y126_CO6;
  wire [0:0] CLBLM_L_X10Y126_SLICE_X13Y126_C_CY;
  wire [0:0] CLBLM_L_X10Y126_SLICE_X13Y126_C_XOR;
  wire [0:0] CLBLM_L_X10Y126_SLICE_X13Y126_D;
  wire [0:0] CLBLM_L_X10Y126_SLICE_X13Y126_D1;
  wire [0:0] CLBLM_L_X10Y126_SLICE_X13Y126_D2;
  wire [0:0] CLBLM_L_X10Y126_SLICE_X13Y126_D3;
  wire [0:0] CLBLM_L_X10Y126_SLICE_X13Y126_D4;
  wire [0:0] CLBLM_L_X10Y126_SLICE_X13Y126_D5;
  wire [0:0] CLBLM_L_X10Y126_SLICE_X13Y126_D6;
  wire [0:0] CLBLM_L_X10Y126_SLICE_X13Y126_DO5;
  wire [0:0] CLBLM_L_X10Y126_SLICE_X13Y126_DO6;
  wire [0:0] CLBLM_L_X10Y126_SLICE_X13Y126_D_CY;
  wire [0:0] CLBLM_L_X10Y126_SLICE_X13Y126_D_XOR;
  wire [0:0] CLBLM_L_X10Y127_SLICE_X12Y127_A;
  wire [0:0] CLBLM_L_X10Y127_SLICE_X12Y127_A1;
  wire [0:0] CLBLM_L_X10Y127_SLICE_X12Y127_A2;
  wire [0:0] CLBLM_L_X10Y127_SLICE_X12Y127_A3;
  wire [0:0] CLBLM_L_X10Y127_SLICE_X12Y127_A4;
  wire [0:0] CLBLM_L_X10Y127_SLICE_X12Y127_A5;
  wire [0:0] CLBLM_L_X10Y127_SLICE_X12Y127_A6;
  wire [0:0] CLBLM_L_X10Y127_SLICE_X12Y127_AO5;
  wire [0:0] CLBLM_L_X10Y127_SLICE_X12Y127_AO6;
  wire [0:0] CLBLM_L_X10Y127_SLICE_X12Y127_AQ;
  wire [0:0] CLBLM_L_X10Y127_SLICE_X12Y127_AX;
  wire [0:0] CLBLM_L_X10Y127_SLICE_X12Y127_A_CY;
  wire [0:0] CLBLM_L_X10Y127_SLICE_X12Y127_A_XOR;
  wire [0:0] CLBLM_L_X10Y127_SLICE_X12Y127_B;
  wire [0:0] CLBLM_L_X10Y127_SLICE_X12Y127_B1;
  wire [0:0] CLBLM_L_X10Y127_SLICE_X12Y127_B2;
  wire [0:0] CLBLM_L_X10Y127_SLICE_X12Y127_B3;
  wire [0:0] CLBLM_L_X10Y127_SLICE_X12Y127_B4;
  wire [0:0] CLBLM_L_X10Y127_SLICE_X12Y127_B5;
  wire [0:0] CLBLM_L_X10Y127_SLICE_X12Y127_B6;
  wire [0:0] CLBLM_L_X10Y127_SLICE_X12Y127_BO5;
  wire [0:0] CLBLM_L_X10Y127_SLICE_X12Y127_BO6;
  wire [0:0] CLBLM_L_X10Y127_SLICE_X12Y127_B_CY;
  wire [0:0] CLBLM_L_X10Y127_SLICE_X12Y127_B_XOR;
  wire [0:0] CLBLM_L_X10Y127_SLICE_X12Y127_C;
  wire [0:0] CLBLM_L_X10Y127_SLICE_X12Y127_C1;
  wire [0:0] CLBLM_L_X10Y127_SLICE_X12Y127_C2;
  wire [0:0] CLBLM_L_X10Y127_SLICE_X12Y127_C3;
  wire [0:0] CLBLM_L_X10Y127_SLICE_X12Y127_C4;
  wire [0:0] CLBLM_L_X10Y127_SLICE_X12Y127_C5;
  wire [0:0] CLBLM_L_X10Y127_SLICE_X12Y127_C6;
  wire [0:0] CLBLM_L_X10Y127_SLICE_X12Y127_CLK;
  wire [0:0] CLBLM_L_X10Y127_SLICE_X12Y127_CO5;
  wire [0:0] CLBLM_L_X10Y127_SLICE_X12Y127_CO6;
  wire [0:0] CLBLM_L_X10Y127_SLICE_X12Y127_C_CY;
  wire [0:0] CLBLM_L_X10Y127_SLICE_X12Y127_C_XOR;
  wire [0:0] CLBLM_L_X10Y127_SLICE_X12Y127_D;
  wire [0:0] CLBLM_L_X10Y127_SLICE_X12Y127_D1;
  wire [0:0] CLBLM_L_X10Y127_SLICE_X12Y127_D2;
  wire [0:0] CLBLM_L_X10Y127_SLICE_X12Y127_D3;
  wire [0:0] CLBLM_L_X10Y127_SLICE_X12Y127_D4;
  wire [0:0] CLBLM_L_X10Y127_SLICE_X12Y127_D5;
  wire [0:0] CLBLM_L_X10Y127_SLICE_X12Y127_D6;
  wire [0:0] CLBLM_L_X10Y127_SLICE_X12Y127_DO5;
  wire [0:0] CLBLM_L_X10Y127_SLICE_X12Y127_DO6;
  wire [0:0] CLBLM_L_X10Y127_SLICE_X12Y127_D_CY;
  wire [0:0] CLBLM_L_X10Y127_SLICE_X12Y127_D_XOR;
  wire [0:0] CLBLM_L_X10Y127_SLICE_X13Y127_A;
  wire [0:0] CLBLM_L_X10Y127_SLICE_X13Y127_A1;
  wire [0:0] CLBLM_L_X10Y127_SLICE_X13Y127_A2;
  wire [0:0] CLBLM_L_X10Y127_SLICE_X13Y127_A3;
  wire [0:0] CLBLM_L_X10Y127_SLICE_X13Y127_A4;
  wire [0:0] CLBLM_L_X10Y127_SLICE_X13Y127_A5;
  wire [0:0] CLBLM_L_X10Y127_SLICE_X13Y127_A6;
  wire [0:0] CLBLM_L_X10Y127_SLICE_X13Y127_AO5;
  wire [0:0] CLBLM_L_X10Y127_SLICE_X13Y127_AO6;
  wire [0:0] CLBLM_L_X10Y127_SLICE_X13Y127_A_CY;
  wire [0:0] CLBLM_L_X10Y127_SLICE_X13Y127_A_XOR;
  wire [0:0] CLBLM_L_X10Y127_SLICE_X13Y127_B;
  wire [0:0] CLBLM_L_X10Y127_SLICE_X13Y127_B1;
  wire [0:0] CLBLM_L_X10Y127_SLICE_X13Y127_B2;
  wire [0:0] CLBLM_L_X10Y127_SLICE_X13Y127_B3;
  wire [0:0] CLBLM_L_X10Y127_SLICE_X13Y127_B4;
  wire [0:0] CLBLM_L_X10Y127_SLICE_X13Y127_B5;
  wire [0:0] CLBLM_L_X10Y127_SLICE_X13Y127_B6;
  wire [0:0] CLBLM_L_X10Y127_SLICE_X13Y127_BO5;
  wire [0:0] CLBLM_L_X10Y127_SLICE_X13Y127_BO6;
  wire [0:0] CLBLM_L_X10Y127_SLICE_X13Y127_B_CY;
  wire [0:0] CLBLM_L_X10Y127_SLICE_X13Y127_B_XOR;
  wire [0:0] CLBLM_L_X10Y127_SLICE_X13Y127_C;
  wire [0:0] CLBLM_L_X10Y127_SLICE_X13Y127_C1;
  wire [0:0] CLBLM_L_X10Y127_SLICE_X13Y127_C2;
  wire [0:0] CLBLM_L_X10Y127_SLICE_X13Y127_C3;
  wire [0:0] CLBLM_L_X10Y127_SLICE_X13Y127_C4;
  wire [0:0] CLBLM_L_X10Y127_SLICE_X13Y127_C5;
  wire [0:0] CLBLM_L_X10Y127_SLICE_X13Y127_C6;
  wire [0:0] CLBLM_L_X10Y127_SLICE_X13Y127_CO5;
  wire [0:0] CLBLM_L_X10Y127_SLICE_X13Y127_CO6;
  wire [0:0] CLBLM_L_X10Y127_SLICE_X13Y127_C_CY;
  wire [0:0] CLBLM_L_X10Y127_SLICE_X13Y127_C_XOR;
  wire [0:0] CLBLM_L_X10Y127_SLICE_X13Y127_D;
  wire [0:0] CLBLM_L_X10Y127_SLICE_X13Y127_D1;
  wire [0:0] CLBLM_L_X10Y127_SLICE_X13Y127_D2;
  wire [0:0] CLBLM_L_X10Y127_SLICE_X13Y127_D3;
  wire [0:0] CLBLM_L_X10Y127_SLICE_X13Y127_D4;
  wire [0:0] CLBLM_L_X10Y127_SLICE_X13Y127_D5;
  wire [0:0] CLBLM_L_X10Y127_SLICE_X13Y127_D6;
  wire [0:0] CLBLM_L_X10Y127_SLICE_X13Y127_DO5;
  wire [0:0] CLBLM_L_X10Y127_SLICE_X13Y127_DO6;
  wire [0:0] CLBLM_L_X10Y127_SLICE_X13Y127_D_CY;
  wire [0:0] CLBLM_L_X10Y127_SLICE_X13Y127_D_XOR;
  wire [0:0] CLBLM_L_X10Y128_SLICE_X12Y128_A;
  wire [0:0] CLBLM_L_X10Y128_SLICE_X12Y128_A1;
  wire [0:0] CLBLM_L_X10Y128_SLICE_X12Y128_A2;
  wire [0:0] CLBLM_L_X10Y128_SLICE_X12Y128_A3;
  wire [0:0] CLBLM_L_X10Y128_SLICE_X12Y128_A4;
  wire [0:0] CLBLM_L_X10Y128_SLICE_X12Y128_A5;
  wire [0:0] CLBLM_L_X10Y128_SLICE_X12Y128_A6;
  wire [0:0] CLBLM_L_X10Y128_SLICE_X12Y128_AO5;
  wire [0:0] CLBLM_L_X10Y128_SLICE_X12Y128_AO6;
  wire [0:0] CLBLM_L_X10Y128_SLICE_X12Y128_A_CY;
  wire [0:0] CLBLM_L_X10Y128_SLICE_X12Y128_A_XOR;
  wire [0:0] CLBLM_L_X10Y128_SLICE_X12Y128_B;
  wire [0:0] CLBLM_L_X10Y128_SLICE_X12Y128_B1;
  wire [0:0] CLBLM_L_X10Y128_SLICE_X12Y128_B2;
  wire [0:0] CLBLM_L_X10Y128_SLICE_X12Y128_B3;
  wire [0:0] CLBLM_L_X10Y128_SLICE_X12Y128_B4;
  wire [0:0] CLBLM_L_X10Y128_SLICE_X12Y128_B5;
  wire [0:0] CLBLM_L_X10Y128_SLICE_X12Y128_B6;
  wire [0:0] CLBLM_L_X10Y128_SLICE_X12Y128_BO5;
  wire [0:0] CLBLM_L_X10Y128_SLICE_X12Y128_BO6;
  wire [0:0] CLBLM_L_X10Y128_SLICE_X12Y128_B_CY;
  wire [0:0] CLBLM_L_X10Y128_SLICE_X12Y128_B_XOR;
  wire [0:0] CLBLM_L_X10Y128_SLICE_X12Y128_C;
  wire [0:0] CLBLM_L_X10Y128_SLICE_X12Y128_C1;
  wire [0:0] CLBLM_L_X10Y128_SLICE_X12Y128_C2;
  wire [0:0] CLBLM_L_X10Y128_SLICE_X12Y128_C3;
  wire [0:0] CLBLM_L_X10Y128_SLICE_X12Y128_C4;
  wire [0:0] CLBLM_L_X10Y128_SLICE_X12Y128_C5;
  wire [0:0] CLBLM_L_X10Y128_SLICE_X12Y128_C6;
  wire [0:0] CLBLM_L_X10Y128_SLICE_X12Y128_CO5;
  wire [0:0] CLBLM_L_X10Y128_SLICE_X12Y128_CO6;
  wire [0:0] CLBLM_L_X10Y128_SLICE_X12Y128_C_CY;
  wire [0:0] CLBLM_L_X10Y128_SLICE_X12Y128_C_XOR;
  wire [0:0] CLBLM_L_X10Y128_SLICE_X12Y128_D;
  wire [0:0] CLBLM_L_X10Y128_SLICE_X12Y128_D1;
  wire [0:0] CLBLM_L_X10Y128_SLICE_X12Y128_D2;
  wire [0:0] CLBLM_L_X10Y128_SLICE_X12Y128_D3;
  wire [0:0] CLBLM_L_X10Y128_SLICE_X12Y128_D4;
  wire [0:0] CLBLM_L_X10Y128_SLICE_X12Y128_D5;
  wire [0:0] CLBLM_L_X10Y128_SLICE_X12Y128_D6;
  wire [0:0] CLBLM_L_X10Y128_SLICE_X12Y128_DO5;
  wire [0:0] CLBLM_L_X10Y128_SLICE_X12Y128_DO6;
  wire [0:0] CLBLM_L_X10Y128_SLICE_X12Y128_D_CY;
  wire [0:0] CLBLM_L_X10Y128_SLICE_X12Y128_D_XOR;
  wire [0:0] CLBLM_L_X10Y128_SLICE_X13Y128_A;
  wire [0:0] CLBLM_L_X10Y128_SLICE_X13Y128_A1;
  wire [0:0] CLBLM_L_X10Y128_SLICE_X13Y128_A2;
  wire [0:0] CLBLM_L_X10Y128_SLICE_X13Y128_A3;
  wire [0:0] CLBLM_L_X10Y128_SLICE_X13Y128_A4;
  wire [0:0] CLBLM_L_X10Y128_SLICE_X13Y128_A5;
  wire [0:0] CLBLM_L_X10Y128_SLICE_X13Y128_A6;
  wire [0:0] CLBLM_L_X10Y128_SLICE_X13Y128_AMUX;
  wire [0:0] CLBLM_L_X10Y128_SLICE_X13Y128_AO5;
  wire [0:0] CLBLM_L_X10Y128_SLICE_X13Y128_AO6;
  wire [0:0] CLBLM_L_X10Y128_SLICE_X13Y128_A_CY;
  wire [0:0] CLBLM_L_X10Y128_SLICE_X13Y128_A_XOR;
  wire [0:0] CLBLM_L_X10Y128_SLICE_X13Y128_B;
  wire [0:0] CLBLM_L_X10Y128_SLICE_X13Y128_B1;
  wire [0:0] CLBLM_L_X10Y128_SLICE_X13Y128_B2;
  wire [0:0] CLBLM_L_X10Y128_SLICE_X13Y128_B3;
  wire [0:0] CLBLM_L_X10Y128_SLICE_X13Y128_B4;
  wire [0:0] CLBLM_L_X10Y128_SLICE_X13Y128_B5;
  wire [0:0] CLBLM_L_X10Y128_SLICE_X13Y128_B6;
  wire [0:0] CLBLM_L_X10Y128_SLICE_X13Y128_BO5;
  wire [0:0] CLBLM_L_X10Y128_SLICE_X13Y128_BO6;
  wire [0:0] CLBLM_L_X10Y128_SLICE_X13Y128_B_CY;
  wire [0:0] CLBLM_L_X10Y128_SLICE_X13Y128_B_XOR;
  wire [0:0] CLBLM_L_X10Y128_SLICE_X13Y128_C;
  wire [0:0] CLBLM_L_X10Y128_SLICE_X13Y128_C1;
  wire [0:0] CLBLM_L_X10Y128_SLICE_X13Y128_C2;
  wire [0:0] CLBLM_L_X10Y128_SLICE_X13Y128_C3;
  wire [0:0] CLBLM_L_X10Y128_SLICE_X13Y128_C4;
  wire [0:0] CLBLM_L_X10Y128_SLICE_X13Y128_C5;
  wire [0:0] CLBLM_L_X10Y128_SLICE_X13Y128_C6;
  wire [0:0] CLBLM_L_X10Y128_SLICE_X13Y128_CO5;
  wire [0:0] CLBLM_L_X10Y128_SLICE_X13Y128_CO6;
  wire [0:0] CLBLM_L_X10Y128_SLICE_X13Y128_C_CY;
  wire [0:0] CLBLM_L_X10Y128_SLICE_X13Y128_C_XOR;
  wire [0:0] CLBLM_L_X10Y128_SLICE_X13Y128_D;
  wire [0:0] CLBLM_L_X10Y128_SLICE_X13Y128_D1;
  wire [0:0] CLBLM_L_X10Y128_SLICE_X13Y128_D2;
  wire [0:0] CLBLM_L_X10Y128_SLICE_X13Y128_D3;
  wire [0:0] CLBLM_L_X10Y128_SLICE_X13Y128_D4;
  wire [0:0] CLBLM_L_X10Y128_SLICE_X13Y128_D5;
  wire [0:0] CLBLM_L_X10Y128_SLICE_X13Y128_D6;
  wire [0:0] CLBLM_L_X10Y128_SLICE_X13Y128_DO5;
  wire [0:0] CLBLM_L_X10Y128_SLICE_X13Y128_DO6;
  wire [0:0] CLBLM_L_X10Y128_SLICE_X13Y128_D_CY;
  wire [0:0] CLBLM_L_X10Y128_SLICE_X13Y128_D_XOR;
  wire [0:0] CLBLM_L_X12Y115_SLICE_X16Y115_A;
  wire [0:0] CLBLM_L_X12Y115_SLICE_X16Y115_A1;
  wire [0:0] CLBLM_L_X12Y115_SLICE_X16Y115_A2;
  wire [0:0] CLBLM_L_X12Y115_SLICE_X16Y115_A3;
  wire [0:0] CLBLM_L_X12Y115_SLICE_X16Y115_A4;
  wire [0:0] CLBLM_L_X12Y115_SLICE_X16Y115_A5;
  wire [0:0] CLBLM_L_X12Y115_SLICE_X16Y115_A6;
  wire [0:0] CLBLM_L_X12Y115_SLICE_X16Y115_AO5;
  wire [0:0] CLBLM_L_X12Y115_SLICE_X16Y115_AO6;
  wire [0:0] CLBLM_L_X12Y115_SLICE_X16Y115_AQ;
  wire [0:0] CLBLM_L_X12Y115_SLICE_X16Y115_A_CY;
  wire [0:0] CLBLM_L_X12Y115_SLICE_X16Y115_A_XOR;
  wire [0:0] CLBLM_L_X12Y115_SLICE_X16Y115_B;
  wire [0:0] CLBLM_L_X12Y115_SLICE_X16Y115_B1;
  wire [0:0] CLBLM_L_X12Y115_SLICE_X16Y115_B2;
  wire [0:0] CLBLM_L_X12Y115_SLICE_X16Y115_B3;
  wire [0:0] CLBLM_L_X12Y115_SLICE_X16Y115_B4;
  wire [0:0] CLBLM_L_X12Y115_SLICE_X16Y115_B5;
  wire [0:0] CLBLM_L_X12Y115_SLICE_X16Y115_B6;
  wire [0:0] CLBLM_L_X12Y115_SLICE_X16Y115_BO5;
  wire [0:0] CLBLM_L_X12Y115_SLICE_X16Y115_BO6;
  wire [0:0] CLBLM_L_X12Y115_SLICE_X16Y115_BQ;
  wire [0:0] CLBLM_L_X12Y115_SLICE_X16Y115_B_CY;
  wire [0:0] CLBLM_L_X12Y115_SLICE_X16Y115_B_XOR;
  wire [0:0] CLBLM_L_X12Y115_SLICE_X16Y115_C;
  wire [0:0] CLBLM_L_X12Y115_SLICE_X16Y115_C1;
  wire [0:0] CLBLM_L_X12Y115_SLICE_X16Y115_C2;
  wire [0:0] CLBLM_L_X12Y115_SLICE_X16Y115_C3;
  wire [0:0] CLBLM_L_X12Y115_SLICE_X16Y115_C4;
  wire [0:0] CLBLM_L_X12Y115_SLICE_X16Y115_C5;
  wire [0:0] CLBLM_L_X12Y115_SLICE_X16Y115_C6;
  wire [0:0] CLBLM_L_X12Y115_SLICE_X16Y115_CLK;
  wire [0:0] CLBLM_L_X12Y115_SLICE_X16Y115_CO5;
  wire [0:0] CLBLM_L_X12Y115_SLICE_X16Y115_CO6;
  wire [0:0] CLBLM_L_X12Y115_SLICE_X16Y115_CQ;
  wire [0:0] CLBLM_L_X12Y115_SLICE_X16Y115_C_CY;
  wire [0:0] CLBLM_L_X12Y115_SLICE_X16Y115_C_XOR;
  wire [0:0] CLBLM_L_X12Y115_SLICE_X16Y115_D;
  wire [0:0] CLBLM_L_X12Y115_SLICE_X16Y115_D1;
  wire [0:0] CLBLM_L_X12Y115_SLICE_X16Y115_D2;
  wire [0:0] CLBLM_L_X12Y115_SLICE_X16Y115_D3;
  wire [0:0] CLBLM_L_X12Y115_SLICE_X16Y115_D4;
  wire [0:0] CLBLM_L_X12Y115_SLICE_X16Y115_D5;
  wire [0:0] CLBLM_L_X12Y115_SLICE_X16Y115_D6;
  wire [0:0] CLBLM_L_X12Y115_SLICE_X16Y115_DO5;
  wire [0:0] CLBLM_L_X12Y115_SLICE_X16Y115_DO6;
  wire [0:0] CLBLM_L_X12Y115_SLICE_X16Y115_DQ;
  wire [0:0] CLBLM_L_X12Y115_SLICE_X16Y115_D_CY;
  wire [0:0] CLBLM_L_X12Y115_SLICE_X16Y115_D_XOR;
  wire [0:0] CLBLM_L_X12Y115_SLICE_X17Y115_A;
  wire [0:0] CLBLM_L_X12Y115_SLICE_X17Y115_A1;
  wire [0:0] CLBLM_L_X12Y115_SLICE_X17Y115_A2;
  wire [0:0] CLBLM_L_X12Y115_SLICE_X17Y115_A3;
  wire [0:0] CLBLM_L_X12Y115_SLICE_X17Y115_A4;
  wire [0:0] CLBLM_L_X12Y115_SLICE_X17Y115_A5;
  wire [0:0] CLBLM_L_X12Y115_SLICE_X17Y115_A6;
  wire [0:0] CLBLM_L_X12Y115_SLICE_X17Y115_AO5;
  wire [0:0] CLBLM_L_X12Y115_SLICE_X17Y115_AO6;
  wire [0:0] CLBLM_L_X12Y115_SLICE_X17Y115_A_CY;
  wire [0:0] CLBLM_L_X12Y115_SLICE_X17Y115_A_XOR;
  wire [0:0] CLBLM_L_X12Y115_SLICE_X17Y115_B;
  wire [0:0] CLBLM_L_X12Y115_SLICE_X17Y115_B1;
  wire [0:0] CLBLM_L_X12Y115_SLICE_X17Y115_B2;
  wire [0:0] CLBLM_L_X12Y115_SLICE_X17Y115_B3;
  wire [0:0] CLBLM_L_X12Y115_SLICE_X17Y115_B4;
  wire [0:0] CLBLM_L_X12Y115_SLICE_X17Y115_B5;
  wire [0:0] CLBLM_L_X12Y115_SLICE_X17Y115_B6;
  wire [0:0] CLBLM_L_X12Y115_SLICE_X17Y115_BO5;
  wire [0:0] CLBLM_L_X12Y115_SLICE_X17Y115_BO6;
  wire [0:0] CLBLM_L_X12Y115_SLICE_X17Y115_B_CY;
  wire [0:0] CLBLM_L_X12Y115_SLICE_X17Y115_B_XOR;
  wire [0:0] CLBLM_L_X12Y115_SLICE_X17Y115_C;
  wire [0:0] CLBLM_L_X12Y115_SLICE_X17Y115_C1;
  wire [0:0] CLBLM_L_X12Y115_SLICE_X17Y115_C2;
  wire [0:0] CLBLM_L_X12Y115_SLICE_X17Y115_C3;
  wire [0:0] CLBLM_L_X12Y115_SLICE_X17Y115_C4;
  wire [0:0] CLBLM_L_X12Y115_SLICE_X17Y115_C5;
  wire [0:0] CLBLM_L_X12Y115_SLICE_X17Y115_C6;
  wire [0:0] CLBLM_L_X12Y115_SLICE_X17Y115_CO5;
  wire [0:0] CLBLM_L_X12Y115_SLICE_X17Y115_CO6;
  wire [0:0] CLBLM_L_X12Y115_SLICE_X17Y115_C_CY;
  wire [0:0] CLBLM_L_X12Y115_SLICE_X17Y115_C_XOR;
  wire [0:0] CLBLM_L_X12Y115_SLICE_X17Y115_D;
  wire [0:0] CLBLM_L_X12Y115_SLICE_X17Y115_D1;
  wire [0:0] CLBLM_L_X12Y115_SLICE_X17Y115_D2;
  wire [0:0] CLBLM_L_X12Y115_SLICE_X17Y115_D3;
  wire [0:0] CLBLM_L_X12Y115_SLICE_X17Y115_D4;
  wire [0:0] CLBLM_L_X12Y115_SLICE_X17Y115_D5;
  wire [0:0] CLBLM_L_X12Y115_SLICE_X17Y115_D6;
  wire [0:0] CLBLM_L_X12Y115_SLICE_X17Y115_DO5;
  wire [0:0] CLBLM_L_X12Y115_SLICE_X17Y115_DO6;
  wire [0:0] CLBLM_L_X12Y115_SLICE_X17Y115_D_CY;
  wire [0:0] CLBLM_L_X12Y115_SLICE_X17Y115_D_XOR;
  wire [0:0] CLBLM_L_X12Y118_SLICE_X16Y118_A;
  wire [0:0] CLBLM_L_X12Y118_SLICE_X16Y118_A1;
  wire [0:0] CLBLM_L_X12Y118_SLICE_X16Y118_A2;
  wire [0:0] CLBLM_L_X12Y118_SLICE_X16Y118_A3;
  wire [0:0] CLBLM_L_X12Y118_SLICE_X16Y118_A4;
  wire [0:0] CLBLM_L_X12Y118_SLICE_X16Y118_A5;
  wire [0:0] CLBLM_L_X12Y118_SLICE_X16Y118_A6;
  wire [0:0] CLBLM_L_X12Y118_SLICE_X16Y118_AO5;
  wire [0:0] CLBLM_L_X12Y118_SLICE_X16Y118_AO6;
  wire [0:0] CLBLM_L_X12Y118_SLICE_X16Y118_AQ;
  wire [0:0] CLBLM_L_X12Y118_SLICE_X16Y118_A_CY;
  wire [0:0] CLBLM_L_X12Y118_SLICE_X16Y118_A_XOR;
  wire [0:0] CLBLM_L_X12Y118_SLICE_X16Y118_B;
  wire [0:0] CLBLM_L_X12Y118_SLICE_X16Y118_B1;
  wire [0:0] CLBLM_L_X12Y118_SLICE_X16Y118_B2;
  wire [0:0] CLBLM_L_X12Y118_SLICE_X16Y118_B3;
  wire [0:0] CLBLM_L_X12Y118_SLICE_X16Y118_B4;
  wire [0:0] CLBLM_L_X12Y118_SLICE_X16Y118_B5;
  wire [0:0] CLBLM_L_X12Y118_SLICE_X16Y118_B6;
  wire [0:0] CLBLM_L_X12Y118_SLICE_X16Y118_BO5;
  wire [0:0] CLBLM_L_X12Y118_SLICE_X16Y118_BO6;
  wire [0:0] CLBLM_L_X12Y118_SLICE_X16Y118_BQ;
  wire [0:0] CLBLM_L_X12Y118_SLICE_X16Y118_B_CY;
  wire [0:0] CLBLM_L_X12Y118_SLICE_X16Y118_B_XOR;
  wire [0:0] CLBLM_L_X12Y118_SLICE_X16Y118_C;
  wire [0:0] CLBLM_L_X12Y118_SLICE_X16Y118_C1;
  wire [0:0] CLBLM_L_X12Y118_SLICE_X16Y118_C2;
  wire [0:0] CLBLM_L_X12Y118_SLICE_X16Y118_C3;
  wire [0:0] CLBLM_L_X12Y118_SLICE_X16Y118_C4;
  wire [0:0] CLBLM_L_X12Y118_SLICE_X16Y118_C5;
  wire [0:0] CLBLM_L_X12Y118_SLICE_X16Y118_C6;
  wire [0:0] CLBLM_L_X12Y118_SLICE_X16Y118_CLK;
  wire [0:0] CLBLM_L_X12Y118_SLICE_X16Y118_CO5;
  wire [0:0] CLBLM_L_X12Y118_SLICE_X16Y118_CO6;
  wire [0:0] CLBLM_L_X12Y118_SLICE_X16Y118_C_CY;
  wire [0:0] CLBLM_L_X12Y118_SLICE_X16Y118_C_XOR;
  wire [0:0] CLBLM_L_X12Y118_SLICE_X16Y118_D;
  wire [0:0] CLBLM_L_X12Y118_SLICE_X16Y118_D1;
  wire [0:0] CLBLM_L_X12Y118_SLICE_X16Y118_D2;
  wire [0:0] CLBLM_L_X12Y118_SLICE_X16Y118_D3;
  wire [0:0] CLBLM_L_X12Y118_SLICE_X16Y118_D4;
  wire [0:0] CLBLM_L_X12Y118_SLICE_X16Y118_D5;
  wire [0:0] CLBLM_L_X12Y118_SLICE_X16Y118_D6;
  wire [0:0] CLBLM_L_X12Y118_SLICE_X16Y118_DO5;
  wire [0:0] CLBLM_L_X12Y118_SLICE_X16Y118_DO6;
  wire [0:0] CLBLM_L_X12Y118_SLICE_X16Y118_D_CY;
  wire [0:0] CLBLM_L_X12Y118_SLICE_X16Y118_D_XOR;
  wire [0:0] CLBLM_L_X12Y118_SLICE_X17Y118_A;
  wire [0:0] CLBLM_L_X12Y118_SLICE_X17Y118_A1;
  wire [0:0] CLBLM_L_X12Y118_SLICE_X17Y118_A2;
  wire [0:0] CLBLM_L_X12Y118_SLICE_X17Y118_A3;
  wire [0:0] CLBLM_L_X12Y118_SLICE_X17Y118_A4;
  wire [0:0] CLBLM_L_X12Y118_SLICE_X17Y118_A5;
  wire [0:0] CLBLM_L_X12Y118_SLICE_X17Y118_A6;
  wire [0:0] CLBLM_L_X12Y118_SLICE_X17Y118_AO5;
  wire [0:0] CLBLM_L_X12Y118_SLICE_X17Y118_AO6;
  wire [0:0] CLBLM_L_X12Y118_SLICE_X17Y118_A_CY;
  wire [0:0] CLBLM_L_X12Y118_SLICE_X17Y118_A_XOR;
  wire [0:0] CLBLM_L_X12Y118_SLICE_X17Y118_B;
  wire [0:0] CLBLM_L_X12Y118_SLICE_X17Y118_B1;
  wire [0:0] CLBLM_L_X12Y118_SLICE_X17Y118_B2;
  wire [0:0] CLBLM_L_X12Y118_SLICE_X17Y118_B3;
  wire [0:0] CLBLM_L_X12Y118_SLICE_X17Y118_B4;
  wire [0:0] CLBLM_L_X12Y118_SLICE_X17Y118_B5;
  wire [0:0] CLBLM_L_X12Y118_SLICE_X17Y118_B6;
  wire [0:0] CLBLM_L_X12Y118_SLICE_X17Y118_BO5;
  wire [0:0] CLBLM_L_X12Y118_SLICE_X17Y118_BO6;
  wire [0:0] CLBLM_L_X12Y118_SLICE_X17Y118_B_CY;
  wire [0:0] CLBLM_L_X12Y118_SLICE_X17Y118_B_XOR;
  wire [0:0] CLBLM_L_X12Y118_SLICE_X17Y118_C;
  wire [0:0] CLBLM_L_X12Y118_SLICE_X17Y118_C1;
  wire [0:0] CLBLM_L_X12Y118_SLICE_X17Y118_C2;
  wire [0:0] CLBLM_L_X12Y118_SLICE_X17Y118_C3;
  wire [0:0] CLBLM_L_X12Y118_SLICE_X17Y118_C4;
  wire [0:0] CLBLM_L_X12Y118_SLICE_X17Y118_C5;
  wire [0:0] CLBLM_L_X12Y118_SLICE_X17Y118_C6;
  wire [0:0] CLBLM_L_X12Y118_SLICE_X17Y118_CO5;
  wire [0:0] CLBLM_L_X12Y118_SLICE_X17Y118_CO6;
  wire [0:0] CLBLM_L_X12Y118_SLICE_X17Y118_C_CY;
  wire [0:0] CLBLM_L_X12Y118_SLICE_X17Y118_C_XOR;
  wire [0:0] CLBLM_L_X12Y118_SLICE_X17Y118_D;
  wire [0:0] CLBLM_L_X12Y118_SLICE_X17Y118_D1;
  wire [0:0] CLBLM_L_X12Y118_SLICE_X17Y118_D2;
  wire [0:0] CLBLM_L_X12Y118_SLICE_X17Y118_D3;
  wire [0:0] CLBLM_L_X12Y118_SLICE_X17Y118_D4;
  wire [0:0] CLBLM_L_X12Y118_SLICE_X17Y118_D5;
  wire [0:0] CLBLM_L_X12Y118_SLICE_X17Y118_D6;
  wire [0:0] CLBLM_L_X12Y118_SLICE_X17Y118_DO5;
  wire [0:0] CLBLM_L_X12Y118_SLICE_X17Y118_DO6;
  wire [0:0] CLBLM_L_X12Y118_SLICE_X17Y118_D_CY;
  wire [0:0] CLBLM_L_X12Y118_SLICE_X17Y118_D_XOR;
  wire [0:0] CLBLM_L_X12Y119_SLICE_X16Y119_A;
  wire [0:0] CLBLM_L_X12Y119_SLICE_X16Y119_A1;
  wire [0:0] CLBLM_L_X12Y119_SLICE_X16Y119_A2;
  wire [0:0] CLBLM_L_X12Y119_SLICE_X16Y119_A3;
  wire [0:0] CLBLM_L_X12Y119_SLICE_X16Y119_A4;
  wire [0:0] CLBLM_L_X12Y119_SLICE_X16Y119_A5;
  wire [0:0] CLBLM_L_X12Y119_SLICE_X16Y119_A6;
  wire [0:0] CLBLM_L_X12Y119_SLICE_X16Y119_AO5;
  wire [0:0] CLBLM_L_X12Y119_SLICE_X16Y119_AO6;
  wire [0:0] CLBLM_L_X12Y119_SLICE_X16Y119_A_CY;
  wire [0:0] CLBLM_L_X12Y119_SLICE_X16Y119_A_XOR;
  wire [0:0] CLBLM_L_X12Y119_SLICE_X16Y119_B;
  wire [0:0] CLBLM_L_X12Y119_SLICE_X16Y119_B1;
  wire [0:0] CLBLM_L_X12Y119_SLICE_X16Y119_B2;
  wire [0:0] CLBLM_L_X12Y119_SLICE_X16Y119_B3;
  wire [0:0] CLBLM_L_X12Y119_SLICE_X16Y119_B4;
  wire [0:0] CLBLM_L_X12Y119_SLICE_X16Y119_B5;
  wire [0:0] CLBLM_L_X12Y119_SLICE_X16Y119_B6;
  wire [0:0] CLBLM_L_X12Y119_SLICE_X16Y119_BO5;
  wire [0:0] CLBLM_L_X12Y119_SLICE_X16Y119_BO6;
  wire [0:0] CLBLM_L_X12Y119_SLICE_X16Y119_B_CY;
  wire [0:0] CLBLM_L_X12Y119_SLICE_X16Y119_B_XOR;
  wire [0:0] CLBLM_L_X12Y119_SLICE_X16Y119_C;
  wire [0:0] CLBLM_L_X12Y119_SLICE_X16Y119_C1;
  wire [0:0] CLBLM_L_X12Y119_SLICE_X16Y119_C2;
  wire [0:0] CLBLM_L_X12Y119_SLICE_X16Y119_C3;
  wire [0:0] CLBLM_L_X12Y119_SLICE_X16Y119_C4;
  wire [0:0] CLBLM_L_X12Y119_SLICE_X16Y119_C5;
  wire [0:0] CLBLM_L_X12Y119_SLICE_X16Y119_C6;
  wire [0:0] CLBLM_L_X12Y119_SLICE_X16Y119_CO5;
  wire [0:0] CLBLM_L_X12Y119_SLICE_X16Y119_CO6;
  wire [0:0] CLBLM_L_X12Y119_SLICE_X16Y119_C_CY;
  wire [0:0] CLBLM_L_X12Y119_SLICE_X16Y119_C_XOR;
  wire [0:0] CLBLM_L_X12Y119_SLICE_X16Y119_D;
  wire [0:0] CLBLM_L_X12Y119_SLICE_X16Y119_D1;
  wire [0:0] CLBLM_L_X12Y119_SLICE_X16Y119_D2;
  wire [0:0] CLBLM_L_X12Y119_SLICE_X16Y119_D3;
  wire [0:0] CLBLM_L_X12Y119_SLICE_X16Y119_D4;
  wire [0:0] CLBLM_L_X12Y119_SLICE_X16Y119_D5;
  wire [0:0] CLBLM_L_X12Y119_SLICE_X16Y119_D6;
  wire [0:0] CLBLM_L_X12Y119_SLICE_X16Y119_DO5;
  wire [0:0] CLBLM_L_X12Y119_SLICE_X16Y119_DO6;
  wire [0:0] CLBLM_L_X12Y119_SLICE_X16Y119_D_CY;
  wire [0:0] CLBLM_L_X12Y119_SLICE_X16Y119_D_XOR;
  wire [0:0] CLBLM_L_X12Y119_SLICE_X17Y119_A;
  wire [0:0] CLBLM_L_X12Y119_SLICE_X17Y119_A1;
  wire [0:0] CLBLM_L_X12Y119_SLICE_X17Y119_A2;
  wire [0:0] CLBLM_L_X12Y119_SLICE_X17Y119_A3;
  wire [0:0] CLBLM_L_X12Y119_SLICE_X17Y119_A4;
  wire [0:0] CLBLM_L_X12Y119_SLICE_X17Y119_A5;
  wire [0:0] CLBLM_L_X12Y119_SLICE_X17Y119_A6;
  wire [0:0] CLBLM_L_X12Y119_SLICE_X17Y119_AMUX;
  wire [0:0] CLBLM_L_X12Y119_SLICE_X17Y119_AO5;
  wire [0:0] CLBLM_L_X12Y119_SLICE_X17Y119_AO6;
  wire [0:0] CLBLM_L_X12Y119_SLICE_X17Y119_A_CY;
  wire [0:0] CLBLM_L_X12Y119_SLICE_X17Y119_A_XOR;
  wire [0:0] CLBLM_L_X12Y119_SLICE_X17Y119_B;
  wire [0:0] CLBLM_L_X12Y119_SLICE_X17Y119_B1;
  wire [0:0] CLBLM_L_X12Y119_SLICE_X17Y119_B2;
  wire [0:0] CLBLM_L_X12Y119_SLICE_X17Y119_B3;
  wire [0:0] CLBLM_L_X12Y119_SLICE_X17Y119_B4;
  wire [0:0] CLBLM_L_X12Y119_SLICE_X17Y119_B5;
  wire [0:0] CLBLM_L_X12Y119_SLICE_X17Y119_B6;
  wire [0:0] CLBLM_L_X12Y119_SLICE_X17Y119_BO5;
  wire [0:0] CLBLM_L_X12Y119_SLICE_X17Y119_BO6;
  wire [0:0] CLBLM_L_X12Y119_SLICE_X17Y119_B_CY;
  wire [0:0] CLBLM_L_X12Y119_SLICE_X17Y119_B_XOR;
  wire [0:0] CLBLM_L_X12Y119_SLICE_X17Y119_C;
  wire [0:0] CLBLM_L_X12Y119_SLICE_X17Y119_C1;
  wire [0:0] CLBLM_L_X12Y119_SLICE_X17Y119_C2;
  wire [0:0] CLBLM_L_X12Y119_SLICE_X17Y119_C3;
  wire [0:0] CLBLM_L_X12Y119_SLICE_X17Y119_C4;
  wire [0:0] CLBLM_L_X12Y119_SLICE_X17Y119_C5;
  wire [0:0] CLBLM_L_X12Y119_SLICE_X17Y119_C6;
  wire [0:0] CLBLM_L_X12Y119_SLICE_X17Y119_CO5;
  wire [0:0] CLBLM_L_X12Y119_SLICE_X17Y119_CO6;
  wire [0:0] CLBLM_L_X12Y119_SLICE_X17Y119_C_CY;
  wire [0:0] CLBLM_L_X12Y119_SLICE_X17Y119_C_XOR;
  wire [0:0] CLBLM_L_X12Y119_SLICE_X17Y119_D;
  wire [0:0] CLBLM_L_X12Y119_SLICE_X17Y119_D1;
  wire [0:0] CLBLM_L_X12Y119_SLICE_X17Y119_D2;
  wire [0:0] CLBLM_L_X12Y119_SLICE_X17Y119_D3;
  wire [0:0] CLBLM_L_X12Y119_SLICE_X17Y119_D4;
  wire [0:0] CLBLM_L_X12Y119_SLICE_X17Y119_D5;
  wire [0:0] CLBLM_L_X12Y119_SLICE_X17Y119_D6;
  wire [0:0] CLBLM_L_X12Y119_SLICE_X17Y119_DO5;
  wire [0:0] CLBLM_L_X12Y119_SLICE_X17Y119_DO6;
  wire [0:0] CLBLM_L_X12Y119_SLICE_X17Y119_D_CY;
  wire [0:0] CLBLM_L_X12Y119_SLICE_X17Y119_D_XOR;
  wire [0:0] CLBLM_L_X12Y120_SLICE_X16Y120_A;
  wire [0:0] CLBLM_L_X12Y120_SLICE_X16Y120_A1;
  wire [0:0] CLBLM_L_X12Y120_SLICE_X16Y120_A2;
  wire [0:0] CLBLM_L_X12Y120_SLICE_X16Y120_A3;
  wire [0:0] CLBLM_L_X12Y120_SLICE_X16Y120_A4;
  wire [0:0] CLBLM_L_X12Y120_SLICE_X16Y120_A5;
  wire [0:0] CLBLM_L_X12Y120_SLICE_X16Y120_A6;
  wire [0:0] CLBLM_L_X12Y120_SLICE_X16Y120_AMUX;
  wire [0:0] CLBLM_L_X12Y120_SLICE_X16Y120_AO5;
  wire [0:0] CLBLM_L_X12Y120_SLICE_X16Y120_AO6;
  wire [0:0] CLBLM_L_X12Y120_SLICE_X16Y120_A_CY;
  wire [0:0] CLBLM_L_X12Y120_SLICE_X16Y120_A_XOR;
  wire [0:0] CLBLM_L_X12Y120_SLICE_X16Y120_B;
  wire [0:0] CLBLM_L_X12Y120_SLICE_X16Y120_B1;
  wire [0:0] CLBLM_L_X12Y120_SLICE_X16Y120_B2;
  wire [0:0] CLBLM_L_X12Y120_SLICE_X16Y120_B3;
  wire [0:0] CLBLM_L_X12Y120_SLICE_X16Y120_B4;
  wire [0:0] CLBLM_L_X12Y120_SLICE_X16Y120_B5;
  wire [0:0] CLBLM_L_X12Y120_SLICE_X16Y120_B6;
  wire [0:0] CLBLM_L_X12Y120_SLICE_X16Y120_BO5;
  wire [0:0] CLBLM_L_X12Y120_SLICE_X16Y120_BO6;
  wire [0:0] CLBLM_L_X12Y120_SLICE_X16Y120_B_CY;
  wire [0:0] CLBLM_L_X12Y120_SLICE_X16Y120_B_XOR;
  wire [0:0] CLBLM_L_X12Y120_SLICE_X16Y120_C;
  wire [0:0] CLBLM_L_X12Y120_SLICE_X16Y120_C1;
  wire [0:0] CLBLM_L_X12Y120_SLICE_X16Y120_C2;
  wire [0:0] CLBLM_L_X12Y120_SLICE_X16Y120_C3;
  wire [0:0] CLBLM_L_X12Y120_SLICE_X16Y120_C4;
  wire [0:0] CLBLM_L_X12Y120_SLICE_X16Y120_C5;
  wire [0:0] CLBLM_L_X12Y120_SLICE_X16Y120_C6;
  wire [0:0] CLBLM_L_X12Y120_SLICE_X16Y120_CO5;
  wire [0:0] CLBLM_L_X12Y120_SLICE_X16Y120_CO6;
  wire [0:0] CLBLM_L_X12Y120_SLICE_X16Y120_C_CY;
  wire [0:0] CLBLM_L_X12Y120_SLICE_X16Y120_C_XOR;
  wire [0:0] CLBLM_L_X12Y120_SLICE_X16Y120_D;
  wire [0:0] CLBLM_L_X12Y120_SLICE_X16Y120_D1;
  wire [0:0] CLBLM_L_X12Y120_SLICE_X16Y120_D2;
  wire [0:0] CLBLM_L_X12Y120_SLICE_X16Y120_D3;
  wire [0:0] CLBLM_L_X12Y120_SLICE_X16Y120_D4;
  wire [0:0] CLBLM_L_X12Y120_SLICE_X16Y120_D5;
  wire [0:0] CLBLM_L_X12Y120_SLICE_X16Y120_D6;
  wire [0:0] CLBLM_L_X12Y120_SLICE_X16Y120_DO5;
  wire [0:0] CLBLM_L_X12Y120_SLICE_X16Y120_DO6;
  wire [0:0] CLBLM_L_X12Y120_SLICE_X16Y120_D_CY;
  wire [0:0] CLBLM_L_X12Y120_SLICE_X16Y120_D_XOR;
  wire [0:0] CLBLM_L_X12Y120_SLICE_X17Y120_A;
  wire [0:0] CLBLM_L_X12Y120_SLICE_X17Y120_A1;
  wire [0:0] CLBLM_L_X12Y120_SLICE_X17Y120_A2;
  wire [0:0] CLBLM_L_X12Y120_SLICE_X17Y120_A3;
  wire [0:0] CLBLM_L_X12Y120_SLICE_X17Y120_A4;
  wire [0:0] CLBLM_L_X12Y120_SLICE_X17Y120_A5;
  wire [0:0] CLBLM_L_X12Y120_SLICE_X17Y120_A6;
  wire [0:0] CLBLM_L_X12Y120_SLICE_X17Y120_AO5;
  wire [0:0] CLBLM_L_X12Y120_SLICE_X17Y120_AO6;
  wire [0:0] CLBLM_L_X12Y120_SLICE_X17Y120_AQ;
  wire [0:0] CLBLM_L_X12Y120_SLICE_X17Y120_A_CY;
  wire [0:0] CLBLM_L_X12Y120_SLICE_X17Y120_A_XOR;
  wire [0:0] CLBLM_L_X12Y120_SLICE_X17Y120_B;
  wire [0:0] CLBLM_L_X12Y120_SLICE_X17Y120_B1;
  wire [0:0] CLBLM_L_X12Y120_SLICE_X17Y120_B2;
  wire [0:0] CLBLM_L_X12Y120_SLICE_X17Y120_B3;
  wire [0:0] CLBLM_L_X12Y120_SLICE_X17Y120_B4;
  wire [0:0] CLBLM_L_X12Y120_SLICE_X17Y120_B5;
  wire [0:0] CLBLM_L_X12Y120_SLICE_X17Y120_B6;
  wire [0:0] CLBLM_L_X12Y120_SLICE_X17Y120_BO5;
  wire [0:0] CLBLM_L_X12Y120_SLICE_X17Y120_BO6;
  wire [0:0] CLBLM_L_X12Y120_SLICE_X17Y120_BQ;
  wire [0:0] CLBLM_L_X12Y120_SLICE_X17Y120_B_CY;
  wire [0:0] CLBLM_L_X12Y120_SLICE_X17Y120_B_XOR;
  wire [0:0] CLBLM_L_X12Y120_SLICE_X17Y120_C;
  wire [0:0] CLBLM_L_X12Y120_SLICE_X17Y120_C1;
  wire [0:0] CLBLM_L_X12Y120_SLICE_X17Y120_C2;
  wire [0:0] CLBLM_L_X12Y120_SLICE_X17Y120_C3;
  wire [0:0] CLBLM_L_X12Y120_SLICE_X17Y120_C4;
  wire [0:0] CLBLM_L_X12Y120_SLICE_X17Y120_C5;
  wire [0:0] CLBLM_L_X12Y120_SLICE_X17Y120_C6;
  wire [0:0] CLBLM_L_X12Y120_SLICE_X17Y120_CLK;
  wire [0:0] CLBLM_L_X12Y120_SLICE_X17Y120_CMUX;
  wire [0:0] CLBLM_L_X12Y120_SLICE_X17Y120_CO5;
  wire [0:0] CLBLM_L_X12Y120_SLICE_X17Y120_CO6;
  wire [0:0] CLBLM_L_X12Y120_SLICE_X17Y120_C_CY;
  wire [0:0] CLBLM_L_X12Y120_SLICE_X17Y120_C_XOR;
  wire [0:0] CLBLM_L_X12Y120_SLICE_X17Y120_D;
  wire [0:0] CLBLM_L_X12Y120_SLICE_X17Y120_D1;
  wire [0:0] CLBLM_L_X12Y120_SLICE_X17Y120_D2;
  wire [0:0] CLBLM_L_X12Y120_SLICE_X17Y120_D3;
  wire [0:0] CLBLM_L_X12Y120_SLICE_X17Y120_D4;
  wire [0:0] CLBLM_L_X12Y120_SLICE_X17Y120_D5;
  wire [0:0] CLBLM_L_X12Y120_SLICE_X17Y120_D6;
  wire [0:0] CLBLM_L_X12Y120_SLICE_X17Y120_DMUX;
  wire [0:0] CLBLM_L_X12Y120_SLICE_X17Y120_DO5;
  wire [0:0] CLBLM_L_X12Y120_SLICE_X17Y120_DO6;
  wire [0:0] CLBLM_L_X12Y120_SLICE_X17Y120_D_CY;
  wire [0:0] CLBLM_L_X12Y120_SLICE_X17Y120_D_XOR;
  wire [0:0] CLBLM_L_X12Y121_SLICE_X16Y121_A;
  wire [0:0] CLBLM_L_X12Y121_SLICE_X16Y121_A1;
  wire [0:0] CLBLM_L_X12Y121_SLICE_X16Y121_A2;
  wire [0:0] CLBLM_L_X12Y121_SLICE_X16Y121_A3;
  wire [0:0] CLBLM_L_X12Y121_SLICE_X16Y121_A4;
  wire [0:0] CLBLM_L_X12Y121_SLICE_X16Y121_A5;
  wire [0:0] CLBLM_L_X12Y121_SLICE_X16Y121_A6;
  wire [0:0] CLBLM_L_X12Y121_SLICE_X16Y121_AO5;
  wire [0:0] CLBLM_L_X12Y121_SLICE_X16Y121_AO6;
  wire [0:0] CLBLM_L_X12Y121_SLICE_X16Y121_AQ;
  wire [0:0] CLBLM_L_X12Y121_SLICE_X16Y121_A_CY;
  wire [0:0] CLBLM_L_X12Y121_SLICE_X16Y121_A_XOR;
  wire [0:0] CLBLM_L_X12Y121_SLICE_X16Y121_B;
  wire [0:0] CLBLM_L_X12Y121_SLICE_X16Y121_B1;
  wire [0:0] CLBLM_L_X12Y121_SLICE_X16Y121_B2;
  wire [0:0] CLBLM_L_X12Y121_SLICE_X16Y121_B3;
  wire [0:0] CLBLM_L_X12Y121_SLICE_X16Y121_B4;
  wire [0:0] CLBLM_L_X12Y121_SLICE_X16Y121_B5;
  wire [0:0] CLBLM_L_X12Y121_SLICE_X16Y121_B6;
  wire [0:0] CLBLM_L_X12Y121_SLICE_X16Y121_BO5;
  wire [0:0] CLBLM_L_X12Y121_SLICE_X16Y121_BO6;
  wire [0:0] CLBLM_L_X12Y121_SLICE_X16Y121_B_CY;
  wire [0:0] CLBLM_L_X12Y121_SLICE_X16Y121_B_XOR;
  wire [0:0] CLBLM_L_X12Y121_SLICE_X16Y121_C;
  wire [0:0] CLBLM_L_X12Y121_SLICE_X16Y121_C1;
  wire [0:0] CLBLM_L_X12Y121_SLICE_X16Y121_C2;
  wire [0:0] CLBLM_L_X12Y121_SLICE_X16Y121_C3;
  wire [0:0] CLBLM_L_X12Y121_SLICE_X16Y121_C4;
  wire [0:0] CLBLM_L_X12Y121_SLICE_X16Y121_C5;
  wire [0:0] CLBLM_L_X12Y121_SLICE_X16Y121_C6;
  wire [0:0] CLBLM_L_X12Y121_SLICE_X16Y121_CLK;
  wire [0:0] CLBLM_L_X12Y121_SLICE_X16Y121_CO5;
  wire [0:0] CLBLM_L_X12Y121_SLICE_X16Y121_CO6;
  wire [0:0] CLBLM_L_X12Y121_SLICE_X16Y121_C_CY;
  wire [0:0] CLBLM_L_X12Y121_SLICE_X16Y121_C_XOR;
  wire [0:0] CLBLM_L_X12Y121_SLICE_X16Y121_D;
  wire [0:0] CLBLM_L_X12Y121_SLICE_X16Y121_D1;
  wire [0:0] CLBLM_L_X12Y121_SLICE_X16Y121_D2;
  wire [0:0] CLBLM_L_X12Y121_SLICE_X16Y121_D3;
  wire [0:0] CLBLM_L_X12Y121_SLICE_X16Y121_D4;
  wire [0:0] CLBLM_L_X12Y121_SLICE_X16Y121_D5;
  wire [0:0] CLBLM_L_X12Y121_SLICE_X16Y121_D6;
  wire [0:0] CLBLM_L_X12Y121_SLICE_X16Y121_DO5;
  wire [0:0] CLBLM_L_X12Y121_SLICE_X16Y121_DO6;
  wire [0:0] CLBLM_L_X12Y121_SLICE_X16Y121_D_CY;
  wire [0:0] CLBLM_L_X12Y121_SLICE_X16Y121_D_XOR;
  wire [0:0] CLBLM_L_X12Y121_SLICE_X17Y121_A;
  wire [0:0] CLBLM_L_X12Y121_SLICE_X17Y121_A1;
  wire [0:0] CLBLM_L_X12Y121_SLICE_X17Y121_A2;
  wire [0:0] CLBLM_L_X12Y121_SLICE_X17Y121_A3;
  wire [0:0] CLBLM_L_X12Y121_SLICE_X17Y121_A4;
  wire [0:0] CLBLM_L_X12Y121_SLICE_X17Y121_A5;
  wire [0:0] CLBLM_L_X12Y121_SLICE_X17Y121_A6;
  wire [0:0] CLBLM_L_X12Y121_SLICE_X17Y121_AO5;
  wire [0:0] CLBLM_L_X12Y121_SLICE_X17Y121_AO6;
  wire [0:0] CLBLM_L_X12Y121_SLICE_X17Y121_A_CY;
  wire [0:0] CLBLM_L_X12Y121_SLICE_X17Y121_A_XOR;
  wire [0:0] CLBLM_L_X12Y121_SLICE_X17Y121_B;
  wire [0:0] CLBLM_L_X12Y121_SLICE_X17Y121_B1;
  wire [0:0] CLBLM_L_X12Y121_SLICE_X17Y121_B2;
  wire [0:0] CLBLM_L_X12Y121_SLICE_X17Y121_B3;
  wire [0:0] CLBLM_L_X12Y121_SLICE_X17Y121_B4;
  wire [0:0] CLBLM_L_X12Y121_SLICE_X17Y121_B5;
  wire [0:0] CLBLM_L_X12Y121_SLICE_X17Y121_B6;
  wire [0:0] CLBLM_L_X12Y121_SLICE_X17Y121_BO5;
  wire [0:0] CLBLM_L_X12Y121_SLICE_X17Y121_BO6;
  wire [0:0] CLBLM_L_X12Y121_SLICE_X17Y121_B_CY;
  wire [0:0] CLBLM_L_X12Y121_SLICE_X17Y121_B_XOR;
  wire [0:0] CLBLM_L_X12Y121_SLICE_X17Y121_C;
  wire [0:0] CLBLM_L_X12Y121_SLICE_X17Y121_C1;
  wire [0:0] CLBLM_L_X12Y121_SLICE_X17Y121_C2;
  wire [0:0] CLBLM_L_X12Y121_SLICE_X17Y121_C3;
  wire [0:0] CLBLM_L_X12Y121_SLICE_X17Y121_C4;
  wire [0:0] CLBLM_L_X12Y121_SLICE_X17Y121_C5;
  wire [0:0] CLBLM_L_X12Y121_SLICE_X17Y121_C6;
  wire [0:0] CLBLM_L_X12Y121_SLICE_X17Y121_CO5;
  wire [0:0] CLBLM_L_X12Y121_SLICE_X17Y121_CO6;
  wire [0:0] CLBLM_L_X12Y121_SLICE_X17Y121_C_CY;
  wire [0:0] CLBLM_L_X12Y121_SLICE_X17Y121_C_XOR;
  wire [0:0] CLBLM_L_X12Y121_SLICE_X17Y121_D;
  wire [0:0] CLBLM_L_X12Y121_SLICE_X17Y121_D1;
  wire [0:0] CLBLM_L_X12Y121_SLICE_X17Y121_D2;
  wire [0:0] CLBLM_L_X12Y121_SLICE_X17Y121_D3;
  wire [0:0] CLBLM_L_X12Y121_SLICE_X17Y121_D4;
  wire [0:0] CLBLM_L_X12Y121_SLICE_X17Y121_D5;
  wire [0:0] CLBLM_L_X12Y121_SLICE_X17Y121_D6;
  wire [0:0] CLBLM_L_X12Y121_SLICE_X17Y121_DO5;
  wire [0:0] CLBLM_L_X12Y121_SLICE_X17Y121_DO6;
  wire [0:0] CLBLM_L_X12Y121_SLICE_X17Y121_D_CY;
  wire [0:0] CLBLM_L_X12Y121_SLICE_X17Y121_D_XOR;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X10Y110_A;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X10Y110_A1;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X10Y110_A2;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X10Y110_A3;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X10Y110_A4;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X10Y110_A5;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X10Y110_A6;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X10Y110_AO5;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X10Y110_AO6;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X10Y110_AQ;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X10Y110_A_CY;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X10Y110_A_XOR;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X10Y110_B;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X10Y110_B1;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X10Y110_B2;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X10Y110_B3;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X10Y110_B4;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X10Y110_B5;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X10Y110_B6;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X10Y110_BO5;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X10Y110_BO6;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X10Y110_BQ;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X10Y110_B_CY;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X10Y110_B_XOR;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X10Y110_C;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X10Y110_C1;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X10Y110_C2;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X10Y110_C3;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X10Y110_C4;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X10Y110_C5;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X10Y110_C6;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X10Y110_CLK;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X10Y110_CO5;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X10Y110_CO6;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X10Y110_C_CY;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X10Y110_C_XOR;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X10Y110_D;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X10Y110_D1;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X10Y110_D2;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X10Y110_D3;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X10Y110_D4;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X10Y110_D5;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X10Y110_D6;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X10Y110_DO5;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X10Y110_DO6;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X10Y110_D_CY;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X10Y110_D_XOR;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X11Y110_A;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X11Y110_A1;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X11Y110_A2;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X11Y110_A3;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X11Y110_A4;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X11Y110_A5;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X11Y110_A6;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X11Y110_AO5;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X11Y110_AO6;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X11Y110_A_CY;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X11Y110_A_XOR;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X11Y110_B;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X11Y110_B1;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X11Y110_B2;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X11Y110_B3;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X11Y110_B4;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X11Y110_B5;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X11Y110_B6;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X11Y110_BO5;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X11Y110_BO6;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X11Y110_B_CY;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X11Y110_B_XOR;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X11Y110_C;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X11Y110_C1;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X11Y110_C2;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X11Y110_C3;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X11Y110_C4;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X11Y110_C5;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X11Y110_C6;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X11Y110_CO5;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X11Y110_CO6;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X11Y110_C_CY;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X11Y110_C_XOR;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X11Y110_D;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X11Y110_D1;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X11Y110_D2;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X11Y110_D3;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X11Y110_D4;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X11Y110_D5;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X11Y110_D6;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X11Y110_DO5;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X11Y110_DO6;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X11Y110_D_CY;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X11Y110_D_XOR;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X10Y111_A;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X10Y111_A1;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X10Y111_A2;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X10Y111_A3;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X10Y111_A4;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X10Y111_A5;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X10Y111_A6;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X10Y111_AO5;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X10Y111_AO6;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X10Y111_AQ;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X10Y111_A_CY;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X10Y111_A_XOR;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X10Y111_B;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X10Y111_B1;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X10Y111_B2;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X10Y111_B3;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X10Y111_B4;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X10Y111_B5;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X10Y111_B6;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X10Y111_BO5;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X10Y111_BO6;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X10Y111_B_CY;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X10Y111_B_XOR;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X10Y111_C;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X10Y111_C1;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X10Y111_C2;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X10Y111_C3;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X10Y111_C4;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X10Y111_C5;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X10Y111_C6;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X10Y111_CLK;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X10Y111_CO5;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X10Y111_CO6;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X10Y111_C_CY;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X10Y111_C_XOR;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X10Y111_D;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X10Y111_D1;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X10Y111_D2;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X10Y111_D3;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X10Y111_D4;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X10Y111_D5;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X10Y111_D6;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X10Y111_DO5;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X10Y111_DO6;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X10Y111_D_CY;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X10Y111_D_XOR;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X11Y111_A;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X11Y111_A1;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X11Y111_A2;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X11Y111_A3;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X11Y111_A4;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X11Y111_A5;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X11Y111_A6;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X11Y111_AO5;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X11Y111_AO6;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X11Y111_A_CY;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X11Y111_A_XOR;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X11Y111_B;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X11Y111_B1;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X11Y111_B2;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X11Y111_B3;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X11Y111_B4;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X11Y111_B5;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X11Y111_B6;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X11Y111_BO5;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X11Y111_BO6;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X11Y111_B_CY;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X11Y111_B_XOR;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X11Y111_C;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X11Y111_C1;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X11Y111_C2;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X11Y111_C3;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X11Y111_C4;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X11Y111_C5;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X11Y111_C6;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X11Y111_CO5;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X11Y111_CO6;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X11Y111_C_CY;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X11Y111_C_XOR;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X11Y111_D;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X11Y111_D1;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X11Y111_D2;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X11Y111_D3;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X11Y111_D4;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X11Y111_D5;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X11Y111_D6;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X11Y111_DO5;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X11Y111_DO6;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X11Y111_D_CY;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X11Y111_D_XOR;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X10Y112_A;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X10Y112_A1;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X10Y112_A2;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X10Y112_A3;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X10Y112_A4;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X10Y112_A5;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X10Y112_A6;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X10Y112_AO5;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X10Y112_AO6;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X10Y112_AQ;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X10Y112_A_CY;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X10Y112_A_XOR;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X10Y112_B;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X10Y112_B1;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X10Y112_B2;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X10Y112_B3;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X10Y112_B4;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X10Y112_B5;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X10Y112_B6;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X10Y112_BO5;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X10Y112_BO6;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X10Y112_BQ;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X10Y112_B_CY;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X10Y112_B_XOR;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X10Y112_C;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X10Y112_C1;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X10Y112_C2;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X10Y112_C3;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X10Y112_C4;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X10Y112_C5;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X10Y112_C6;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X10Y112_CLK;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X10Y112_CO5;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X10Y112_CO6;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X10Y112_CQ;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X10Y112_C_CY;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X10Y112_C_XOR;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X10Y112_D;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X10Y112_D1;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X10Y112_D2;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X10Y112_D3;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X10Y112_D4;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X10Y112_D5;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X10Y112_D6;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X10Y112_DO5;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X10Y112_DO6;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X10Y112_DQ;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X10Y112_D_CY;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X10Y112_D_XOR;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X11Y112_A;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X11Y112_A1;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X11Y112_A2;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X11Y112_A3;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X11Y112_A4;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X11Y112_A5;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X11Y112_A6;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X11Y112_AO5;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X11Y112_AO6;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X11Y112_AQ;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X11Y112_A_CY;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X11Y112_A_XOR;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X11Y112_B;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X11Y112_B1;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X11Y112_B2;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X11Y112_B3;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X11Y112_B4;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X11Y112_B5;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X11Y112_B6;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X11Y112_BMUX;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X11Y112_BO5;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X11Y112_BO6;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X11Y112_B_CY;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X11Y112_B_XOR;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X11Y112_C;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X11Y112_C1;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X11Y112_C2;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X11Y112_C3;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X11Y112_C4;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X11Y112_C5;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X11Y112_C6;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X11Y112_CLK;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X11Y112_CO5;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X11Y112_CO6;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X11Y112_C_CY;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X11Y112_C_XOR;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X11Y112_D;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X11Y112_D1;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X11Y112_D2;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X11Y112_D3;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X11Y112_D4;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X11Y112_D5;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X11Y112_D6;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X11Y112_DO5;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X11Y112_DO6;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X11Y112_D_CY;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X11Y112_D_XOR;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X10Y113_A;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X10Y113_A1;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X10Y113_A2;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X10Y113_A3;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X10Y113_A4;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X10Y113_A5;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X10Y113_A6;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X10Y113_AO5;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X10Y113_AO6;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X10Y113_A_CY;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X10Y113_A_XOR;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X10Y113_B;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X10Y113_B1;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X10Y113_B2;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X10Y113_B3;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X10Y113_B4;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X10Y113_B5;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X10Y113_B6;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X10Y113_BO5;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X10Y113_BO6;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X10Y113_B_CY;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X10Y113_B_XOR;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X10Y113_C;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X10Y113_C1;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X10Y113_C2;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X10Y113_C3;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X10Y113_C4;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X10Y113_C5;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X10Y113_C6;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X10Y113_CO5;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X10Y113_CO6;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X10Y113_C_CY;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X10Y113_C_XOR;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X10Y113_D;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X10Y113_D1;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X10Y113_D2;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X10Y113_D3;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X10Y113_D4;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X10Y113_D5;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X10Y113_D6;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X10Y113_DO5;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X10Y113_DO6;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X10Y113_D_CY;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X10Y113_D_XOR;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X11Y113_A;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X11Y113_A1;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X11Y113_A2;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X11Y113_A3;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X11Y113_A4;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X11Y113_A5;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X11Y113_A6;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X11Y113_AO5;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X11Y113_AO6;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X11Y113_AQ;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X11Y113_A_CY;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X11Y113_A_XOR;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X11Y113_B;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X11Y113_B1;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X11Y113_B2;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X11Y113_B3;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X11Y113_B4;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X11Y113_B5;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X11Y113_B6;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X11Y113_BO5;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X11Y113_BO6;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X11Y113_BQ;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X11Y113_B_CY;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X11Y113_B_XOR;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X11Y113_C;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X11Y113_C1;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X11Y113_C2;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X11Y113_C3;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X11Y113_C4;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X11Y113_C5;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X11Y113_C6;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X11Y113_CLK;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X11Y113_CO5;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X11Y113_CO6;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X11Y113_CQ;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X11Y113_C_CY;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X11Y113_C_XOR;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X11Y113_D;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X11Y113_D1;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X11Y113_D2;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X11Y113_D3;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X11Y113_D4;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X11Y113_D5;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X11Y113_D6;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X11Y113_DO5;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X11Y113_DO6;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X11Y113_D_CY;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X11Y113_D_XOR;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X10Y114_A;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X10Y114_A1;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X10Y114_A2;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X10Y114_A3;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X10Y114_A4;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X10Y114_A5;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X10Y114_A6;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X10Y114_AO5;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X10Y114_AO6;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X10Y114_AQ;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X10Y114_A_CY;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X10Y114_A_XOR;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X10Y114_B;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X10Y114_B1;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X10Y114_B2;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X10Y114_B3;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X10Y114_B4;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X10Y114_B5;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X10Y114_B5Q;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X10Y114_B6;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X10Y114_BMUX;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X10Y114_BO5;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X10Y114_BO6;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X10Y114_BQ;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X10Y114_B_CY;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X10Y114_B_XOR;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X10Y114_C;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X10Y114_C1;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X10Y114_C2;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X10Y114_C3;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X10Y114_C4;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X10Y114_C5;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X10Y114_C5Q;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X10Y114_C6;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X10Y114_CLK;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X10Y114_CMUX;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X10Y114_CO5;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X10Y114_CO6;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X10Y114_CQ;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X10Y114_C_CY;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X10Y114_C_XOR;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X10Y114_D;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X10Y114_D1;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X10Y114_D2;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X10Y114_D3;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X10Y114_D4;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X10Y114_D5;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X10Y114_D6;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X10Y114_DO5;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X10Y114_DO6;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X10Y114_DQ;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X10Y114_D_CY;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X10Y114_D_XOR;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X11Y114_A;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X11Y114_A1;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X11Y114_A2;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X11Y114_A3;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X11Y114_A4;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X11Y114_A5;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X11Y114_A6;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X11Y114_AO5;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X11Y114_AO6;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X11Y114_AQ;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X11Y114_A_CY;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X11Y114_A_XOR;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X11Y114_B;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X11Y114_B1;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X11Y114_B2;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X11Y114_B3;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X11Y114_B4;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X11Y114_B5;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X11Y114_B6;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X11Y114_BO5;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X11Y114_BO6;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X11Y114_BQ;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X11Y114_B_CY;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X11Y114_B_XOR;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X11Y114_C;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X11Y114_C1;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X11Y114_C2;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X11Y114_C3;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X11Y114_C4;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X11Y114_C5;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X11Y114_C6;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X11Y114_CLK;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X11Y114_CO5;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X11Y114_CO6;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X11Y114_CQ;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X11Y114_C_CY;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X11Y114_C_XOR;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X11Y114_D;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X11Y114_D1;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X11Y114_D2;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X11Y114_D3;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X11Y114_D4;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X11Y114_D5;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X11Y114_D6;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X11Y114_DO5;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X11Y114_DO6;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X11Y114_D_CY;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X11Y114_D_XOR;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X10Y115_A;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X10Y115_A1;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X10Y115_A2;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X10Y115_A3;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X10Y115_A4;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X10Y115_A5;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X10Y115_A6;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X10Y115_AO5;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X10Y115_AO6;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X10Y115_AQ;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X10Y115_A_CY;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X10Y115_A_XOR;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X10Y115_B;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X10Y115_B1;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X10Y115_B2;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X10Y115_B3;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X10Y115_B4;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X10Y115_B5;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X10Y115_B6;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X10Y115_BMUX;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X10Y115_BO5;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X10Y115_BO6;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X10Y115_B_CY;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X10Y115_B_XOR;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X10Y115_C;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X10Y115_C1;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X10Y115_C2;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X10Y115_C3;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X10Y115_C4;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X10Y115_C5;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X10Y115_C5Q;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X10Y115_C6;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X10Y115_CLK;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X10Y115_CMUX;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X10Y115_CO5;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X10Y115_CO6;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X10Y115_CQ;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X10Y115_C_CY;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X10Y115_C_XOR;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X10Y115_D;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X10Y115_D1;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X10Y115_D2;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X10Y115_D3;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X10Y115_D4;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X10Y115_D5;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X10Y115_D6;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X10Y115_DO5;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X10Y115_DO6;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X10Y115_DQ;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X10Y115_D_CY;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X10Y115_D_XOR;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X11Y115_A;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X11Y115_A1;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X11Y115_A2;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X11Y115_A3;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X11Y115_A4;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X11Y115_A5;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X11Y115_A6;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X11Y115_AO5;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X11Y115_AO6;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X11Y115_AQ;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X11Y115_A_CY;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X11Y115_A_XOR;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X11Y115_B;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X11Y115_B1;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X11Y115_B2;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X11Y115_B3;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X11Y115_B4;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X11Y115_B5;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X11Y115_B6;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X11Y115_BO5;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X11Y115_BO6;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X11Y115_BQ;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X11Y115_B_CY;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X11Y115_B_XOR;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X11Y115_C;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X11Y115_C1;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X11Y115_C2;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X11Y115_C3;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X11Y115_C4;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X11Y115_C5;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X11Y115_C5Q;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X11Y115_C6;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X11Y115_CLK;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X11Y115_CMUX;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X11Y115_CO5;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X11Y115_CO6;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X11Y115_CQ;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X11Y115_C_CY;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X11Y115_C_XOR;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X11Y115_D;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X11Y115_D1;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X11Y115_D2;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X11Y115_D3;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X11Y115_D4;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X11Y115_D5;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X11Y115_D6;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X11Y115_DO5;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X11Y115_DO6;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X11Y115_DQ;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X11Y115_D_CY;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X11Y115_D_XOR;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X10Y116_A;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X10Y116_A1;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X10Y116_A2;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X10Y116_A3;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X10Y116_A4;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X10Y116_A5;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X10Y116_A6;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X10Y116_AO5;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X10Y116_AO6;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X10Y116_AQ;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X10Y116_AX;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X10Y116_A_CY;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X10Y116_A_XOR;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X10Y116_B;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X10Y116_B1;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X10Y116_B2;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X10Y116_B3;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X10Y116_B4;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X10Y116_B5;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X10Y116_B6;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X10Y116_BO5;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X10Y116_BO6;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X10Y116_B_CY;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X10Y116_B_XOR;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X10Y116_C;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X10Y116_C1;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X10Y116_C2;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X10Y116_C3;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X10Y116_C4;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X10Y116_C5;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X10Y116_C6;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X10Y116_CE;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X10Y116_CLK;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X10Y116_CO5;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X10Y116_CO6;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X10Y116_C_CY;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X10Y116_C_XOR;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X10Y116_D;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X10Y116_D1;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X10Y116_D2;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X10Y116_D3;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X10Y116_D4;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X10Y116_D5;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X10Y116_D6;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X10Y116_DO5;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X10Y116_DO6;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X10Y116_D_CY;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X10Y116_D_XOR;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X10Y116_SR;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X11Y116_A;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X11Y116_A1;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X11Y116_A2;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X11Y116_A3;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X11Y116_A4;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X11Y116_A5;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X11Y116_A5Q;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X11Y116_A6;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X11Y116_AMUX;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X11Y116_AO5;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X11Y116_AO6;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X11Y116_AQ;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X11Y116_AX;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X11Y116_A_CY;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X11Y116_A_XOR;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X11Y116_B;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X11Y116_B1;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X11Y116_B2;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X11Y116_B3;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X11Y116_B4;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X11Y116_B5;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X11Y116_B6;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X11Y116_BO5;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X11Y116_BO6;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X11Y116_BQ;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X11Y116_B_CY;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X11Y116_B_XOR;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X11Y116_C;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X11Y116_C1;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X11Y116_C2;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X11Y116_C3;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X11Y116_C4;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X11Y116_C5;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X11Y116_C6;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X11Y116_CLK;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X11Y116_CMUX;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X11Y116_CO5;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X11Y116_CO6;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X11Y116_C_CY;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X11Y116_C_XOR;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X11Y116_D;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X11Y116_D1;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X11Y116_D2;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X11Y116_D3;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X11Y116_D4;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X11Y116_D5;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X11Y116_D6;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X11Y116_DO5;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X11Y116_DO6;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X11Y116_DQ;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X11Y116_D_CY;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X11Y116_D_XOR;
  wire [0:0] CLBLM_L_X8Y117_SLICE_X10Y117_A;
  wire [0:0] CLBLM_L_X8Y117_SLICE_X10Y117_A1;
  wire [0:0] CLBLM_L_X8Y117_SLICE_X10Y117_A2;
  wire [0:0] CLBLM_L_X8Y117_SLICE_X10Y117_A3;
  wire [0:0] CLBLM_L_X8Y117_SLICE_X10Y117_A4;
  wire [0:0] CLBLM_L_X8Y117_SLICE_X10Y117_A5;
  wire [0:0] CLBLM_L_X8Y117_SLICE_X10Y117_A6;
  wire [0:0] CLBLM_L_X8Y117_SLICE_X10Y117_AO5;
  wire [0:0] CLBLM_L_X8Y117_SLICE_X10Y117_AO6;
  wire [0:0] CLBLM_L_X8Y117_SLICE_X10Y117_AQ;
  wire [0:0] CLBLM_L_X8Y117_SLICE_X10Y117_A_CY;
  wire [0:0] CLBLM_L_X8Y117_SLICE_X10Y117_A_XOR;
  wire [0:0] CLBLM_L_X8Y117_SLICE_X10Y117_B;
  wire [0:0] CLBLM_L_X8Y117_SLICE_X10Y117_B1;
  wire [0:0] CLBLM_L_X8Y117_SLICE_X10Y117_B2;
  wire [0:0] CLBLM_L_X8Y117_SLICE_X10Y117_B3;
  wire [0:0] CLBLM_L_X8Y117_SLICE_X10Y117_B4;
  wire [0:0] CLBLM_L_X8Y117_SLICE_X10Y117_B5;
  wire [0:0] CLBLM_L_X8Y117_SLICE_X10Y117_B6;
  wire [0:0] CLBLM_L_X8Y117_SLICE_X10Y117_BO5;
  wire [0:0] CLBLM_L_X8Y117_SLICE_X10Y117_BO6;
  wire [0:0] CLBLM_L_X8Y117_SLICE_X10Y117_BQ;
  wire [0:0] CLBLM_L_X8Y117_SLICE_X10Y117_B_CY;
  wire [0:0] CLBLM_L_X8Y117_SLICE_X10Y117_B_XOR;
  wire [0:0] CLBLM_L_X8Y117_SLICE_X10Y117_C;
  wire [0:0] CLBLM_L_X8Y117_SLICE_X10Y117_C1;
  wire [0:0] CLBLM_L_X8Y117_SLICE_X10Y117_C2;
  wire [0:0] CLBLM_L_X8Y117_SLICE_X10Y117_C3;
  wire [0:0] CLBLM_L_X8Y117_SLICE_X10Y117_C4;
  wire [0:0] CLBLM_L_X8Y117_SLICE_X10Y117_C5;
  wire [0:0] CLBLM_L_X8Y117_SLICE_X10Y117_C6;
  wire [0:0] CLBLM_L_X8Y117_SLICE_X10Y117_CLK;
  wire [0:0] CLBLM_L_X8Y117_SLICE_X10Y117_CO5;
  wire [0:0] CLBLM_L_X8Y117_SLICE_X10Y117_CO6;
  wire [0:0] CLBLM_L_X8Y117_SLICE_X10Y117_CQ;
  wire [0:0] CLBLM_L_X8Y117_SLICE_X10Y117_C_CY;
  wire [0:0] CLBLM_L_X8Y117_SLICE_X10Y117_C_XOR;
  wire [0:0] CLBLM_L_X8Y117_SLICE_X10Y117_D;
  wire [0:0] CLBLM_L_X8Y117_SLICE_X10Y117_D1;
  wire [0:0] CLBLM_L_X8Y117_SLICE_X10Y117_D2;
  wire [0:0] CLBLM_L_X8Y117_SLICE_X10Y117_D3;
  wire [0:0] CLBLM_L_X8Y117_SLICE_X10Y117_D4;
  wire [0:0] CLBLM_L_X8Y117_SLICE_X10Y117_D5;
  wire [0:0] CLBLM_L_X8Y117_SLICE_X10Y117_D6;
  wire [0:0] CLBLM_L_X8Y117_SLICE_X10Y117_DMUX;
  wire [0:0] CLBLM_L_X8Y117_SLICE_X10Y117_DO5;
  wire [0:0] CLBLM_L_X8Y117_SLICE_X10Y117_DO6;
  wire [0:0] CLBLM_L_X8Y117_SLICE_X10Y117_D_CY;
  wire [0:0] CLBLM_L_X8Y117_SLICE_X10Y117_D_XOR;
  wire [0:0] CLBLM_L_X8Y117_SLICE_X11Y117_A;
  wire [0:0] CLBLM_L_X8Y117_SLICE_X11Y117_A1;
  wire [0:0] CLBLM_L_X8Y117_SLICE_X11Y117_A2;
  wire [0:0] CLBLM_L_X8Y117_SLICE_X11Y117_A3;
  wire [0:0] CLBLM_L_X8Y117_SLICE_X11Y117_A4;
  wire [0:0] CLBLM_L_X8Y117_SLICE_X11Y117_A5;
  wire [0:0] CLBLM_L_X8Y117_SLICE_X11Y117_A6;
  wire [0:0] CLBLM_L_X8Y117_SLICE_X11Y117_AO5;
  wire [0:0] CLBLM_L_X8Y117_SLICE_X11Y117_AO6;
  wire [0:0] CLBLM_L_X8Y117_SLICE_X11Y117_AQ;
  wire [0:0] CLBLM_L_X8Y117_SLICE_X11Y117_A_CY;
  wire [0:0] CLBLM_L_X8Y117_SLICE_X11Y117_A_XOR;
  wire [0:0] CLBLM_L_X8Y117_SLICE_X11Y117_B;
  wire [0:0] CLBLM_L_X8Y117_SLICE_X11Y117_B1;
  wire [0:0] CLBLM_L_X8Y117_SLICE_X11Y117_B2;
  wire [0:0] CLBLM_L_X8Y117_SLICE_X11Y117_B3;
  wire [0:0] CLBLM_L_X8Y117_SLICE_X11Y117_B4;
  wire [0:0] CLBLM_L_X8Y117_SLICE_X11Y117_B5;
  wire [0:0] CLBLM_L_X8Y117_SLICE_X11Y117_B6;
  wire [0:0] CLBLM_L_X8Y117_SLICE_X11Y117_BO5;
  wire [0:0] CLBLM_L_X8Y117_SLICE_X11Y117_BO6;
  wire [0:0] CLBLM_L_X8Y117_SLICE_X11Y117_BQ;
  wire [0:0] CLBLM_L_X8Y117_SLICE_X11Y117_B_CY;
  wire [0:0] CLBLM_L_X8Y117_SLICE_X11Y117_B_XOR;
  wire [0:0] CLBLM_L_X8Y117_SLICE_X11Y117_C;
  wire [0:0] CLBLM_L_X8Y117_SLICE_X11Y117_C1;
  wire [0:0] CLBLM_L_X8Y117_SLICE_X11Y117_C2;
  wire [0:0] CLBLM_L_X8Y117_SLICE_X11Y117_C3;
  wire [0:0] CLBLM_L_X8Y117_SLICE_X11Y117_C4;
  wire [0:0] CLBLM_L_X8Y117_SLICE_X11Y117_C5;
  wire [0:0] CLBLM_L_X8Y117_SLICE_X11Y117_C6;
  wire [0:0] CLBLM_L_X8Y117_SLICE_X11Y117_CLK;
  wire [0:0] CLBLM_L_X8Y117_SLICE_X11Y117_CO5;
  wire [0:0] CLBLM_L_X8Y117_SLICE_X11Y117_CO6;
  wire [0:0] CLBLM_L_X8Y117_SLICE_X11Y117_CQ;
  wire [0:0] CLBLM_L_X8Y117_SLICE_X11Y117_C_CY;
  wire [0:0] CLBLM_L_X8Y117_SLICE_X11Y117_C_XOR;
  wire [0:0] CLBLM_L_X8Y117_SLICE_X11Y117_D;
  wire [0:0] CLBLM_L_X8Y117_SLICE_X11Y117_D1;
  wire [0:0] CLBLM_L_X8Y117_SLICE_X11Y117_D2;
  wire [0:0] CLBLM_L_X8Y117_SLICE_X11Y117_D3;
  wire [0:0] CLBLM_L_X8Y117_SLICE_X11Y117_D4;
  wire [0:0] CLBLM_L_X8Y117_SLICE_X11Y117_D5;
  wire [0:0] CLBLM_L_X8Y117_SLICE_X11Y117_D6;
  wire [0:0] CLBLM_L_X8Y117_SLICE_X11Y117_DO5;
  wire [0:0] CLBLM_L_X8Y117_SLICE_X11Y117_DO6;
  wire [0:0] CLBLM_L_X8Y117_SLICE_X11Y117_DQ;
  wire [0:0] CLBLM_L_X8Y117_SLICE_X11Y117_D_CY;
  wire [0:0] CLBLM_L_X8Y117_SLICE_X11Y117_D_XOR;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X10Y118_A;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X10Y118_A1;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X10Y118_A2;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X10Y118_A3;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X10Y118_A4;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X10Y118_A5;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X10Y118_A6;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X10Y118_AO5;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X10Y118_AO6;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X10Y118_AQ;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X10Y118_A_CY;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X10Y118_A_XOR;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X10Y118_B;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X10Y118_B1;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X10Y118_B2;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X10Y118_B3;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X10Y118_B4;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X10Y118_B5;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X10Y118_B6;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X10Y118_BO5;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X10Y118_BO6;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X10Y118_BQ;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X10Y118_B_CY;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X10Y118_B_XOR;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X10Y118_C;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X10Y118_C1;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X10Y118_C2;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X10Y118_C3;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X10Y118_C4;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X10Y118_C5;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X10Y118_C6;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X10Y118_CLK;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X10Y118_CO5;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X10Y118_CO6;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X10Y118_CQ;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X10Y118_C_CY;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X10Y118_C_XOR;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X10Y118_D;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X10Y118_D1;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X10Y118_D2;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X10Y118_D3;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X10Y118_D4;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X10Y118_D5;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X10Y118_D5Q;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X10Y118_D6;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X10Y118_DMUX;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X10Y118_DO5;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X10Y118_DO6;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X10Y118_DQ;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X10Y118_D_CY;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X10Y118_D_XOR;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X11Y118_A;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X11Y118_A1;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X11Y118_A2;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X11Y118_A3;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X11Y118_A4;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X11Y118_A5;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X11Y118_A6;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X11Y118_AO5;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X11Y118_AO6;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X11Y118_AQ;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X11Y118_A_CY;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X11Y118_A_XOR;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X11Y118_B;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X11Y118_B1;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X11Y118_B2;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X11Y118_B3;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X11Y118_B4;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X11Y118_B5;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X11Y118_B6;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X11Y118_BMUX;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X11Y118_BO5;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X11Y118_BO6;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X11Y118_B_CY;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X11Y118_B_XOR;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X11Y118_C;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X11Y118_C1;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X11Y118_C2;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X11Y118_C3;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X11Y118_C4;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X11Y118_C5;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X11Y118_C6;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X11Y118_CLK;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X11Y118_CO5;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X11Y118_CO6;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X11Y118_C_CY;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X11Y118_C_XOR;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X11Y118_D;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X11Y118_D1;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X11Y118_D2;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X11Y118_D3;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X11Y118_D4;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X11Y118_D5;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X11Y118_D6;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X11Y118_DO5;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X11Y118_DO6;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X11Y118_D_CY;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X11Y118_D_XOR;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X10Y119_A;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X10Y119_A1;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X10Y119_A2;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X10Y119_A3;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X10Y119_A4;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X10Y119_A5;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X10Y119_A5Q;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X10Y119_A6;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X10Y119_AMUX;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X10Y119_AO5;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X10Y119_AO6;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X10Y119_AQ;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X10Y119_AX;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X10Y119_A_CY;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X10Y119_A_XOR;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X10Y119_B;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X10Y119_B1;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X10Y119_B2;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X10Y119_B3;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X10Y119_B4;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X10Y119_B5;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X10Y119_B6;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X10Y119_BO5;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X10Y119_BO6;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X10Y119_BQ;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X10Y119_B_CY;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X10Y119_B_XOR;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X10Y119_C;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X10Y119_C1;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X10Y119_C2;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X10Y119_C3;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X10Y119_C4;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X10Y119_C5;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X10Y119_C6;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X10Y119_CLK;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X10Y119_CO5;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X10Y119_CO6;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X10Y119_CQ;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X10Y119_C_CY;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X10Y119_C_XOR;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X10Y119_D;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X10Y119_D1;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X10Y119_D2;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X10Y119_D3;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X10Y119_D4;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X10Y119_D5;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X10Y119_D6;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X10Y119_DMUX;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X10Y119_DO5;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X10Y119_DO6;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X10Y119_D_CY;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X10Y119_D_XOR;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X11Y119_A;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X11Y119_A1;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X11Y119_A2;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X11Y119_A3;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X11Y119_A4;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X11Y119_A5;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X11Y119_A6;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X11Y119_AO5;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X11Y119_AO6;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X11Y119_AQ;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X11Y119_A_CY;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X11Y119_A_XOR;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X11Y119_B;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X11Y119_B1;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X11Y119_B2;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X11Y119_B3;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X11Y119_B4;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X11Y119_B5;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X11Y119_B6;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X11Y119_BO5;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X11Y119_BO6;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X11Y119_BQ;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X11Y119_B_CY;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X11Y119_B_XOR;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X11Y119_C;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X11Y119_C1;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X11Y119_C2;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X11Y119_C3;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X11Y119_C4;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X11Y119_C5;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X11Y119_C5Q;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X11Y119_C6;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X11Y119_CLK;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X11Y119_CMUX;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X11Y119_CO5;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X11Y119_CO6;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X11Y119_CQ;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X11Y119_C_CY;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X11Y119_C_XOR;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X11Y119_D;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X11Y119_D1;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X11Y119_D2;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X11Y119_D3;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X11Y119_D4;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X11Y119_D5;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X11Y119_D6;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X11Y119_DO5;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X11Y119_DO6;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X11Y119_DQ;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X11Y119_D_CY;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X11Y119_D_XOR;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X10Y120_A;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X10Y120_A1;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X10Y120_A2;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X10Y120_A3;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X10Y120_A4;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X10Y120_A5;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X10Y120_A5Q;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X10Y120_A6;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X10Y120_AMUX;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X10Y120_AO5;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X10Y120_AO6;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X10Y120_AQ;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X10Y120_A_CY;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X10Y120_A_XOR;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X10Y120_B;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X10Y120_B1;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X10Y120_B2;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X10Y120_B3;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X10Y120_B4;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X10Y120_B5;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X10Y120_B6;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X10Y120_BO5;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X10Y120_BO6;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X10Y120_BQ;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X10Y120_B_CY;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X10Y120_B_XOR;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X10Y120_C;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X10Y120_C1;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X10Y120_C2;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X10Y120_C3;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X10Y120_C4;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X10Y120_C5;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X10Y120_C6;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X10Y120_CLK;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X10Y120_CO5;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X10Y120_CO6;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X10Y120_CQ;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X10Y120_C_CY;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X10Y120_C_XOR;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X10Y120_D;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X10Y120_D1;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X10Y120_D2;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X10Y120_D3;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X10Y120_D4;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X10Y120_D5;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X10Y120_D5Q;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X10Y120_D6;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X10Y120_DMUX;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X10Y120_DO5;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X10Y120_DO6;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X10Y120_DQ;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X10Y120_D_CY;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X10Y120_D_XOR;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X11Y120_A;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X11Y120_A1;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X11Y120_A2;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X11Y120_A3;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X11Y120_A4;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X11Y120_A5;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X11Y120_A6;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X11Y120_AO5;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X11Y120_AO6;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X11Y120_AQ;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X11Y120_A_CY;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X11Y120_A_XOR;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X11Y120_B;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X11Y120_B1;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X11Y120_B2;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X11Y120_B3;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X11Y120_B4;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X11Y120_B5;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X11Y120_B6;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X11Y120_BO5;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X11Y120_BO6;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X11Y120_BQ;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X11Y120_B_CY;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X11Y120_B_XOR;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X11Y120_C;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X11Y120_C1;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X11Y120_C2;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X11Y120_C3;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X11Y120_C4;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X11Y120_C5;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X11Y120_C5Q;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X11Y120_C6;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X11Y120_CLK;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X11Y120_CMUX;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X11Y120_CO5;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X11Y120_CO6;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X11Y120_CQ;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X11Y120_C_CY;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X11Y120_C_XOR;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X11Y120_D;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X11Y120_D1;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X11Y120_D2;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X11Y120_D3;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X11Y120_D4;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X11Y120_D5;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X11Y120_D6;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X11Y120_DO5;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X11Y120_DO6;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X11Y120_D_CY;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X11Y120_D_XOR;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X10Y121_A;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X10Y121_A1;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X10Y121_A2;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X10Y121_A3;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X10Y121_A4;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X10Y121_A5;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X10Y121_A6;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X10Y121_AO5;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X10Y121_AO6;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X10Y121_AQ;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X10Y121_A_CY;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X10Y121_A_XOR;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X10Y121_B;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X10Y121_B1;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X10Y121_B2;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X10Y121_B3;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X10Y121_B4;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X10Y121_B5;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X10Y121_B6;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X10Y121_BO5;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X10Y121_BO6;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X10Y121_BQ;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X10Y121_B_CY;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X10Y121_B_XOR;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X10Y121_C;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X10Y121_C1;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X10Y121_C2;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X10Y121_C3;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X10Y121_C4;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X10Y121_C5;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X10Y121_C6;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X10Y121_CLK;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X10Y121_CO5;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X10Y121_CO6;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X10Y121_CQ;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X10Y121_C_CY;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X10Y121_C_XOR;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X10Y121_D;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X10Y121_D1;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X10Y121_D2;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X10Y121_D3;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X10Y121_D4;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X10Y121_D5;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X10Y121_D6;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X10Y121_DO5;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X10Y121_DO6;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X10Y121_D_CY;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X10Y121_D_XOR;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X11Y121_A;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X11Y121_A1;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X11Y121_A2;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X11Y121_A3;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X11Y121_A4;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X11Y121_A5;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X11Y121_A6;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X11Y121_AO5;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X11Y121_AO6;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X11Y121_AQ;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X11Y121_A_CY;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X11Y121_A_XOR;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X11Y121_B;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X11Y121_B1;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X11Y121_B2;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X11Y121_B3;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X11Y121_B4;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X11Y121_B5;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X11Y121_B6;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X11Y121_BO5;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X11Y121_BO6;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X11Y121_BQ;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X11Y121_B_CY;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X11Y121_B_XOR;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X11Y121_C;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X11Y121_C1;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X11Y121_C2;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X11Y121_C3;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X11Y121_C4;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X11Y121_C5;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X11Y121_C6;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X11Y121_CLK;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X11Y121_CO5;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X11Y121_CO6;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X11Y121_CQ;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X11Y121_C_CY;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X11Y121_C_XOR;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X11Y121_D;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X11Y121_D1;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X11Y121_D2;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X11Y121_D3;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X11Y121_D4;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X11Y121_D5;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X11Y121_D6;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X11Y121_DO5;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X11Y121_DO6;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X11Y121_DQ;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X11Y121_D_CY;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X11Y121_D_XOR;
  wire [0:0] CLBLM_L_X8Y122_SLICE_X10Y122_A;
  wire [0:0] CLBLM_L_X8Y122_SLICE_X10Y122_A1;
  wire [0:0] CLBLM_L_X8Y122_SLICE_X10Y122_A2;
  wire [0:0] CLBLM_L_X8Y122_SLICE_X10Y122_A3;
  wire [0:0] CLBLM_L_X8Y122_SLICE_X10Y122_A4;
  wire [0:0] CLBLM_L_X8Y122_SLICE_X10Y122_A5;
  wire [0:0] CLBLM_L_X8Y122_SLICE_X10Y122_A6;
  wire [0:0] CLBLM_L_X8Y122_SLICE_X10Y122_AMUX;
  wire [0:0] CLBLM_L_X8Y122_SLICE_X10Y122_AO5;
  wire [0:0] CLBLM_L_X8Y122_SLICE_X10Y122_AO6;
  wire [0:0] CLBLM_L_X8Y122_SLICE_X10Y122_AQ;
  wire [0:0] CLBLM_L_X8Y122_SLICE_X10Y122_AX;
  wire [0:0] CLBLM_L_X8Y122_SLICE_X10Y122_A_CY;
  wire [0:0] CLBLM_L_X8Y122_SLICE_X10Y122_A_XOR;
  wire [0:0] CLBLM_L_X8Y122_SLICE_X10Y122_B;
  wire [0:0] CLBLM_L_X8Y122_SLICE_X10Y122_B1;
  wire [0:0] CLBLM_L_X8Y122_SLICE_X10Y122_B2;
  wire [0:0] CLBLM_L_X8Y122_SLICE_X10Y122_B3;
  wire [0:0] CLBLM_L_X8Y122_SLICE_X10Y122_B4;
  wire [0:0] CLBLM_L_X8Y122_SLICE_X10Y122_B5;
  wire [0:0] CLBLM_L_X8Y122_SLICE_X10Y122_B6;
  wire [0:0] CLBLM_L_X8Y122_SLICE_X10Y122_BMUX;
  wire [0:0] CLBLM_L_X8Y122_SLICE_X10Y122_BO5;
  wire [0:0] CLBLM_L_X8Y122_SLICE_X10Y122_BO6;
  wire [0:0] CLBLM_L_X8Y122_SLICE_X10Y122_B_CY;
  wire [0:0] CLBLM_L_X8Y122_SLICE_X10Y122_B_XOR;
  wire [0:0] CLBLM_L_X8Y122_SLICE_X10Y122_C;
  wire [0:0] CLBLM_L_X8Y122_SLICE_X10Y122_C1;
  wire [0:0] CLBLM_L_X8Y122_SLICE_X10Y122_C2;
  wire [0:0] CLBLM_L_X8Y122_SLICE_X10Y122_C3;
  wire [0:0] CLBLM_L_X8Y122_SLICE_X10Y122_C4;
  wire [0:0] CLBLM_L_X8Y122_SLICE_X10Y122_C5;
  wire [0:0] CLBLM_L_X8Y122_SLICE_X10Y122_C6;
  wire [0:0] CLBLM_L_X8Y122_SLICE_X10Y122_CE;
  wire [0:0] CLBLM_L_X8Y122_SLICE_X10Y122_CLK;
  wire [0:0] CLBLM_L_X8Y122_SLICE_X10Y122_CO5;
  wire [0:0] CLBLM_L_X8Y122_SLICE_X10Y122_CO6;
  wire [0:0] CLBLM_L_X8Y122_SLICE_X10Y122_C_CY;
  wire [0:0] CLBLM_L_X8Y122_SLICE_X10Y122_C_XOR;
  wire [0:0] CLBLM_L_X8Y122_SLICE_X10Y122_D;
  wire [0:0] CLBLM_L_X8Y122_SLICE_X10Y122_D1;
  wire [0:0] CLBLM_L_X8Y122_SLICE_X10Y122_D2;
  wire [0:0] CLBLM_L_X8Y122_SLICE_X10Y122_D3;
  wire [0:0] CLBLM_L_X8Y122_SLICE_X10Y122_D4;
  wire [0:0] CLBLM_L_X8Y122_SLICE_X10Y122_D5;
  wire [0:0] CLBLM_L_X8Y122_SLICE_X10Y122_D6;
  wire [0:0] CLBLM_L_X8Y122_SLICE_X10Y122_DO5;
  wire [0:0] CLBLM_L_X8Y122_SLICE_X10Y122_DO6;
  wire [0:0] CLBLM_L_X8Y122_SLICE_X10Y122_D_CY;
  wire [0:0] CLBLM_L_X8Y122_SLICE_X10Y122_D_XOR;
  wire [0:0] CLBLM_L_X8Y122_SLICE_X10Y122_SR;
  wire [0:0] CLBLM_L_X8Y122_SLICE_X11Y122_A;
  wire [0:0] CLBLM_L_X8Y122_SLICE_X11Y122_A1;
  wire [0:0] CLBLM_L_X8Y122_SLICE_X11Y122_A2;
  wire [0:0] CLBLM_L_X8Y122_SLICE_X11Y122_A3;
  wire [0:0] CLBLM_L_X8Y122_SLICE_X11Y122_A4;
  wire [0:0] CLBLM_L_X8Y122_SLICE_X11Y122_A5;
  wire [0:0] CLBLM_L_X8Y122_SLICE_X11Y122_A5Q;
  wire [0:0] CLBLM_L_X8Y122_SLICE_X11Y122_A6;
  wire [0:0] CLBLM_L_X8Y122_SLICE_X11Y122_AMUX;
  wire [0:0] CLBLM_L_X8Y122_SLICE_X11Y122_AO5;
  wire [0:0] CLBLM_L_X8Y122_SLICE_X11Y122_AO6;
  wire [0:0] CLBLM_L_X8Y122_SLICE_X11Y122_AQ;
  wire [0:0] CLBLM_L_X8Y122_SLICE_X11Y122_AX;
  wire [0:0] CLBLM_L_X8Y122_SLICE_X11Y122_A_CY;
  wire [0:0] CLBLM_L_X8Y122_SLICE_X11Y122_A_XOR;
  wire [0:0] CLBLM_L_X8Y122_SLICE_X11Y122_B;
  wire [0:0] CLBLM_L_X8Y122_SLICE_X11Y122_B1;
  wire [0:0] CLBLM_L_X8Y122_SLICE_X11Y122_B2;
  wire [0:0] CLBLM_L_X8Y122_SLICE_X11Y122_B3;
  wire [0:0] CLBLM_L_X8Y122_SLICE_X11Y122_B4;
  wire [0:0] CLBLM_L_X8Y122_SLICE_X11Y122_B5;
  wire [0:0] CLBLM_L_X8Y122_SLICE_X11Y122_B6;
  wire [0:0] CLBLM_L_X8Y122_SLICE_X11Y122_BO5;
  wire [0:0] CLBLM_L_X8Y122_SLICE_X11Y122_BO6;
  wire [0:0] CLBLM_L_X8Y122_SLICE_X11Y122_BQ;
  wire [0:0] CLBLM_L_X8Y122_SLICE_X11Y122_B_CY;
  wire [0:0] CLBLM_L_X8Y122_SLICE_X11Y122_B_XOR;
  wire [0:0] CLBLM_L_X8Y122_SLICE_X11Y122_C;
  wire [0:0] CLBLM_L_X8Y122_SLICE_X11Y122_C1;
  wire [0:0] CLBLM_L_X8Y122_SLICE_X11Y122_C2;
  wire [0:0] CLBLM_L_X8Y122_SLICE_X11Y122_C3;
  wire [0:0] CLBLM_L_X8Y122_SLICE_X11Y122_C4;
  wire [0:0] CLBLM_L_X8Y122_SLICE_X11Y122_C5;
  wire [0:0] CLBLM_L_X8Y122_SLICE_X11Y122_C6;
  wire [0:0] CLBLM_L_X8Y122_SLICE_X11Y122_CLK;
  wire [0:0] CLBLM_L_X8Y122_SLICE_X11Y122_CO5;
  wire [0:0] CLBLM_L_X8Y122_SLICE_X11Y122_CO6;
  wire [0:0] CLBLM_L_X8Y122_SLICE_X11Y122_C_CY;
  wire [0:0] CLBLM_L_X8Y122_SLICE_X11Y122_C_XOR;
  wire [0:0] CLBLM_L_X8Y122_SLICE_X11Y122_D;
  wire [0:0] CLBLM_L_X8Y122_SLICE_X11Y122_D1;
  wire [0:0] CLBLM_L_X8Y122_SLICE_X11Y122_D2;
  wire [0:0] CLBLM_L_X8Y122_SLICE_X11Y122_D3;
  wire [0:0] CLBLM_L_X8Y122_SLICE_X11Y122_D4;
  wire [0:0] CLBLM_L_X8Y122_SLICE_X11Y122_D5;
  wire [0:0] CLBLM_L_X8Y122_SLICE_X11Y122_D6;
  wire [0:0] CLBLM_L_X8Y122_SLICE_X11Y122_DO5;
  wire [0:0] CLBLM_L_X8Y122_SLICE_X11Y122_DO6;
  wire [0:0] CLBLM_L_X8Y122_SLICE_X11Y122_D_CY;
  wire [0:0] CLBLM_L_X8Y122_SLICE_X11Y122_D_XOR;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X10Y123_A;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X10Y123_A1;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X10Y123_A2;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X10Y123_A3;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X10Y123_A4;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X10Y123_A5;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X10Y123_A5Q;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X10Y123_A6;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X10Y123_AMUX;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X10Y123_AO5;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X10Y123_AO6;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X10Y123_AQ;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X10Y123_A_CY;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X10Y123_A_XOR;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X10Y123_B;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X10Y123_B1;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X10Y123_B2;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X10Y123_B3;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X10Y123_B4;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X10Y123_B5;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X10Y123_B5Q;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X10Y123_B6;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X10Y123_BMUX;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X10Y123_BO5;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X10Y123_BO6;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X10Y123_BQ;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X10Y123_B_CY;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X10Y123_B_XOR;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X10Y123_C;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X10Y123_C1;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X10Y123_C2;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X10Y123_C3;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X10Y123_C4;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X10Y123_C5;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X10Y123_C6;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X10Y123_CLK;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X10Y123_CO5;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X10Y123_CO6;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X10Y123_C_CY;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X10Y123_C_XOR;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X10Y123_D;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X10Y123_D1;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X10Y123_D2;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X10Y123_D3;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X10Y123_D4;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X10Y123_D5;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X10Y123_D6;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X10Y123_DO5;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X10Y123_DO6;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X10Y123_D_CY;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X10Y123_D_XOR;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X11Y123_A;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X11Y123_A1;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X11Y123_A2;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X11Y123_A3;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X11Y123_A4;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X11Y123_A5;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X11Y123_A5Q;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X11Y123_A6;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X11Y123_AMUX;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X11Y123_AO5;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X11Y123_AO6;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X11Y123_AQ;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X11Y123_A_CY;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X11Y123_A_XOR;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X11Y123_B;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X11Y123_B1;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X11Y123_B2;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X11Y123_B3;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X11Y123_B4;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X11Y123_B5;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X11Y123_B6;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X11Y123_BO5;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X11Y123_BO6;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X11Y123_B_CY;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X11Y123_B_XOR;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X11Y123_C;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X11Y123_C1;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X11Y123_C2;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X11Y123_C3;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X11Y123_C4;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X11Y123_C5;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X11Y123_C6;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X11Y123_CLK;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X11Y123_CO5;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X11Y123_CO6;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X11Y123_C_CY;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X11Y123_C_XOR;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X11Y123_D;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X11Y123_D1;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X11Y123_D2;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X11Y123_D3;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X11Y123_D4;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X11Y123_D5;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X11Y123_D6;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X11Y123_DO5;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X11Y123_DO6;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X11Y123_D_CY;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X11Y123_D_XOR;
  wire [0:0] CLBLM_L_X8Y128_SLICE_X10Y128_A;
  wire [0:0] CLBLM_L_X8Y128_SLICE_X10Y128_A1;
  wire [0:0] CLBLM_L_X8Y128_SLICE_X10Y128_A2;
  wire [0:0] CLBLM_L_X8Y128_SLICE_X10Y128_A3;
  wire [0:0] CLBLM_L_X8Y128_SLICE_X10Y128_A4;
  wire [0:0] CLBLM_L_X8Y128_SLICE_X10Y128_A5;
  wire [0:0] CLBLM_L_X8Y128_SLICE_X10Y128_A6;
  wire [0:0] CLBLM_L_X8Y128_SLICE_X10Y128_AMUX;
  wire [0:0] CLBLM_L_X8Y128_SLICE_X10Y128_AO5;
  wire [0:0] CLBLM_L_X8Y128_SLICE_X10Y128_AO6;
  wire [0:0] CLBLM_L_X8Y128_SLICE_X10Y128_A_CY;
  wire [0:0] CLBLM_L_X8Y128_SLICE_X10Y128_A_XOR;
  wire [0:0] CLBLM_L_X8Y128_SLICE_X10Y128_B;
  wire [0:0] CLBLM_L_X8Y128_SLICE_X10Y128_B1;
  wire [0:0] CLBLM_L_X8Y128_SLICE_X10Y128_B2;
  wire [0:0] CLBLM_L_X8Y128_SLICE_X10Y128_B3;
  wire [0:0] CLBLM_L_X8Y128_SLICE_X10Y128_B4;
  wire [0:0] CLBLM_L_X8Y128_SLICE_X10Y128_B5;
  wire [0:0] CLBLM_L_X8Y128_SLICE_X10Y128_B6;
  wire [0:0] CLBLM_L_X8Y128_SLICE_X10Y128_BO5;
  wire [0:0] CLBLM_L_X8Y128_SLICE_X10Y128_BO6;
  wire [0:0] CLBLM_L_X8Y128_SLICE_X10Y128_B_CY;
  wire [0:0] CLBLM_L_X8Y128_SLICE_X10Y128_B_XOR;
  wire [0:0] CLBLM_L_X8Y128_SLICE_X10Y128_C;
  wire [0:0] CLBLM_L_X8Y128_SLICE_X10Y128_C1;
  wire [0:0] CLBLM_L_X8Y128_SLICE_X10Y128_C2;
  wire [0:0] CLBLM_L_X8Y128_SLICE_X10Y128_C3;
  wire [0:0] CLBLM_L_X8Y128_SLICE_X10Y128_C4;
  wire [0:0] CLBLM_L_X8Y128_SLICE_X10Y128_C5;
  wire [0:0] CLBLM_L_X8Y128_SLICE_X10Y128_C6;
  wire [0:0] CLBLM_L_X8Y128_SLICE_X10Y128_CO5;
  wire [0:0] CLBLM_L_X8Y128_SLICE_X10Y128_CO6;
  wire [0:0] CLBLM_L_X8Y128_SLICE_X10Y128_C_CY;
  wire [0:0] CLBLM_L_X8Y128_SLICE_X10Y128_C_XOR;
  wire [0:0] CLBLM_L_X8Y128_SLICE_X10Y128_D;
  wire [0:0] CLBLM_L_X8Y128_SLICE_X10Y128_D1;
  wire [0:0] CLBLM_L_X8Y128_SLICE_X10Y128_D2;
  wire [0:0] CLBLM_L_X8Y128_SLICE_X10Y128_D3;
  wire [0:0] CLBLM_L_X8Y128_SLICE_X10Y128_D4;
  wire [0:0] CLBLM_L_X8Y128_SLICE_X10Y128_D5;
  wire [0:0] CLBLM_L_X8Y128_SLICE_X10Y128_D6;
  wire [0:0] CLBLM_L_X8Y128_SLICE_X10Y128_DO5;
  wire [0:0] CLBLM_L_X8Y128_SLICE_X10Y128_DO6;
  wire [0:0] CLBLM_L_X8Y128_SLICE_X10Y128_D_CY;
  wire [0:0] CLBLM_L_X8Y128_SLICE_X10Y128_D_XOR;
  wire [0:0] CLBLM_L_X8Y128_SLICE_X11Y128_A;
  wire [0:0] CLBLM_L_X8Y128_SLICE_X11Y128_A1;
  wire [0:0] CLBLM_L_X8Y128_SLICE_X11Y128_A2;
  wire [0:0] CLBLM_L_X8Y128_SLICE_X11Y128_A3;
  wire [0:0] CLBLM_L_X8Y128_SLICE_X11Y128_A4;
  wire [0:0] CLBLM_L_X8Y128_SLICE_X11Y128_A5;
  wire [0:0] CLBLM_L_X8Y128_SLICE_X11Y128_A6;
  wire [0:0] CLBLM_L_X8Y128_SLICE_X11Y128_AO5;
  wire [0:0] CLBLM_L_X8Y128_SLICE_X11Y128_AO6;
  wire [0:0] CLBLM_L_X8Y128_SLICE_X11Y128_A_CY;
  wire [0:0] CLBLM_L_X8Y128_SLICE_X11Y128_A_XOR;
  wire [0:0] CLBLM_L_X8Y128_SLICE_X11Y128_B;
  wire [0:0] CLBLM_L_X8Y128_SLICE_X11Y128_B1;
  wire [0:0] CLBLM_L_X8Y128_SLICE_X11Y128_B2;
  wire [0:0] CLBLM_L_X8Y128_SLICE_X11Y128_B3;
  wire [0:0] CLBLM_L_X8Y128_SLICE_X11Y128_B4;
  wire [0:0] CLBLM_L_X8Y128_SLICE_X11Y128_B5;
  wire [0:0] CLBLM_L_X8Y128_SLICE_X11Y128_B6;
  wire [0:0] CLBLM_L_X8Y128_SLICE_X11Y128_BO5;
  wire [0:0] CLBLM_L_X8Y128_SLICE_X11Y128_BO6;
  wire [0:0] CLBLM_L_X8Y128_SLICE_X11Y128_B_CY;
  wire [0:0] CLBLM_L_X8Y128_SLICE_X11Y128_B_XOR;
  wire [0:0] CLBLM_L_X8Y128_SLICE_X11Y128_C;
  wire [0:0] CLBLM_L_X8Y128_SLICE_X11Y128_C1;
  wire [0:0] CLBLM_L_X8Y128_SLICE_X11Y128_C2;
  wire [0:0] CLBLM_L_X8Y128_SLICE_X11Y128_C3;
  wire [0:0] CLBLM_L_X8Y128_SLICE_X11Y128_C4;
  wire [0:0] CLBLM_L_X8Y128_SLICE_X11Y128_C5;
  wire [0:0] CLBLM_L_X8Y128_SLICE_X11Y128_C6;
  wire [0:0] CLBLM_L_X8Y128_SLICE_X11Y128_CO5;
  wire [0:0] CLBLM_L_X8Y128_SLICE_X11Y128_CO6;
  wire [0:0] CLBLM_L_X8Y128_SLICE_X11Y128_C_CY;
  wire [0:0] CLBLM_L_X8Y128_SLICE_X11Y128_C_XOR;
  wire [0:0] CLBLM_L_X8Y128_SLICE_X11Y128_D;
  wire [0:0] CLBLM_L_X8Y128_SLICE_X11Y128_D1;
  wire [0:0] CLBLM_L_X8Y128_SLICE_X11Y128_D2;
  wire [0:0] CLBLM_L_X8Y128_SLICE_X11Y128_D3;
  wire [0:0] CLBLM_L_X8Y128_SLICE_X11Y128_D4;
  wire [0:0] CLBLM_L_X8Y128_SLICE_X11Y128_D5;
  wire [0:0] CLBLM_L_X8Y128_SLICE_X11Y128_D6;
  wire [0:0] CLBLM_L_X8Y128_SLICE_X11Y128_DO5;
  wire [0:0] CLBLM_L_X8Y128_SLICE_X11Y128_DO6;
  wire [0:0] CLBLM_L_X8Y128_SLICE_X11Y128_D_CY;
  wire [0:0] CLBLM_L_X8Y128_SLICE_X11Y128_D_XOR;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X10Y133_A;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X10Y133_A1;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X10Y133_A2;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X10Y133_A3;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X10Y133_A4;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X10Y133_A5;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X10Y133_A6;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X10Y133_AO5;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X10Y133_AO6;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X10Y133_A_CY;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X10Y133_A_XOR;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X10Y133_B;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X10Y133_B1;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X10Y133_B2;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X10Y133_B3;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X10Y133_B4;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X10Y133_B5;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X10Y133_B6;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X10Y133_BO5;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X10Y133_BO6;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X10Y133_B_CY;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X10Y133_B_XOR;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X10Y133_C;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X10Y133_C1;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X10Y133_C2;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X10Y133_C3;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X10Y133_C4;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X10Y133_C5;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X10Y133_C6;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X10Y133_CO5;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X10Y133_CO6;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X10Y133_C_CY;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X10Y133_C_XOR;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X10Y133_D;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X10Y133_D1;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X10Y133_D2;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X10Y133_D3;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X10Y133_D4;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X10Y133_D5;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X10Y133_D6;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X10Y133_DO5;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X10Y133_DO6;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X10Y133_D_CY;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X10Y133_D_XOR;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X11Y133_A;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X11Y133_A1;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X11Y133_A2;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X11Y133_A3;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X11Y133_A4;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X11Y133_A5;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X11Y133_A6;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X11Y133_AMUX;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X11Y133_AO5;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X11Y133_AO6;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X11Y133_A_CY;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X11Y133_A_XOR;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X11Y133_B;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X11Y133_B1;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X11Y133_B2;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X11Y133_B3;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X11Y133_B4;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X11Y133_B5;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X11Y133_B6;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X11Y133_BO5;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X11Y133_BO6;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X11Y133_B_CY;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X11Y133_B_XOR;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X11Y133_C;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X11Y133_C1;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X11Y133_C2;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X11Y133_C3;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X11Y133_C4;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X11Y133_C5;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X11Y133_C6;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X11Y133_CO5;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X11Y133_CO6;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X11Y133_C_CY;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X11Y133_C_XOR;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X11Y133_D;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X11Y133_D1;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X11Y133_D2;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X11Y133_D3;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X11Y133_D4;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X11Y133_D5;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X11Y133_D6;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X11Y133_DO5;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X11Y133_DO6;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X11Y133_D_CY;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X11Y133_D_XOR;
  wire [0:0] CLBLM_R_X103Y138_SLICE_X162Y138_A;
  wire [0:0] CLBLM_R_X103Y138_SLICE_X162Y138_A1;
  wire [0:0] CLBLM_R_X103Y138_SLICE_X162Y138_A2;
  wire [0:0] CLBLM_R_X103Y138_SLICE_X162Y138_A3;
  wire [0:0] CLBLM_R_X103Y138_SLICE_X162Y138_A4;
  wire [0:0] CLBLM_R_X103Y138_SLICE_X162Y138_A5;
  wire [0:0] CLBLM_R_X103Y138_SLICE_X162Y138_A6;
  wire [0:0] CLBLM_R_X103Y138_SLICE_X162Y138_AO5;
  wire [0:0] CLBLM_R_X103Y138_SLICE_X162Y138_AO6;
  wire [0:0] CLBLM_R_X103Y138_SLICE_X162Y138_A_CY;
  wire [0:0] CLBLM_R_X103Y138_SLICE_X162Y138_A_XOR;
  wire [0:0] CLBLM_R_X103Y138_SLICE_X162Y138_B;
  wire [0:0] CLBLM_R_X103Y138_SLICE_X162Y138_B1;
  wire [0:0] CLBLM_R_X103Y138_SLICE_X162Y138_B2;
  wire [0:0] CLBLM_R_X103Y138_SLICE_X162Y138_B3;
  wire [0:0] CLBLM_R_X103Y138_SLICE_X162Y138_B4;
  wire [0:0] CLBLM_R_X103Y138_SLICE_X162Y138_B5;
  wire [0:0] CLBLM_R_X103Y138_SLICE_X162Y138_B6;
  wire [0:0] CLBLM_R_X103Y138_SLICE_X162Y138_BO5;
  wire [0:0] CLBLM_R_X103Y138_SLICE_X162Y138_BO6;
  wire [0:0] CLBLM_R_X103Y138_SLICE_X162Y138_B_CY;
  wire [0:0] CLBLM_R_X103Y138_SLICE_X162Y138_B_XOR;
  wire [0:0] CLBLM_R_X103Y138_SLICE_X162Y138_C;
  wire [0:0] CLBLM_R_X103Y138_SLICE_X162Y138_C1;
  wire [0:0] CLBLM_R_X103Y138_SLICE_X162Y138_C2;
  wire [0:0] CLBLM_R_X103Y138_SLICE_X162Y138_C3;
  wire [0:0] CLBLM_R_X103Y138_SLICE_X162Y138_C4;
  wire [0:0] CLBLM_R_X103Y138_SLICE_X162Y138_C5;
  wire [0:0] CLBLM_R_X103Y138_SLICE_X162Y138_C6;
  wire [0:0] CLBLM_R_X103Y138_SLICE_X162Y138_CO5;
  wire [0:0] CLBLM_R_X103Y138_SLICE_X162Y138_CO6;
  wire [0:0] CLBLM_R_X103Y138_SLICE_X162Y138_C_CY;
  wire [0:0] CLBLM_R_X103Y138_SLICE_X162Y138_C_XOR;
  wire [0:0] CLBLM_R_X103Y138_SLICE_X162Y138_D;
  wire [0:0] CLBLM_R_X103Y138_SLICE_X162Y138_D1;
  wire [0:0] CLBLM_R_X103Y138_SLICE_X162Y138_D2;
  wire [0:0] CLBLM_R_X103Y138_SLICE_X162Y138_D3;
  wire [0:0] CLBLM_R_X103Y138_SLICE_X162Y138_D4;
  wire [0:0] CLBLM_R_X103Y138_SLICE_X162Y138_D5;
  wire [0:0] CLBLM_R_X103Y138_SLICE_X162Y138_D6;
  wire [0:0] CLBLM_R_X103Y138_SLICE_X162Y138_DO5;
  wire [0:0] CLBLM_R_X103Y138_SLICE_X162Y138_DO6;
  wire [0:0] CLBLM_R_X103Y138_SLICE_X162Y138_D_CY;
  wire [0:0] CLBLM_R_X103Y138_SLICE_X162Y138_D_XOR;
  wire [0:0] CLBLM_R_X103Y138_SLICE_X163Y138_A;
  wire [0:0] CLBLM_R_X103Y138_SLICE_X163Y138_A1;
  wire [0:0] CLBLM_R_X103Y138_SLICE_X163Y138_A2;
  wire [0:0] CLBLM_R_X103Y138_SLICE_X163Y138_A3;
  wire [0:0] CLBLM_R_X103Y138_SLICE_X163Y138_A4;
  wire [0:0] CLBLM_R_X103Y138_SLICE_X163Y138_A5;
  wire [0:0] CLBLM_R_X103Y138_SLICE_X163Y138_A6;
  wire [0:0] CLBLM_R_X103Y138_SLICE_X163Y138_AO5;
  wire [0:0] CLBLM_R_X103Y138_SLICE_X163Y138_AO6;
  wire [0:0] CLBLM_R_X103Y138_SLICE_X163Y138_A_CY;
  wire [0:0] CLBLM_R_X103Y138_SLICE_X163Y138_A_XOR;
  wire [0:0] CLBLM_R_X103Y138_SLICE_X163Y138_B;
  wire [0:0] CLBLM_R_X103Y138_SLICE_X163Y138_B1;
  wire [0:0] CLBLM_R_X103Y138_SLICE_X163Y138_B2;
  wire [0:0] CLBLM_R_X103Y138_SLICE_X163Y138_B3;
  wire [0:0] CLBLM_R_X103Y138_SLICE_X163Y138_B4;
  wire [0:0] CLBLM_R_X103Y138_SLICE_X163Y138_B5;
  wire [0:0] CLBLM_R_X103Y138_SLICE_X163Y138_B6;
  wire [0:0] CLBLM_R_X103Y138_SLICE_X163Y138_BO5;
  wire [0:0] CLBLM_R_X103Y138_SLICE_X163Y138_BO6;
  wire [0:0] CLBLM_R_X103Y138_SLICE_X163Y138_B_CY;
  wire [0:0] CLBLM_R_X103Y138_SLICE_X163Y138_B_XOR;
  wire [0:0] CLBLM_R_X103Y138_SLICE_X163Y138_C;
  wire [0:0] CLBLM_R_X103Y138_SLICE_X163Y138_C1;
  wire [0:0] CLBLM_R_X103Y138_SLICE_X163Y138_C2;
  wire [0:0] CLBLM_R_X103Y138_SLICE_X163Y138_C3;
  wire [0:0] CLBLM_R_X103Y138_SLICE_X163Y138_C4;
  wire [0:0] CLBLM_R_X103Y138_SLICE_X163Y138_C5;
  wire [0:0] CLBLM_R_X103Y138_SLICE_X163Y138_C6;
  wire [0:0] CLBLM_R_X103Y138_SLICE_X163Y138_CO5;
  wire [0:0] CLBLM_R_X103Y138_SLICE_X163Y138_CO6;
  wire [0:0] CLBLM_R_X103Y138_SLICE_X163Y138_C_CY;
  wire [0:0] CLBLM_R_X103Y138_SLICE_X163Y138_C_XOR;
  wire [0:0] CLBLM_R_X103Y138_SLICE_X163Y138_D;
  wire [0:0] CLBLM_R_X103Y138_SLICE_X163Y138_D1;
  wire [0:0] CLBLM_R_X103Y138_SLICE_X163Y138_D2;
  wire [0:0] CLBLM_R_X103Y138_SLICE_X163Y138_D3;
  wire [0:0] CLBLM_R_X103Y138_SLICE_X163Y138_D4;
  wire [0:0] CLBLM_R_X103Y138_SLICE_X163Y138_D5;
  wire [0:0] CLBLM_R_X103Y138_SLICE_X163Y138_D6;
  wire [0:0] CLBLM_R_X103Y138_SLICE_X163Y138_DO5;
  wire [0:0] CLBLM_R_X103Y138_SLICE_X163Y138_DO6;
  wire [0:0] CLBLM_R_X103Y138_SLICE_X163Y138_D_CY;
  wire [0:0] CLBLM_R_X103Y138_SLICE_X163Y138_D_XOR;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X162Y169_A;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X162Y169_A1;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X162Y169_A2;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X162Y169_A3;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X162Y169_A4;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X162Y169_A5;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X162Y169_A6;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X162Y169_AO5;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X162Y169_AO6;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X162Y169_A_CY;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X162Y169_A_XOR;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X162Y169_B;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X162Y169_B1;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X162Y169_B2;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X162Y169_B3;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X162Y169_B4;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X162Y169_B5;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X162Y169_B6;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X162Y169_BO5;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X162Y169_BO6;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X162Y169_B_CY;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X162Y169_B_XOR;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X162Y169_C;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X162Y169_C1;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X162Y169_C2;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X162Y169_C3;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X162Y169_C4;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X162Y169_C5;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X162Y169_C6;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X162Y169_CO5;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X162Y169_CO6;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X162Y169_C_CY;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X162Y169_C_XOR;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X162Y169_D;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X162Y169_D1;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X162Y169_D2;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X162Y169_D3;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X162Y169_D4;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X162Y169_D5;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X162Y169_D6;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X162Y169_DO5;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X162Y169_DO6;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X162Y169_D_CY;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X162Y169_D_XOR;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X163Y169_A;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X163Y169_A1;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X163Y169_A2;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X163Y169_A3;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X163Y169_A4;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X163Y169_A5;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X163Y169_A6;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X163Y169_AMUX;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X163Y169_AO5;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X163Y169_AO6;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X163Y169_A_CY;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X163Y169_A_XOR;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X163Y169_B;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X163Y169_B1;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X163Y169_B2;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X163Y169_B3;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X163Y169_B4;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X163Y169_B5;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X163Y169_B6;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X163Y169_BO5;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X163Y169_BO6;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X163Y169_B_CY;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X163Y169_B_XOR;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X163Y169_C;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X163Y169_C1;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X163Y169_C2;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X163Y169_C3;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X163Y169_C4;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X163Y169_C5;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X163Y169_C6;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X163Y169_CO5;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X163Y169_CO6;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X163Y169_C_CY;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X163Y169_C_XOR;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X163Y169_D;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X163Y169_D1;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X163Y169_D2;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X163Y169_D3;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X163Y169_D4;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X163Y169_D5;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X163Y169_D6;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X163Y169_DO5;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X163Y169_DO6;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X163Y169_D_CY;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X163Y169_D_XOR;
  wire [0:0] CLBLM_R_X103Y172_SLICE_X162Y172_A;
  wire [0:0] CLBLM_R_X103Y172_SLICE_X162Y172_A1;
  wire [0:0] CLBLM_R_X103Y172_SLICE_X162Y172_A2;
  wire [0:0] CLBLM_R_X103Y172_SLICE_X162Y172_A3;
  wire [0:0] CLBLM_R_X103Y172_SLICE_X162Y172_A4;
  wire [0:0] CLBLM_R_X103Y172_SLICE_X162Y172_A5;
  wire [0:0] CLBLM_R_X103Y172_SLICE_X162Y172_A6;
  wire [0:0] CLBLM_R_X103Y172_SLICE_X162Y172_AO5;
  wire [0:0] CLBLM_R_X103Y172_SLICE_X162Y172_AO6;
  wire [0:0] CLBLM_R_X103Y172_SLICE_X162Y172_A_CY;
  wire [0:0] CLBLM_R_X103Y172_SLICE_X162Y172_A_XOR;
  wire [0:0] CLBLM_R_X103Y172_SLICE_X162Y172_B;
  wire [0:0] CLBLM_R_X103Y172_SLICE_X162Y172_B1;
  wire [0:0] CLBLM_R_X103Y172_SLICE_X162Y172_B2;
  wire [0:0] CLBLM_R_X103Y172_SLICE_X162Y172_B3;
  wire [0:0] CLBLM_R_X103Y172_SLICE_X162Y172_B4;
  wire [0:0] CLBLM_R_X103Y172_SLICE_X162Y172_B5;
  wire [0:0] CLBLM_R_X103Y172_SLICE_X162Y172_B6;
  wire [0:0] CLBLM_R_X103Y172_SLICE_X162Y172_BO5;
  wire [0:0] CLBLM_R_X103Y172_SLICE_X162Y172_BO6;
  wire [0:0] CLBLM_R_X103Y172_SLICE_X162Y172_B_CY;
  wire [0:0] CLBLM_R_X103Y172_SLICE_X162Y172_B_XOR;
  wire [0:0] CLBLM_R_X103Y172_SLICE_X162Y172_C;
  wire [0:0] CLBLM_R_X103Y172_SLICE_X162Y172_C1;
  wire [0:0] CLBLM_R_X103Y172_SLICE_X162Y172_C2;
  wire [0:0] CLBLM_R_X103Y172_SLICE_X162Y172_C3;
  wire [0:0] CLBLM_R_X103Y172_SLICE_X162Y172_C4;
  wire [0:0] CLBLM_R_X103Y172_SLICE_X162Y172_C5;
  wire [0:0] CLBLM_R_X103Y172_SLICE_X162Y172_C6;
  wire [0:0] CLBLM_R_X103Y172_SLICE_X162Y172_CO5;
  wire [0:0] CLBLM_R_X103Y172_SLICE_X162Y172_CO6;
  wire [0:0] CLBLM_R_X103Y172_SLICE_X162Y172_C_CY;
  wire [0:0] CLBLM_R_X103Y172_SLICE_X162Y172_C_XOR;
  wire [0:0] CLBLM_R_X103Y172_SLICE_X162Y172_D;
  wire [0:0] CLBLM_R_X103Y172_SLICE_X162Y172_D1;
  wire [0:0] CLBLM_R_X103Y172_SLICE_X162Y172_D2;
  wire [0:0] CLBLM_R_X103Y172_SLICE_X162Y172_D3;
  wire [0:0] CLBLM_R_X103Y172_SLICE_X162Y172_D4;
  wire [0:0] CLBLM_R_X103Y172_SLICE_X162Y172_D5;
  wire [0:0] CLBLM_R_X103Y172_SLICE_X162Y172_D6;
  wire [0:0] CLBLM_R_X103Y172_SLICE_X162Y172_DO5;
  wire [0:0] CLBLM_R_X103Y172_SLICE_X162Y172_DO6;
  wire [0:0] CLBLM_R_X103Y172_SLICE_X162Y172_D_CY;
  wire [0:0] CLBLM_R_X103Y172_SLICE_X162Y172_D_XOR;
  wire [0:0] CLBLM_R_X103Y172_SLICE_X163Y172_A;
  wire [0:0] CLBLM_R_X103Y172_SLICE_X163Y172_A1;
  wire [0:0] CLBLM_R_X103Y172_SLICE_X163Y172_A2;
  wire [0:0] CLBLM_R_X103Y172_SLICE_X163Y172_A3;
  wire [0:0] CLBLM_R_X103Y172_SLICE_X163Y172_A4;
  wire [0:0] CLBLM_R_X103Y172_SLICE_X163Y172_A5;
  wire [0:0] CLBLM_R_X103Y172_SLICE_X163Y172_A6;
  wire [0:0] CLBLM_R_X103Y172_SLICE_X163Y172_AMUX;
  wire [0:0] CLBLM_R_X103Y172_SLICE_X163Y172_AO5;
  wire [0:0] CLBLM_R_X103Y172_SLICE_X163Y172_AO6;
  wire [0:0] CLBLM_R_X103Y172_SLICE_X163Y172_A_CY;
  wire [0:0] CLBLM_R_X103Y172_SLICE_X163Y172_A_XOR;
  wire [0:0] CLBLM_R_X103Y172_SLICE_X163Y172_B;
  wire [0:0] CLBLM_R_X103Y172_SLICE_X163Y172_B1;
  wire [0:0] CLBLM_R_X103Y172_SLICE_X163Y172_B2;
  wire [0:0] CLBLM_R_X103Y172_SLICE_X163Y172_B3;
  wire [0:0] CLBLM_R_X103Y172_SLICE_X163Y172_B4;
  wire [0:0] CLBLM_R_X103Y172_SLICE_X163Y172_B5;
  wire [0:0] CLBLM_R_X103Y172_SLICE_X163Y172_B6;
  wire [0:0] CLBLM_R_X103Y172_SLICE_X163Y172_BO5;
  wire [0:0] CLBLM_R_X103Y172_SLICE_X163Y172_BO6;
  wire [0:0] CLBLM_R_X103Y172_SLICE_X163Y172_B_CY;
  wire [0:0] CLBLM_R_X103Y172_SLICE_X163Y172_B_XOR;
  wire [0:0] CLBLM_R_X103Y172_SLICE_X163Y172_C;
  wire [0:0] CLBLM_R_X103Y172_SLICE_X163Y172_C1;
  wire [0:0] CLBLM_R_X103Y172_SLICE_X163Y172_C2;
  wire [0:0] CLBLM_R_X103Y172_SLICE_X163Y172_C3;
  wire [0:0] CLBLM_R_X103Y172_SLICE_X163Y172_C4;
  wire [0:0] CLBLM_R_X103Y172_SLICE_X163Y172_C5;
  wire [0:0] CLBLM_R_X103Y172_SLICE_X163Y172_C6;
  wire [0:0] CLBLM_R_X103Y172_SLICE_X163Y172_CO5;
  wire [0:0] CLBLM_R_X103Y172_SLICE_X163Y172_CO6;
  wire [0:0] CLBLM_R_X103Y172_SLICE_X163Y172_C_CY;
  wire [0:0] CLBLM_R_X103Y172_SLICE_X163Y172_C_XOR;
  wire [0:0] CLBLM_R_X103Y172_SLICE_X163Y172_D;
  wire [0:0] CLBLM_R_X103Y172_SLICE_X163Y172_D1;
  wire [0:0] CLBLM_R_X103Y172_SLICE_X163Y172_D2;
  wire [0:0] CLBLM_R_X103Y172_SLICE_X163Y172_D3;
  wire [0:0] CLBLM_R_X103Y172_SLICE_X163Y172_D4;
  wire [0:0] CLBLM_R_X103Y172_SLICE_X163Y172_D5;
  wire [0:0] CLBLM_R_X103Y172_SLICE_X163Y172_D6;
  wire [0:0] CLBLM_R_X103Y172_SLICE_X163Y172_DO5;
  wire [0:0] CLBLM_R_X103Y172_SLICE_X163Y172_DO6;
  wire [0:0] CLBLM_R_X103Y172_SLICE_X163Y172_D_CY;
  wire [0:0] CLBLM_R_X103Y172_SLICE_X163Y172_D_XOR;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X162Y174_A;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X162Y174_A1;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X162Y174_A2;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X162Y174_A3;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X162Y174_A4;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X162Y174_A5;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X162Y174_A6;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X162Y174_AO5;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X162Y174_AO6;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X162Y174_A_CY;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X162Y174_A_XOR;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X162Y174_B;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X162Y174_B1;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X162Y174_B2;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X162Y174_B3;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X162Y174_B4;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X162Y174_B5;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X162Y174_B6;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X162Y174_BO5;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X162Y174_BO6;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X162Y174_B_CY;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X162Y174_B_XOR;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X162Y174_C;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X162Y174_C1;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X162Y174_C2;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X162Y174_C3;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X162Y174_C4;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X162Y174_C5;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X162Y174_C6;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X162Y174_CO5;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X162Y174_CO6;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X162Y174_C_CY;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X162Y174_C_XOR;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X162Y174_D;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X162Y174_D1;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X162Y174_D2;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X162Y174_D3;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X162Y174_D4;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X162Y174_D5;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X162Y174_D6;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X162Y174_DO5;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X162Y174_DO6;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X162Y174_D_CY;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X162Y174_D_XOR;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X163Y174_A;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X163Y174_A1;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X163Y174_A2;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X163Y174_A3;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X163Y174_A4;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X163Y174_A5;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X163Y174_A6;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X163Y174_AMUX;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X163Y174_AO5;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X163Y174_AO6;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X163Y174_A_CY;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X163Y174_A_XOR;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X163Y174_B;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X163Y174_B1;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X163Y174_B2;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X163Y174_B3;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X163Y174_B4;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X163Y174_B5;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X163Y174_B6;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X163Y174_BO5;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X163Y174_BO6;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X163Y174_B_CY;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X163Y174_B_XOR;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X163Y174_C;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X163Y174_C1;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X163Y174_C2;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X163Y174_C3;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X163Y174_C4;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X163Y174_C5;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X163Y174_C6;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X163Y174_CO5;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X163Y174_CO6;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X163Y174_C_CY;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X163Y174_C_XOR;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X163Y174_D;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X163Y174_D1;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X163Y174_D2;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X163Y174_D3;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X163Y174_D4;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X163Y174_D5;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X163Y174_D6;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X163Y174_DO5;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X163Y174_DO6;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X163Y174_D_CY;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X163Y174_D_XOR;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X162Y177_A;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X162Y177_A1;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X162Y177_A2;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X162Y177_A3;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X162Y177_A4;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X162Y177_A5;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X162Y177_A6;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X162Y177_AO5;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X162Y177_AO6;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X162Y177_A_CY;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X162Y177_A_XOR;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X162Y177_B;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X162Y177_B1;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X162Y177_B2;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X162Y177_B3;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X162Y177_B4;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X162Y177_B5;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X162Y177_B6;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X162Y177_BO5;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X162Y177_BO6;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X162Y177_B_CY;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X162Y177_B_XOR;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X162Y177_C;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X162Y177_C1;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X162Y177_C2;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X162Y177_C3;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X162Y177_C4;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X162Y177_C5;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X162Y177_C6;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X162Y177_CO5;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X162Y177_CO6;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X162Y177_C_CY;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X162Y177_C_XOR;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X162Y177_D;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X162Y177_D1;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X162Y177_D2;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X162Y177_D3;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X162Y177_D4;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X162Y177_D5;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X162Y177_D6;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X162Y177_DO5;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X162Y177_DO6;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X162Y177_D_CY;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X162Y177_D_XOR;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X163Y177_A;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X163Y177_A1;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X163Y177_A2;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X163Y177_A3;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X163Y177_A4;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X163Y177_A5;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X163Y177_A6;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X163Y177_AMUX;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X163Y177_AO5;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X163Y177_AO6;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X163Y177_A_CY;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X163Y177_A_XOR;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X163Y177_B;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X163Y177_B1;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X163Y177_B2;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X163Y177_B3;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X163Y177_B4;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X163Y177_B5;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X163Y177_B6;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X163Y177_BO5;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X163Y177_BO6;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X163Y177_B_CY;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X163Y177_B_XOR;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X163Y177_C;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X163Y177_C1;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X163Y177_C2;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X163Y177_C3;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X163Y177_C4;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X163Y177_C5;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X163Y177_C6;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X163Y177_CO5;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X163Y177_CO6;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X163Y177_C_CY;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X163Y177_C_XOR;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X163Y177_D;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X163Y177_D1;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X163Y177_D2;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X163Y177_D3;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X163Y177_D4;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X163Y177_D5;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X163Y177_D6;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X163Y177_DO5;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X163Y177_DO6;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X163Y177_D_CY;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X163Y177_D_XOR;
  wire [0:0] CLBLM_R_X11Y113_SLICE_X14Y113_A;
  wire [0:0] CLBLM_R_X11Y113_SLICE_X14Y113_A1;
  wire [0:0] CLBLM_R_X11Y113_SLICE_X14Y113_A2;
  wire [0:0] CLBLM_R_X11Y113_SLICE_X14Y113_A3;
  wire [0:0] CLBLM_R_X11Y113_SLICE_X14Y113_A4;
  wire [0:0] CLBLM_R_X11Y113_SLICE_X14Y113_A5;
  wire [0:0] CLBLM_R_X11Y113_SLICE_X14Y113_A6;
  wire [0:0] CLBLM_R_X11Y113_SLICE_X14Y113_AO5;
  wire [0:0] CLBLM_R_X11Y113_SLICE_X14Y113_AO6;
  wire [0:0] CLBLM_R_X11Y113_SLICE_X14Y113_AQ;
  wire [0:0] CLBLM_R_X11Y113_SLICE_X14Y113_A_CY;
  wire [0:0] CLBLM_R_X11Y113_SLICE_X14Y113_A_XOR;
  wire [0:0] CLBLM_R_X11Y113_SLICE_X14Y113_B;
  wire [0:0] CLBLM_R_X11Y113_SLICE_X14Y113_B1;
  wire [0:0] CLBLM_R_X11Y113_SLICE_X14Y113_B2;
  wire [0:0] CLBLM_R_X11Y113_SLICE_X14Y113_B3;
  wire [0:0] CLBLM_R_X11Y113_SLICE_X14Y113_B4;
  wire [0:0] CLBLM_R_X11Y113_SLICE_X14Y113_B5;
  wire [0:0] CLBLM_R_X11Y113_SLICE_X14Y113_B6;
  wire [0:0] CLBLM_R_X11Y113_SLICE_X14Y113_BO5;
  wire [0:0] CLBLM_R_X11Y113_SLICE_X14Y113_BO6;
  wire [0:0] CLBLM_R_X11Y113_SLICE_X14Y113_BQ;
  wire [0:0] CLBLM_R_X11Y113_SLICE_X14Y113_B_CY;
  wire [0:0] CLBLM_R_X11Y113_SLICE_X14Y113_B_XOR;
  wire [0:0] CLBLM_R_X11Y113_SLICE_X14Y113_C;
  wire [0:0] CLBLM_R_X11Y113_SLICE_X14Y113_C1;
  wire [0:0] CLBLM_R_X11Y113_SLICE_X14Y113_C2;
  wire [0:0] CLBLM_R_X11Y113_SLICE_X14Y113_C3;
  wire [0:0] CLBLM_R_X11Y113_SLICE_X14Y113_C4;
  wire [0:0] CLBLM_R_X11Y113_SLICE_X14Y113_C5;
  wire [0:0] CLBLM_R_X11Y113_SLICE_X14Y113_C6;
  wire [0:0] CLBLM_R_X11Y113_SLICE_X14Y113_CLK;
  wire [0:0] CLBLM_R_X11Y113_SLICE_X14Y113_CO5;
  wire [0:0] CLBLM_R_X11Y113_SLICE_X14Y113_CO6;
  wire [0:0] CLBLM_R_X11Y113_SLICE_X14Y113_C_CY;
  wire [0:0] CLBLM_R_X11Y113_SLICE_X14Y113_C_XOR;
  wire [0:0] CLBLM_R_X11Y113_SLICE_X14Y113_D;
  wire [0:0] CLBLM_R_X11Y113_SLICE_X14Y113_D1;
  wire [0:0] CLBLM_R_X11Y113_SLICE_X14Y113_D2;
  wire [0:0] CLBLM_R_X11Y113_SLICE_X14Y113_D3;
  wire [0:0] CLBLM_R_X11Y113_SLICE_X14Y113_D4;
  wire [0:0] CLBLM_R_X11Y113_SLICE_X14Y113_D5;
  wire [0:0] CLBLM_R_X11Y113_SLICE_X14Y113_D6;
  wire [0:0] CLBLM_R_X11Y113_SLICE_X14Y113_DO5;
  wire [0:0] CLBLM_R_X11Y113_SLICE_X14Y113_DO6;
  wire [0:0] CLBLM_R_X11Y113_SLICE_X14Y113_D_CY;
  wire [0:0] CLBLM_R_X11Y113_SLICE_X14Y113_D_XOR;
  wire [0:0] CLBLM_R_X11Y113_SLICE_X15Y113_A;
  wire [0:0] CLBLM_R_X11Y113_SLICE_X15Y113_A1;
  wire [0:0] CLBLM_R_X11Y113_SLICE_X15Y113_A2;
  wire [0:0] CLBLM_R_X11Y113_SLICE_X15Y113_A3;
  wire [0:0] CLBLM_R_X11Y113_SLICE_X15Y113_A4;
  wire [0:0] CLBLM_R_X11Y113_SLICE_X15Y113_A5;
  wire [0:0] CLBLM_R_X11Y113_SLICE_X15Y113_A6;
  wire [0:0] CLBLM_R_X11Y113_SLICE_X15Y113_AO5;
  wire [0:0] CLBLM_R_X11Y113_SLICE_X15Y113_AO6;
  wire [0:0] CLBLM_R_X11Y113_SLICE_X15Y113_AQ;
  wire [0:0] CLBLM_R_X11Y113_SLICE_X15Y113_A_CY;
  wire [0:0] CLBLM_R_X11Y113_SLICE_X15Y113_A_XOR;
  wire [0:0] CLBLM_R_X11Y113_SLICE_X15Y113_B;
  wire [0:0] CLBLM_R_X11Y113_SLICE_X15Y113_B1;
  wire [0:0] CLBLM_R_X11Y113_SLICE_X15Y113_B2;
  wire [0:0] CLBLM_R_X11Y113_SLICE_X15Y113_B3;
  wire [0:0] CLBLM_R_X11Y113_SLICE_X15Y113_B4;
  wire [0:0] CLBLM_R_X11Y113_SLICE_X15Y113_B5;
  wire [0:0] CLBLM_R_X11Y113_SLICE_X15Y113_B6;
  wire [0:0] CLBLM_R_X11Y113_SLICE_X15Y113_BO5;
  wire [0:0] CLBLM_R_X11Y113_SLICE_X15Y113_BO6;
  wire [0:0] CLBLM_R_X11Y113_SLICE_X15Y113_BQ;
  wire [0:0] CLBLM_R_X11Y113_SLICE_X15Y113_B_CY;
  wire [0:0] CLBLM_R_X11Y113_SLICE_X15Y113_B_XOR;
  wire [0:0] CLBLM_R_X11Y113_SLICE_X15Y113_C;
  wire [0:0] CLBLM_R_X11Y113_SLICE_X15Y113_C1;
  wire [0:0] CLBLM_R_X11Y113_SLICE_X15Y113_C2;
  wire [0:0] CLBLM_R_X11Y113_SLICE_X15Y113_C3;
  wire [0:0] CLBLM_R_X11Y113_SLICE_X15Y113_C4;
  wire [0:0] CLBLM_R_X11Y113_SLICE_X15Y113_C5;
  wire [0:0] CLBLM_R_X11Y113_SLICE_X15Y113_C6;
  wire [0:0] CLBLM_R_X11Y113_SLICE_X15Y113_CLK;
  wire [0:0] CLBLM_R_X11Y113_SLICE_X15Y113_CO5;
  wire [0:0] CLBLM_R_X11Y113_SLICE_X15Y113_CO6;
  wire [0:0] CLBLM_R_X11Y113_SLICE_X15Y113_C_CY;
  wire [0:0] CLBLM_R_X11Y113_SLICE_X15Y113_C_XOR;
  wire [0:0] CLBLM_R_X11Y113_SLICE_X15Y113_D;
  wire [0:0] CLBLM_R_X11Y113_SLICE_X15Y113_D1;
  wire [0:0] CLBLM_R_X11Y113_SLICE_X15Y113_D2;
  wire [0:0] CLBLM_R_X11Y113_SLICE_X15Y113_D3;
  wire [0:0] CLBLM_R_X11Y113_SLICE_X15Y113_D4;
  wire [0:0] CLBLM_R_X11Y113_SLICE_X15Y113_D5;
  wire [0:0] CLBLM_R_X11Y113_SLICE_X15Y113_D6;
  wire [0:0] CLBLM_R_X11Y113_SLICE_X15Y113_DO5;
  wire [0:0] CLBLM_R_X11Y113_SLICE_X15Y113_DO6;
  wire [0:0] CLBLM_R_X11Y113_SLICE_X15Y113_D_CY;
  wire [0:0] CLBLM_R_X11Y113_SLICE_X15Y113_D_XOR;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X14Y114_A;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X14Y114_A1;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X14Y114_A2;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X14Y114_A3;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X14Y114_A4;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X14Y114_A5;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X14Y114_A6;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X14Y114_AO5;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X14Y114_AO6;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X14Y114_AQ;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X14Y114_A_CY;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X14Y114_A_XOR;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X14Y114_B;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X14Y114_B1;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X14Y114_B2;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X14Y114_B3;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X14Y114_B4;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X14Y114_B5;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X14Y114_B6;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X14Y114_BO5;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X14Y114_BO6;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X14Y114_BQ;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X14Y114_B_CY;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X14Y114_B_XOR;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X14Y114_C;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X14Y114_C1;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X14Y114_C2;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X14Y114_C3;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X14Y114_C4;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X14Y114_C5;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X14Y114_C6;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X14Y114_CLK;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X14Y114_CO5;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X14Y114_CO6;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X14Y114_CQ;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X14Y114_C_CY;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X14Y114_C_XOR;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X14Y114_D;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X14Y114_D1;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X14Y114_D2;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X14Y114_D3;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X14Y114_D4;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X14Y114_D5;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X14Y114_D5Q;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X14Y114_D6;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X14Y114_DMUX;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X14Y114_DO5;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X14Y114_DO6;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X14Y114_DQ;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X14Y114_D_CY;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X14Y114_D_XOR;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X15Y114_A;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X15Y114_A1;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X15Y114_A2;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X15Y114_A3;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X15Y114_A4;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X15Y114_A5;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X15Y114_A6;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X15Y114_AO5;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X15Y114_AO6;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X15Y114_A_CY;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X15Y114_A_XOR;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X15Y114_B;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X15Y114_B1;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X15Y114_B2;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X15Y114_B3;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X15Y114_B4;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X15Y114_B5;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X15Y114_B6;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X15Y114_BO5;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X15Y114_BO6;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X15Y114_B_CY;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X15Y114_B_XOR;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X15Y114_C;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X15Y114_C1;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X15Y114_C2;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X15Y114_C3;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X15Y114_C4;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X15Y114_C5;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X15Y114_C6;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X15Y114_CO5;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X15Y114_CO6;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X15Y114_C_CY;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X15Y114_C_XOR;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X15Y114_D;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X15Y114_D1;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X15Y114_D2;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X15Y114_D3;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X15Y114_D4;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X15Y114_D5;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X15Y114_D6;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X15Y114_DO5;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X15Y114_DO6;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X15Y114_D_CY;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X15Y114_D_XOR;
  wire [0:0] CLBLM_R_X11Y115_SLICE_X14Y115_A;
  wire [0:0] CLBLM_R_X11Y115_SLICE_X14Y115_A1;
  wire [0:0] CLBLM_R_X11Y115_SLICE_X14Y115_A2;
  wire [0:0] CLBLM_R_X11Y115_SLICE_X14Y115_A3;
  wire [0:0] CLBLM_R_X11Y115_SLICE_X14Y115_A4;
  wire [0:0] CLBLM_R_X11Y115_SLICE_X14Y115_A5;
  wire [0:0] CLBLM_R_X11Y115_SLICE_X14Y115_A6;
  wire [0:0] CLBLM_R_X11Y115_SLICE_X14Y115_AO5;
  wire [0:0] CLBLM_R_X11Y115_SLICE_X14Y115_AO6;
  wire [0:0] CLBLM_R_X11Y115_SLICE_X14Y115_AQ;
  wire [0:0] CLBLM_R_X11Y115_SLICE_X14Y115_A_CY;
  wire [0:0] CLBLM_R_X11Y115_SLICE_X14Y115_A_XOR;
  wire [0:0] CLBLM_R_X11Y115_SLICE_X14Y115_B;
  wire [0:0] CLBLM_R_X11Y115_SLICE_X14Y115_B1;
  wire [0:0] CLBLM_R_X11Y115_SLICE_X14Y115_B2;
  wire [0:0] CLBLM_R_X11Y115_SLICE_X14Y115_B3;
  wire [0:0] CLBLM_R_X11Y115_SLICE_X14Y115_B4;
  wire [0:0] CLBLM_R_X11Y115_SLICE_X14Y115_B5;
  wire [0:0] CLBLM_R_X11Y115_SLICE_X14Y115_B6;
  wire [0:0] CLBLM_R_X11Y115_SLICE_X14Y115_BO5;
  wire [0:0] CLBLM_R_X11Y115_SLICE_X14Y115_BO6;
  wire [0:0] CLBLM_R_X11Y115_SLICE_X14Y115_BQ;
  wire [0:0] CLBLM_R_X11Y115_SLICE_X14Y115_B_CY;
  wire [0:0] CLBLM_R_X11Y115_SLICE_X14Y115_B_XOR;
  wire [0:0] CLBLM_R_X11Y115_SLICE_X14Y115_C;
  wire [0:0] CLBLM_R_X11Y115_SLICE_X14Y115_C1;
  wire [0:0] CLBLM_R_X11Y115_SLICE_X14Y115_C2;
  wire [0:0] CLBLM_R_X11Y115_SLICE_X14Y115_C3;
  wire [0:0] CLBLM_R_X11Y115_SLICE_X14Y115_C4;
  wire [0:0] CLBLM_R_X11Y115_SLICE_X14Y115_C5;
  wire [0:0] CLBLM_R_X11Y115_SLICE_X14Y115_C6;
  wire [0:0] CLBLM_R_X11Y115_SLICE_X14Y115_CLK;
  wire [0:0] CLBLM_R_X11Y115_SLICE_X14Y115_CO5;
  wire [0:0] CLBLM_R_X11Y115_SLICE_X14Y115_CO6;
  wire [0:0] CLBLM_R_X11Y115_SLICE_X14Y115_CQ;
  wire [0:0] CLBLM_R_X11Y115_SLICE_X14Y115_C_CY;
  wire [0:0] CLBLM_R_X11Y115_SLICE_X14Y115_C_XOR;
  wire [0:0] CLBLM_R_X11Y115_SLICE_X14Y115_D;
  wire [0:0] CLBLM_R_X11Y115_SLICE_X14Y115_D1;
  wire [0:0] CLBLM_R_X11Y115_SLICE_X14Y115_D2;
  wire [0:0] CLBLM_R_X11Y115_SLICE_X14Y115_D3;
  wire [0:0] CLBLM_R_X11Y115_SLICE_X14Y115_D4;
  wire [0:0] CLBLM_R_X11Y115_SLICE_X14Y115_D5;
  wire [0:0] CLBLM_R_X11Y115_SLICE_X14Y115_D6;
  wire [0:0] CLBLM_R_X11Y115_SLICE_X14Y115_DO5;
  wire [0:0] CLBLM_R_X11Y115_SLICE_X14Y115_DO6;
  wire [0:0] CLBLM_R_X11Y115_SLICE_X14Y115_DQ;
  wire [0:0] CLBLM_R_X11Y115_SLICE_X14Y115_D_CY;
  wire [0:0] CLBLM_R_X11Y115_SLICE_X14Y115_D_XOR;
  wire [0:0] CLBLM_R_X11Y115_SLICE_X15Y115_A;
  wire [0:0] CLBLM_R_X11Y115_SLICE_X15Y115_A1;
  wire [0:0] CLBLM_R_X11Y115_SLICE_X15Y115_A2;
  wire [0:0] CLBLM_R_X11Y115_SLICE_X15Y115_A3;
  wire [0:0] CLBLM_R_X11Y115_SLICE_X15Y115_A4;
  wire [0:0] CLBLM_R_X11Y115_SLICE_X15Y115_A5;
  wire [0:0] CLBLM_R_X11Y115_SLICE_X15Y115_A6;
  wire [0:0] CLBLM_R_X11Y115_SLICE_X15Y115_AO5;
  wire [0:0] CLBLM_R_X11Y115_SLICE_X15Y115_AO6;
  wire [0:0] CLBLM_R_X11Y115_SLICE_X15Y115_AQ;
  wire [0:0] CLBLM_R_X11Y115_SLICE_X15Y115_A_CY;
  wire [0:0] CLBLM_R_X11Y115_SLICE_X15Y115_A_XOR;
  wire [0:0] CLBLM_R_X11Y115_SLICE_X15Y115_B;
  wire [0:0] CLBLM_R_X11Y115_SLICE_X15Y115_B1;
  wire [0:0] CLBLM_R_X11Y115_SLICE_X15Y115_B2;
  wire [0:0] CLBLM_R_X11Y115_SLICE_X15Y115_B3;
  wire [0:0] CLBLM_R_X11Y115_SLICE_X15Y115_B4;
  wire [0:0] CLBLM_R_X11Y115_SLICE_X15Y115_B5;
  wire [0:0] CLBLM_R_X11Y115_SLICE_X15Y115_B6;
  wire [0:0] CLBLM_R_X11Y115_SLICE_X15Y115_BO5;
  wire [0:0] CLBLM_R_X11Y115_SLICE_X15Y115_BO6;
  wire [0:0] CLBLM_R_X11Y115_SLICE_X15Y115_BQ;
  wire [0:0] CLBLM_R_X11Y115_SLICE_X15Y115_B_CY;
  wire [0:0] CLBLM_R_X11Y115_SLICE_X15Y115_B_XOR;
  wire [0:0] CLBLM_R_X11Y115_SLICE_X15Y115_C;
  wire [0:0] CLBLM_R_X11Y115_SLICE_X15Y115_C1;
  wire [0:0] CLBLM_R_X11Y115_SLICE_X15Y115_C2;
  wire [0:0] CLBLM_R_X11Y115_SLICE_X15Y115_C3;
  wire [0:0] CLBLM_R_X11Y115_SLICE_X15Y115_C4;
  wire [0:0] CLBLM_R_X11Y115_SLICE_X15Y115_C5;
  wire [0:0] CLBLM_R_X11Y115_SLICE_X15Y115_C6;
  wire [0:0] CLBLM_R_X11Y115_SLICE_X15Y115_CLK;
  wire [0:0] CLBLM_R_X11Y115_SLICE_X15Y115_CO5;
  wire [0:0] CLBLM_R_X11Y115_SLICE_X15Y115_CO6;
  wire [0:0] CLBLM_R_X11Y115_SLICE_X15Y115_CQ;
  wire [0:0] CLBLM_R_X11Y115_SLICE_X15Y115_C_CY;
  wire [0:0] CLBLM_R_X11Y115_SLICE_X15Y115_C_XOR;
  wire [0:0] CLBLM_R_X11Y115_SLICE_X15Y115_D;
  wire [0:0] CLBLM_R_X11Y115_SLICE_X15Y115_D1;
  wire [0:0] CLBLM_R_X11Y115_SLICE_X15Y115_D2;
  wire [0:0] CLBLM_R_X11Y115_SLICE_X15Y115_D3;
  wire [0:0] CLBLM_R_X11Y115_SLICE_X15Y115_D4;
  wire [0:0] CLBLM_R_X11Y115_SLICE_X15Y115_D5;
  wire [0:0] CLBLM_R_X11Y115_SLICE_X15Y115_D6;
  wire [0:0] CLBLM_R_X11Y115_SLICE_X15Y115_DO5;
  wire [0:0] CLBLM_R_X11Y115_SLICE_X15Y115_DO6;
  wire [0:0] CLBLM_R_X11Y115_SLICE_X15Y115_DQ;
  wire [0:0] CLBLM_R_X11Y115_SLICE_X15Y115_D_CY;
  wire [0:0] CLBLM_R_X11Y115_SLICE_X15Y115_D_XOR;
  wire [0:0] CLBLM_R_X11Y116_SLICE_X14Y116_A;
  wire [0:0] CLBLM_R_X11Y116_SLICE_X14Y116_A1;
  wire [0:0] CLBLM_R_X11Y116_SLICE_X14Y116_A2;
  wire [0:0] CLBLM_R_X11Y116_SLICE_X14Y116_A3;
  wire [0:0] CLBLM_R_X11Y116_SLICE_X14Y116_A4;
  wire [0:0] CLBLM_R_X11Y116_SLICE_X14Y116_A5;
  wire [0:0] CLBLM_R_X11Y116_SLICE_X14Y116_A6;
  wire [0:0] CLBLM_R_X11Y116_SLICE_X14Y116_AO5;
  wire [0:0] CLBLM_R_X11Y116_SLICE_X14Y116_AO6;
  wire [0:0] CLBLM_R_X11Y116_SLICE_X14Y116_AQ;
  wire [0:0] CLBLM_R_X11Y116_SLICE_X14Y116_A_CY;
  wire [0:0] CLBLM_R_X11Y116_SLICE_X14Y116_A_XOR;
  wire [0:0] CLBLM_R_X11Y116_SLICE_X14Y116_B;
  wire [0:0] CLBLM_R_X11Y116_SLICE_X14Y116_B1;
  wire [0:0] CLBLM_R_X11Y116_SLICE_X14Y116_B2;
  wire [0:0] CLBLM_R_X11Y116_SLICE_X14Y116_B3;
  wire [0:0] CLBLM_R_X11Y116_SLICE_X14Y116_B4;
  wire [0:0] CLBLM_R_X11Y116_SLICE_X14Y116_B5;
  wire [0:0] CLBLM_R_X11Y116_SLICE_X14Y116_B6;
  wire [0:0] CLBLM_R_X11Y116_SLICE_X14Y116_BMUX;
  wire [0:0] CLBLM_R_X11Y116_SLICE_X14Y116_BO5;
  wire [0:0] CLBLM_R_X11Y116_SLICE_X14Y116_BO6;
  wire [0:0] CLBLM_R_X11Y116_SLICE_X14Y116_B_CY;
  wire [0:0] CLBLM_R_X11Y116_SLICE_X14Y116_B_XOR;
  wire [0:0] CLBLM_R_X11Y116_SLICE_X14Y116_C;
  wire [0:0] CLBLM_R_X11Y116_SLICE_X14Y116_C1;
  wire [0:0] CLBLM_R_X11Y116_SLICE_X14Y116_C2;
  wire [0:0] CLBLM_R_X11Y116_SLICE_X14Y116_C3;
  wire [0:0] CLBLM_R_X11Y116_SLICE_X14Y116_C4;
  wire [0:0] CLBLM_R_X11Y116_SLICE_X14Y116_C5;
  wire [0:0] CLBLM_R_X11Y116_SLICE_X14Y116_C6;
  wire [0:0] CLBLM_R_X11Y116_SLICE_X14Y116_CLK;
  wire [0:0] CLBLM_R_X11Y116_SLICE_X14Y116_CO5;
  wire [0:0] CLBLM_R_X11Y116_SLICE_X14Y116_CO6;
  wire [0:0] CLBLM_R_X11Y116_SLICE_X14Y116_CQ;
  wire [0:0] CLBLM_R_X11Y116_SLICE_X14Y116_C_CY;
  wire [0:0] CLBLM_R_X11Y116_SLICE_X14Y116_C_XOR;
  wire [0:0] CLBLM_R_X11Y116_SLICE_X14Y116_D;
  wire [0:0] CLBLM_R_X11Y116_SLICE_X14Y116_D1;
  wire [0:0] CLBLM_R_X11Y116_SLICE_X14Y116_D2;
  wire [0:0] CLBLM_R_X11Y116_SLICE_X14Y116_D3;
  wire [0:0] CLBLM_R_X11Y116_SLICE_X14Y116_D4;
  wire [0:0] CLBLM_R_X11Y116_SLICE_X14Y116_D5;
  wire [0:0] CLBLM_R_X11Y116_SLICE_X14Y116_D6;
  wire [0:0] CLBLM_R_X11Y116_SLICE_X14Y116_DO5;
  wire [0:0] CLBLM_R_X11Y116_SLICE_X14Y116_DO6;
  wire [0:0] CLBLM_R_X11Y116_SLICE_X14Y116_DQ;
  wire [0:0] CLBLM_R_X11Y116_SLICE_X14Y116_D_CY;
  wire [0:0] CLBLM_R_X11Y116_SLICE_X14Y116_D_XOR;
  wire [0:0] CLBLM_R_X11Y116_SLICE_X15Y116_A;
  wire [0:0] CLBLM_R_X11Y116_SLICE_X15Y116_A1;
  wire [0:0] CLBLM_R_X11Y116_SLICE_X15Y116_A2;
  wire [0:0] CLBLM_R_X11Y116_SLICE_X15Y116_A3;
  wire [0:0] CLBLM_R_X11Y116_SLICE_X15Y116_A4;
  wire [0:0] CLBLM_R_X11Y116_SLICE_X15Y116_A5;
  wire [0:0] CLBLM_R_X11Y116_SLICE_X15Y116_A6;
  wire [0:0] CLBLM_R_X11Y116_SLICE_X15Y116_AO5;
  wire [0:0] CLBLM_R_X11Y116_SLICE_X15Y116_AO6;
  wire [0:0] CLBLM_R_X11Y116_SLICE_X15Y116_AQ;
  wire [0:0] CLBLM_R_X11Y116_SLICE_X15Y116_A_CY;
  wire [0:0] CLBLM_R_X11Y116_SLICE_X15Y116_A_XOR;
  wire [0:0] CLBLM_R_X11Y116_SLICE_X15Y116_B;
  wire [0:0] CLBLM_R_X11Y116_SLICE_X15Y116_B1;
  wire [0:0] CLBLM_R_X11Y116_SLICE_X15Y116_B2;
  wire [0:0] CLBLM_R_X11Y116_SLICE_X15Y116_B3;
  wire [0:0] CLBLM_R_X11Y116_SLICE_X15Y116_B4;
  wire [0:0] CLBLM_R_X11Y116_SLICE_X15Y116_B5;
  wire [0:0] CLBLM_R_X11Y116_SLICE_X15Y116_B6;
  wire [0:0] CLBLM_R_X11Y116_SLICE_X15Y116_BO5;
  wire [0:0] CLBLM_R_X11Y116_SLICE_X15Y116_BO6;
  wire [0:0] CLBLM_R_X11Y116_SLICE_X15Y116_B_CY;
  wire [0:0] CLBLM_R_X11Y116_SLICE_X15Y116_B_XOR;
  wire [0:0] CLBLM_R_X11Y116_SLICE_X15Y116_C;
  wire [0:0] CLBLM_R_X11Y116_SLICE_X15Y116_C1;
  wire [0:0] CLBLM_R_X11Y116_SLICE_X15Y116_C2;
  wire [0:0] CLBLM_R_X11Y116_SLICE_X15Y116_C3;
  wire [0:0] CLBLM_R_X11Y116_SLICE_X15Y116_C4;
  wire [0:0] CLBLM_R_X11Y116_SLICE_X15Y116_C5;
  wire [0:0] CLBLM_R_X11Y116_SLICE_X15Y116_C6;
  wire [0:0] CLBLM_R_X11Y116_SLICE_X15Y116_CLK;
  wire [0:0] CLBLM_R_X11Y116_SLICE_X15Y116_CO5;
  wire [0:0] CLBLM_R_X11Y116_SLICE_X15Y116_CO6;
  wire [0:0] CLBLM_R_X11Y116_SLICE_X15Y116_C_CY;
  wire [0:0] CLBLM_R_X11Y116_SLICE_X15Y116_C_XOR;
  wire [0:0] CLBLM_R_X11Y116_SLICE_X15Y116_D;
  wire [0:0] CLBLM_R_X11Y116_SLICE_X15Y116_D1;
  wire [0:0] CLBLM_R_X11Y116_SLICE_X15Y116_D2;
  wire [0:0] CLBLM_R_X11Y116_SLICE_X15Y116_D3;
  wire [0:0] CLBLM_R_X11Y116_SLICE_X15Y116_D4;
  wire [0:0] CLBLM_R_X11Y116_SLICE_X15Y116_D5;
  wire [0:0] CLBLM_R_X11Y116_SLICE_X15Y116_D6;
  wire [0:0] CLBLM_R_X11Y116_SLICE_X15Y116_DO5;
  wire [0:0] CLBLM_R_X11Y116_SLICE_X15Y116_DO6;
  wire [0:0] CLBLM_R_X11Y116_SLICE_X15Y116_D_CY;
  wire [0:0] CLBLM_R_X11Y116_SLICE_X15Y116_D_XOR;
  wire [0:0] CLBLM_R_X11Y117_SLICE_X14Y117_A;
  wire [0:0] CLBLM_R_X11Y117_SLICE_X14Y117_A1;
  wire [0:0] CLBLM_R_X11Y117_SLICE_X14Y117_A2;
  wire [0:0] CLBLM_R_X11Y117_SLICE_X14Y117_A3;
  wire [0:0] CLBLM_R_X11Y117_SLICE_X14Y117_A4;
  wire [0:0] CLBLM_R_X11Y117_SLICE_X14Y117_A5;
  wire [0:0] CLBLM_R_X11Y117_SLICE_X14Y117_A6;
  wire [0:0] CLBLM_R_X11Y117_SLICE_X14Y117_AO5;
  wire [0:0] CLBLM_R_X11Y117_SLICE_X14Y117_AO6;
  wire [0:0] CLBLM_R_X11Y117_SLICE_X14Y117_AQ;
  wire [0:0] CLBLM_R_X11Y117_SLICE_X14Y117_A_CY;
  wire [0:0] CLBLM_R_X11Y117_SLICE_X14Y117_A_XOR;
  wire [0:0] CLBLM_R_X11Y117_SLICE_X14Y117_B;
  wire [0:0] CLBLM_R_X11Y117_SLICE_X14Y117_B1;
  wire [0:0] CLBLM_R_X11Y117_SLICE_X14Y117_B2;
  wire [0:0] CLBLM_R_X11Y117_SLICE_X14Y117_B3;
  wire [0:0] CLBLM_R_X11Y117_SLICE_X14Y117_B4;
  wire [0:0] CLBLM_R_X11Y117_SLICE_X14Y117_B5;
  wire [0:0] CLBLM_R_X11Y117_SLICE_X14Y117_B6;
  wire [0:0] CLBLM_R_X11Y117_SLICE_X14Y117_BO5;
  wire [0:0] CLBLM_R_X11Y117_SLICE_X14Y117_BO6;
  wire [0:0] CLBLM_R_X11Y117_SLICE_X14Y117_BQ;
  wire [0:0] CLBLM_R_X11Y117_SLICE_X14Y117_B_CY;
  wire [0:0] CLBLM_R_X11Y117_SLICE_X14Y117_B_XOR;
  wire [0:0] CLBLM_R_X11Y117_SLICE_X14Y117_C;
  wire [0:0] CLBLM_R_X11Y117_SLICE_X14Y117_C1;
  wire [0:0] CLBLM_R_X11Y117_SLICE_X14Y117_C2;
  wire [0:0] CLBLM_R_X11Y117_SLICE_X14Y117_C3;
  wire [0:0] CLBLM_R_X11Y117_SLICE_X14Y117_C4;
  wire [0:0] CLBLM_R_X11Y117_SLICE_X14Y117_C5;
  wire [0:0] CLBLM_R_X11Y117_SLICE_X14Y117_C6;
  wire [0:0] CLBLM_R_X11Y117_SLICE_X14Y117_CLK;
  wire [0:0] CLBLM_R_X11Y117_SLICE_X14Y117_CO5;
  wire [0:0] CLBLM_R_X11Y117_SLICE_X14Y117_CO6;
  wire [0:0] CLBLM_R_X11Y117_SLICE_X14Y117_CQ;
  wire [0:0] CLBLM_R_X11Y117_SLICE_X14Y117_C_CY;
  wire [0:0] CLBLM_R_X11Y117_SLICE_X14Y117_C_XOR;
  wire [0:0] CLBLM_R_X11Y117_SLICE_X14Y117_D;
  wire [0:0] CLBLM_R_X11Y117_SLICE_X14Y117_D1;
  wire [0:0] CLBLM_R_X11Y117_SLICE_X14Y117_D2;
  wire [0:0] CLBLM_R_X11Y117_SLICE_X14Y117_D3;
  wire [0:0] CLBLM_R_X11Y117_SLICE_X14Y117_D4;
  wire [0:0] CLBLM_R_X11Y117_SLICE_X14Y117_D5;
  wire [0:0] CLBLM_R_X11Y117_SLICE_X14Y117_D6;
  wire [0:0] CLBLM_R_X11Y117_SLICE_X14Y117_DMUX;
  wire [0:0] CLBLM_R_X11Y117_SLICE_X14Y117_DO5;
  wire [0:0] CLBLM_R_X11Y117_SLICE_X14Y117_DO6;
  wire [0:0] CLBLM_R_X11Y117_SLICE_X14Y117_D_CY;
  wire [0:0] CLBLM_R_X11Y117_SLICE_X14Y117_D_XOR;
  wire [0:0] CLBLM_R_X11Y117_SLICE_X15Y117_A;
  wire [0:0] CLBLM_R_X11Y117_SLICE_X15Y117_A1;
  wire [0:0] CLBLM_R_X11Y117_SLICE_X15Y117_A2;
  wire [0:0] CLBLM_R_X11Y117_SLICE_X15Y117_A3;
  wire [0:0] CLBLM_R_X11Y117_SLICE_X15Y117_A4;
  wire [0:0] CLBLM_R_X11Y117_SLICE_X15Y117_A5;
  wire [0:0] CLBLM_R_X11Y117_SLICE_X15Y117_A6;
  wire [0:0] CLBLM_R_X11Y117_SLICE_X15Y117_AO5;
  wire [0:0] CLBLM_R_X11Y117_SLICE_X15Y117_AO6;
  wire [0:0] CLBLM_R_X11Y117_SLICE_X15Y117_AQ;
  wire [0:0] CLBLM_R_X11Y117_SLICE_X15Y117_A_CY;
  wire [0:0] CLBLM_R_X11Y117_SLICE_X15Y117_A_XOR;
  wire [0:0] CLBLM_R_X11Y117_SLICE_X15Y117_B;
  wire [0:0] CLBLM_R_X11Y117_SLICE_X15Y117_B1;
  wire [0:0] CLBLM_R_X11Y117_SLICE_X15Y117_B2;
  wire [0:0] CLBLM_R_X11Y117_SLICE_X15Y117_B3;
  wire [0:0] CLBLM_R_X11Y117_SLICE_X15Y117_B4;
  wire [0:0] CLBLM_R_X11Y117_SLICE_X15Y117_B5;
  wire [0:0] CLBLM_R_X11Y117_SLICE_X15Y117_B6;
  wire [0:0] CLBLM_R_X11Y117_SLICE_X15Y117_BO5;
  wire [0:0] CLBLM_R_X11Y117_SLICE_X15Y117_BO6;
  wire [0:0] CLBLM_R_X11Y117_SLICE_X15Y117_B_CY;
  wire [0:0] CLBLM_R_X11Y117_SLICE_X15Y117_B_XOR;
  wire [0:0] CLBLM_R_X11Y117_SLICE_X15Y117_C;
  wire [0:0] CLBLM_R_X11Y117_SLICE_X15Y117_C1;
  wire [0:0] CLBLM_R_X11Y117_SLICE_X15Y117_C2;
  wire [0:0] CLBLM_R_X11Y117_SLICE_X15Y117_C3;
  wire [0:0] CLBLM_R_X11Y117_SLICE_X15Y117_C4;
  wire [0:0] CLBLM_R_X11Y117_SLICE_X15Y117_C5;
  wire [0:0] CLBLM_R_X11Y117_SLICE_X15Y117_C6;
  wire [0:0] CLBLM_R_X11Y117_SLICE_X15Y117_CLK;
  wire [0:0] CLBLM_R_X11Y117_SLICE_X15Y117_CO5;
  wire [0:0] CLBLM_R_X11Y117_SLICE_X15Y117_CO6;
  wire [0:0] CLBLM_R_X11Y117_SLICE_X15Y117_C_CY;
  wire [0:0] CLBLM_R_X11Y117_SLICE_X15Y117_C_XOR;
  wire [0:0] CLBLM_R_X11Y117_SLICE_X15Y117_D;
  wire [0:0] CLBLM_R_X11Y117_SLICE_X15Y117_D1;
  wire [0:0] CLBLM_R_X11Y117_SLICE_X15Y117_D2;
  wire [0:0] CLBLM_R_X11Y117_SLICE_X15Y117_D3;
  wire [0:0] CLBLM_R_X11Y117_SLICE_X15Y117_D4;
  wire [0:0] CLBLM_R_X11Y117_SLICE_X15Y117_D5;
  wire [0:0] CLBLM_R_X11Y117_SLICE_X15Y117_D6;
  wire [0:0] CLBLM_R_X11Y117_SLICE_X15Y117_DO5;
  wire [0:0] CLBLM_R_X11Y117_SLICE_X15Y117_DO6;
  wire [0:0] CLBLM_R_X11Y117_SLICE_X15Y117_D_CY;
  wire [0:0] CLBLM_R_X11Y117_SLICE_X15Y117_D_XOR;
  wire [0:0] CLBLM_R_X11Y118_SLICE_X14Y118_A;
  wire [0:0] CLBLM_R_X11Y118_SLICE_X14Y118_A1;
  wire [0:0] CLBLM_R_X11Y118_SLICE_X14Y118_A2;
  wire [0:0] CLBLM_R_X11Y118_SLICE_X14Y118_A3;
  wire [0:0] CLBLM_R_X11Y118_SLICE_X14Y118_A4;
  wire [0:0] CLBLM_R_X11Y118_SLICE_X14Y118_A5;
  wire [0:0] CLBLM_R_X11Y118_SLICE_X14Y118_A6;
  wire [0:0] CLBLM_R_X11Y118_SLICE_X14Y118_AO5;
  wire [0:0] CLBLM_R_X11Y118_SLICE_X14Y118_AO6;
  wire [0:0] CLBLM_R_X11Y118_SLICE_X14Y118_AQ;
  wire [0:0] CLBLM_R_X11Y118_SLICE_X14Y118_A_CY;
  wire [0:0] CLBLM_R_X11Y118_SLICE_X14Y118_A_XOR;
  wire [0:0] CLBLM_R_X11Y118_SLICE_X14Y118_B;
  wire [0:0] CLBLM_R_X11Y118_SLICE_X14Y118_B1;
  wire [0:0] CLBLM_R_X11Y118_SLICE_X14Y118_B2;
  wire [0:0] CLBLM_R_X11Y118_SLICE_X14Y118_B3;
  wire [0:0] CLBLM_R_X11Y118_SLICE_X14Y118_B4;
  wire [0:0] CLBLM_R_X11Y118_SLICE_X14Y118_B5;
  wire [0:0] CLBLM_R_X11Y118_SLICE_X14Y118_B6;
  wire [0:0] CLBLM_R_X11Y118_SLICE_X14Y118_BO5;
  wire [0:0] CLBLM_R_X11Y118_SLICE_X14Y118_BO6;
  wire [0:0] CLBLM_R_X11Y118_SLICE_X14Y118_BQ;
  wire [0:0] CLBLM_R_X11Y118_SLICE_X14Y118_B_CY;
  wire [0:0] CLBLM_R_X11Y118_SLICE_X14Y118_B_XOR;
  wire [0:0] CLBLM_R_X11Y118_SLICE_X14Y118_C;
  wire [0:0] CLBLM_R_X11Y118_SLICE_X14Y118_C1;
  wire [0:0] CLBLM_R_X11Y118_SLICE_X14Y118_C2;
  wire [0:0] CLBLM_R_X11Y118_SLICE_X14Y118_C3;
  wire [0:0] CLBLM_R_X11Y118_SLICE_X14Y118_C4;
  wire [0:0] CLBLM_R_X11Y118_SLICE_X14Y118_C5;
  wire [0:0] CLBLM_R_X11Y118_SLICE_X14Y118_C6;
  wire [0:0] CLBLM_R_X11Y118_SLICE_X14Y118_CLK;
  wire [0:0] CLBLM_R_X11Y118_SLICE_X14Y118_CO5;
  wire [0:0] CLBLM_R_X11Y118_SLICE_X14Y118_CO6;
  wire [0:0] CLBLM_R_X11Y118_SLICE_X14Y118_CQ;
  wire [0:0] CLBLM_R_X11Y118_SLICE_X14Y118_C_CY;
  wire [0:0] CLBLM_R_X11Y118_SLICE_X14Y118_C_XOR;
  wire [0:0] CLBLM_R_X11Y118_SLICE_X14Y118_D;
  wire [0:0] CLBLM_R_X11Y118_SLICE_X14Y118_D1;
  wire [0:0] CLBLM_R_X11Y118_SLICE_X14Y118_D2;
  wire [0:0] CLBLM_R_X11Y118_SLICE_X14Y118_D3;
  wire [0:0] CLBLM_R_X11Y118_SLICE_X14Y118_D4;
  wire [0:0] CLBLM_R_X11Y118_SLICE_X14Y118_D5;
  wire [0:0] CLBLM_R_X11Y118_SLICE_X14Y118_D6;
  wire [0:0] CLBLM_R_X11Y118_SLICE_X14Y118_DMUX;
  wire [0:0] CLBLM_R_X11Y118_SLICE_X14Y118_DO5;
  wire [0:0] CLBLM_R_X11Y118_SLICE_X14Y118_DO6;
  wire [0:0] CLBLM_R_X11Y118_SLICE_X14Y118_D_CY;
  wire [0:0] CLBLM_R_X11Y118_SLICE_X14Y118_D_XOR;
  wire [0:0] CLBLM_R_X11Y118_SLICE_X15Y118_A;
  wire [0:0] CLBLM_R_X11Y118_SLICE_X15Y118_A1;
  wire [0:0] CLBLM_R_X11Y118_SLICE_X15Y118_A2;
  wire [0:0] CLBLM_R_X11Y118_SLICE_X15Y118_A3;
  wire [0:0] CLBLM_R_X11Y118_SLICE_X15Y118_A4;
  wire [0:0] CLBLM_R_X11Y118_SLICE_X15Y118_A5;
  wire [0:0] CLBLM_R_X11Y118_SLICE_X15Y118_A6;
  wire [0:0] CLBLM_R_X11Y118_SLICE_X15Y118_AO5;
  wire [0:0] CLBLM_R_X11Y118_SLICE_X15Y118_AO6;
  wire [0:0] CLBLM_R_X11Y118_SLICE_X15Y118_AQ;
  wire [0:0] CLBLM_R_X11Y118_SLICE_X15Y118_A_CY;
  wire [0:0] CLBLM_R_X11Y118_SLICE_X15Y118_A_XOR;
  wire [0:0] CLBLM_R_X11Y118_SLICE_X15Y118_B;
  wire [0:0] CLBLM_R_X11Y118_SLICE_X15Y118_B1;
  wire [0:0] CLBLM_R_X11Y118_SLICE_X15Y118_B2;
  wire [0:0] CLBLM_R_X11Y118_SLICE_X15Y118_B3;
  wire [0:0] CLBLM_R_X11Y118_SLICE_X15Y118_B4;
  wire [0:0] CLBLM_R_X11Y118_SLICE_X15Y118_B5;
  wire [0:0] CLBLM_R_X11Y118_SLICE_X15Y118_B6;
  wire [0:0] CLBLM_R_X11Y118_SLICE_X15Y118_BO5;
  wire [0:0] CLBLM_R_X11Y118_SLICE_X15Y118_BO6;
  wire [0:0] CLBLM_R_X11Y118_SLICE_X15Y118_BQ;
  wire [0:0] CLBLM_R_X11Y118_SLICE_X15Y118_B_CY;
  wire [0:0] CLBLM_R_X11Y118_SLICE_X15Y118_B_XOR;
  wire [0:0] CLBLM_R_X11Y118_SLICE_X15Y118_C;
  wire [0:0] CLBLM_R_X11Y118_SLICE_X15Y118_C1;
  wire [0:0] CLBLM_R_X11Y118_SLICE_X15Y118_C2;
  wire [0:0] CLBLM_R_X11Y118_SLICE_X15Y118_C3;
  wire [0:0] CLBLM_R_X11Y118_SLICE_X15Y118_C4;
  wire [0:0] CLBLM_R_X11Y118_SLICE_X15Y118_C5;
  wire [0:0] CLBLM_R_X11Y118_SLICE_X15Y118_C6;
  wire [0:0] CLBLM_R_X11Y118_SLICE_X15Y118_CLK;
  wire [0:0] CLBLM_R_X11Y118_SLICE_X15Y118_CO5;
  wire [0:0] CLBLM_R_X11Y118_SLICE_X15Y118_CO6;
  wire [0:0] CLBLM_R_X11Y118_SLICE_X15Y118_CQ;
  wire [0:0] CLBLM_R_X11Y118_SLICE_X15Y118_C_CY;
  wire [0:0] CLBLM_R_X11Y118_SLICE_X15Y118_C_XOR;
  wire [0:0] CLBLM_R_X11Y118_SLICE_X15Y118_D;
  wire [0:0] CLBLM_R_X11Y118_SLICE_X15Y118_D1;
  wire [0:0] CLBLM_R_X11Y118_SLICE_X15Y118_D2;
  wire [0:0] CLBLM_R_X11Y118_SLICE_X15Y118_D3;
  wire [0:0] CLBLM_R_X11Y118_SLICE_X15Y118_D4;
  wire [0:0] CLBLM_R_X11Y118_SLICE_X15Y118_D5;
  wire [0:0] CLBLM_R_X11Y118_SLICE_X15Y118_D6;
  wire [0:0] CLBLM_R_X11Y118_SLICE_X15Y118_DO5;
  wire [0:0] CLBLM_R_X11Y118_SLICE_X15Y118_DO6;
  wire [0:0] CLBLM_R_X11Y118_SLICE_X15Y118_D_CY;
  wire [0:0] CLBLM_R_X11Y118_SLICE_X15Y118_D_XOR;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X14Y119_A;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X14Y119_A1;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X14Y119_A2;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X14Y119_A3;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X14Y119_A4;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X14Y119_A5;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X14Y119_A6;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X14Y119_AMUX;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X14Y119_AO5;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X14Y119_AO6;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X14Y119_AQ;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X14Y119_AX;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X14Y119_A_CY;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X14Y119_A_XOR;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X14Y119_B;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X14Y119_B1;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X14Y119_B2;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X14Y119_B3;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X14Y119_B4;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X14Y119_B5;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X14Y119_B6;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X14Y119_BMUX;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X14Y119_BO5;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X14Y119_BO6;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X14Y119_B_CY;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X14Y119_B_XOR;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X14Y119_C;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X14Y119_C1;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X14Y119_C2;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X14Y119_C3;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X14Y119_C4;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X14Y119_C5;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X14Y119_C6;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X14Y119_CE;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X14Y119_CLK;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X14Y119_CMUX;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X14Y119_CO5;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X14Y119_CO6;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X14Y119_C_CY;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X14Y119_C_XOR;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X14Y119_D;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X14Y119_D1;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X14Y119_D2;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X14Y119_D3;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X14Y119_D4;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X14Y119_D5;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X14Y119_D6;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X14Y119_DO5;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X14Y119_DO6;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X14Y119_D_CY;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X14Y119_D_XOR;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X14Y119_SR;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X15Y119_A;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X15Y119_A1;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X15Y119_A2;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X15Y119_A3;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X15Y119_A4;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X15Y119_A5;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X15Y119_A6;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X15Y119_AO5;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X15Y119_AO6;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X15Y119_AQ;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X15Y119_A_CY;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X15Y119_A_XOR;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X15Y119_B;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X15Y119_B1;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X15Y119_B2;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X15Y119_B3;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X15Y119_B4;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X15Y119_B5;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X15Y119_B6;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X15Y119_BO5;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X15Y119_BO6;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X15Y119_BQ;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X15Y119_B_CY;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X15Y119_B_XOR;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X15Y119_C;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X15Y119_C1;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X15Y119_C2;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X15Y119_C3;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X15Y119_C4;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X15Y119_C5;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X15Y119_C6;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X15Y119_CLK;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X15Y119_CO5;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X15Y119_CO6;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X15Y119_CQ;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X15Y119_C_CY;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X15Y119_C_XOR;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X15Y119_D;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X15Y119_D1;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X15Y119_D2;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X15Y119_D3;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X15Y119_D4;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X15Y119_D5;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X15Y119_D6;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X15Y119_DO5;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X15Y119_DO6;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X15Y119_D_CY;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X15Y119_D_XOR;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X14Y120_A;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X14Y120_A1;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X14Y120_A2;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X14Y120_A3;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X14Y120_A4;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X14Y120_A5;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X14Y120_A6;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X14Y120_AMUX;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X14Y120_AO5;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X14Y120_AO6;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X14Y120_AQ;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X14Y120_AX;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X14Y120_A_CY;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X14Y120_A_XOR;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X14Y120_B;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X14Y120_B1;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X14Y120_B2;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X14Y120_B3;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X14Y120_B4;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X14Y120_B5;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X14Y120_B6;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X14Y120_BMUX;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X14Y120_BO5;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X14Y120_BO6;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X14Y120_B_CY;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X14Y120_B_XOR;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X14Y120_C;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X14Y120_C1;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X14Y120_C2;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X14Y120_C3;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X14Y120_C4;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X14Y120_C5;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X14Y120_C6;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X14Y120_CE;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X14Y120_CLK;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X14Y120_CO5;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X14Y120_CO6;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X14Y120_C_CY;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X14Y120_C_XOR;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X14Y120_D;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X14Y120_D1;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X14Y120_D2;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X14Y120_D3;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X14Y120_D4;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X14Y120_D5;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X14Y120_D6;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X14Y120_DO5;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X14Y120_DO6;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X14Y120_D_CY;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X14Y120_D_XOR;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X14Y120_SR;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X15Y120_A;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X15Y120_A1;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X15Y120_A2;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X15Y120_A3;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X15Y120_A4;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X15Y120_A5;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X15Y120_A6;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X15Y120_AO5;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X15Y120_AO6;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X15Y120_AQ;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X15Y120_A_CY;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X15Y120_A_XOR;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X15Y120_B;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X15Y120_B1;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X15Y120_B2;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X15Y120_B3;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X15Y120_B4;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X15Y120_B5;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X15Y120_B6;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X15Y120_BO5;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X15Y120_BO6;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X15Y120_BQ;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X15Y120_B_CY;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X15Y120_B_XOR;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X15Y120_C;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X15Y120_C1;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X15Y120_C2;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X15Y120_C3;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X15Y120_C4;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X15Y120_C5;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X15Y120_C6;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X15Y120_CLK;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X15Y120_CO5;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X15Y120_CO6;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X15Y120_CQ;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X15Y120_C_CY;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X15Y120_C_XOR;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X15Y120_D;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X15Y120_D1;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X15Y120_D2;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X15Y120_D3;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X15Y120_D4;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X15Y120_D5;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X15Y120_D6;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X15Y120_DO5;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X15Y120_DO6;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X15Y120_D_CY;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X15Y120_D_XOR;
  wire [0:0] CLBLM_R_X11Y121_SLICE_X14Y121_A;
  wire [0:0] CLBLM_R_X11Y121_SLICE_X14Y121_A1;
  wire [0:0] CLBLM_R_X11Y121_SLICE_X14Y121_A2;
  wire [0:0] CLBLM_R_X11Y121_SLICE_X14Y121_A3;
  wire [0:0] CLBLM_R_X11Y121_SLICE_X14Y121_A4;
  wire [0:0] CLBLM_R_X11Y121_SLICE_X14Y121_A5;
  wire [0:0] CLBLM_R_X11Y121_SLICE_X14Y121_A6;
  wire [0:0] CLBLM_R_X11Y121_SLICE_X14Y121_AO5;
  wire [0:0] CLBLM_R_X11Y121_SLICE_X14Y121_AO6;
  wire [0:0] CLBLM_R_X11Y121_SLICE_X14Y121_AQ;
  wire [0:0] CLBLM_R_X11Y121_SLICE_X14Y121_A_CY;
  wire [0:0] CLBLM_R_X11Y121_SLICE_X14Y121_A_XOR;
  wire [0:0] CLBLM_R_X11Y121_SLICE_X14Y121_B;
  wire [0:0] CLBLM_R_X11Y121_SLICE_X14Y121_B1;
  wire [0:0] CLBLM_R_X11Y121_SLICE_X14Y121_B2;
  wire [0:0] CLBLM_R_X11Y121_SLICE_X14Y121_B3;
  wire [0:0] CLBLM_R_X11Y121_SLICE_X14Y121_B4;
  wire [0:0] CLBLM_R_X11Y121_SLICE_X14Y121_B5;
  wire [0:0] CLBLM_R_X11Y121_SLICE_X14Y121_B6;
  wire [0:0] CLBLM_R_X11Y121_SLICE_X14Y121_BMUX;
  wire [0:0] CLBLM_R_X11Y121_SLICE_X14Y121_BO5;
  wire [0:0] CLBLM_R_X11Y121_SLICE_X14Y121_BO6;
  wire [0:0] CLBLM_R_X11Y121_SLICE_X14Y121_B_CY;
  wire [0:0] CLBLM_R_X11Y121_SLICE_X14Y121_B_XOR;
  wire [0:0] CLBLM_R_X11Y121_SLICE_X14Y121_C;
  wire [0:0] CLBLM_R_X11Y121_SLICE_X14Y121_C1;
  wire [0:0] CLBLM_R_X11Y121_SLICE_X14Y121_C2;
  wire [0:0] CLBLM_R_X11Y121_SLICE_X14Y121_C3;
  wire [0:0] CLBLM_R_X11Y121_SLICE_X14Y121_C4;
  wire [0:0] CLBLM_R_X11Y121_SLICE_X14Y121_C5;
  wire [0:0] CLBLM_R_X11Y121_SLICE_X14Y121_C6;
  wire [0:0] CLBLM_R_X11Y121_SLICE_X14Y121_CLK;
  wire [0:0] CLBLM_R_X11Y121_SLICE_X14Y121_CO5;
  wire [0:0] CLBLM_R_X11Y121_SLICE_X14Y121_CO6;
  wire [0:0] CLBLM_R_X11Y121_SLICE_X14Y121_C_CY;
  wire [0:0] CLBLM_R_X11Y121_SLICE_X14Y121_C_XOR;
  wire [0:0] CLBLM_R_X11Y121_SLICE_X14Y121_D;
  wire [0:0] CLBLM_R_X11Y121_SLICE_X14Y121_D1;
  wire [0:0] CLBLM_R_X11Y121_SLICE_X14Y121_D2;
  wire [0:0] CLBLM_R_X11Y121_SLICE_X14Y121_D3;
  wire [0:0] CLBLM_R_X11Y121_SLICE_X14Y121_D4;
  wire [0:0] CLBLM_R_X11Y121_SLICE_X14Y121_D5;
  wire [0:0] CLBLM_R_X11Y121_SLICE_X14Y121_D6;
  wire [0:0] CLBLM_R_X11Y121_SLICE_X14Y121_DO5;
  wire [0:0] CLBLM_R_X11Y121_SLICE_X14Y121_DO6;
  wire [0:0] CLBLM_R_X11Y121_SLICE_X14Y121_D_CY;
  wire [0:0] CLBLM_R_X11Y121_SLICE_X14Y121_D_XOR;
  wire [0:0] CLBLM_R_X11Y121_SLICE_X15Y121_A;
  wire [0:0] CLBLM_R_X11Y121_SLICE_X15Y121_A1;
  wire [0:0] CLBLM_R_X11Y121_SLICE_X15Y121_A2;
  wire [0:0] CLBLM_R_X11Y121_SLICE_X15Y121_A3;
  wire [0:0] CLBLM_R_X11Y121_SLICE_X15Y121_A4;
  wire [0:0] CLBLM_R_X11Y121_SLICE_X15Y121_A5;
  wire [0:0] CLBLM_R_X11Y121_SLICE_X15Y121_A6;
  wire [0:0] CLBLM_R_X11Y121_SLICE_X15Y121_AMUX;
  wire [0:0] CLBLM_R_X11Y121_SLICE_X15Y121_AO5;
  wire [0:0] CLBLM_R_X11Y121_SLICE_X15Y121_AO6;
  wire [0:0] CLBLM_R_X11Y121_SLICE_X15Y121_A_CY;
  wire [0:0] CLBLM_R_X11Y121_SLICE_X15Y121_A_XOR;
  wire [0:0] CLBLM_R_X11Y121_SLICE_X15Y121_B;
  wire [0:0] CLBLM_R_X11Y121_SLICE_X15Y121_B1;
  wire [0:0] CLBLM_R_X11Y121_SLICE_X15Y121_B2;
  wire [0:0] CLBLM_R_X11Y121_SLICE_X15Y121_B3;
  wire [0:0] CLBLM_R_X11Y121_SLICE_X15Y121_B4;
  wire [0:0] CLBLM_R_X11Y121_SLICE_X15Y121_B5;
  wire [0:0] CLBLM_R_X11Y121_SLICE_X15Y121_B6;
  wire [0:0] CLBLM_R_X11Y121_SLICE_X15Y121_BO5;
  wire [0:0] CLBLM_R_X11Y121_SLICE_X15Y121_BO6;
  wire [0:0] CLBLM_R_X11Y121_SLICE_X15Y121_B_CY;
  wire [0:0] CLBLM_R_X11Y121_SLICE_X15Y121_B_XOR;
  wire [0:0] CLBLM_R_X11Y121_SLICE_X15Y121_C;
  wire [0:0] CLBLM_R_X11Y121_SLICE_X15Y121_C1;
  wire [0:0] CLBLM_R_X11Y121_SLICE_X15Y121_C2;
  wire [0:0] CLBLM_R_X11Y121_SLICE_X15Y121_C3;
  wire [0:0] CLBLM_R_X11Y121_SLICE_X15Y121_C4;
  wire [0:0] CLBLM_R_X11Y121_SLICE_X15Y121_C5;
  wire [0:0] CLBLM_R_X11Y121_SLICE_X15Y121_C6;
  wire [0:0] CLBLM_R_X11Y121_SLICE_X15Y121_CO5;
  wire [0:0] CLBLM_R_X11Y121_SLICE_X15Y121_CO6;
  wire [0:0] CLBLM_R_X11Y121_SLICE_X15Y121_C_CY;
  wire [0:0] CLBLM_R_X11Y121_SLICE_X15Y121_C_XOR;
  wire [0:0] CLBLM_R_X11Y121_SLICE_X15Y121_D;
  wire [0:0] CLBLM_R_X11Y121_SLICE_X15Y121_D1;
  wire [0:0] CLBLM_R_X11Y121_SLICE_X15Y121_D2;
  wire [0:0] CLBLM_R_X11Y121_SLICE_X15Y121_D3;
  wire [0:0] CLBLM_R_X11Y121_SLICE_X15Y121_D4;
  wire [0:0] CLBLM_R_X11Y121_SLICE_X15Y121_D5;
  wire [0:0] CLBLM_R_X11Y121_SLICE_X15Y121_D6;
  wire [0:0] CLBLM_R_X11Y121_SLICE_X15Y121_DO5;
  wire [0:0] CLBLM_R_X11Y121_SLICE_X15Y121_DO6;
  wire [0:0] CLBLM_R_X11Y121_SLICE_X15Y121_D_CY;
  wire [0:0] CLBLM_R_X11Y121_SLICE_X15Y121_D_XOR;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X14Y122_A;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X14Y122_A1;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X14Y122_A2;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X14Y122_A3;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X14Y122_A4;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X14Y122_A5;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X14Y122_A6;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X14Y122_AO5;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X14Y122_AO6;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X14Y122_AQ;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X14Y122_A_CY;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X14Y122_A_XOR;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X14Y122_B;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X14Y122_B1;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X14Y122_B2;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X14Y122_B3;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X14Y122_B4;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X14Y122_B5;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X14Y122_B6;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X14Y122_BO5;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X14Y122_BO6;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X14Y122_B_CY;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X14Y122_B_XOR;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X14Y122_C;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X14Y122_C1;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X14Y122_C2;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X14Y122_C3;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X14Y122_C4;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X14Y122_C5;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X14Y122_C6;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X14Y122_CLK;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X14Y122_CO5;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X14Y122_CO6;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X14Y122_C_CY;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X14Y122_C_XOR;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X14Y122_D;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X14Y122_D1;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X14Y122_D2;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X14Y122_D3;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X14Y122_D4;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X14Y122_D5;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X14Y122_D6;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X14Y122_DO5;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X14Y122_DO6;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X14Y122_D_CY;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X14Y122_D_XOR;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X15Y122_A;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X15Y122_A1;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X15Y122_A2;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X15Y122_A3;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X15Y122_A4;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X15Y122_A5;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X15Y122_A6;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X15Y122_AO5;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X15Y122_AO6;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X15Y122_A_CY;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X15Y122_A_XOR;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X15Y122_B;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X15Y122_B1;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X15Y122_B2;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X15Y122_B3;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X15Y122_B4;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X15Y122_B5;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X15Y122_B6;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X15Y122_BO5;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X15Y122_BO6;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X15Y122_B_CY;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X15Y122_B_XOR;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X15Y122_C;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X15Y122_C1;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X15Y122_C2;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X15Y122_C3;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X15Y122_C4;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X15Y122_C5;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X15Y122_C6;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X15Y122_CO5;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X15Y122_CO6;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X15Y122_C_CY;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X15Y122_C_XOR;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X15Y122_D;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X15Y122_D1;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X15Y122_D2;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X15Y122_D3;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X15Y122_D4;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X15Y122_D5;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X15Y122_D6;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X15Y122_DO5;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X15Y122_DO6;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X15Y122_D_CY;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X15Y122_D_XOR;
  wire [0:0] CLBLM_R_X11Y123_SLICE_X14Y123_A;
  wire [0:0] CLBLM_R_X11Y123_SLICE_X14Y123_A1;
  wire [0:0] CLBLM_R_X11Y123_SLICE_X14Y123_A2;
  wire [0:0] CLBLM_R_X11Y123_SLICE_X14Y123_A3;
  wire [0:0] CLBLM_R_X11Y123_SLICE_X14Y123_A4;
  wire [0:0] CLBLM_R_X11Y123_SLICE_X14Y123_A5;
  wire [0:0] CLBLM_R_X11Y123_SLICE_X14Y123_A6;
  wire [0:0] CLBLM_R_X11Y123_SLICE_X14Y123_AMUX;
  wire [0:0] CLBLM_R_X11Y123_SLICE_X14Y123_AO5;
  wire [0:0] CLBLM_R_X11Y123_SLICE_X14Y123_AO6;
  wire [0:0] CLBLM_R_X11Y123_SLICE_X14Y123_A_CY;
  wire [0:0] CLBLM_R_X11Y123_SLICE_X14Y123_A_XOR;
  wire [0:0] CLBLM_R_X11Y123_SLICE_X14Y123_B;
  wire [0:0] CLBLM_R_X11Y123_SLICE_X14Y123_B1;
  wire [0:0] CLBLM_R_X11Y123_SLICE_X14Y123_B2;
  wire [0:0] CLBLM_R_X11Y123_SLICE_X14Y123_B3;
  wire [0:0] CLBLM_R_X11Y123_SLICE_X14Y123_B4;
  wire [0:0] CLBLM_R_X11Y123_SLICE_X14Y123_B5;
  wire [0:0] CLBLM_R_X11Y123_SLICE_X14Y123_B6;
  wire [0:0] CLBLM_R_X11Y123_SLICE_X14Y123_BMUX;
  wire [0:0] CLBLM_R_X11Y123_SLICE_X14Y123_BO5;
  wire [0:0] CLBLM_R_X11Y123_SLICE_X14Y123_BO6;
  wire [0:0] CLBLM_R_X11Y123_SLICE_X14Y123_B_CY;
  wire [0:0] CLBLM_R_X11Y123_SLICE_X14Y123_B_XOR;
  wire [0:0] CLBLM_R_X11Y123_SLICE_X14Y123_C;
  wire [0:0] CLBLM_R_X11Y123_SLICE_X14Y123_C1;
  wire [0:0] CLBLM_R_X11Y123_SLICE_X14Y123_C2;
  wire [0:0] CLBLM_R_X11Y123_SLICE_X14Y123_C3;
  wire [0:0] CLBLM_R_X11Y123_SLICE_X14Y123_C4;
  wire [0:0] CLBLM_R_X11Y123_SLICE_X14Y123_C5;
  wire [0:0] CLBLM_R_X11Y123_SLICE_X14Y123_C6;
  wire [0:0] CLBLM_R_X11Y123_SLICE_X14Y123_CO5;
  wire [0:0] CLBLM_R_X11Y123_SLICE_X14Y123_CO6;
  wire [0:0] CLBLM_R_X11Y123_SLICE_X14Y123_C_CY;
  wire [0:0] CLBLM_R_X11Y123_SLICE_X14Y123_C_XOR;
  wire [0:0] CLBLM_R_X11Y123_SLICE_X14Y123_D;
  wire [0:0] CLBLM_R_X11Y123_SLICE_X14Y123_D1;
  wire [0:0] CLBLM_R_X11Y123_SLICE_X14Y123_D2;
  wire [0:0] CLBLM_R_X11Y123_SLICE_X14Y123_D3;
  wire [0:0] CLBLM_R_X11Y123_SLICE_X14Y123_D4;
  wire [0:0] CLBLM_R_X11Y123_SLICE_X14Y123_D5;
  wire [0:0] CLBLM_R_X11Y123_SLICE_X14Y123_D6;
  wire [0:0] CLBLM_R_X11Y123_SLICE_X14Y123_DO5;
  wire [0:0] CLBLM_R_X11Y123_SLICE_X14Y123_DO6;
  wire [0:0] CLBLM_R_X11Y123_SLICE_X14Y123_D_CY;
  wire [0:0] CLBLM_R_X11Y123_SLICE_X14Y123_D_XOR;
  wire [0:0] CLBLM_R_X11Y123_SLICE_X15Y123_A;
  wire [0:0] CLBLM_R_X11Y123_SLICE_X15Y123_A1;
  wire [0:0] CLBLM_R_X11Y123_SLICE_X15Y123_A2;
  wire [0:0] CLBLM_R_X11Y123_SLICE_X15Y123_A3;
  wire [0:0] CLBLM_R_X11Y123_SLICE_X15Y123_A4;
  wire [0:0] CLBLM_R_X11Y123_SLICE_X15Y123_A5;
  wire [0:0] CLBLM_R_X11Y123_SLICE_X15Y123_A6;
  wire [0:0] CLBLM_R_X11Y123_SLICE_X15Y123_AO5;
  wire [0:0] CLBLM_R_X11Y123_SLICE_X15Y123_AO6;
  wire [0:0] CLBLM_R_X11Y123_SLICE_X15Y123_A_CY;
  wire [0:0] CLBLM_R_X11Y123_SLICE_X15Y123_A_XOR;
  wire [0:0] CLBLM_R_X11Y123_SLICE_X15Y123_B;
  wire [0:0] CLBLM_R_X11Y123_SLICE_X15Y123_B1;
  wire [0:0] CLBLM_R_X11Y123_SLICE_X15Y123_B2;
  wire [0:0] CLBLM_R_X11Y123_SLICE_X15Y123_B3;
  wire [0:0] CLBLM_R_X11Y123_SLICE_X15Y123_B4;
  wire [0:0] CLBLM_R_X11Y123_SLICE_X15Y123_B5;
  wire [0:0] CLBLM_R_X11Y123_SLICE_X15Y123_B6;
  wire [0:0] CLBLM_R_X11Y123_SLICE_X15Y123_BO5;
  wire [0:0] CLBLM_R_X11Y123_SLICE_X15Y123_BO6;
  wire [0:0] CLBLM_R_X11Y123_SLICE_X15Y123_B_CY;
  wire [0:0] CLBLM_R_X11Y123_SLICE_X15Y123_B_XOR;
  wire [0:0] CLBLM_R_X11Y123_SLICE_X15Y123_C;
  wire [0:0] CLBLM_R_X11Y123_SLICE_X15Y123_C1;
  wire [0:0] CLBLM_R_X11Y123_SLICE_X15Y123_C2;
  wire [0:0] CLBLM_R_X11Y123_SLICE_X15Y123_C3;
  wire [0:0] CLBLM_R_X11Y123_SLICE_X15Y123_C4;
  wire [0:0] CLBLM_R_X11Y123_SLICE_X15Y123_C5;
  wire [0:0] CLBLM_R_X11Y123_SLICE_X15Y123_C6;
  wire [0:0] CLBLM_R_X11Y123_SLICE_X15Y123_CO5;
  wire [0:0] CLBLM_R_X11Y123_SLICE_X15Y123_CO6;
  wire [0:0] CLBLM_R_X11Y123_SLICE_X15Y123_C_CY;
  wire [0:0] CLBLM_R_X11Y123_SLICE_X15Y123_C_XOR;
  wire [0:0] CLBLM_R_X11Y123_SLICE_X15Y123_D;
  wire [0:0] CLBLM_R_X11Y123_SLICE_X15Y123_D1;
  wire [0:0] CLBLM_R_X11Y123_SLICE_X15Y123_D2;
  wire [0:0] CLBLM_R_X11Y123_SLICE_X15Y123_D3;
  wire [0:0] CLBLM_R_X11Y123_SLICE_X15Y123_D4;
  wire [0:0] CLBLM_R_X11Y123_SLICE_X15Y123_D5;
  wire [0:0] CLBLM_R_X11Y123_SLICE_X15Y123_D6;
  wire [0:0] CLBLM_R_X11Y123_SLICE_X15Y123_DO5;
  wire [0:0] CLBLM_R_X11Y123_SLICE_X15Y123_DO6;
  wire [0:0] CLBLM_R_X11Y123_SLICE_X15Y123_D_CY;
  wire [0:0] CLBLM_R_X11Y123_SLICE_X15Y123_D_XOR;
  wire [0:0] CLBLM_R_X11Y128_SLICE_X14Y128_A;
  wire [0:0] CLBLM_R_X11Y128_SLICE_X14Y128_A1;
  wire [0:0] CLBLM_R_X11Y128_SLICE_X14Y128_A2;
  wire [0:0] CLBLM_R_X11Y128_SLICE_X14Y128_A3;
  wire [0:0] CLBLM_R_X11Y128_SLICE_X14Y128_A4;
  wire [0:0] CLBLM_R_X11Y128_SLICE_X14Y128_A5;
  wire [0:0] CLBLM_R_X11Y128_SLICE_X14Y128_A6;
  wire [0:0] CLBLM_R_X11Y128_SLICE_X14Y128_AMUX;
  wire [0:0] CLBLM_R_X11Y128_SLICE_X14Y128_AO5;
  wire [0:0] CLBLM_R_X11Y128_SLICE_X14Y128_AO6;
  wire [0:0] CLBLM_R_X11Y128_SLICE_X14Y128_A_CY;
  wire [0:0] CLBLM_R_X11Y128_SLICE_X14Y128_A_XOR;
  wire [0:0] CLBLM_R_X11Y128_SLICE_X14Y128_B;
  wire [0:0] CLBLM_R_X11Y128_SLICE_X14Y128_B1;
  wire [0:0] CLBLM_R_X11Y128_SLICE_X14Y128_B2;
  wire [0:0] CLBLM_R_X11Y128_SLICE_X14Y128_B3;
  wire [0:0] CLBLM_R_X11Y128_SLICE_X14Y128_B4;
  wire [0:0] CLBLM_R_X11Y128_SLICE_X14Y128_B5;
  wire [0:0] CLBLM_R_X11Y128_SLICE_X14Y128_B6;
  wire [0:0] CLBLM_R_X11Y128_SLICE_X14Y128_BO5;
  wire [0:0] CLBLM_R_X11Y128_SLICE_X14Y128_BO6;
  wire [0:0] CLBLM_R_X11Y128_SLICE_X14Y128_B_CY;
  wire [0:0] CLBLM_R_X11Y128_SLICE_X14Y128_B_XOR;
  wire [0:0] CLBLM_R_X11Y128_SLICE_X14Y128_C;
  wire [0:0] CLBLM_R_X11Y128_SLICE_X14Y128_C1;
  wire [0:0] CLBLM_R_X11Y128_SLICE_X14Y128_C2;
  wire [0:0] CLBLM_R_X11Y128_SLICE_X14Y128_C3;
  wire [0:0] CLBLM_R_X11Y128_SLICE_X14Y128_C4;
  wire [0:0] CLBLM_R_X11Y128_SLICE_X14Y128_C5;
  wire [0:0] CLBLM_R_X11Y128_SLICE_X14Y128_C6;
  wire [0:0] CLBLM_R_X11Y128_SLICE_X14Y128_CO5;
  wire [0:0] CLBLM_R_X11Y128_SLICE_X14Y128_CO6;
  wire [0:0] CLBLM_R_X11Y128_SLICE_X14Y128_C_CY;
  wire [0:0] CLBLM_R_X11Y128_SLICE_X14Y128_C_XOR;
  wire [0:0] CLBLM_R_X11Y128_SLICE_X14Y128_D;
  wire [0:0] CLBLM_R_X11Y128_SLICE_X14Y128_D1;
  wire [0:0] CLBLM_R_X11Y128_SLICE_X14Y128_D2;
  wire [0:0] CLBLM_R_X11Y128_SLICE_X14Y128_D3;
  wire [0:0] CLBLM_R_X11Y128_SLICE_X14Y128_D4;
  wire [0:0] CLBLM_R_X11Y128_SLICE_X14Y128_D5;
  wire [0:0] CLBLM_R_X11Y128_SLICE_X14Y128_D6;
  wire [0:0] CLBLM_R_X11Y128_SLICE_X14Y128_DO5;
  wire [0:0] CLBLM_R_X11Y128_SLICE_X14Y128_DO6;
  wire [0:0] CLBLM_R_X11Y128_SLICE_X14Y128_D_CY;
  wire [0:0] CLBLM_R_X11Y128_SLICE_X14Y128_D_XOR;
  wire [0:0] CLBLM_R_X11Y128_SLICE_X15Y128_A;
  wire [0:0] CLBLM_R_X11Y128_SLICE_X15Y128_A1;
  wire [0:0] CLBLM_R_X11Y128_SLICE_X15Y128_A2;
  wire [0:0] CLBLM_R_X11Y128_SLICE_X15Y128_A3;
  wire [0:0] CLBLM_R_X11Y128_SLICE_X15Y128_A4;
  wire [0:0] CLBLM_R_X11Y128_SLICE_X15Y128_A5;
  wire [0:0] CLBLM_R_X11Y128_SLICE_X15Y128_A6;
  wire [0:0] CLBLM_R_X11Y128_SLICE_X15Y128_AO5;
  wire [0:0] CLBLM_R_X11Y128_SLICE_X15Y128_AO6;
  wire [0:0] CLBLM_R_X11Y128_SLICE_X15Y128_AQ;
  wire [0:0] CLBLM_R_X11Y128_SLICE_X15Y128_A_CY;
  wire [0:0] CLBLM_R_X11Y128_SLICE_X15Y128_A_XOR;
  wire [0:0] CLBLM_R_X11Y128_SLICE_X15Y128_B;
  wire [0:0] CLBLM_R_X11Y128_SLICE_X15Y128_B1;
  wire [0:0] CLBLM_R_X11Y128_SLICE_X15Y128_B2;
  wire [0:0] CLBLM_R_X11Y128_SLICE_X15Y128_B3;
  wire [0:0] CLBLM_R_X11Y128_SLICE_X15Y128_B4;
  wire [0:0] CLBLM_R_X11Y128_SLICE_X15Y128_B5;
  wire [0:0] CLBLM_R_X11Y128_SLICE_X15Y128_B6;
  wire [0:0] CLBLM_R_X11Y128_SLICE_X15Y128_BO5;
  wire [0:0] CLBLM_R_X11Y128_SLICE_X15Y128_BO6;
  wire [0:0] CLBLM_R_X11Y128_SLICE_X15Y128_B_CY;
  wire [0:0] CLBLM_R_X11Y128_SLICE_X15Y128_B_XOR;
  wire [0:0] CLBLM_R_X11Y128_SLICE_X15Y128_C;
  wire [0:0] CLBLM_R_X11Y128_SLICE_X15Y128_C1;
  wire [0:0] CLBLM_R_X11Y128_SLICE_X15Y128_C2;
  wire [0:0] CLBLM_R_X11Y128_SLICE_X15Y128_C3;
  wire [0:0] CLBLM_R_X11Y128_SLICE_X15Y128_C4;
  wire [0:0] CLBLM_R_X11Y128_SLICE_X15Y128_C5;
  wire [0:0] CLBLM_R_X11Y128_SLICE_X15Y128_C6;
  wire [0:0] CLBLM_R_X11Y128_SLICE_X15Y128_CLK;
  wire [0:0] CLBLM_R_X11Y128_SLICE_X15Y128_CO5;
  wire [0:0] CLBLM_R_X11Y128_SLICE_X15Y128_CO6;
  wire [0:0] CLBLM_R_X11Y128_SLICE_X15Y128_C_CY;
  wire [0:0] CLBLM_R_X11Y128_SLICE_X15Y128_C_XOR;
  wire [0:0] CLBLM_R_X11Y128_SLICE_X15Y128_D;
  wire [0:0] CLBLM_R_X11Y128_SLICE_X15Y128_D1;
  wire [0:0] CLBLM_R_X11Y128_SLICE_X15Y128_D2;
  wire [0:0] CLBLM_R_X11Y128_SLICE_X15Y128_D3;
  wire [0:0] CLBLM_R_X11Y128_SLICE_X15Y128_D4;
  wire [0:0] CLBLM_R_X11Y128_SLICE_X15Y128_D5;
  wire [0:0] CLBLM_R_X11Y128_SLICE_X15Y128_D6;
  wire [0:0] CLBLM_R_X11Y128_SLICE_X15Y128_DO5;
  wire [0:0] CLBLM_R_X11Y128_SLICE_X15Y128_DO6;
  wire [0:0] CLBLM_R_X11Y128_SLICE_X15Y128_D_CY;
  wire [0:0] CLBLM_R_X11Y128_SLICE_X15Y128_D_XOR;
  wire [0:0] CLBLM_R_X13Y119_SLICE_X18Y119_A;
  wire [0:0] CLBLM_R_X13Y119_SLICE_X18Y119_A1;
  wire [0:0] CLBLM_R_X13Y119_SLICE_X18Y119_A2;
  wire [0:0] CLBLM_R_X13Y119_SLICE_X18Y119_A3;
  wire [0:0] CLBLM_R_X13Y119_SLICE_X18Y119_A4;
  wire [0:0] CLBLM_R_X13Y119_SLICE_X18Y119_A5;
  wire [0:0] CLBLM_R_X13Y119_SLICE_X18Y119_A6;
  wire [0:0] CLBLM_R_X13Y119_SLICE_X18Y119_AO5;
  wire [0:0] CLBLM_R_X13Y119_SLICE_X18Y119_AO6;
  wire [0:0] CLBLM_R_X13Y119_SLICE_X18Y119_AQ;
  wire [0:0] CLBLM_R_X13Y119_SLICE_X18Y119_A_CY;
  wire [0:0] CLBLM_R_X13Y119_SLICE_X18Y119_A_XOR;
  wire [0:0] CLBLM_R_X13Y119_SLICE_X18Y119_B;
  wire [0:0] CLBLM_R_X13Y119_SLICE_X18Y119_B1;
  wire [0:0] CLBLM_R_X13Y119_SLICE_X18Y119_B2;
  wire [0:0] CLBLM_R_X13Y119_SLICE_X18Y119_B3;
  wire [0:0] CLBLM_R_X13Y119_SLICE_X18Y119_B4;
  wire [0:0] CLBLM_R_X13Y119_SLICE_X18Y119_B5;
  wire [0:0] CLBLM_R_X13Y119_SLICE_X18Y119_B6;
  wire [0:0] CLBLM_R_X13Y119_SLICE_X18Y119_BO5;
  wire [0:0] CLBLM_R_X13Y119_SLICE_X18Y119_BO6;
  wire [0:0] CLBLM_R_X13Y119_SLICE_X18Y119_BQ;
  wire [0:0] CLBLM_R_X13Y119_SLICE_X18Y119_B_CY;
  wire [0:0] CLBLM_R_X13Y119_SLICE_X18Y119_B_XOR;
  wire [0:0] CLBLM_R_X13Y119_SLICE_X18Y119_C;
  wire [0:0] CLBLM_R_X13Y119_SLICE_X18Y119_C1;
  wire [0:0] CLBLM_R_X13Y119_SLICE_X18Y119_C2;
  wire [0:0] CLBLM_R_X13Y119_SLICE_X18Y119_C3;
  wire [0:0] CLBLM_R_X13Y119_SLICE_X18Y119_C4;
  wire [0:0] CLBLM_R_X13Y119_SLICE_X18Y119_C5;
  wire [0:0] CLBLM_R_X13Y119_SLICE_X18Y119_C6;
  wire [0:0] CLBLM_R_X13Y119_SLICE_X18Y119_CLK;
  wire [0:0] CLBLM_R_X13Y119_SLICE_X18Y119_CO5;
  wire [0:0] CLBLM_R_X13Y119_SLICE_X18Y119_CO6;
  wire [0:0] CLBLM_R_X13Y119_SLICE_X18Y119_CQ;
  wire [0:0] CLBLM_R_X13Y119_SLICE_X18Y119_C_CY;
  wire [0:0] CLBLM_R_X13Y119_SLICE_X18Y119_C_XOR;
  wire [0:0] CLBLM_R_X13Y119_SLICE_X18Y119_D;
  wire [0:0] CLBLM_R_X13Y119_SLICE_X18Y119_D1;
  wire [0:0] CLBLM_R_X13Y119_SLICE_X18Y119_D2;
  wire [0:0] CLBLM_R_X13Y119_SLICE_X18Y119_D3;
  wire [0:0] CLBLM_R_X13Y119_SLICE_X18Y119_D4;
  wire [0:0] CLBLM_R_X13Y119_SLICE_X18Y119_D5;
  wire [0:0] CLBLM_R_X13Y119_SLICE_X18Y119_D6;
  wire [0:0] CLBLM_R_X13Y119_SLICE_X18Y119_DO5;
  wire [0:0] CLBLM_R_X13Y119_SLICE_X18Y119_DO6;
  wire [0:0] CLBLM_R_X13Y119_SLICE_X18Y119_D_CY;
  wire [0:0] CLBLM_R_X13Y119_SLICE_X18Y119_D_XOR;
  wire [0:0] CLBLM_R_X13Y119_SLICE_X19Y119_A;
  wire [0:0] CLBLM_R_X13Y119_SLICE_X19Y119_A1;
  wire [0:0] CLBLM_R_X13Y119_SLICE_X19Y119_A2;
  wire [0:0] CLBLM_R_X13Y119_SLICE_X19Y119_A3;
  wire [0:0] CLBLM_R_X13Y119_SLICE_X19Y119_A4;
  wire [0:0] CLBLM_R_X13Y119_SLICE_X19Y119_A5;
  wire [0:0] CLBLM_R_X13Y119_SLICE_X19Y119_A6;
  wire [0:0] CLBLM_R_X13Y119_SLICE_X19Y119_AO5;
  wire [0:0] CLBLM_R_X13Y119_SLICE_X19Y119_AO6;
  wire [0:0] CLBLM_R_X13Y119_SLICE_X19Y119_A_CY;
  wire [0:0] CLBLM_R_X13Y119_SLICE_X19Y119_A_XOR;
  wire [0:0] CLBLM_R_X13Y119_SLICE_X19Y119_B;
  wire [0:0] CLBLM_R_X13Y119_SLICE_X19Y119_B1;
  wire [0:0] CLBLM_R_X13Y119_SLICE_X19Y119_B2;
  wire [0:0] CLBLM_R_X13Y119_SLICE_X19Y119_B3;
  wire [0:0] CLBLM_R_X13Y119_SLICE_X19Y119_B4;
  wire [0:0] CLBLM_R_X13Y119_SLICE_X19Y119_B5;
  wire [0:0] CLBLM_R_X13Y119_SLICE_X19Y119_B6;
  wire [0:0] CLBLM_R_X13Y119_SLICE_X19Y119_BO5;
  wire [0:0] CLBLM_R_X13Y119_SLICE_X19Y119_BO6;
  wire [0:0] CLBLM_R_X13Y119_SLICE_X19Y119_B_CY;
  wire [0:0] CLBLM_R_X13Y119_SLICE_X19Y119_B_XOR;
  wire [0:0] CLBLM_R_X13Y119_SLICE_X19Y119_C;
  wire [0:0] CLBLM_R_X13Y119_SLICE_X19Y119_C1;
  wire [0:0] CLBLM_R_X13Y119_SLICE_X19Y119_C2;
  wire [0:0] CLBLM_R_X13Y119_SLICE_X19Y119_C3;
  wire [0:0] CLBLM_R_X13Y119_SLICE_X19Y119_C4;
  wire [0:0] CLBLM_R_X13Y119_SLICE_X19Y119_C5;
  wire [0:0] CLBLM_R_X13Y119_SLICE_X19Y119_C6;
  wire [0:0] CLBLM_R_X13Y119_SLICE_X19Y119_CO5;
  wire [0:0] CLBLM_R_X13Y119_SLICE_X19Y119_CO6;
  wire [0:0] CLBLM_R_X13Y119_SLICE_X19Y119_C_CY;
  wire [0:0] CLBLM_R_X13Y119_SLICE_X19Y119_C_XOR;
  wire [0:0] CLBLM_R_X13Y119_SLICE_X19Y119_D;
  wire [0:0] CLBLM_R_X13Y119_SLICE_X19Y119_D1;
  wire [0:0] CLBLM_R_X13Y119_SLICE_X19Y119_D2;
  wire [0:0] CLBLM_R_X13Y119_SLICE_X19Y119_D3;
  wire [0:0] CLBLM_R_X13Y119_SLICE_X19Y119_D4;
  wire [0:0] CLBLM_R_X13Y119_SLICE_X19Y119_D5;
  wire [0:0] CLBLM_R_X13Y119_SLICE_X19Y119_D6;
  wire [0:0] CLBLM_R_X13Y119_SLICE_X19Y119_DO5;
  wire [0:0] CLBLM_R_X13Y119_SLICE_X19Y119_DO6;
  wire [0:0] CLBLM_R_X13Y119_SLICE_X19Y119_D_CY;
  wire [0:0] CLBLM_R_X13Y119_SLICE_X19Y119_D_XOR;
  wire [0:0] CLBLM_R_X13Y120_SLICE_X18Y120_A;
  wire [0:0] CLBLM_R_X13Y120_SLICE_X18Y120_A1;
  wire [0:0] CLBLM_R_X13Y120_SLICE_X18Y120_A2;
  wire [0:0] CLBLM_R_X13Y120_SLICE_X18Y120_A3;
  wire [0:0] CLBLM_R_X13Y120_SLICE_X18Y120_A4;
  wire [0:0] CLBLM_R_X13Y120_SLICE_X18Y120_A5;
  wire [0:0] CLBLM_R_X13Y120_SLICE_X18Y120_A6;
  wire [0:0] CLBLM_R_X13Y120_SLICE_X18Y120_AO5;
  wire [0:0] CLBLM_R_X13Y120_SLICE_X18Y120_AO6;
  wire [0:0] CLBLM_R_X13Y120_SLICE_X18Y120_A_CY;
  wire [0:0] CLBLM_R_X13Y120_SLICE_X18Y120_A_XOR;
  wire [0:0] CLBLM_R_X13Y120_SLICE_X18Y120_B;
  wire [0:0] CLBLM_R_X13Y120_SLICE_X18Y120_B1;
  wire [0:0] CLBLM_R_X13Y120_SLICE_X18Y120_B2;
  wire [0:0] CLBLM_R_X13Y120_SLICE_X18Y120_B3;
  wire [0:0] CLBLM_R_X13Y120_SLICE_X18Y120_B4;
  wire [0:0] CLBLM_R_X13Y120_SLICE_X18Y120_B5;
  wire [0:0] CLBLM_R_X13Y120_SLICE_X18Y120_B6;
  wire [0:0] CLBLM_R_X13Y120_SLICE_X18Y120_BO5;
  wire [0:0] CLBLM_R_X13Y120_SLICE_X18Y120_BO6;
  wire [0:0] CLBLM_R_X13Y120_SLICE_X18Y120_B_CY;
  wire [0:0] CLBLM_R_X13Y120_SLICE_X18Y120_B_XOR;
  wire [0:0] CLBLM_R_X13Y120_SLICE_X18Y120_C;
  wire [0:0] CLBLM_R_X13Y120_SLICE_X18Y120_C1;
  wire [0:0] CLBLM_R_X13Y120_SLICE_X18Y120_C2;
  wire [0:0] CLBLM_R_X13Y120_SLICE_X18Y120_C3;
  wire [0:0] CLBLM_R_X13Y120_SLICE_X18Y120_C4;
  wire [0:0] CLBLM_R_X13Y120_SLICE_X18Y120_C5;
  wire [0:0] CLBLM_R_X13Y120_SLICE_X18Y120_C6;
  wire [0:0] CLBLM_R_X13Y120_SLICE_X18Y120_CO5;
  wire [0:0] CLBLM_R_X13Y120_SLICE_X18Y120_CO6;
  wire [0:0] CLBLM_R_X13Y120_SLICE_X18Y120_C_CY;
  wire [0:0] CLBLM_R_X13Y120_SLICE_X18Y120_C_XOR;
  wire [0:0] CLBLM_R_X13Y120_SLICE_X18Y120_D;
  wire [0:0] CLBLM_R_X13Y120_SLICE_X18Y120_D1;
  wire [0:0] CLBLM_R_X13Y120_SLICE_X18Y120_D2;
  wire [0:0] CLBLM_R_X13Y120_SLICE_X18Y120_D3;
  wire [0:0] CLBLM_R_X13Y120_SLICE_X18Y120_D4;
  wire [0:0] CLBLM_R_X13Y120_SLICE_X18Y120_D5;
  wire [0:0] CLBLM_R_X13Y120_SLICE_X18Y120_D6;
  wire [0:0] CLBLM_R_X13Y120_SLICE_X18Y120_DO5;
  wire [0:0] CLBLM_R_X13Y120_SLICE_X18Y120_DO6;
  wire [0:0] CLBLM_R_X13Y120_SLICE_X18Y120_D_CY;
  wire [0:0] CLBLM_R_X13Y120_SLICE_X18Y120_D_XOR;
  wire [0:0] CLBLM_R_X13Y120_SLICE_X19Y120_A;
  wire [0:0] CLBLM_R_X13Y120_SLICE_X19Y120_A1;
  wire [0:0] CLBLM_R_X13Y120_SLICE_X19Y120_A2;
  wire [0:0] CLBLM_R_X13Y120_SLICE_X19Y120_A3;
  wire [0:0] CLBLM_R_X13Y120_SLICE_X19Y120_A4;
  wire [0:0] CLBLM_R_X13Y120_SLICE_X19Y120_A5;
  wire [0:0] CLBLM_R_X13Y120_SLICE_X19Y120_A6;
  wire [0:0] CLBLM_R_X13Y120_SLICE_X19Y120_AO5;
  wire [0:0] CLBLM_R_X13Y120_SLICE_X19Y120_AO6;
  wire [0:0] CLBLM_R_X13Y120_SLICE_X19Y120_A_CY;
  wire [0:0] CLBLM_R_X13Y120_SLICE_X19Y120_A_XOR;
  wire [0:0] CLBLM_R_X13Y120_SLICE_X19Y120_B;
  wire [0:0] CLBLM_R_X13Y120_SLICE_X19Y120_B1;
  wire [0:0] CLBLM_R_X13Y120_SLICE_X19Y120_B2;
  wire [0:0] CLBLM_R_X13Y120_SLICE_X19Y120_B3;
  wire [0:0] CLBLM_R_X13Y120_SLICE_X19Y120_B4;
  wire [0:0] CLBLM_R_X13Y120_SLICE_X19Y120_B5;
  wire [0:0] CLBLM_R_X13Y120_SLICE_X19Y120_B6;
  wire [0:0] CLBLM_R_X13Y120_SLICE_X19Y120_BO5;
  wire [0:0] CLBLM_R_X13Y120_SLICE_X19Y120_BO6;
  wire [0:0] CLBLM_R_X13Y120_SLICE_X19Y120_B_CY;
  wire [0:0] CLBLM_R_X13Y120_SLICE_X19Y120_B_XOR;
  wire [0:0] CLBLM_R_X13Y120_SLICE_X19Y120_C;
  wire [0:0] CLBLM_R_X13Y120_SLICE_X19Y120_C1;
  wire [0:0] CLBLM_R_X13Y120_SLICE_X19Y120_C2;
  wire [0:0] CLBLM_R_X13Y120_SLICE_X19Y120_C3;
  wire [0:0] CLBLM_R_X13Y120_SLICE_X19Y120_C4;
  wire [0:0] CLBLM_R_X13Y120_SLICE_X19Y120_C5;
  wire [0:0] CLBLM_R_X13Y120_SLICE_X19Y120_C6;
  wire [0:0] CLBLM_R_X13Y120_SLICE_X19Y120_CO5;
  wire [0:0] CLBLM_R_X13Y120_SLICE_X19Y120_CO6;
  wire [0:0] CLBLM_R_X13Y120_SLICE_X19Y120_C_CY;
  wire [0:0] CLBLM_R_X13Y120_SLICE_X19Y120_C_XOR;
  wire [0:0] CLBLM_R_X13Y120_SLICE_X19Y120_D;
  wire [0:0] CLBLM_R_X13Y120_SLICE_X19Y120_D1;
  wire [0:0] CLBLM_R_X13Y120_SLICE_X19Y120_D2;
  wire [0:0] CLBLM_R_X13Y120_SLICE_X19Y120_D3;
  wire [0:0] CLBLM_R_X13Y120_SLICE_X19Y120_D4;
  wire [0:0] CLBLM_R_X13Y120_SLICE_X19Y120_D5;
  wire [0:0] CLBLM_R_X13Y120_SLICE_X19Y120_D6;
  wire [0:0] CLBLM_R_X13Y120_SLICE_X19Y120_DO5;
  wire [0:0] CLBLM_R_X13Y120_SLICE_X19Y120_DO6;
  wire [0:0] CLBLM_R_X13Y120_SLICE_X19Y120_D_CY;
  wire [0:0] CLBLM_R_X13Y120_SLICE_X19Y120_D_XOR;
  wire [0:0] CLBLM_R_X37Y119_SLICE_X56Y119_A;
  wire [0:0] CLBLM_R_X37Y119_SLICE_X56Y119_A1;
  wire [0:0] CLBLM_R_X37Y119_SLICE_X56Y119_A2;
  wire [0:0] CLBLM_R_X37Y119_SLICE_X56Y119_A3;
  wire [0:0] CLBLM_R_X37Y119_SLICE_X56Y119_A4;
  wire [0:0] CLBLM_R_X37Y119_SLICE_X56Y119_A5;
  wire [0:0] CLBLM_R_X37Y119_SLICE_X56Y119_A6;
  wire [0:0] CLBLM_R_X37Y119_SLICE_X56Y119_AO5;
  wire [0:0] CLBLM_R_X37Y119_SLICE_X56Y119_AO6;
  wire [0:0] CLBLM_R_X37Y119_SLICE_X56Y119_A_CY;
  wire [0:0] CLBLM_R_X37Y119_SLICE_X56Y119_A_XOR;
  wire [0:0] CLBLM_R_X37Y119_SLICE_X56Y119_B;
  wire [0:0] CLBLM_R_X37Y119_SLICE_X56Y119_B1;
  wire [0:0] CLBLM_R_X37Y119_SLICE_X56Y119_B2;
  wire [0:0] CLBLM_R_X37Y119_SLICE_X56Y119_B3;
  wire [0:0] CLBLM_R_X37Y119_SLICE_X56Y119_B4;
  wire [0:0] CLBLM_R_X37Y119_SLICE_X56Y119_B5;
  wire [0:0] CLBLM_R_X37Y119_SLICE_X56Y119_B6;
  wire [0:0] CLBLM_R_X37Y119_SLICE_X56Y119_BO5;
  wire [0:0] CLBLM_R_X37Y119_SLICE_X56Y119_BO6;
  wire [0:0] CLBLM_R_X37Y119_SLICE_X56Y119_B_CY;
  wire [0:0] CLBLM_R_X37Y119_SLICE_X56Y119_B_XOR;
  wire [0:0] CLBLM_R_X37Y119_SLICE_X56Y119_C;
  wire [0:0] CLBLM_R_X37Y119_SLICE_X56Y119_C1;
  wire [0:0] CLBLM_R_X37Y119_SLICE_X56Y119_C2;
  wire [0:0] CLBLM_R_X37Y119_SLICE_X56Y119_C3;
  wire [0:0] CLBLM_R_X37Y119_SLICE_X56Y119_C4;
  wire [0:0] CLBLM_R_X37Y119_SLICE_X56Y119_C5;
  wire [0:0] CLBLM_R_X37Y119_SLICE_X56Y119_C6;
  wire [0:0] CLBLM_R_X37Y119_SLICE_X56Y119_CO5;
  wire [0:0] CLBLM_R_X37Y119_SLICE_X56Y119_CO6;
  wire [0:0] CLBLM_R_X37Y119_SLICE_X56Y119_C_CY;
  wire [0:0] CLBLM_R_X37Y119_SLICE_X56Y119_C_XOR;
  wire [0:0] CLBLM_R_X37Y119_SLICE_X56Y119_D;
  wire [0:0] CLBLM_R_X37Y119_SLICE_X56Y119_D1;
  wire [0:0] CLBLM_R_X37Y119_SLICE_X56Y119_D2;
  wire [0:0] CLBLM_R_X37Y119_SLICE_X56Y119_D3;
  wire [0:0] CLBLM_R_X37Y119_SLICE_X56Y119_D4;
  wire [0:0] CLBLM_R_X37Y119_SLICE_X56Y119_D5;
  wire [0:0] CLBLM_R_X37Y119_SLICE_X56Y119_D6;
  wire [0:0] CLBLM_R_X37Y119_SLICE_X56Y119_DO5;
  wire [0:0] CLBLM_R_X37Y119_SLICE_X56Y119_DO6;
  wire [0:0] CLBLM_R_X37Y119_SLICE_X56Y119_D_CY;
  wire [0:0] CLBLM_R_X37Y119_SLICE_X56Y119_D_XOR;
  wire [0:0] CLBLM_R_X37Y119_SLICE_X57Y119_A;
  wire [0:0] CLBLM_R_X37Y119_SLICE_X57Y119_A1;
  wire [0:0] CLBLM_R_X37Y119_SLICE_X57Y119_A2;
  wire [0:0] CLBLM_R_X37Y119_SLICE_X57Y119_A3;
  wire [0:0] CLBLM_R_X37Y119_SLICE_X57Y119_A4;
  wire [0:0] CLBLM_R_X37Y119_SLICE_X57Y119_A5;
  wire [0:0] CLBLM_R_X37Y119_SLICE_X57Y119_A6;
  wire [0:0] CLBLM_R_X37Y119_SLICE_X57Y119_AO5;
  wire [0:0] CLBLM_R_X37Y119_SLICE_X57Y119_AO6;
  wire [0:0] CLBLM_R_X37Y119_SLICE_X57Y119_A_CY;
  wire [0:0] CLBLM_R_X37Y119_SLICE_X57Y119_A_XOR;
  wire [0:0] CLBLM_R_X37Y119_SLICE_X57Y119_B;
  wire [0:0] CLBLM_R_X37Y119_SLICE_X57Y119_B1;
  wire [0:0] CLBLM_R_X37Y119_SLICE_X57Y119_B2;
  wire [0:0] CLBLM_R_X37Y119_SLICE_X57Y119_B3;
  wire [0:0] CLBLM_R_X37Y119_SLICE_X57Y119_B4;
  wire [0:0] CLBLM_R_X37Y119_SLICE_X57Y119_B5;
  wire [0:0] CLBLM_R_X37Y119_SLICE_X57Y119_B6;
  wire [0:0] CLBLM_R_X37Y119_SLICE_X57Y119_BO5;
  wire [0:0] CLBLM_R_X37Y119_SLICE_X57Y119_BO6;
  wire [0:0] CLBLM_R_X37Y119_SLICE_X57Y119_B_CY;
  wire [0:0] CLBLM_R_X37Y119_SLICE_X57Y119_B_XOR;
  wire [0:0] CLBLM_R_X37Y119_SLICE_X57Y119_C;
  wire [0:0] CLBLM_R_X37Y119_SLICE_X57Y119_C1;
  wire [0:0] CLBLM_R_X37Y119_SLICE_X57Y119_C2;
  wire [0:0] CLBLM_R_X37Y119_SLICE_X57Y119_C3;
  wire [0:0] CLBLM_R_X37Y119_SLICE_X57Y119_C4;
  wire [0:0] CLBLM_R_X37Y119_SLICE_X57Y119_C5;
  wire [0:0] CLBLM_R_X37Y119_SLICE_X57Y119_C6;
  wire [0:0] CLBLM_R_X37Y119_SLICE_X57Y119_CO5;
  wire [0:0] CLBLM_R_X37Y119_SLICE_X57Y119_CO6;
  wire [0:0] CLBLM_R_X37Y119_SLICE_X57Y119_C_CY;
  wire [0:0] CLBLM_R_X37Y119_SLICE_X57Y119_C_XOR;
  wire [0:0] CLBLM_R_X37Y119_SLICE_X57Y119_D;
  wire [0:0] CLBLM_R_X37Y119_SLICE_X57Y119_D1;
  wire [0:0] CLBLM_R_X37Y119_SLICE_X57Y119_D2;
  wire [0:0] CLBLM_R_X37Y119_SLICE_X57Y119_D3;
  wire [0:0] CLBLM_R_X37Y119_SLICE_X57Y119_D4;
  wire [0:0] CLBLM_R_X37Y119_SLICE_X57Y119_D5;
  wire [0:0] CLBLM_R_X37Y119_SLICE_X57Y119_D6;
  wire [0:0] CLBLM_R_X37Y119_SLICE_X57Y119_DO5;
  wire [0:0] CLBLM_R_X37Y119_SLICE_X57Y119_DO6;
  wire [0:0] CLBLM_R_X37Y119_SLICE_X57Y119_D_CY;
  wire [0:0] CLBLM_R_X37Y119_SLICE_X57Y119_D_XOR;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X2Y110_A;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X2Y110_A1;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X2Y110_A2;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X2Y110_A3;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X2Y110_A4;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X2Y110_A5;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X2Y110_A6;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X2Y110_AO5;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X2Y110_AO6;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X2Y110_AQ;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X2Y110_AX;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X2Y110_A_CY;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X2Y110_A_XOR;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X2Y110_B;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X2Y110_B1;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X2Y110_B2;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X2Y110_B3;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X2Y110_B4;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X2Y110_B5;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X2Y110_B6;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X2Y110_BO5;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X2Y110_BO6;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X2Y110_B_CY;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X2Y110_B_XOR;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X2Y110_C;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X2Y110_C1;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X2Y110_C2;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X2Y110_C3;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X2Y110_C4;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X2Y110_C5;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X2Y110_C6;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X2Y110_CLK;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X2Y110_CO5;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X2Y110_CO6;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X2Y110_C_CY;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X2Y110_C_XOR;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X2Y110_D;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X2Y110_D1;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X2Y110_D2;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X2Y110_D3;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X2Y110_D4;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X2Y110_D5;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X2Y110_D6;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X2Y110_DO5;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X2Y110_DO6;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X2Y110_D_CY;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X2Y110_D_XOR;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X3Y110_A;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X3Y110_A1;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X3Y110_A2;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X3Y110_A3;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X3Y110_A4;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X3Y110_A5;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X3Y110_A6;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X3Y110_AO5;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X3Y110_AO6;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X3Y110_AQ;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X3Y110_A_CY;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X3Y110_A_XOR;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X3Y110_B;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X3Y110_B1;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X3Y110_B2;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X3Y110_B3;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X3Y110_B4;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X3Y110_B5;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X3Y110_B6;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X3Y110_BO5;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X3Y110_BO6;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X3Y110_BQ;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X3Y110_B_CY;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X3Y110_B_XOR;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X3Y110_C;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X3Y110_C1;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X3Y110_C2;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X3Y110_C3;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X3Y110_C4;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X3Y110_C5;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X3Y110_C6;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X3Y110_CLK;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X3Y110_CO5;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X3Y110_CO6;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X3Y110_C_CY;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X3Y110_C_XOR;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X3Y110_D;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X3Y110_D1;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X3Y110_D2;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X3Y110_D3;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X3Y110_D4;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X3Y110_D5;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X3Y110_D6;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X3Y110_DO5;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X3Y110_DO6;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X3Y110_D_CY;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X3Y110_D_XOR;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X2Y111_A;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X2Y111_A1;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X2Y111_A2;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X2Y111_A3;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X2Y111_A4;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X2Y111_A5;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X2Y111_A6;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X2Y111_AO5;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X2Y111_AO6;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X2Y111_AQ;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X2Y111_A_CY;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X2Y111_A_XOR;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X2Y111_B;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X2Y111_B1;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X2Y111_B2;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X2Y111_B3;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X2Y111_B4;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X2Y111_B5;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X2Y111_B6;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X2Y111_BMUX;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X2Y111_BO5;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X2Y111_BO6;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X2Y111_B_CY;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X2Y111_B_XOR;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X2Y111_C;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X2Y111_C1;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X2Y111_C2;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X2Y111_C3;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X2Y111_C4;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X2Y111_C5;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X2Y111_C6;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X2Y111_CLK;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X2Y111_CO5;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X2Y111_CO6;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X2Y111_C_CY;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X2Y111_C_XOR;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X2Y111_D;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X2Y111_D1;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X2Y111_D2;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X2Y111_D3;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X2Y111_D4;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X2Y111_D5;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X2Y111_D6;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X2Y111_DO5;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X2Y111_DO6;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X2Y111_D_CY;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X2Y111_D_XOR;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X3Y111_A;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X3Y111_A1;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X3Y111_A2;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X3Y111_A3;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X3Y111_A4;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X3Y111_A5;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X3Y111_A6;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X3Y111_AMUX;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X3Y111_AO5;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X3Y111_AO6;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X3Y111_AQ;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X3Y111_A_CY;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X3Y111_A_XOR;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X3Y111_B;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X3Y111_B1;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X3Y111_B2;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X3Y111_B3;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X3Y111_B4;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X3Y111_B5;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X3Y111_B6;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X3Y111_BO5;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X3Y111_BO6;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X3Y111_BQ;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X3Y111_B_CY;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X3Y111_B_XOR;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X3Y111_C;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X3Y111_C1;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X3Y111_C2;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X3Y111_C3;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X3Y111_C4;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X3Y111_C5;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X3Y111_C6;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X3Y111_CLK;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X3Y111_CMUX;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X3Y111_CO5;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X3Y111_CO6;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X3Y111_C_CY;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X3Y111_C_XOR;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X3Y111_D;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X3Y111_D1;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X3Y111_D2;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X3Y111_D3;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X3Y111_D4;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X3Y111_D5;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X3Y111_D6;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X3Y111_DO5;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X3Y111_DO6;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X3Y111_D_CY;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X3Y111_D_XOR;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X2Y112_A;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X2Y112_A1;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X2Y112_A2;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X2Y112_A3;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X2Y112_A4;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X2Y112_A5;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X2Y112_A6;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X2Y112_AO5;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X2Y112_AO6;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X2Y112_AQ;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X2Y112_A_CY;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X2Y112_A_XOR;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X2Y112_B;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X2Y112_B1;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X2Y112_B2;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X2Y112_B3;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X2Y112_B4;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X2Y112_B5;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X2Y112_B6;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X2Y112_BO5;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X2Y112_BO6;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X2Y112_BQ;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X2Y112_B_CY;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X2Y112_B_XOR;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X2Y112_C;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X2Y112_C1;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X2Y112_C2;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X2Y112_C3;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X2Y112_C4;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X2Y112_C5;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X2Y112_C6;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X2Y112_CLK;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X2Y112_CO5;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X2Y112_CO6;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X2Y112_C_CY;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X2Y112_C_XOR;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X2Y112_D;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X2Y112_D1;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X2Y112_D2;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X2Y112_D3;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X2Y112_D4;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X2Y112_D5;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X2Y112_D6;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X2Y112_DO5;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X2Y112_DO6;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X2Y112_D_CY;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X2Y112_D_XOR;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X3Y112_A;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X3Y112_A1;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X3Y112_A2;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X3Y112_A3;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X3Y112_A4;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X3Y112_A5;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X3Y112_A6;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X3Y112_AO5;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X3Y112_AO6;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X3Y112_AQ;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X3Y112_A_CY;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X3Y112_A_XOR;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X3Y112_B;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X3Y112_B1;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X3Y112_B2;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X3Y112_B3;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X3Y112_B4;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X3Y112_B5;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X3Y112_B5Q;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X3Y112_B6;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X3Y112_BMUX;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X3Y112_BO5;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X3Y112_BO6;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X3Y112_BQ;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X3Y112_B_CY;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X3Y112_B_XOR;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X3Y112_C;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X3Y112_C1;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X3Y112_C2;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X3Y112_C3;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X3Y112_C4;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X3Y112_C5;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X3Y112_C5Q;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X3Y112_C6;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X3Y112_CLK;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X3Y112_CMUX;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X3Y112_CO5;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X3Y112_CO6;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X3Y112_CQ;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X3Y112_C_CY;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X3Y112_C_XOR;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X3Y112_D;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X3Y112_D1;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X3Y112_D2;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X3Y112_D3;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X3Y112_D4;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X3Y112_D5;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X3Y112_D6;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X3Y112_DO5;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X3Y112_DO6;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X3Y112_D_CY;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X3Y112_D_XOR;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X2Y113_A;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X2Y113_A1;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X2Y113_A2;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X2Y113_A3;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X2Y113_A4;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X2Y113_A5;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X2Y113_A6;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X2Y113_AO5;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X2Y113_AO6;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X2Y113_AQ;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X2Y113_A_CY;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X2Y113_A_XOR;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X2Y113_B;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X2Y113_B1;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X2Y113_B2;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X2Y113_B3;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X2Y113_B4;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X2Y113_B5;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X2Y113_B6;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X2Y113_BO5;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X2Y113_BO6;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X2Y113_BQ;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X2Y113_B_CY;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X2Y113_B_XOR;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X2Y113_C;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X2Y113_C1;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X2Y113_C2;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X2Y113_C3;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X2Y113_C4;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X2Y113_C5;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X2Y113_C6;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X2Y113_CLK;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X2Y113_CMUX;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X2Y113_CO5;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X2Y113_CO6;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X2Y113_C_CY;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X2Y113_C_XOR;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X2Y113_D;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X2Y113_D1;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X2Y113_D2;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X2Y113_D3;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X2Y113_D4;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X2Y113_D5;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X2Y113_D6;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X2Y113_DMUX;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X2Y113_DO5;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X2Y113_DO6;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X2Y113_D_CY;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X2Y113_D_XOR;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X3Y113_A;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X3Y113_A1;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X3Y113_A2;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X3Y113_A3;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X3Y113_A4;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X3Y113_A5;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X3Y113_A6;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X3Y113_AO5;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X3Y113_AO6;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X3Y113_AQ;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X3Y113_A_CY;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X3Y113_A_XOR;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X3Y113_B;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X3Y113_B1;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X3Y113_B2;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X3Y113_B3;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X3Y113_B4;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X3Y113_B5;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X3Y113_B6;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X3Y113_BMUX;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X3Y113_BO5;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X3Y113_BO6;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X3Y113_B_CY;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X3Y113_B_XOR;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X3Y113_C;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X3Y113_C1;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X3Y113_C2;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X3Y113_C3;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X3Y113_C4;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X3Y113_C5;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X3Y113_C6;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X3Y113_CLK;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X3Y113_CO5;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X3Y113_CO6;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X3Y113_C_CY;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X3Y113_C_XOR;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X3Y113_D;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X3Y113_D1;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X3Y113_D2;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X3Y113_D3;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X3Y113_D4;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X3Y113_D5;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X3Y113_D6;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X3Y113_DO5;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X3Y113_DO6;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X3Y113_D_CY;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X3Y113_D_XOR;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X2Y114_A;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X2Y114_A1;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X2Y114_A2;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X2Y114_A3;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X2Y114_A4;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X2Y114_A5;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X2Y114_A6;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X2Y114_AMUX;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X2Y114_AO5;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X2Y114_AO6;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X2Y114_AQ;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X2Y114_A_CY;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X2Y114_A_XOR;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X2Y114_B;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X2Y114_B1;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X2Y114_B2;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X2Y114_B3;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X2Y114_B4;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X2Y114_B5;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X2Y114_B6;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X2Y114_BO5;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X2Y114_BO6;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X2Y114_BQ;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X2Y114_B_CY;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X2Y114_B_XOR;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X2Y114_C;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X2Y114_C1;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X2Y114_C2;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X2Y114_C3;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X2Y114_C4;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X2Y114_C5;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X2Y114_C6;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X2Y114_CLK;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X2Y114_CO5;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X2Y114_CO6;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X2Y114_CQ;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X2Y114_C_CY;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X2Y114_C_XOR;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X2Y114_D;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X2Y114_D1;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X2Y114_D2;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X2Y114_D3;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X2Y114_D4;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X2Y114_D5;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X2Y114_D6;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X2Y114_DO5;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X2Y114_DO6;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X2Y114_DQ;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X2Y114_D_CY;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X2Y114_D_XOR;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X3Y114_A;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X3Y114_A1;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X3Y114_A2;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X3Y114_A3;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X3Y114_A4;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X3Y114_A5;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X3Y114_A6;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X3Y114_AO5;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X3Y114_AO6;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X3Y114_AQ;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X3Y114_A_CY;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X3Y114_A_XOR;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X3Y114_B;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X3Y114_B1;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X3Y114_B2;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X3Y114_B3;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X3Y114_B4;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X3Y114_B5;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X3Y114_B6;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X3Y114_BO5;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X3Y114_BO6;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X3Y114_BQ;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X3Y114_B_CY;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X3Y114_B_XOR;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X3Y114_C;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X3Y114_C1;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X3Y114_C2;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X3Y114_C3;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X3Y114_C4;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X3Y114_C5;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X3Y114_C6;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X3Y114_CLK;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X3Y114_CO5;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X3Y114_CO6;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X3Y114_CQ;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X3Y114_C_CY;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X3Y114_C_XOR;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X3Y114_D;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X3Y114_D1;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X3Y114_D2;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X3Y114_D3;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X3Y114_D4;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X3Y114_D5;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X3Y114_D6;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X3Y114_DO5;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X3Y114_DO6;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X3Y114_D_CY;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X3Y114_D_XOR;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X2Y115_A;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X2Y115_A1;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X2Y115_A2;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X2Y115_A3;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X2Y115_A4;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X2Y115_A5;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X2Y115_A6;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X2Y115_AO5;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X2Y115_AO6;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X2Y115_AQ;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X2Y115_A_CY;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X2Y115_A_XOR;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X2Y115_B;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X2Y115_B1;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X2Y115_B2;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X2Y115_B3;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X2Y115_B4;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X2Y115_B5;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X2Y115_B6;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X2Y115_BO5;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X2Y115_BO6;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X2Y115_BQ;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X2Y115_B_CY;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X2Y115_B_XOR;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X2Y115_C;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X2Y115_C1;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X2Y115_C2;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X2Y115_C3;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X2Y115_C4;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X2Y115_C5;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X2Y115_C6;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X2Y115_CLK;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X2Y115_CO5;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X2Y115_CO6;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X2Y115_CQ;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X2Y115_C_CY;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X2Y115_C_XOR;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X2Y115_D;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X2Y115_D1;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X2Y115_D2;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X2Y115_D3;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X2Y115_D4;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X2Y115_D5;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X2Y115_D6;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X2Y115_DO5;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X2Y115_DO6;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X2Y115_DQ;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X2Y115_D_CY;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X2Y115_D_XOR;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X3Y115_A;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X3Y115_A1;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X3Y115_A2;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X3Y115_A3;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X3Y115_A4;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X3Y115_A5;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X3Y115_A6;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X3Y115_AO5;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X3Y115_AO6;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X3Y115_AQ;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X3Y115_A_CY;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X3Y115_A_XOR;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X3Y115_B;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X3Y115_B1;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X3Y115_B2;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X3Y115_B3;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X3Y115_B4;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X3Y115_B5;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X3Y115_B6;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X3Y115_BO5;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X3Y115_BO6;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X3Y115_BQ;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X3Y115_B_CY;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X3Y115_B_XOR;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X3Y115_C;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X3Y115_C1;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X3Y115_C2;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X3Y115_C3;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X3Y115_C4;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X3Y115_C5;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X3Y115_C6;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X3Y115_CLK;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X3Y115_CO5;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X3Y115_CO6;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X3Y115_CQ;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X3Y115_C_CY;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X3Y115_C_XOR;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X3Y115_D;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X3Y115_D1;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X3Y115_D2;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X3Y115_D3;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X3Y115_D4;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X3Y115_D5;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X3Y115_D6;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X3Y115_DO5;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X3Y115_DO6;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X3Y115_DQ;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X3Y115_D_CY;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X3Y115_D_XOR;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X2Y116_A;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X2Y116_A1;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X2Y116_A2;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X2Y116_A3;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X2Y116_A4;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X2Y116_A5;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X2Y116_A6;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X2Y116_AO5;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X2Y116_AO6;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X2Y116_AQ;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X2Y116_A_CY;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X2Y116_A_XOR;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X2Y116_B;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X2Y116_B1;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X2Y116_B2;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X2Y116_B3;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X2Y116_B4;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X2Y116_B5;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X2Y116_B6;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X2Y116_BO5;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X2Y116_BO6;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X2Y116_BQ;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X2Y116_B_CY;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X2Y116_B_XOR;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X2Y116_C;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X2Y116_C1;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X2Y116_C2;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X2Y116_C3;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X2Y116_C4;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X2Y116_C5;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X2Y116_C6;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X2Y116_CLK;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X2Y116_CO5;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X2Y116_CO6;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X2Y116_C_CY;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X2Y116_C_XOR;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X2Y116_D;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X2Y116_D1;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X2Y116_D2;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X2Y116_D3;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X2Y116_D4;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X2Y116_D5;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X2Y116_D6;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X2Y116_DO5;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X2Y116_DO6;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X2Y116_D_CY;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X2Y116_D_XOR;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X3Y116_A;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X3Y116_A1;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X3Y116_A2;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X3Y116_A3;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X3Y116_A4;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X3Y116_A5;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X3Y116_A5Q;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X3Y116_A6;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X3Y116_AMUX;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X3Y116_AO5;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X3Y116_AO6;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X3Y116_AQ;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X3Y116_AX;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X3Y116_A_CY;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X3Y116_A_XOR;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X3Y116_B;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X3Y116_B1;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X3Y116_B2;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X3Y116_B3;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X3Y116_B4;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X3Y116_B5;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X3Y116_B6;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X3Y116_BO5;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X3Y116_BO6;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X3Y116_BQ;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X3Y116_B_CY;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X3Y116_B_XOR;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X3Y116_C;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X3Y116_C1;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X3Y116_C2;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X3Y116_C3;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X3Y116_C4;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X3Y116_C5;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X3Y116_C6;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X3Y116_CLK;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X3Y116_CO5;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X3Y116_CO6;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X3Y116_CQ;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X3Y116_C_CY;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X3Y116_C_XOR;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X3Y116_D;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X3Y116_D1;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X3Y116_D2;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X3Y116_D3;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X3Y116_D4;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X3Y116_D5;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X3Y116_D6;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X3Y116_DO5;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X3Y116_DO6;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X3Y116_D_CY;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X3Y116_D_XOR;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X2Y117_A;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X2Y117_A1;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X2Y117_A2;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X2Y117_A3;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X2Y117_A4;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X2Y117_A5;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X2Y117_A6;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X2Y117_AO5;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X2Y117_AO6;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X2Y117_AQ;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X2Y117_A_CY;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X2Y117_A_XOR;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X2Y117_B;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X2Y117_B1;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X2Y117_B2;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X2Y117_B3;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X2Y117_B4;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X2Y117_B5;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X2Y117_B6;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X2Y117_BMUX;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X2Y117_BO5;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X2Y117_BO6;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X2Y117_B_CY;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X2Y117_B_XOR;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X2Y117_C;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X2Y117_C1;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X2Y117_C2;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X2Y117_C3;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X2Y117_C4;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X2Y117_C5;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X2Y117_C6;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X2Y117_CLK;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X2Y117_CO5;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X2Y117_CO6;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X2Y117_C_CY;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X2Y117_C_XOR;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X2Y117_D;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X2Y117_D1;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X2Y117_D2;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X2Y117_D3;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X2Y117_D4;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X2Y117_D5;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X2Y117_D6;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X2Y117_DO5;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X2Y117_DO6;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X2Y117_D_CY;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X2Y117_D_XOR;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X3Y117_A;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X3Y117_A1;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X3Y117_A2;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X3Y117_A3;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X3Y117_A4;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X3Y117_A5;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X3Y117_A5Q;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X3Y117_A6;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X3Y117_AMUX;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X3Y117_AO5;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X3Y117_AO6;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X3Y117_AQ;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X3Y117_A_CY;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X3Y117_A_XOR;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X3Y117_B;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X3Y117_B1;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X3Y117_B2;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X3Y117_B3;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X3Y117_B4;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X3Y117_B5;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X3Y117_B5Q;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X3Y117_B6;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X3Y117_BMUX;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X3Y117_BO5;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X3Y117_BO6;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X3Y117_BQ;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X3Y117_B_CY;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X3Y117_B_XOR;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X3Y117_C;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X3Y117_C1;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X3Y117_C2;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X3Y117_C3;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X3Y117_C4;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X3Y117_C5;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X3Y117_C5Q;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X3Y117_C6;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X3Y117_CLK;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X3Y117_CMUX;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X3Y117_CO5;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X3Y117_CO6;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X3Y117_CQ;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X3Y117_C_CY;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X3Y117_C_XOR;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X3Y117_D;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X3Y117_D1;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X3Y117_D2;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X3Y117_D3;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X3Y117_D4;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X3Y117_D5;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X3Y117_D6;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X3Y117_DO5;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X3Y117_DO6;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X3Y117_D_CY;
  wire [0:0] CLBLM_R_X3Y117_SLICE_X3Y117_D_XOR;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X2Y118_A;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X2Y118_A1;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X2Y118_A2;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X2Y118_A3;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X2Y118_A4;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X2Y118_A5;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X2Y118_A6;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X2Y118_AO5;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X2Y118_AO6;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X2Y118_AQ;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X2Y118_A_CY;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X2Y118_A_XOR;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X2Y118_B;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X2Y118_B1;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X2Y118_B2;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X2Y118_B3;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X2Y118_B4;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X2Y118_B5;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X2Y118_B6;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X2Y118_BO5;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X2Y118_BO6;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X2Y118_B_CY;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X2Y118_B_XOR;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X2Y118_C;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X2Y118_C1;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X2Y118_C2;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X2Y118_C3;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X2Y118_C4;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X2Y118_C5;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X2Y118_C6;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X2Y118_CLK;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X2Y118_CO5;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X2Y118_CO6;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X2Y118_C_CY;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X2Y118_C_XOR;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X2Y118_D;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X2Y118_D1;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X2Y118_D2;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X2Y118_D3;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X2Y118_D4;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X2Y118_D5;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X2Y118_D6;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X2Y118_DO5;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X2Y118_DO6;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X2Y118_D_CY;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X2Y118_D_XOR;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X3Y118_A;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X3Y118_A1;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X3Y118_A2;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X3Y118_A3;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X3Y118_A4;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X3Y118_A5;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X3Y118_A6;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X3Y118_AO5;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X3Y118_AO6;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X3Y118_AQ;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X3Y118_A_CY;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X3Y118_A_XOR;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X3Y118_B;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X3Y118_B1;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X3Y118_B2;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X3Y118_B3;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X3Y118_B4;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X3Y118_B5;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X3Y118_B6;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X3Y118_BO5;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X3Y118_BO6;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X3Y118_B_CY;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X3Y118_B_XOR;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X3Y118_C;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X3Y118_C1;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X3Y118_C2;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X3Y118_C3;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X3Y118_C4;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X3Y118_C5;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X3Y118_C6;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X3Y118_CLK;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X3Y118_CO5;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X3Y118_CO6;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X3Y118_C_CY;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X3Y118_C_XOR;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X3Y118_D;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X3Y118_D1;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X3Y118_D2;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X3Y118_D3;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X3Y118_D4;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X3Y118_D5;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X3Y118_D6;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X3Y118_DO5;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X3Y118_DO6;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X3Y118_D_CY;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X3Y118_D_XOR;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X2Y119_A;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X2Y119_A1;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X2Y119_A2;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X2Y119_A3;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X2Y119_A4;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X2Y119_A5;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X2Y119_A6;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X2Y119_AO5;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X2Y119_AO6;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X2Y119_A_CY;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X2Y119_A_XOR;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X2Y119_B;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X2Y119_B1;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X2Y119_B2;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X2Y119_B3;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X2Y119_B4;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X2Y119_B5;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X2Y119_B6;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X2Y119_BO5;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X2Y119_BO6;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X2Y119_B_CY;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X2Y119_B_XOR;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X2Y119_C;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X2Y119_C1;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X2Y119_C2;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X2Y119_C3;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X2Y119_C4;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X2Y119_C5;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X2Y119_C6;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X2Y119_CO5;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X2Y119_CO6;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X2Y119_C_CY;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X2Y119_C_XOR;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X2Y119_D;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X2Y119_D1;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X2Y119_D2;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X2Y119_D3;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X2Y119_D4;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X2Y119_D5;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X2Y119_D6;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X2Y119_DO5;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X2Y119_DO6;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X2Y119_D_CY;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X2Y119_D_XOR;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X3Y119_A;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X3Y119_A1;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X3Y119_A2;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X3Y119_A3;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X3Y119_A4;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X3Y119_A5;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X3Y119_A6;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X3Y119_AO5;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X3Y119_AO6;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X3Y119_AQ;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X3Y119_A_CY;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X3Y119_A_XOR;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X3Y119_B;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X3Y119_B1;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X3Y119_B2;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X3Y119_B3;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X3Y119_B4;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X3Y119_B5;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X3Y119_B6;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X3Y119_BO5;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X3Y119_BO6;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X3Y119_B_CY;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X3Y119_B_XOR;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X3Y119_C;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X3Y119_C1;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X3Y119_C2;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X3Y119_C3;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X3Y119_C4;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X3Y119_C5;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X3Y119_C6;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X3Y119_CLK;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X3Y119_CO5;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X3Y119_CO6;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X3Y119_C_CY;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X3Y119_C_XOR;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X3Y119_D;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X3Y119_D1;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X3Y119_D2;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X3Y119_D3;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X3Y119_D4;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X3Y119_D5;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X3Y119_D6;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X3Y119_DO5;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X3Y119_DO6;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X3Y119_D_CY;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X3Y119_D_XOR;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X2Y120_A;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X2Y120_A1;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X2Y120_A2;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X2Y120_A3;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X2Y120_A4;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X2Y120_A5;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X2Y120_A6;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X2Y120_AO5;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X2Y120_AO6;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X2Y120_A_CY;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X2Y120_A_XOR;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X2Y120_B;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X2Y120_B1;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X2Y120_B2;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X2Y120_B3;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X2Y120_B4;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X2Y120_B5;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X2Y120_B6;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X2Y120_BO5;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X2Y120_BO6;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X2Y120_B_CY;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X2Y120_B_XOR;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X2Y120_C;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X2Y120_C1;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X2Y120_C2;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X2Y120_C3;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X2Y120_C4;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X2Y120_C5;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X2Y120_C6;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X2Y120_CO5;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X2Y120_CO6;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X2Y120_C_CY;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X2Y120_C_XOR;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X2Y120_D;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X2Y120_D1;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X2Y120_D2;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X2Y120_D3;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X2Y120_D4;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X2Y120_D5;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X2Y120_D6;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X2Y120_DO5;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X2Y120_DO6;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X2Y120_D_CY;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X2Y120_D_XOR;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X3Y120_A;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X3Y120_A1;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X3Y120_A2;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X3Y120_A3;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X3Y120_A4;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X3Y120_A5;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X3Y120_A6;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X3Y120_AO5;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X3Y120_AO6;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X3Y120_A_CY;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X3Y120_A_XOR;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X3Y120_B;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X3Y120_B1;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X3Y120_B2;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X3Y120_B3;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X3Y120_B4;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X3Y120_B5;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X3Y120_B6;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X3Y120_BMUX;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X3Y120_BO5;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X3Y120_BO6;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X3Y120_B_CY;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X3Y120_B_XOR;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X3Y120_C;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X3Y120_C1;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X3Y120_C2;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X3Y120_C3;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X3Y120_C4;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X3Y120_C5;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X3Y120_C6;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X3Y120_CO5;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X3Y120_CO6;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X3Y120_C_CY;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X3Y120_C_XOR;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X3Y120_D;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X3Y120_D1;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X3Y120_D2;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X3Y120_D3;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X3Y120_D4;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X3Y120_D5;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X3Y120_D6;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X3Y120_DMUX;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X3Y120_DO5;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X3Y120_DO6;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X3Y120_D_CY;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X3Y120_D_XOR;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X2Y121_A;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X2Y121_A1;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X2Y121_A2;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X2Y121_A3;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X2Y121_A4;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X2Y121_A5;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X2Y121_A6;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X2Y121_AMUX;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X2Y121_AO5;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X2Y121_AO6;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X2Y121_A_CY;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X2Y121_A_XOR;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X2Y121_B;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X2Y121_B1;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X2Y121_B2;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X2Y121_B3;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X2Y121_B4;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X2Y121_B5;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X2Y121_B6;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X2Y121_BO5;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X2Y121_BO6;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X2Y121_B_CY;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X2Y121_B_XOR;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X2Y121_C;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X2Y121_C1;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X2Y121_C2;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X2Y121_C3;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X2Y121_C4;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X2Y121_C5;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X2Y121_C6;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X2Y121_CMUX;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X2Y121_CO5;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X2Y121_CO6;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X2Y121_C_CY;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X2Y121_C_XOR;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X2Y121_D;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X2Y121_D1;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X2Y121_D2;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X2Y121_D3;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X2Y121_D4;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X2Y121_D5;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X2Y121_D6;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X2Y121_DO5;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X2Y121_DO6;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X2Y121_D_CY;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X2Y121_D_XOR;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X3Y121_A;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X3Y121_A1;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X3Y121_A2;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X3Y121_A3;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X3Y121_A4;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X3Y121_A5;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X3Y121_A6;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X3Y121_AMUX;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X3Y121_AO5;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X3Y121_AO6;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X3Y121_A_CY;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X3Y121_A_XOR;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X3Y121_B;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X3Y121_B1;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X3Y121_B2;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X3Y121_B3;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X3Y121_B4;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X3Y121_B5;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X3Y121_B6;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X3Y121_BO5;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X3Y121_BO6;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X3Y121_B_CY;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X3Y121_B_XOR;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X3Y121_C;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X3Y121_C1;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X3Y121_C2;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X3Y121_C3;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X3Y121_C4;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X3Y121_C5;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X3Y121_C6;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X3Y121_CO5;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X3Y121_CO6;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X3Y121_C_CY;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X3Y121_C_XOR;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X3Y121_D;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X3Y121_D1;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X3Y121_D2;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X3Y121_D3;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X3Y121_D4;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X3Y121_D5;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X3Y121_D6;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X3Y121_DMUX;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X3Y121_DO5;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X3Y121_DO6;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X3Y121_D_CY;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X3Y121_D_XOR;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X2Y122_A;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X2Y122_A1;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X2Y122_A2;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X2Y122_A3;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X2Y122_A4;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X2Y122_A5;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X2Y122_A6;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X2Y122_AMUX;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X2Y122_AO5;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X2Y122_AO6;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X2Y122_A_CY;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X2Y122_A_XOR;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X2Y122_B;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X2Y122_B1;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X2Y122_B2;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X2Y122_B3;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X2Y122_B4;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X2Y122_B5;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X2Y122_B6;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X2Y122_BMUX;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X2Y122_BO5;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X2Y122_BO6;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X2Y122_B_CY;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X2Y122_B_XOR;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X2Y122_C;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X2Y122_C1;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X2Y122_C2;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X2Y122_C3;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X2Y122_C4;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X2Y122_C5;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X2Y122_C6;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X2Y122_CO5;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X2Y122_CO6;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X2Y122_C_CY;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X2Y122_C_XOR;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X2Y122_D;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X2Y122_D1;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X2Y122_D2;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X2Y122_D3;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X2Y122_D4;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X2Y122_D5;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X2Y122_D6;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X2Y122_DMUX;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X2Y122_DO5;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X2Y122_DO6;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X2Y122_D_CY;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X2Y122_D_XOR;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X3Y122_A;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X3Y122_A1;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X3Y122_A2;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X3Y122_A3;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X3Y122_A4;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X3Y122_A5;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X3Y122_A6;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X3Y122_AMUX;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X3Y122_AO5;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X3Y122_AO6;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X3Y122_A_CY;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X3Y122_A_XOR;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X3Y122_B;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X3Y122_B1;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X3Y122_B2;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X3Y122_B3;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X3Y122_B4;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X3Y122_B5;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X3Y122_B6;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X3Y122_BO5;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X3Y122_BO6;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X3Y122_B_CY;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X3Y122_B_XOR;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X3Y122_C;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X3Y122_C1;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X3Y122_C2;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X3Y122_C3;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X3Y122_C4;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X3Y122_C5;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X3Y122_C6;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X3Y122_CO5;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X3Y122_CO6;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X3Y122_C_CY;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X3Y122_C_XOR;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X3Y122_D;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X3Y122_D1;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X3Y122_D2;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X3Y122_D3;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X3Y122_D4;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X3Y122_D5;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X3Y122_D6;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X3Y122_DO5;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X3Y122_DO6;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X3Y122_D_CY;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X3Y122_D_XOR;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X2Y123_A;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X2Y123_A1;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X2Y123_A2;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X2Y123_A3;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X2Y123_A4;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X2Y123_A5;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X2Y123_A6;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X2Y123_AO5;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X2Y123_AO6;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X2Y123_A_CY;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X2Y123_A_XOR;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X2Y123_B;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X2Y123_B1;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X2Y123_B2;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X2Y123_B3;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X2Y123_B4;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X2Y123_B5;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X2Y123_B6;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X2Y123_BO5;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X2Y123_BO6;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X2Y123_B_CY;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X2Y123_B_XOR;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X2Y123_C;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X2Y123_C1;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X2Y123_C2;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X2Y123_C3;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X2Y123_C4;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X2Y123_C5;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X2Y123_C6;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X2Y123_CO5;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X2Y123_CO6;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X2Y123_C_CY;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X2Y123_C_XOR;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X2Y123_D;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X2Y123_D1;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X2Y123_D2;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X2Y123_D3;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X2Y123_D4;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X2Y123_D5;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X2Y123_D6;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X2Y123_DO5;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X2Y123_DO6;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X2Y123_D_CY;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X2Y123_D_XOR;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X3Y123_A;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X3Y123_A1;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X3Y123_A2;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X3Y123_A3;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X3Y123_A4;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X3Y123_A5;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X3Y123_A6;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X3Y123_AO5;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X3Y123_AO6;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X3Y123_AQ;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X3Y123_A_CY;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X3Y123_A_XOR;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X3Y123_B;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X3Y123_B1;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X3Y123_B2;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X3Y123_B3;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X3Y123_B4;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X3Y123_B5;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X3Y123_B6;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X3Y123_BMUX;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X3Y123_BO5;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X3Y123_BO6;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X3Y123_B_CY;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X3Y123_B_XOR;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X3Y123_C;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X3Y123_C1;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X3Y123_C2;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X3Y123_C3;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X3Y123_C4;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X3Y123_C5;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X3Y123_C6;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X3Y123_CLK;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X3Y123_CO5;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X3Y123_CO6;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X3Y123_C_CY;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X3Y123_C_XOR;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X3Y123_D;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X3Y123_D1;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X3Y123_D2;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X3Y123_D3;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X3Y123_D4;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X3Y123_D5;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X3Y123_D6;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X3Y123_DO5;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X3Y123_DO6;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X3Y123_D_CY;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X3Y123_D_XOR;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X2Y124_A;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X2Y124_A1;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X2Y124_A2;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X2Y124_A3;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X2Y124_A4;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X2Y124_A5;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X2Y124_A6;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X2Y124_AMUX;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X2Y124_AO5;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X2Y124_AO6;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X2Y124_A_CY;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X2Y124_A_XOR;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X2Y124_B;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X2Y124_B1;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X2Y124_B2;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X2Y124_B3;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X2Y124_B4;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X2Y124_B5;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X2Y124_B6;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X2Y124_BMUX;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X2Y124_BO5;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X2Y124_BO6;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X2Y124_B_CY;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X2Y124_B_XOR;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X2Y124_C;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X2Y124_C1;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X2Y124_C2;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X2Y124_C3;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X2Y124_C4;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X2Y124_C5;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X2Y124_C6;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X2Y124_CO5;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X2Y124_CO6;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X2Y124_C_CY;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X2Y124_C_XOR;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X2Y124_D;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X2Y124_D1;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X2Y124_D2;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X2Y124_D3;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X2Y124_D4;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X2Y124_D5;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X2Y124_D6;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X2Y124_DO5;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X2Y124_DO6;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X2Y124_D_CY;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X2Y124_D_XOR;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X3Y124_A;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X3Y124_A1;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X3Y124_A2;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X3Y124_A3;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X3Y124_A4;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X3Y124_A5;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X3Y124_A6;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X3Y124_AO5;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X3Y124_AO6;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X3Y124_A_CY;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X3Y124_A_XOR;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X3Y124_B;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X3Y124_B1;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X3Y124_B2;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X3Y124_B3;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X3Y124_B4;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X3Y124_B5;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X3Y124_B6;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X3Y124_BO5;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X3Y124_BO6;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X3Y124_B_CY;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X3Y124_B_XOR;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X3Y124_C;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X3Y124_C1;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X3Y124_C2;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X3Y124_C3;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X3Y124_C4;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X3Y124_C5;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X3Y124_C6;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X3Y124_CO5;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X3Y124_CO6;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X3Y124_C_CY;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X3Y124_C_XOR;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X3Y124_D;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X3Y124_D1;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X3Y124_D2;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X3Y124_D3;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X3Y124_D4;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X3Y124_D5;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X3Y124_D6;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X3Y124_DO5;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X3Y124_DO6;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X3Y124_D_CY;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X3Y124_D_XOR;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X6Y109_A;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X6Y109_A1;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X6Y109_A2;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X6Y109_A3;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X6Y109_A4;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X6Y109_A5;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X6Y109_A6;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X6Y109_AO5;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X6Y109_AO6;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X6Y109_AQ;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X6Y109_A_CY;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X6Y109_A_XOR;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X6Y109_B;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X6Y109_B1;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X6Y109_B2;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X6Y109_B3;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X6Y109_B4;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X6Y109_B5;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X6Y109_B6;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X6Y109_BO5;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X6Y109_BO6;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X6Y109_BQ;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X6Y109_B_CY;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X6Y109_B_XOR;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X6Y109_C;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X6Y109_C1;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X6Y109_C2;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X6Y109_C3;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X6Y109_C4;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X6Y109_C5;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X6Y109_C6;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X6Y109_CLK;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X6Y109_CO5;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X6Y109_CO6;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X6Y109_CQ;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X6Y109_C_CY;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X6Y109_C_XOR;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X6Y109_D;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X6Y109_D1;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X6Y109_D2;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X6Y109_D3;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X6Y109_D4;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X6Y109_D5;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X6Y109_D6;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X6Y109_DO5;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X6Y109_DO6;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X6Y109_D_CY;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X6Y109_D_XOR;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X7Y109_A;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X7Y109_A1;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X7Y109_A2;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X7Y109_A3;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X7Y109_A4;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X7Y109_A5;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X7Y109_A6;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X7Y109_AO5;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X7Y109_AO6;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X7Y109_AQ;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X7Y109_A_CY;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X7Y109_A_XOR;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X7Y109_B;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X7Y109_B1;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X7Y109_B2;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X7Y109_B3;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X7Y109_B4;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X7Y109_B5;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X7Y109_B6;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X7Y109_BO5;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X7Y109_BO6;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X7Y109_B_CY;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X7Y109_B_XOR;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X7Y109_C;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X7Y109_C1;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X7Y109_C2;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X7Y109_C3;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X7Y109_C4;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X7Y109_C5;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X7Y109_C6;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X7Y109_CLK;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X7Y109_CO5;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X7Y109_CO6;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X7Y109_C_CY;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X7Y109_C_XOR;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X7Y109_D;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X7Y109_D1;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X7Y109_D2;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X7Y109_D3;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X7Y109_D4;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X7Y109_D5;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X7Y109_D6;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X7Y109_DO5;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X7Y109_DO6;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X7Y109_D_CY;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X7Y109_D_XOR;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X6Y110_A;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X6Y110_A1;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X6Y110_A2;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X6Y110_A3;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X6Y110_A4;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X6Y110_A5;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X6Y110_A6;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X6Y110_AO5;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X6Y110_AO6;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X6Y110_AQ;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X6Y110_A_CY;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X6Y110_A_XOR;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X6Y110_B;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X6Y110_B1;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X6Y110_B2;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X6Y110_B3;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X6Y110_B4;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X6Y110_B5;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X6Y110_B6;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X6Y110_BO5;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X6Y110_BO6;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X6Y110_B_CY;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X6Y110_B_XOR;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X6Y110_C;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X6Y110_C1;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X6Y110_C2;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X6Y110_C3;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X6Y110_C4;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X6Y110_C5;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X6Y110_C6;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X6Y110_CLK;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X6Y110_CO5;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X6Y110_CO6;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X6Y110_C_CY;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X6Y110_C_XOR;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X6Y110_D;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X6Y110_D1;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X6Y110_D2;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X6Y110_D3;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X6Y110_D4;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X6Y110_D5;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X6Y110_D6;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X6Y110_DO5;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X6Y110_DO6;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X6Y110_D_CY;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X6Y110_D_XOR;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X7Y110_A;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X7Y110_A1;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X7Y110_A2;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X7Y110_A3;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X7Y110_A4;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X7Y110_A5;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X7Y110_A6;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X7Y110_AMUX;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X7Y110_AO5;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X7Y110_AO6;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X7Y110_AQ;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X7Y110_A_CY;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X7Y110_A_XOR;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X7Y110_B;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X7Y110_B1;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X7Y110_B2;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X7Y110_B3;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X7Y110_B4;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X7Y110_B5;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X7Y110_B6;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X7Y110_BO5;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X7Y110_BO6;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X7Y110_BQ;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X7Y110_B_CY;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X7Y110_B_XOR;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X7Y110_C;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X7Y110_C1;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X7Y110_C2;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X7Y110_C3;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X7Y110_C4;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X7Y110_C5;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X7Y110_C6;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X7Y110_CLK;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X7Y110_CO5;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X7Y110_CO6;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X7Y110_CQ;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X7Y110_C_CY;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X7Y110_C_XOR;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X7Y110_D;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X7Y110_D1;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X7Y110_D2;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X7Y110_D3;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X7Y110_D4;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X7Y110_D5;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X7Y110_D6;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X7Y110_DMUX;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X7Y110_DO5;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X7Y110_DO6;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X7Y110_D_CY;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X7Y110_D_XOR;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X6Y111_A;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X6Y111_A1;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X6Y111_A2;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X6Y111_A3;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X6Y111_A4;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X6Y111_A5;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X6Y111_A6;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X6Y111_AO5;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X6Y111_AO6;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X6Y111_AQ;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X6Y111_A_CY;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X6Y111_A_XOR;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X6Y111_B;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X6Y111_B1;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X6Y111_B2;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X6Y111_B3;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X6Y111_B4;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X6Y111_B5;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X6Y111_B6;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X6Y111_BO5;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X6Y111_BO6;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X6Y111_BQ;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X6Y111_B_CY;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X6Y111_B_XOR;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X6Y111_C;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X6Y111_C1;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X6Y111_C2;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X6Y111_C3;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X6Y111_C4;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X6Y111_C5;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X6Y111_C5Q;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X6Y111_C6;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X6Y111_CLK;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X6Y111_CMUX;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X6Y111_CO5;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X6Y111_CO6;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X6Y111_CQ;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X6Y111_C_CY;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X6Y111_C_XOR;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X6Y111_D;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X6Y111_D1;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X6Y111_D2;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X6Y111_D3;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X6Y111_D4;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X6Y111_D5;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X6Y111_D6;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X6Y111_DO5;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X6Y111_DO6;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X6Y111_D_CY;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X6Y111_D_XOR;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X7Y111_A;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X7Y111_A1;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X7Y111_A2;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X7Y111_A3;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X7Y111_A4;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X7Y111_A5;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X7Y111_A6;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X7Y111_AO5;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X7Y111_AO6;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X7Y111_AQ;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X7Y111_A_CY;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X7Y111_A_XOR;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X7Y111_B;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X7Y111_B1;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X7Y111_B2;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X7Y111_B3;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X7Y111_B4;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X7Y111_B5;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X7Y111_B6;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X7Y111_BO5;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X7Y111_BO6;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X7Y111_BQ;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X7Y111_B_CY;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X7Y111_B_XOR;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X7Y111_C;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X7Y111_C1;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X7Y111_C2;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X7Y111_C3;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X7Y111_C4;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X7Y111_C5;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X7Y111_C6;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X7Y111_CLK;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X7Y111_CMUX;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X7Y111_CO5;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X7Y111_CO6;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X7Y111_C_CY;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X7Y111_C_XOR;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X7Y111_D;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X7Y111_D1;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X7Y111_D2;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X7Y111_D3;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X7Y111_D4;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X7Y111_D5;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X7Y111_D6;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X7Y111_DO5;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X7Y111_DO6;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X7Y111_D_CY;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X7Y111_D_XOR;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X6Y112_A;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X6Y112_A1;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X6Y112_A2;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X6Y112_A3;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X6Y112_A4;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X6Y112_A5;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X6Y112_A6;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X6Y112_AO5;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X6Y112_AO6;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X6Y112_AQ;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X6Y112_A_CY;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X6Y112_A_XOR;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X6Y112_B;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X6Y112_B1;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X6Y112_B2;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X6Y112_B3;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X6Y112_B4;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X6Y112_B5;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X6Y112_B6;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X6Y112_BMUX;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X6Y112_BO5;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X6Y112_BO6;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X6Y112_B_CY;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X6Y112_B_XOR;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X6Y112_C;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X6Y112_C1;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X6Y112_C2;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X6Y112_C3;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X6Y112_C4;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X6Y112_C5;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X6Y112_C6;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X6Y112_CLK;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X6Y112_CO5;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X6Y112_CO6;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X6Y112_C_CY;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X6Y112_C_XOR;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X6Y112_D;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X6Y112_D1;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X6Y112_D2;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X6Y112_D3;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X6Y112_D4;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X6Y112_D5;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X6Y112_D6;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X6Y112_DO5;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X6Y112_DO6;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X6Y112_D_CY;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X6Y112_D_XOR;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X7Y112_A;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X7Y112_A1;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X7Y112_A2;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X7Y112_A3;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X7Y112_A4;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X7Y112_A5;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X7Y112_A6;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X7Y112_AMUX;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X7Y112_AO5;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X7Y112_AO6;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X7Y112_A_CY;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X7Y112_A_XOR;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X7Y112_B;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X7Y112_B1;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X7Y112_B2;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X7Y112_B3;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X7Y112_B4;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X7Y112_B5;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X7Y112_B6;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X7Y112_BO5;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X7Y112_BO6;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X7Y112_B_CY;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X7Y112_B_XOR;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X7Y112_C;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X7Y112_C1;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X7Y112_C2;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X7Y112_C3;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X7Y112_C4;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X7Y112_C5;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X7Y112_C6;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X7Y112_CO5;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X7Y112_CO6;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X7Y112_C_CY;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X7Y112_C_XOR;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X7Y112_D;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X7Y112_D1;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X7Y112_D2;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X7Y112_D3;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X7Y112_D4;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X7Y112_D5;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X7Y112_D6;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X7Y112_DO5;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X7Y112_DO6;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X7Y112_D_CY;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X7Y112_D_XOR;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X6Y113_A;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X6Y113_A1;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X6Y113_A2;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X6Y113_A3;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X6Y113_A4;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X6Y113_A5;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X6Y113_A6;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X6Y113_AO5;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X6Y113_AO6;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X6Y113_AQ;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X6Y113_A_CY;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X6Y113_A_XOR;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X6Y113_B;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X6Y113_B1;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X6Y113_B2;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X6Y113_B3;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X6Y113_B4;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X6Y113_B5;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X6Y113_B6;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X6Y113_BO5;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X6Y113_BO6;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X6Y113_BQ;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X6Y113_B_CY;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X6Y113_B_XOR;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X6Y113_C;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X6Y113_C1;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X6Y113_C2;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X6Y113_C3;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X6Y113_C4;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X6Y113_C5;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X6Y113_C6;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X6Y113_CLK;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X6Y113_CO5;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X6Y113_CO6;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X6Y113_CQ;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X6Y113_C_CY;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X6Y113_C_XOR;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X6Y113_D;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X6Y113_D1;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X6Y113_D2;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X6Y113_D3;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X6Y113_D4;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X6Y113_D5;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X6Y113_D6;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X6Y113_DMUX;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X6Y113_DO5;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X6Y113_DO6;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X6Y113_D_CY;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X6Y113_D_XOR;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X7Y113_A;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X7Y113_A1;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X7Y113_A2;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X7Y113_A3;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X7Y113_A4;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X7Y113_A5;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X7Y113_A5Q;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X7Y113_A6;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X7Y113_AMUX;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X7Y113_AO5;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X7Y113_AO6;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X7Y113_AQ;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X7Y113_A_CY;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X7Y113_A_XOR;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X7Y113_B;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X7Y113_B1;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X7Y113_B2;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X7Y113_B3;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X7Y113_B4;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X7Y113_B5;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X7Y113_B6;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X7Y113_BMUX;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X7Y113_BO5;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X7Y113_BO6;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X7Y113_B_CY;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X7Y113_B_XOR;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X7Y113_C;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X7Y113_C1;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X7Y113_C2;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X7Y113_C3;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X7Y113_C4;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X7Y113_C5;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X7Y113_C6;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X7Y113_CLK;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X7Y113_CO5;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X7Y113_CO6;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X7Y113_C_CY;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X7Y113_C_XOR;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X7Y113_D;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X7Y113_D1;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X7Y113_D2;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X7Y113_D3;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X7Y113_D4;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X7Y113_D5;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X7Y113_D6;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X7Y113_DO5;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X7Y113_DO6;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X7Y113_D_CY;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X7Y113_D_XOR;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X6Y114_A;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X6Y114_A1;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X6Y114_A2;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X6Y114_A3;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X6Y114_A4;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X6Y114_A5;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X6Y114_A6;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X6Y114_AO5;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X6Y114_AO6;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X6Y114_AQ;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X6Y114_A_CY;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X6Y114_A_XOR;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X6Y114_B;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X6Y114_B1;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X6Y114_B2;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X6Y114_B3;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X6Y114_B4;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X6Y114_B5;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X6Y114_B6;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X6Y114_BO5;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X6Y114_BO6;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X6Y114_BQ;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X6Y114_B_CY;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X6Y114_B_XOR;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X6Y114_C;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X6Y114_C1;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X6Y114_C2;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X6Y114_C3;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X6Y114_C4;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X6Y114_C5;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X6Y114_C6;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X6Y114_CLK;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X6Y114_CO5;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X6Y114_CO6;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X6Y114_CQ;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X6Y114_C_CY;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X6Y114_C_XOR;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X6Y114_D;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X6Y114_D1;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X6Y114_D2;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X6Y114_D3;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X6Y114_D4;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X6Y114_D5;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X6Y114_D6;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X6Y114_DO5;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X6Y114_DO6;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X6Y114_DQ;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X6Y114_D_CY;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X6Y114_D_XOR;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X7Y114_A;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X7Y114_A1;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X7Y114_A2;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X7Y114_A3;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X7Y114_A4;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X7Y114_A5;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X7Y114_A6;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X7Y114_AO5;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X7Y114_AO6;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X7Y114_AQ;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X7Y114_A_CY;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X7Y114_A_XOR;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X7Y114_B;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X7Y114_B1;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X7Y114_B2;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X7Y114_B3;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X7Y114_B4;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X7Y114_B5;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X7Y114_B6;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X7Y114_BMUX;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X7Y114_BO5;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X7Y114_BO6;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X7Y114_B_CY;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X7Y114_B_XOR;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X7Y114_C;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X7Y114_C1;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X7Y114_C2;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X7Y114_C3;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X7Y114_C4;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X7Y114_C5;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X7Y114_C6;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X7Y114_CLK;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X7Y114_CO5;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X7Y114_CO6;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X7Y114_C_CY;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X7Y114_C_XOR;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X7Y114_D;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X7Y114_D1;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X7Y114_D2;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X7Y114_D3;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X7Y114_D4;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X7Y114_D5;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X7Y114_D6;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X7Y114_DO5;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X7Y114_DO6;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X7Y114_D_CY;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X7Y114_D_XOR;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X6Y115_A;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X6Y115_A1;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X6Y115_A2;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X6Y115_A3;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X6Y115_A4;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X6Y115_A5;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X6Y115_A6;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X6Y115_AO5;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X6Y115_AO6;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X6Y115_AQ;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X6Y115_A_CY;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X6Y115_A_XOR;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X6Y115_B;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X6Y115_B1;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X6Y115_B2;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X6Y115_B3;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X6Y115_B4;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X6Y115_B5;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X6Y115_B6;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X6Y115_BO5;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X6Y115_BO6;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X6Y115_BQ;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X6Y115_B_CY;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X6Y115_B_XOR;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X6Y115_C;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X6Y115_C1;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X6Y115_C2;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X6Y115_C3;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X6Y115_C4;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X6Y115_C5;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X6Y115_C6;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X6Y115_CLK;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X6Y115_CMUX;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X6Y115_CO5;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X6Y115_CO6;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X6Y115_C_CY;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X6Y115_C_XOR;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X6Y115_D;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X6Y115_D1;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X6Y115_D2;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X6Y115_D3;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X6Y115_D4;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X6Y115_D5;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X6Y115_D6;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X6Y115_DO5;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X6Y115_DO6;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X6Y115_D_CY;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X6Y115_D_XOR;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X7Y115_A;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X7Y115_A1;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X7Y115_A2;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X7Y115_A3;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X7Y115_A4;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X7Y115_A5;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X7Y115_A5Q;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X7Y115_A6;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X7Y115_AMUX;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X7Y115_AO5;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X7Y115_AO6;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X7Y115_AQ;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X7Y115_A_CY;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X7Y115_A_XOR;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X7Y115_B;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X7Y115_B1;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X7Y115_B2;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X7Y115_B3;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X7Y115_B4;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X7Y115_B5;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X7Y115_B6;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X7Y115_BO5;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X7Y115_BO6;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X7Y115_BQ;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X7Y115_B_CY;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X7Y115_B_XOR;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X7Y115_C;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X7Y115_C1;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X7Y115_C2;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X7Y115_C3;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X7Y115_C4;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X7Y115_C5;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X7Y115_C6;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X7Y115_CLK;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X7Y115_CMUX;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X7Y115_CO5;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X7Y115_CO6;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X7Y115_C_CY;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X7Y115_C_XOR;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X7Y115_D;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X7Y115_D1;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X7Y115_D2;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X7Y115_D3;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X7Y115_D4;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X7Y115_D5;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X7Y115_D6;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X7Y115_DO5;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X7Y115_DO6;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X7Y115_D_CY;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X7Y115_D_XOR;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X6Y116_A;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X6Y116_A1;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X6Y116_A2;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X6Y116_A3;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X6Y116_A4;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X6Y116_A5;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X6Y116_A5Q;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X6Y116_A6;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X6Y116_AMUX;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X6Y116_AO5;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X6Y116_AO6;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X6Y116_AQ;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X6Y116_AX;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X6Y116_A_CY;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X6Y116_A_XOR;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X6Y116_B;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X6Y116_B1;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X6Y116_B2;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X6Y116_B3;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X6Y116_B4;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X6Y116_B5;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X6Y116_B6;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X6Y116_BO5;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X6Y116_BO6;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X6Y116_BQ;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X6Y116_B_CY;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X6Y116_B_XOR;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X6Y116_C;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X6Y116_C1;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X6Y116_C2;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X6Y116_C3;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X6Y116_C4;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X6Y116_C5;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X6Y116_C6;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X6Y116_CLK;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X6Y116_CMUX;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X6Y116_CO5;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X6Y116_CO6;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X6Y116_C_CY;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X6Y116_C_XOR;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X6Y116_D;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X6Y116_D1;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X6Y116_D2;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X6Y116_D3;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X6Y116_D4;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X6Y116_D5;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X6Y116_D6;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X6Y116_DO5;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X6Y116_DO6;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X6Y116_DQ;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X6Y116_D_CY;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X6Y116_D_XOR;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X7Y116_A;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X7Y116_A1;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X7Y116_A2;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X7Y116_A3;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X7Y116_A4;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X7Y116_A5;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X7Y116_A5Q;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X7Y116_A6;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X7Y116_AMUX;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X7Y116_AO5;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X7Y116_AO6;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X7Y116_AQ;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X7Y116_AX;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X7Y116_A_CY;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X7Y116_A_XOR;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X7Y116_B;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X7Y116_B1;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X7Y116_B2;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X7Y116_B3;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X7Y116_B4;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X7Y116_B5;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X7Y116_B6;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X7Y116_BMUX;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X7Y116_BO5;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X7Y116_BO6;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X7Y116_B_CY;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X7Y116_B_XOR;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X7Y116_C;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X7Y116_C1;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X7Y116_C2;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X7Y116_C3;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X7Y116_C4;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X7Y116_C5;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X7Y116_C6;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X7Y116_CLK;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X7Y116_CO5;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X7Y116_CO6;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X7Y116_CQ;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X7Y116_C_CY;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X7Y116_C_XOR;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X7Y116_D;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X7Y116_D1;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X7Y116_D2;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X7Y116_D3;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X7Y116_D4;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X7Y116_D5;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X7Y116_D6;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X7Y116_DO5;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X7Y116_DO6;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X7Y116_D_CY;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X7Y116_D_XOR;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X6Y117_A;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X6Y117_A1;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X6Y117_A2;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X6Y117_A3;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X6Y117_A4;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X6Y117_A5;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X6Y117_A6;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X6Y117_AO5;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X6Y117_AO6;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X6Y117_AQ;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X6Y117_A_CY;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X6Y117_A_XOR;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X6Y117_B;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X6Y117_B1;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X6Y117_B2;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X6Y117_B3;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X6Y117_B4;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X6Y117_B5;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X6Y117_B6;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X6Y117_BO5;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X6Y117_BO6;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X6Y117_BQ;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X6Y117_B_CY;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X6Y117_B_XOR;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X6Y117_C;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X6Y117_C1;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X6Y117_C2;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X6Y117_C3;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X6Y117_C4;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X6Y117_C5;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X6Y117_C6;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X6Y117_CLK;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X6Y117_CO5;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X6Y117_CO6;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X6Y117_CQ;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X6Y117_C_CY;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X6Y117_C_XOR;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X6Y117_D;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X6Y117_D1;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X6Y117_D2;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X6Y117_D3;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X6Y117_D4;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X6Y117_D5;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X6Y117_D5Q;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X6Y117_D6;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X6Y117_DMUX;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X6Y117_DO5;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X6Y117_DO6;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X6Y117_DQ;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X6Y117_D_CY;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X6Y117_D_XOR;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X7Y117_A;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X7Y117_A1;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X7Y117_A2;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X7Y117_A3;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X7Y117_A4;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X7Y117_A5;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X7Y117_A6;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X7Y117_AO5;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X7Y117_AO6;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X7Y117_AQ;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X7Y117_A_CY;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X7Y117_A_XOR;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X7Y117_B;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X7Y117_B1;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X7Y117_B2;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X7Y117_B3;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X7Y117_B4;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X7Y117_B5;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X7Y117_B6;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X7Y117_BO5;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X7Y117_BO6;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X7Y117_BQ;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X7Y117_B_CY;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X7Y117_B_XOR;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X7Y117_C;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X7Y117_C1;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X7Y117_C2;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X7Y117_C3;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X7Y117_C4;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X7Y117_C5;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X7Y117_C6;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X7Y117_CLK;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X7Y117_CO5;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X7Y117_CO6;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X7Y117_C_CY;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X7Y117_C_XOR;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X7Y117_D;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X7Y117_D1;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X7Y117_D2;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X7Y117_D3;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X7Y117_D4;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X7Y117_D5;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X7Y117_D6;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X7Y117_DO5;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X7Y117_DO6;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X7Y117_D_CY;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X7Y117_D_XOR;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X6Y118_A;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X6Y118_A1;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X6Y118_A2;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X6Y118_A3;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X6Y118_A4;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X6Y118_A5;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X6Y118_A6;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X6Y118_AO5;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X6Y118_AO6;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X6Y118_AQ;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X6Y118_A_CY;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X6Y118_A_XOR;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X6Y118_B;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X6Y118_B1;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X6Y118_B2;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X6Y118_B3;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X6Y118_B4;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X6Y118_B5;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X6Y118_B6;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X6Y118_BO5;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X6Y118_BO6;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X6Y118_BQ;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X6Y118_B_CY;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X6Y118_B_XOR;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X6Y118_C;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X6Y118_C1;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X6Y118_C2;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X6Y118_C3;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X6Y118_C4;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X6Y118_C5;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X6Y118_C6;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X6Y118_CLK;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X6Y118_CO5;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X6Y118_CO6;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X6Y118_CQ;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X6Y118_C_CY;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X6Y118_C_XOR;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X6Y118_D;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X6Y118_D1;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X6Y118_D2;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X6Y118_D3;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X6Y118_D4;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X6Y118_D5;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X6Y118_D6;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X6Y118_DO5;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X6Y118_DO6;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X6Y118_D_CY;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X6Y118_D_XOR;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X7Y118_A;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X7Y118_A1;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X7Y118_A2;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X7Y118_A3;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X7Y118_A4;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X7Y118_A5;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X7Y118_A6;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X7Y118_AO5;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X7Y118_AO6;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X7Y118_AQ;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X7Y118_A_CY;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X7Y118_A_XOR;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X7Y118_B;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X7Y118_B1;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X7Y118_B2;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X7Y118_B3;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X7Y118_B4;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X7Y118_B5;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X7Y118_B6;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X7Y118_BMUX;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X7Y118_BO5;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X7Y118_BO6;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X7Y118_B_CY;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X7Y118_B_XOR;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X7Y118_C;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X7Y118_C1;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X7Y118_C2;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X7Y118_C3;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X7Y118_C4;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X7Y118_C5;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X7Y118_C6;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X7Y118_CLK;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X7Y118_CO5;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X7Y118_CO6;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X7Y118_C_CY;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X7Y118_C_XOR;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X7Y118_D;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X7Y118_D1;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X7Y118_D2;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X7Y118_D3;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X7Y118_D4;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X7Y118_D5;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X7Y118_D6;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X7Y118_DO5;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X7Y118_DO6;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X7Y118_D_CY;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X7Y118_D_XOR;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X6Y119_A;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X6Y119_A1;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X6Y119_A2;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X6Y119_A3;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X6Y119_A4;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X6Y119_A5;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X6Y119_A6;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X6Y119_AO5;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X6Y119_AO6;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X6Y119_AQ;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X6Y119_A_CY;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X6Y119_A_XOR;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X6Y119_B;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X6Y119_B1;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X6Y119_B2;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X6Y119_B3;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X6Y119_B4;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X6Y119_B5;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X6Y119_B5Q;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X6Y119_B6;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X6Y119_BMUX;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X6Y119_BO5;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X6Y119_BO6;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X6Y119_BQ;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X6Y119_B_CY;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X6Y119_B_XOR;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X6Y119_C;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X6Y119_C1;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X6Y119_C2;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X6Y119_C3;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X6Y119_C4;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X6Y119_C5;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X6Y119_C6;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X6Y119_CLK;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X6Y119_CO5;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X6Y119_CO6;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X6Y119_CQ;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X6Y119_C_CY;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X6Y119_C_XOR;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X6Y119_D;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X6Y119_D1;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X6Y119_D2;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X6Y119_D3;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X6Y119_D4;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X6Y119_D5;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X6Y119_D6;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X6Y119_DO5;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X6Y119_DO6;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X6Y119_D_CY;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X6Y119_D_XOR;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X7Y119_A;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X7Y119_A1;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X7Y119_A2;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X7Y119_A3;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X7Y119_A4;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X7Y119_A5;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X7Y119_A6;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X7Y119_AO5;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X7Y119_AO6;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X7Y119_A_CY;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X7Y119_A_XOR;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X7Y119_B;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X7Y119_B1;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X7Y119_B2;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X7Y119_B3;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X7Y119_B4;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X7Y119_B5;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X7Y119_B6;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X7Y119_BO5;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X7Y119_BO6;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X7Y119_B_CY;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X7Y119_B_XOR;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X7Y119_C;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X7Y119_C1;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X7Y119_C2;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X7Y119_C3;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X7Y119_C4;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X7Y119_C5;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X7Y119_C6;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X7Y119_CO5;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X7Y119_CO6;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X7Y119_C_CY;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X7Y119_C_XOR;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X7Y119_D;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X7Y119_D1;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X7Y119_D2;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X7Y119_D3;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X7Y119_D4;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X7Y119_D5;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X7Y119_D6;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X7Y119_DO5;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X7Y119_DO6;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X7Y119_D_CY;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X7Y119_D_XOR;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X6Y120_A;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X6Y120_A1;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X6Y120_A2;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X6Y120_A3;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X6Y120_A4;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X6Y120_A5;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X6Y120_A5Q;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X6Y120_A6;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X6Y120_AMUX;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X6Y120_AO5;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X6Y120_AO6;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X6Y120_AQ;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X6Y120_A_CY;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X6Y120_A_XOR;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X6Y120_B;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X6Y120_B1;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X6Y120_B2;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X6Y120_B3;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X6Y120_B4;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X6Y120_B5;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X6Y120_B6;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X6Y120_BO5;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X6Y120_BO6;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X6Y120_BQ;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X6Y120_B_CY;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X6Y120_B_XOR;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X6Y120_C;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X6Y120_C1;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X6Y120_C2;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X6Y120_C3;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X6Y120_C4;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X6Y120_C5;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X6Y120_C6;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X6Y120_CLK;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X6Y120_CMUX;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X6Y120_CO5;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X6Y120_CO6;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X6Y120_C_CY;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X6Y120_C_XOR;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X6Y120_D;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X6Y120_D1;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X6Y120_D2;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X6Y120_D3;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X6Y120_D4;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X6Y120_D5;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X6Y120_D6;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X6Y120_DO5;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X6Y120_DO6;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X6Y120_D_CY;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X6Y120_D_XOR;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X7Y120_A;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X7Y120_A1;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X7Y120_A2;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X7Y120_A3;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X7Y120_A4;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X7Y120_A5;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X7Y120_A6;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X7Y120_AO5;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X7Y120_AO6;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X7Y120_AQ;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X7Y120_A_CY;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X7Y120_A_XOR;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X7Y120_B;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X7Y120_B1;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X7Y120_B2;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X7Y120_B3;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X7Y120_B4;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X7Y120_B5;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X7Y120_B6;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X7Y120_BO5;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X7Y120_BO6;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X7Y120_BQ;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X7Y120_B_CY;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X7Y120_B_XOR;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X7Y120_C;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X7Y120_C1;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X7Y120_C2;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X7Y120_C3;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X7Y120_C4;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X7Y120_C5;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X7Y120_C6;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X7Y120_CLK;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X7Y120_CO5;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X7Y120_CO6;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X7Y120_CQ;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X7Y120_C_CY;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X7Y120_C_XOR;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X7Y120_D;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X7Y120_D1;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X7Y120_D2;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X7Y120_D3;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X7Y120_D4;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X7Y120_D5;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X7Y120_D6;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X7Y120_DMUX;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X7Y120_DO5;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X7Y120_DO6;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X7Y120_D_CY;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X7Y120_D_XOR;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X6Y121_A;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X6Y121_A1;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X6Y121_A2;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X6Y121_A3;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X6Y121_A4;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X6Y121_A5;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X6Y121_A5Q;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X6Y121_A6;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X6Y121_AMUX;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X6Y121_AO5;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X6Y121_AO6;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X6Y121_AQ;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X6Y121_AX;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X6Y121_A_CY;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X6Y121_A_XOR;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X6Y121_B;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X6Y121_B1;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X6Y121_B2;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X6Y121_B3;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X6Y121_B4;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X6Y121_B5;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X6Y121_B5Q;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X6Y121_B6;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X6Y121_BMUX;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X6Y121_BO5;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X6Y121_BO6;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X6Y121_BQ;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X6Y121_BX;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X6Y121_B_CY;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X6Y121_B_XOR;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X6Y121_C;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X6Y121_C1;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X6Y121_C2;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X6Y121_C3;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X6Y121_C4;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X6Y121_C5;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X6Y121_C6;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X6Y121_CLK;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X6Y121_CMUX;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X6Y121_CO5;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X6Y121_CO6;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X6Y121_C_CY;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X6Y121_C_XOR;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X6Y121_D;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X6Y121_D1;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X6Y121_D2;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X6Y121_D3;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X6Y121_D4;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X6Y121_D5;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X6Y121_D6;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X6Y121_DO5;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X6Y121_DO6;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X6Y121_D_CY;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X6Y121_D_XOR;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X7Y121_A;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X7Y121_A1;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X7Y121_A2;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X7Y121_A3;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X7Y121_A4;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X7Y121_A5;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X7Y121_A5Q;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X7Y121_A6;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X7Y121_AMUX;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X7Y121_AO5;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X7Y121_AO6;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X7Y121_AQ;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X7Y121_A_CY;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X7Y121_A_XOR;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X7Y121_B;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X7Y121_B1;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X7Y121_B2;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X7Y121_B3;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X7Y121_B4;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X7Y121_B5;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X7Y121_B6;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X7Y121_BO5;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X7Y121_BO6;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X7Y121_B_CY;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X7Y121_B_XOR;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X7Y121_C;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X7Y121_C1;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X7Y121_C2;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X7Y121_C3;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X7Y121_C4;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X7Y121_C5;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X7Y121_C6;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X7Y121_CLK;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X7Y121_CO5;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X7Y121_CO6;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X7Y121_C_CY;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X7Y121_C_XOR;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X7Y121_D;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X7Y121_D1;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X7Y121_D2;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X7Y121_D3;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X7Y121_D4;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X7Y121_D5;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X7Y121_D6;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X7Y121_DO5;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X7Y121_DO6;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X7Y121_D_CY;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X7Y121_D_XOR;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X6Y122_A;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X6Y122_A1;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X6Y122_A2;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X6Y122_A3;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X6Y122_A4;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X6Y122_A5;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X6Y122_A6;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X6Y122_AMUX;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X6Y122_AO5;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X6Y122_AO6;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X6Y122_AQ;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X6Y122_A_CY;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X6Y122_A_XOR;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X6Y122_B;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X6Y122_B1;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X6Y122_B2;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X6Y122_B3;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X6Y122_B4;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X6Y122_B5;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X6Y122_B6;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X6Y122_BO5;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X6Y122_BO6;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X6Y122_BQ;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X6Y122_B_CY;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X6Y122_B_XOR;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X6Y122_C;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X6Y122_C1;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X6Y122_C2;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X6Y122_C3;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X6Y122_C4;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X6Y122_C5;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X6Y122_C6;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X6Y122_CLK;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X6Y122_CMUX;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X6Y122_CO5;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X6Y122_CO6;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X6Y122_C_CY;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X6Y122_C_XOR;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X6Y122_D;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X6Y122_D1;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X6Y122_D2;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X6Y122_D3;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X6Y122_D4;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X6Y122_D5;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X6Y122_D6;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X6Y122_DO5;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X6Y122_DO6;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X6Y122_D_CY;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X6Y122_D_XOR;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X7Y122_A;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X7Y122_A1;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X7Y122_A2;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X7Y122_A3;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X7Y122_A4;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X7Y122_A5;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X7Y122_A5Q;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X7Y122_A6;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X7Y122_AMUX;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X7Y122_AO5;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X7Y122_AO6;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X7Y122_AQ;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X7Y122_A_CY;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X7Y122_A_XOR;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X7Y122_B;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X7Y122_B1;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X7Y122_B2;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X7Y122_B3;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X7Y122_B4;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X7Y122_B5;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X7Y122_B6;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X7Y122_BO5;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X7Y122_BO6;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X7Y122_BQ;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X7Y122_B_CY;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X7Y122_B_XOR;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X7Y122_C;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X7Y122_C1;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X7Y122_C2;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X7Y122_C3;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X7Y122_C4;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X7Y122_C5;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X7Y122_C6;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X7Y122_CLK;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X7Y122_CO5;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X7Y122_CO6;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X7Y122_CQ;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X7Y122_C_CY;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X7Y122_C_XOR;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X7Y122_D;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X7Y122_D1;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X7Y122_D2;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X7Y122_D3;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X7Y122_D4;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X7Y122_D5;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X7Y122_D6;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X7Y122_DO5;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X7Y122_DO6;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X7Y122_DQ;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X7Y122_D_CY;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X7Y122_D_XOR;
  wire [0:0] CLBLM_R_X5Y123_SLICE_X6Y123_A;
  wire [0:0] CLBLM_R_X5Y123_SLICE_X6Y123_A1;
  wire [0:0] CLBLM_R_X5Y123_SLICE_X6Y123_A2;
  wire [0:0] CLBLM_R_X5Y123_SLICE_X6Y123_A3;
  wire [0:0] CLBLM_R_X5Y123_SLICE_X6Y123_A4;
  wire [0:0] CLBLM_R_X5Y123_SLICE_X6Y123_A5;
  wire [0:0] CLBLM_R_X5Y123_SLICE_X6Y123_A6;
  wire [0:0] CLBLM_R_X5Y123_SLICE_X6Y123_AO5;
  wire [0:0] CLBLM_R_X5Y123_SLICE_X6Y123_AO6;
  wire [0:0] CLBLM_R_X5Y123_SLICE_X6Y123_AQ;
  wire [0:0] CLBLM_R_X5Y123_SLICE_X6Y123_A_CY;
  wire [0:0] CLBLM_R_X5Y123_SLICE_X6Y123_A_XOR;
  wire [0:0] CLBLM_R_X5Y123_SLICE_X6Y123_B;
  wire [0:0] CLBLM_R_X5Y123_SLICE_X6Y123_B1;
  wire [0:0] CLBLM_R_X5Y123_SLICE_X6Y123_B2;
  wire [0:0] CLBLM_R_X5Y123_SLICE_X6Y123_B3;
  wire [0:0] CLBLM_R_X5Y123_SLICE_X6Y123_B4;
  wire [0:0] CLBLM_R_X5Y123_SLICE_X6Y123_B5;
  wire [0:0] CLBLM_R_X5Y123_SLICE_X6Y123_B6;
  wire [0:0] CLBLM_R_X5Y123_SLICE_X6Y123_BO5;
  wire [0:0] CLBLM_R_X5Y123_SLICE_X6Y123_BO6;
  wire [0:0] CLBLM_R_X5Y123_SLICE_X6Y123_BQ;
  wire [0:0] CLBLM_R_X5Y123_SLICE_X6Y123_B_CY;
  wire [0:0] CLBLM_R_X5Y123_SLICE_X6Y123_B_XOR;
  wire [0:0] CLBLM_R_X5Y123_SLICE_X6Y123_C;
  wire [0:0] CLBLM_R_X5Y123_SLICE_X6Y123_C1;
  wire [0:0] CLBLM_R_X5Y123_SLICE_X6Y123_C2;
  wire [0:0] CLBLM_R_X5Y123_SLICE_X6Y123_C3;
  wire [0:0] CLBLM_R_X5Y123_SLICE_X6Y123_C4;
  wire [0:0] CLBLM_R_X5Y123_SLICE_X6Y123_C5;
  wire [0:0] CLBLM_R_X5Y123_SLICE_X6Y123_C6;
  wire [0:0] CLBLM_R_X5Y123_SLICE_X6Y123_CLK;
  wire [0:0] CLBLM_R_X5Y123_SLICE_X6Y123_CO5;
  wire [0:0] CLBLM_R_X5Y123_SLICE_X6Y123_CO6;
  wire [0:0] CLBLM_R_X5Y123_SLICE_X6Y123_CQ;
  wire [0:0] CLBLM_R_X5Y123_SLICE_X6Y123_C_CY;
  wire [0:0] CLBLM_R_X5Y123_SLICE_X6Y123_C_XOR;
  wire [0:0] CLBLM_R_X5Y123_SLICE_X6Y123_D;
  wire [0:0] CLBLM_R_X5Y123_SLICE_X6Y123_D1;
  wire [0:0] CLBLM_R_X5Y123_SLICE_X6Y123_D2;
  wire [0:0] CLBLM_R_X5Y123_SLICE_X6Y123_D3;
  wire [0:0] CLBLM_R_X5Y123_SLICE_X6Y123_D4;
  wire [0:0] CLBLM_R_X5Y123_SLICE_X6Y123_D5;
  wire [0:0] CLBLM_R_X5Y123_SLICE_X6Y123_D6;
  wire [0:0] CLBLM_R_X5Y123_SLICE_X6Y123_DMUX;
  wire [0:0] CLBLM_R_X5Y123_SLICE_X6Y123_DO5;
  wire [0:0] CLBLM_R_X5Y123_SLICE_X6Y123_DO6;
  wire [0:0] CLBLM_R_X5Y123_SLICE_X6Y123_D_CY;
  wire [0:0] CLBLM_R_X5Y123_SLICE_X6Y123_D_XOR;
  wire [0:0] CLBLM_R_X5Y123_SLICE_X7Y123_A;
  wire [0:0] CLBLM_R_X5Y123_SLICE_X7Y123_A1;
  wire [0:0] CLBLM_R_X5Y123_SLICE_X7Y123_A2;
  wire [0:0] CLBLM_R_X5Y123_SLICE_X7Y123_A3;
  wire [0:0] CLBLM_R_X5Y123_SLICE_X7Y123_A4;
  wire [0:0] CLBLM_R_X5Y123_SLICE_X7Y123_A5;
  wire [0:0] CLBLM_R_X5Y123_SLICE_X7Y123_A6;
  wire [0:0] CLBLM_R_X5Y123_SLICE_X7Y123_AO5;
  wire [0:0] CLBLM_R_X5Y123_SLICE_X7Y123_AO6;
  wire [0:0] CLBLM_R_X5Y123_SLICE_X7Y123_AQ;
  wire [0:0] CLBLM_R_X5Y123_SLICE_X7Y123_A_CY;
  wire [0:0] CLBLM_R_X5Y123_SLICE_X7Y123_A_XOR;
  wire [0:0] CLBLM_R_X5Y123_SLICE_X7Y123_B;
  wire [0:0] CLBLM_R_X5Y123_SLICE_X7Y123_B1;
  wire [0:0] CLBLM_R_X5Y123_SLICE_X7Y123_B2;
  wire [0:0] CLBLM_R_X5Y123_SLICE_X7Y123_B3;
  wire [0:0] CLBLM_R_X5Y123_SLICE_X7Y123_B4;
  wire [0:0] CLBLM_R_X5Y123_SLICE_X7Y123_B5;
  wire [0:0] CLBLM_R_X5Y123_SLICE_X7Y123_B6;
  wire [0:0] CLBLM_R_X5Y123_SLICE_X7Y123_BO5;
  wire [0:0] CLBLM_R_X5Y123_SLICE_X7Y123_BO6;
  wire [0:0] CLBLM_R_X5Y123_SLICE_X7Y123_B_CY;
  wire [0:0] CLBLM_R_X5Y123_SLICE_X7Y123_B_XOR;
  wire [0:0] CLBLM_R_X5Y123_SLICE_X7Y123_C;
  wire [0:0] CLBLM_R_X5Y123_SLICE_X7Y123_C1;
  wire [0:0] CLBLM_R_X5Y123_SLICE_X7Y123_C2;
  wire [0:0] CLBLM_R_X5Y123_SLICE_X7Y123_C3;
  wire [0:0] CLBLM_R_X5Y123_SLICE_X7Y123_C4;
  wire [0:0] CLBLM_R_X5Y123_SLICE_X7Y123_C5;
  wire [0:0] CLBLM_R_X5Y123_SLICE_X7Y123_C6;
  wire [0:0] CLBLM_R_X5Y123_SLICE_X7Y123_CLK;
  wire [0:0] CLBLM_R_X5Y123_SLICE_X7Y123_CO5;
  wire [0:0] CLBLM_R_X5Y123_SLICE_X7Y123_CO6;
  wire [0:0] CLBLM_R_X5Y123_SLICE_X7Y123_C_CY;
  wire [0:0] CLBLM_R_X5Y123_SLICE_X7Y123_C_XOR;
  wire [0:0] CLBLM_R_X5Y123_SLICE_X7Y123_D;
  wire [0:0] CLBLM_R_X5Y123_SLICE_X7Y123_D1;
  wire [0:0] CLBLM_R_X5Y123_SLICE_X7Y123_D2;
  wire [0:0] CLBLM_R_X5Y123_SLICE_X7Y123_D3;
  wire [0:0] CLBLM_R_X5Y123_SLICE_X7Y123_D4;
  wire [0:0] CLBLM_R_X5Y123_SLICE_X7Y123_D5;
  wire [0:0] CLBLM_R_X5Y123_SLICE_X7Y123_D6;
  wire [0:0] CLBLM_R_X5Y123_SLICE_X7Y123_DO5;
  wire [0:0] CLBLM_R_X5Y123_SLICE_X7Y123_DO6;
  wire [0:0] CLBLM_R_X5Y123_SLICE_X7Y123_D_CY;
  wire [0:0] CLBLM_R_X5Y123_SLICE_X7Y123_D_XOR;
  wire [0:0] CLBLM_R_X5Y124_SLICE_X6Y124_A;
  wire [0:0] CLBLM_R_X5Y124_SLICE_X6Y124_A1;
  wire [0:0] CLBLM_R_X5Y124_SLICE_X6Y124_A2;
  wire [0:0] CLBLM_R_X5Y124_SLICE_X6Y124_A3;
  wire [0:0] CLBLM_R_X5Y124_SLICE_X6Y124_A4;
  wire [0:0] CLBLM_R_X5Y124_SLICE_X6Y124_A5;
  wire [0:0] CLBLM_R_X5Y124_SLICE_X6Y124_A6;
  wire [0:0] CLBLM_R_X5Y124_SLICE_X6Y124_AO5;
  wire [0:0] CLBLM_R_X5Y124_SLICE_X6Y124_AO6;
  wire [0:0] CLBLM_R_X5Y124_SLICE_X6Y124_AQ;
  wire [0:0] CLBLM_R_X5Y124_SLICE_X6Y124_A_CY;
  wire [0:0] CLBLM_R_X5Y124_SLICE_X6Y124_A_XOR;
  wire [0:0] CLBLM_R_X5Y124_SLICE_X6Y124_B;
  wire [0:0] CLBLM_R_X5Y124_SLICE_X6Y124_B1;
  wire [0:0] CLBLM_R_X5Y124_SLICE_X6Y124_B2;
  wire [0:0] CLBLM_R_X5Y124_SLICE_X6Y124_B3;
  wire [0:0] CLBLM_R_X5Y124_SLICE_X6Y124_B4;
  wire [0:0] CLBLM_R_X5Y124_SLICE_X6Y124_B5;
  wire [0:0] CLBLM_R_X5Y124_SLICE_X6Y124_B6;
  wire [0:0] CLBLM_R_X5Y124_SLICE_X6Y124_BO5;
  wire [0:0] CLBLM_R_X5Y124_SLICE_X6Y124_BO6;
  wire [0:0] CLBLM_R_X5Y124_SLICE_X6Y124_BQ;
  wire [0:0] CLBLM_R_X5Y124_SLICE_X6Y124_B_CY;
  wire [0:0] CLBLM_R_X5Y124_SLICE_X6Y124_B_XOR;
  wire [0:0] CLBLM_R_X5Y124_SLICE_X6Y124_C;
  wire [0:0] CLBLM_R_X5Y124_SLICE_X6Y124_C1;
  wire [0:0] CLBLM_R_X5Y124_SLICE_X6Y124_C2;
  wire [0:0] CLBLM_R_X5Y124_SLICE_X6Y124_C3;
  wire [0:0] CLBLM_R_X5Y124_SLICE_X6Y124_C4;
  wire [0:0] CLBLM_R_X5Y124_SLICE_X6Y124_C5;
  wire [0:0] CLBLM_R_X5Y124_SLICE_X6Y124_C6;
  wire [0:0] CLBLM_R_X5Y124_SLICE_X6Y124_CLK;
  wire [0:0] CLBLM_R_X5Y124_SLICE_X6Y124_CO5;
  wire [0:0] CLBLM_R_X5Y124_SLICE_X6Y124_CO6;
  wire [0:0] CLBLM_R_X5Y124_SLICE_X6Y124_CQ;
  wire [0:0] CLBLM_R_X5Y124_SLICE_X6Y124_C_CY;
  wire [0:0] CLBLM_R_X5Y124_SLICE_X6Y124_C_XOR;
  wire [0:0] CLBLM_R_X5Y124_SLICE_X6Y124_D;
  wire [0:0] CLBLM_R_X5Y124_SLICE_X6Y124_D1;
  wire [0:0] CLBLM_R_X5Y124_SLICE_X6Y124_D2;
  wire [0:0] CLBLM_R_X5Y124_SLICE_X6Y124_D3;
  wire [0:0] CLBLM_R_X5Y124_SLICE_X6Y124_D4;
  wire [0:0] CLBLM_R_X5Y124_SLICE_X6Y124_D5;
  wire [0:0] CLBLM_R_X5Y124_SLICE_X6Y124_D6;
  wire [0:0] CLBLM_R_X5Y124_SLICE_X6Y124_DO5;
  wire [0:0] CLBLM_R_X5Y124_SLICE_X6Y124_DO6;
  wire [0:0] CLBLM_R_X5Y124_SLICE_X6Y124_D_CY;
  wire [0:0] CLBLM_R_X5Y124_SLICE_X6Y124_D_XOR;
  wire [0:0] CLBLM_R_X5Y124_SLICE_X7Y124_A;
  wire [0:0] CLBLM_R_X5Y124_SLICE_X7Y124_A1;
  wire [0:0] CLBLM_R_X5Y124_SLICE_X7Y124_A2;
  wire [0:0] CLBLM_R_X5Y124_SLICE_X7Y124_A3;
  wire [0:0] CLBLM_R_X5Y124_SLICE_X7Y124_A4;
  wire [0:0] CLBLM_R_X5Y124_SLICE_X7Y124_A5;
  wire [0:0] CLBLM_R_X5Y124_SLICE_X7Y124_A6;
  wire [0:0] CLBLM_R_X5Y124_SLICE_X7Y124_AO5;
  wire [0:0] CLBLM_R_X5Y124_SLICE_X7Y124_AO6;
  wire [0:0] CLBLM_R_X5Y124_SLICE_X7Y124_A_CY;
  wire [0:0] CLBLM_R_X5Y124_SLICE_X7Y124_A_XOR;
  wire [0:0] CLBLM_R_X5Y124_SLICE_X7Y124_B;
  wire [0:0] CLBLM_R_X5Y124_SLICE_X7Y124_B1;
  wire [0:0] CLBLM_R_X5Y124_SLICE_X7Y124_B2;
  wire [0:0] CLBLM_R_X5Y124_SLICE_X7Y124_B3;
  wire [0:0] CLBLM_R_X5Y124_SLICE_X7Y124_B4;
  wire [0:0] CLBLM_R_X5Y124_SLICE_X7Y124_B5;
  wire [0:0] CLBLM_R_X5Y124_SLICE_X7Y124_B6;
  wire [0:0] CLBLM_R_X5Y124_SLICE_X7Y124_BO5;
  wire [0:0] CLBLM_R_X5Y124_SLICE_X7Y124_BO6;
  wire [0:0] CLBLM_R_X5Y124_SLICE_X7Y124_B_CY;
  wire [0:0] CLBLM_R_X5Y124_SLICE_X7Y124_B_XOR;
  wire [0:0] CLBLM_R_X5Y124_SLICE_X7Y124_C;
  wire [0:0] CLBLM_R_X5Y124_SLICE_X7Y124_C1;
  wire [0:0] CLBLM_R_X5Y124_SLICE_X7Y124_C2;
  wire [0:0] CLBLM_R_X5Y124_SLICE_X7Y124_C3;
  wire [0:0] CLBLM_R_X5Y124_SLICE_X7Y124_C4;
  wire [0:0] CLBLM_R_X5Y124_SLICE_X7Y124_C5;
  wire [0:0] CLBLM_R_X5Y124_SLICE_X7Y124_C6;
  wire [0:0] CLBLM_R_X5Y124_SLICE_X7Y124_CO5;
  wire [0:0] CLBLM_R_X5Y124_SLICE_X7Y124_CO6;
  wire [0:0] CLBLM_R_X5Y124_SLICE_X7Y124_C_CY;
  wire [0:0] CLBLM_R_X5Y124_SLICE_X7Y124_C_XOR;
  wire [0:0] CLBLM_R_X5Y124_SLICE_X7Y124_D;
  wire [0:0] CLBLM_R_X5Y124_SLICE_X7Y124_D1;
  wire [0:0] CLBLM_R_X5Y124_SLICE_X7Y124_D2;
  wire [0:0] CLBLM_R_X5Y124_SLICE_X7Y124_D3;
  wire [0:0] CLBLM_R_X5Y124_SLICE_X7Y124_D4;
  wire [0:0] CLBLM_R_X5Y124_SLICE_X7Y124_D5;
  wire [0:0] CLBLM_R_X5Y124_SLICE_X7Y124_D6;
  wire [0:0] CLBLM_R_X5Y124_SLICE_X7Y124_DO5;
  wire [0:0] CLBLM_R_X5Y124_SLICE_X7Y124_DO6;
  wire [0:0] CLBLM_R_X5Y124_SLICE_X7Y124_D_CY;
  wire [0:0] CLBLM_R_X5Y124_SLICE_X7Y124_D_XOR;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X6Y125_A;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X6Y125_A1;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X6Y125_A2;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X6Y125_A3;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X6Y125_A4;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X6Y125_A5;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X6Y125_A5Q;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X6Y125_A6;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X6Y125_AMUX;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X6Y125_AO5;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X6Y125_AO6;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X6Y125_AQ;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X6Y125_AX;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X6Y125_A_CY;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X6Y125_A_XOR;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X6Y125_B;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X6Y125_B1;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X6Y125_B2;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X6Y125_B3;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X6Y125_B4;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X6Y125_B5;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X6Y125_B6;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X6Y125_BMUX;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X6Y125_BO5;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X6Y125_BO6;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X6Y125_B_CY;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X6Y125_B_XOR;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X6Y125_C;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X6Y125_C1;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X6Y125_C2;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X6Y125_C3;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X6Y125_C4;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X6Y125_C5;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X6Y125_C6;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X6Y125_CLK;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X6Y125_CMUX;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X6Y125_CO5;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X6Y125_CO6;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X6Y125_C_CY;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X6Y125_C_XOR;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X6Y125_D;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X6Y125_D1;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X6Y125_D2;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X6Y125_D3;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X6Y125_D4;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X6Y125_D5;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X6Y125_D6;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X6Y125_DO5;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X6Y125_DO6;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X6Y125_D_CY;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X6Y125_D_XOR;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X7Y125_A;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X7Y125_A1;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X7Y125_A2;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X7Y125_A3;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X7Y125_A4;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X7Y125_A5;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X7Y125_A6;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X7Y125_AO5;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X7Y125_AO6;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X7Y125_A_CY;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X7Y125_A_XOR;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X7Y125_B;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X7Y125_B1;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X7Y125_B2;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X7Y125_B3;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X7Y125_B4;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X7Y125_B5;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X7Y125_B6;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X7Y125_BO5;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X7Y125_BO6;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X7Y125_B_CY;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X7Y125_B_XOR;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X7Y125_C;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X7Y125_C1;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X7Y125_C2;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X7Y125_C3;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X7Y125_C4;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X7Y125_C5;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X7Y125_C6;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X7Y125_CO5;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X7Y125_CO6;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X7Y125_C_CY;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X7Y125_C_XOR;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X7Y125_D;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X7Y125_D1;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X7Y125_D2;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X7Y125_D3;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X7Y125_D4;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X7Y125_D5;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X7Y125_D6;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X7Y125_DO5;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X7Y125_DO6;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X7Y125_D_CY;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X7Y125_D_XOR;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X8Y109_A;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X8Y109_A1;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X8Y109_A2;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X8Y109_A3;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X8Y109_A4;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X8Y109_A5;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X8Y109_A6;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X8Y109_AO5;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X8Y109_AO6;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X8Y109_AQ;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X8Y109_A_CY;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X8Y109_A_XOR;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X8Y109_B;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X8Y109_B1;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X8Y109_B2;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X8Y109_B3;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X8Y109_B4;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X8Y109_B5;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X8Y109_B6;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X8Y109_BO5;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X8Y109_BO6;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X8Y109_BQ;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X8Y109_B_CY;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X8Y109_B_XOR;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X8Y109_C;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X8Y109_C1;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X8Y109_C2;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X8Y109_C3;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X8Y109_C4;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X8Y109_C5;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X8Y109_C6;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X8Y109_CLK;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X8Y109_CO5;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X8Y109_CO6;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X8Y109_CQ;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X8Y109_C_CY;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X8Y109_C_XOR;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X8Y109_D;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X8Y109_D1;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X8Y109_D2;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X8Y109_D3;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X8Y109_D4;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X8Y109_D5;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X8Y109_D6;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X8Y109_DO5;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X8Y109_DO6;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X8Y109_D_CY;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X8Y109_D_XOR;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X9Y109_A;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X9Y109_A1;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X9Y109_A2;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X9Y109_A3;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X9Y109_A4;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X9Y109_A5;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X9Y109_A6;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X9Y109_AO5;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X9Y109_AO6;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X9Y109_A_CY;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X9Y109_A_XOR;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X9Y109_B;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X9Y109_B1;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X9Y109_B2;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X9Y109_B3;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X9Y109_B4;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X9Y109_B5;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X9Y109_B6;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X9Y109_BO5;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X9Y109_BO6;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X9Y109_B_CY;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X9Y109_B_XOR;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X9Y109_C;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X9Y109_C1;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X9Y109_C2;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X9Y109_C3;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X9Y109_C4;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X9Y109_C5;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X9Y109_C6;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X9Y109_CO5;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X9Y109_CO6;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X9Y109_C_CY;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X9Y109_C_XOR;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X9Y109_D;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X9Y109_D1;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X9Y109_D2;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X9Y109_D3;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X9Y109_D4;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X9Y109_D5;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X9Y109_D6;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X9Y109_DO5;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X9Y109_DO6;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X9Y109_D_CY;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X9Y109_D_XOR;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X8Y110_A;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X8Y110_A1;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X8Y110_A2;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X8Y110_A3;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X8Y110_A4;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X8Y110_A5;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X8Y110_A6;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X8Y110_AO5;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X8Y110_AO6;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X8Y110_AQ;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X8Y110_A_CY;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X8Y110_A_XOR;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X8Y110_B;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X8Y110_B1;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X8Y110_B2;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X8Y110_B3;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X8Y110_B4;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X8Y110_B5;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X8Y110_B6;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X8Y110_BO5;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X8Y110_BO6;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X8Y110_BQ;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X8Y110_B_CY;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X8Y110_B_XOR;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X8Y110_C;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X8Y110_C1;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X8Y110_C2;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X8Y110_C3;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X8Y110_C4;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X8Y110_C5;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X8Y110_C6;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X8Y110_CLK;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X8Y110_CO5;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X8Y110_CO6;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X8Y110_CQ;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X8Y110_C_CY;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X8Y110_C_XOR;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X8Y110_D;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X8Y110_D1;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X8Y110_D2;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X8Y110_D3;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X8Y110_D4;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X8Y110_D5;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X8Y110_D6;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X8Y110_DMUX;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X8Y110_DO5;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X8Y110_DO6;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X8Y110_D_CY;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X8Y110_D_XOR;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X9Y110_A;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X9Y110_A1;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X9Y110_A2;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X9Y110_A3;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X9Y110_A4;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X9Y110_A5;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X9Y110_A6;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X9Y110_AO5;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X9Y110_AO6;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X9Y110_AQ;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X9Y110_A_CY;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X9Y110_A_XOR;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X9Y110_B;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X9Y110_B1;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X9Y110_B2;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X9Y110_B3;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X9Y110_B4;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X9Y110_B5;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X9Y110_B6;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X9Y110_BO5;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X9Y110_BO6;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X9Y110_BQ;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X9Y110_B_CY;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X9Y110_B_XOR;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X9Y110_C;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X9Y110_C1;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X9Y110_C2;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X9Y110_C3;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X9Y110_C4;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X9Y110_C5;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X9Y110_C6;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X9Y110_CLK;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X9Y110_CO5;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X9Y110_CO6;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X9Y110_CQ;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X9Y110_C_CY;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X9Y110_C_XOR;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X9Y110_D;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X9Y110_D1;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X9Y110_D2;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X9Y110_D3;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X9Y110_D4;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X9Y110_D5;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X9Y110_D6;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X9Y110_DO5;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X9Y110_DO6;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X9Y110_D_CY;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X9Y110_D_XOR;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X8Y111_A;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X8Y111_A1;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X8Y111_A2;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X8Y111_A3;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X8Y111_A4;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X8Y111_A5;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X8Y111_A6;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X8Y111_AO5;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X8Y111_AO6;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X8Y111_AQ;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X8Y111_A_CY;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X8Y111_A_XOR;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X8Y111_B;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X8Y111_B1;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X8Y111_B2;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X8Y111_B3;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X8Y111_B4;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X8Y111_B5;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X8Y111_B6;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X8Y111_BO5;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X8Y111_BO6;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X8Y111_BQ;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X8Y111_B_CY;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X8Y111_B_XOR;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X8Y111_C;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X8Y111_C1;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X8Y111_C2;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X8Y111_C3;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X8Y111_C4;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X8Y111_C5;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X8Y111_C6;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X8Y111_CLK;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X8Y111_CO5;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X8Y111_CO6;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X8Y111_CQ;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X8Y111_C_CY;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X8Y111_C_XOR;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X8Y111_D;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X8Y111_D1;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X8Y111_D2;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X8Y111_D3;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X8Y111_D4;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X8Y111_D5;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X8Y111_D6;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X8Y111_DO5;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X8Y111_DO6;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X8Y111_D_CY;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X8Y111_D_XOR;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X9Y111_A;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X9Y111_A1;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X9Y111_A2;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X9Y111_A3;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X9Y111_A4;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X9Y111_A5;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X9Y111_A6;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X9Y111_AMUX;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X9Y111_AO5;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X9Y111_AO6;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X9Y111_A_CY;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X9Y111_A_XOR;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X9Y111_B;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X9Y111_B1;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X9Y111_B2;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X9Y111_B3;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X9Y111_B4;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X9Y111_B5;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X9Y111_B6;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X9Y111_BMUX;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X9Y111_BO5;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X9Y111_BO6;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X9Y111_B_CY;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X9Y111_B_XOR;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X9Y111_C;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X9Y111_C1;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X9Y111_C2;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X9Y111_C3;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X9Y111_C4;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X9Y111_C5;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X9Y111_C6;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X9Y111_CO5;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X9Y111_CO6;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X9Y111_C_CY;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X9Y111_C_XOR;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X9Y111_D;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X9Y111_D1;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X9Y111_D2;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X9Y111_D3;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X9Y111_D4;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X9Y111_D5;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X9Y111_D6;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X9Y111_DO5;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X9Y111_DO6;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X9Y111_D_CY;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X9Y111_D_XOR;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X8Y112_A;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X8Y112_A1;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X8Y112_A2;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X8Y112_A3;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X8Y112_A4;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X8Y112_A5;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X8Y112_A6;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X8Y112_AO5;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X8Y112_AO6;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X8Y112_AQ;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X8Y112_A_CY;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X8Y112_A_XOR;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X8Y112_B;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X8Y112_B1;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X8Y112_B2;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X8Y112_B3;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X8Y112_B4;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X8Y112_B5;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X8Y112_B6;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X8Y112_BO5;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X8Y112_BO6;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X8Y112_BQ;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X8Y112_B_CY;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X8Y112_B_XOR;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X8Y112_C;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X8Y112_C1;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X8Y112_C2;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X8Y112_C3;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X8Y112_C4;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X8Y112_C5;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X8Y112_C6;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X8Y112_CLK;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X8Y112_CO5;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X8Y112_CO6;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X8Y112_CQ;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X8Y112_C_CY;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X8Y112_C_XOR;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X8Y112_D;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X8Y112_D1;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X8Y112_D2;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X8Y112_D3;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X8Y112_D4;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X8Y112_D5;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X8Y112_D6;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X8Y112_DO5;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X8Y112_DO6;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X8Y112_D_CY;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X8Y112_D_XOR;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X9Y112_A;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X9Y112_A1;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X9Y112_A2;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X9Y112_A3;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X9Y112_A4;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X9Y112_A5;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X9Y112_A6;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X9Y112_AO5;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X9Y112_AO6;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X9Y112_AQ;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X9Y112_A_CY;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X9Y112_A_XOR;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X9Y112_B;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X9Y112_B1;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X9Y112_B2;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X9Y112_B3;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X9Y112_B4;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X9Y112_B5;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X9Y112_B6;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X9Y112_BO5;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X9Y112_BO6;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X9Y112_BQ;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X9Y112_B_CY;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X9Y112_B_XOR;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X9Y112_C;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X9Y112_C1;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X9Y112_C2;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X9Y112_C3;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X9Y112_C4;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X9Y112_C5;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X9Y112_C6;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X9Y112_CLK;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X9Y112_CO5;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X9Y112_CO6;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X9Y112_CQ;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X9Y112_C_CY;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X9Y112_C_XOR;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X9Y112_D;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X9Y112_D1;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X9Y112_D2;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X9Y112_D3;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X9Y112_D4;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X9Y112_D5;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X9Y112_D6;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X9Y112_DO5;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X9Y112_DO6;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X9Y112_D_CY;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X9Y112_D_XOR;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X8Y113_A;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X8Y113_A1;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X8Y113_A2;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X8Y113_A3;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X8Y113_A4;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X8Y113_A5;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X8Y113_A6;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X8Y113_AO5;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X8Y113_AO6;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X8Y113_AQ;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X8Y113_A_CY;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X8Y113_A_XOR;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X8Y113_B;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X8Y113_B1;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X8Y113_B2;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X8Y113_B3;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X8Y113_B4;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X8Y113_B5;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X8Y113_B6;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X8Y113_BMUX;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X8Y113_BO5;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X8Y113_BO6;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X8Y113_B_CY;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X8Y113_B_XOR;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X8Y113_C;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X8Y113_C1;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X8Y113_C2;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X8Y113_C3;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X8Y113_C4;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X8Y113_C5;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X8Y113_C6;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X8Y113_CLK;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X8Y113_CO5;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X8Y113_CO6;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X8Y113_C_CY;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X8Y113_C_XOR;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X8Y113_D;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X8Y113_D1;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X8Y113_D2;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X8Y113_D3;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X8Y113_D4;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X8Y113_D5;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X8Y113_D6;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X8Y113_DO5;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X8Y113_DO6;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X8Y113_D_CY;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X8Y113_D_XOR;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X9Y113_A;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X9Y113_A1;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X9Y113_A2;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X9Y113_A3;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X9Y113_A4;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X9Y113_A5;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X9Y113_A5Q;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X9Y113_A6;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X9Y113_AMUX;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X9Y113_AO5;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X9Y113_AO6;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X9Y113_AQ;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X9Y113_A_CY;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X9Y113_A_XOR;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X9Y113_B;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X9Y113_B1;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X9Y113_B2;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X9Y113_B3;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X9Y113_B4;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X9Y113_B5;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X9Y113_B6;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X9Y113_BO5;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X9Y113_BO6;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X9Y113_BQ;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X9Y113_B_CY;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X9Y113_B_XOR;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X9Y113_C;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X9Y113_C1;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X9Y113_C2;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X9Y113_C3;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X9Y113_C4;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X9Y113_C5;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X9Y113_C6;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X9Y113_CLK;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X9Y113_CO5;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X9Y113_CO6;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X9Y113_C_CY;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X9Y113_C_XOR;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X9Y113_D;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X9Y113_D1;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X9Y113_D2;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X9Y113_D3;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X9Y113_D4;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X9Y113_D5;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X9Y113_D6;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X9Y113_DO5;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X9Y113_DO6;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X9Y113_D_CY;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X9Y113_D_XOR;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X8Y114_A;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X8Y114_A1;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X8Y114_A2;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X8Y114_A3;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X8Y114_A4;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X8Y114_A5;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X8Y114_A6;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X8Y114_AO5;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X8Y114_AO6;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X8Y114_AQ;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X8Y114_A_CY;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X8Y114_A_XOR;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X8Y114_B;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X8Y114_B1;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X8Y114_B2;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X8Y114_B3;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X8Y114_B4;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X8Y114_B5;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X8Y114_B6;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X8Y114_BO5;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X8Y114_BO6;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X8Y114_BQ;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X8Y114_B_CY;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X8Y114_B_XOR;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X8Y114_C;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X8Y114_C1;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X8Y114_C2;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X8Y114_C3;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X8Y114_C4;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X8Y114_C5;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X8Y114_C6;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X8Y114_CLK;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X8Y114_CO5;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X8Y114_CO6;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X8Y114_C_CY;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X8Y114_C_XOR;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X8Y114_D;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X8Y114_D1;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X8Y114_D2;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X8Y114_D3;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X8Y114_D4;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X8Y114_D5;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X8Y114_D6;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X8Y114_DO5;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X8Y114_DO6;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X8Y114_D_CY;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X8Y114_D_XOR;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X9Y114_A;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X9Y114_A1;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X9Y114_A2;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X9Y114_A3;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X9Y114_A4;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X9Y114_A5;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X9Y114_A6;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X9Y114_AO5;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X9Y114_AO6;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X9Y114_A_CY;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X9Y114_A_XOR;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X9Y114_B;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X9Y114_B1;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X9Y114_B2;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X9Y114_B3;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X9Y114_B4;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X9Y114_B5;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X9Y114_B6;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X9Y114_BO5;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X9Y114_BO6;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X9Y114_B_CY;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X9Y114_B_XOR;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X9Y114_C;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X9Y114_C1;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X9Y114_C2;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X9Y114_C3;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X9Y114_C4;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X9Y114_C5;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X9Y114_C6;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X9Y114_CO5;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X9Y114_CO6;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X9Y114_C_CY;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X9Y114_C_XOR;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X9Y114_D;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X9Y114_D1;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X9Y114_D2;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X9Y114_D3;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X9Y114_D4;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X9Y114_D5;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X9Y114_D6;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X9Y114_DO5;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X9Y114_DO6;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X9Y114_D_CY;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X9Y114_D_XOR;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X8Y115_A;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X8Y115_A1;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X8Y115_A2;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X8Y115_A3;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X8Y115_A4;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X8Y115_A5;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X8Y115_A5Q;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X8Y115_A6;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X8Y115_AMUX;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X8Y115_AO5;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X8Y115_AO6;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X8Y115_AQ;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X8Y115_AX;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X8Y115_A_CY;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X8Y115_A_XOR;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X8Y115_B;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X8Y115_B1;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X8Y115_B2;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X8Y115_B3;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X8Y115_B4;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X8Y115_B5;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X8Y115_B6;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X8Y115_BO5;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X8Y115_BO6;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X8Y115_BQ;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X8Y115_B_CY;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X8Y115_B_XOR;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X8Y115_C;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X8Y115_C1;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X8Y115_C2;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X8Y115_C3;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X8Y115_C4;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X8Y115_C5;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X8Y115_C6;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X8Y115_CLK;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X8Y115_CO5;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X8Y115_CO6;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X8Y115_CQ;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X8Y115_C_CY;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X8Y115_C_XOR;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X8Y115_D;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X8Y115_D1;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X8Y115_D2;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X8Y115_D3;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X8Y115_D4;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X8Y115_D5;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X8Y115_D6;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X8Y115_DMUX;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X8Y115_DO5;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X8Y115_DO6;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X8Y115_D_CY;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X8Y115_D_XOR;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X9Y115_A;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X9Y115_A1;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X9Y115_A2;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X9Y115_A3;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X9Y115_A4;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X9Y115_A5;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X9Y115_A6;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X9Y115_AO5;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X9Y115_AO6;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X9Y115_AQ;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X9Y115_A_CY;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X9Y115_A_XOR;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X9Y115_B;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X9Y115_B1;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X9Y115_B2;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X9Y115_B3;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X9Y115_B4;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X9Y115_B5;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X9Y115_B5Q;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X9Y115_B6;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X9Y115_BMUX;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X9Y115_BO5;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X9Y115_BO6;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X9Y115_BQ;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X9Y115_B_CY;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X9Y115_B_XOR;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X9Y115_C;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X9Y115_C1;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X9Y115_C2;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X9Y115_C3;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X9Y115_C4;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X9Y115_C5;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X9Y115_C5Q;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X9Y115_C6;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X9Y115_CLK;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X9Y115_CMUX;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X9Y115_CO5;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X9Y115_CO6;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X9Y115_CQ;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X9Y115_C_CY;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X9Y115_C_XOR;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X9Y115_D;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X9Y115_D1;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X9Y115_D2;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X9Y115_D3;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X9Y115_D4;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X9Y115_D5;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X9Y115_D6;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X9Y115_DO5;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X9Y115_DO6;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X9Y115_DQ;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X9Y115_D_CY;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X9Y115_D_XOR;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X8Y116_A;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X8Y116_A1;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X8Y116_A2;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X8Y116_A3;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X8Y116_A4;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X8Y116_A5;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X8Y116_A6;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X8Y116_AO5;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X8Y116_AO6;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X8Y116_AQ;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X8Y116_A_CY;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X8Y116_A_XOR;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X8Y116_B;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X8Y116_B1;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X8Y116_B2;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X8Y116_B3;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X8Y116_B4;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X8Y116_B5;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X8Y116_B6;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X8Y116_BO5;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X8Y116_BO6;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X8Y116_BQ;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X8Y116_B_CY;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X8Y116_B_XOR;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X8Y116_C;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X8Y116_C1;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X8Y116_C2;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X8Y116_C3;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X8Y116_C4;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X8Y116_C5;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X8Y116_C6;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X8Y116_CLK;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X8Y116_CO5;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X8Y116_CO6;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X8Y116_CQ;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X8Y116_C_CY;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X8Y116_C_XOR;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X8Y116_D;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X8Y116_D1;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X8Y116_D2;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X8Y116_D3;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X8Y116_D4;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X8Y116_D5;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X8Y116_D6;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X8Y116_DO5;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X8Y116_DO6;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X8Y116_D_CY;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X8Y116_D_XOR;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X9Y116_A;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X9Y116_A1;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X9Y116_A2;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X9Y116_A3;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X9Y116_A4;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X9Y116_A5;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X9Y116_A6;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X9Y116_AO5;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X9Y116_AO6;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X9Y116_AQ;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X9Y116_A_CY;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X9Y116_A_XOR;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X9Y116_B;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X9Y116_B1;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X9Y116_B2;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X9Y116_B3;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X9Y116_B4;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X9Y116_B5;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X9Y116_B6;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X9Y116_BO5;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X9Y116_BO6;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X9Y116_B_CY;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X9Y116_B_XOR;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X9Y116_C;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X9Y116_C1;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X9Y116_C2;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X9Y116_C3;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X9Y116_C4;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X9Y116_C5;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X9Y116_C6;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X9Y116_CLK;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X9Y116_CO5;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X9Y116_CO6;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X9Y116_C_CY;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X9Y116_C_XOR;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X9Y116_D;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X9Y116_D1;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X9Y116_D2;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X9Y116_D3;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X9Y116_D4;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X9Y116_D5;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X9Y116_D6;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X9Y116_DO5;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X9Y116_DO6;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X9Y116_D_CY;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X9Y116_D_XOR;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X8Y117_A;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X8Y117_A1;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X8Y117_A2;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X8Y117_A3;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X8Y117_A4;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X8Y117_A5;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X8Y117_A5Q;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X8Y117_A6;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X8Y117_AMUX;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X8Y117_AO5;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X8Y117_AO6;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X8Y117_AQ;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X8Y117_AX;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X8Y117_A_CY;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X8Y117_A_XOR;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X8Y117_B;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X8Y117_B1;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X8Y117_B2;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X8Y117_B3;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X8Y117_B4;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X8Y117_B5;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X8Y117_B6;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X8Y117_BO5;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X8Y117_BO6;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X8Y117_BQ;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X8Y117_B_CY;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X8Y117_B_XOR;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X8Y117_C;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X8Y117_C1;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X8Y117_C2;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X8Y117_C3;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X8Y117_C4;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X8Y117_C5;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X8Y117_C6;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X8Y117_CLK;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X8Y117_CO5;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X8Y117_CO6;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X8Y117_CQ;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X8Y117_C_CY;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X8Y117_C_XOR;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X8Y117_D;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X8Y117_D1;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X8Y117_D2;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X8Y117_D3;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X8Y117_D4;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X8Y117_D5;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X8Y117_D6;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X8Y117_DMUX;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X8Y117_DO5;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X8Y117_DO6;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X8Y117_D_CY;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X8Y117_D_XOR;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X9Y117_A;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X9Y117_A1;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X9Y117_A2;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X9Y117_A3;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X9Y117_A4;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X9Y117_A5;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X9Y117_A6;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X9Y117_AO5;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X9Y117_AO6;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X9Y117_AQ;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X9Y117_A_CY;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X9Y117_A_XOR;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X9Y117_B;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X9Y117_B1;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X9Y117_B2;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X9Y117_B3;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X9Y117_B4;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X9Y117_B5;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X9Y117_B6;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X9Y117_BO5;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X9Y117_BO6;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X9Y117_BQ;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X9Y117_B_CY;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X9Y117_B_XOR;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X9Y117_C;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X9Y117_C1;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X9Y117_C2;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X9Y117_C3;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X9Y117_C4;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X9Y117_C5;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X9Y117_C6;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X9Y117_CLK;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X9Y117_CO5;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X9Y117_CO6;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X9Y117_CQ;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X9Y117_C_CY;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X9Y117_C_XOR;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X9Y117_D;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X9Y117_D1;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X9Y117_D2;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X9Y117_D3;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X9Y117_D4;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X9Y117_D5;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X9Y117_D6;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X9Y117_DO5;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X9Y117_DO6;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X9Y117_DQ;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X9Y117_D_CY;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X9Y117_D_XOR;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X8Y118_A;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X8Y118_A1;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X8Y118_A2;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X8Y118_A3;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X8Y118_A4;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X8Y118_A5;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X8Y118_A6;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X8Y118_AO5;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X8Y118_AO6;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X8Y118_AQ;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X8Y118_A_CY;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X8Y118_A_XOR;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X8Y118_B;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X8Y118_B1;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X8Y118_B2;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X8Y118_B3;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X8Y118_B4;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X8Y118_B5;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X8Y118_B6;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X8Y118_BO5;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X8Y118_BO6;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X8Y118_BQ;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X8Y118_B_CY;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X8Y118_B_XOR;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X8Y118_C;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X8Y118_C1;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X8Y118_C2;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X8Y118_C3;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X8Y118_C4;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X8Y118_C5;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X8Y118_C6;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X8Y118_CLK;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X8Y118_CO5;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X8Y118_CO6;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X8Y118_CQ;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X8Y118_C_CY;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X8Y118_C_XOR;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X8Y118_D;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X8Y118_D1;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X8Y118_D2;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X8Y118_D3;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X8Y118_D4;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X8Y118_D5;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X8Y118_D6;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X8Y118_DO5;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X8Y118_DO6;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X8Y118_DQ;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X8Y118_D_CY;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X8Y118_D_XOR;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X9Y118_A;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X9Y118_A1;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X9Y118_A2;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X9Y118_A3;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X9Y118_A4;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X9Y118_A5;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X9Y118_A6;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X9Y118_AO5;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X9Y118_AO6;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X9Y118_AQ;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X9Y118_A_CY;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X9Y118_A_XOR;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X9Y118_B;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X9Y118_B1;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X9Y118_B2;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X9Y118_B3;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X9Y118_B4;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X9Y118_B5;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X9Y118_B6;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X9Y118_BO5;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X9Y118_BO6;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X9Y118_BQ;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X9Y118_B_CY;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X9Y118_B_XOR;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X9Y118_C;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X9Y118_C1;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X9Y118_C2;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X9Y118_C3;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X9Y118_C4;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X9Y118_C5;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X9Y118_C6;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X9Y118_CLK;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X9Y118_CO5;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X9Y118_CO6;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X9Y118_CQ;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X9Y118_C_CY;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X9Y118_C_XOR;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X9Y118_D;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X9Y118_D1;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X9Y118_D2;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X9Y118_D3;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X9Y118_D4;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X9Y118_D5;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X9Y118_D6;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X9Y118_DO5;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X9Y118_DO6;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X9Y118_D_CY;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X9Y118_D_XOR;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X8Y119_A;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X8Y119_A1;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X8Y119_A2;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X8Y119_A3;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X8Y119_A4;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X8Y119_A5;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X8Y119_A6;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X8Y119_AO5;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X8Y119_AO6;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X8Y119_AQ;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X8Y119_A_CY;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X8Y119_A_XOR;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X8Y119_B;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X8Y119_B1;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X8Y119_B2;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X8Y119_B3;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X8Y119_B4;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X8Y119_B5;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X8Y119_B6;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X8Y119_BO5;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X8Y119_BO6;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X8Y119_BQ;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X8Y119_B_CY;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X8Y119_B_XOR;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X8Y119_C;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X8Y119_C1;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X8Y119_C2;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X8Y119_C3;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X8Y119_C4;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X8Y119_C5;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X8Y119_C5Q;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X8Y119_C6;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X8Y119_CLK;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X8Y119_CMUX;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X8Y119_CO5;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X8Y119_CO6;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X8Y119_CQ;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X8Y119_C_CY;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X8Y119_C_XOR;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X8Y119_D;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X8Y119_D1;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X8Y119_D2;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X8Y119_D3;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X8Y119_D4;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X8Y119_D5;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X8Y119_D5Q;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X8Y119_D6;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X8Y119_DMUX;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X8Y119_DO5;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X8Y119_DO6;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X8Y119_DQ;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X8Y119_D_CY;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X8Y119_D_XOR;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X9Y119_A;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X9Y119_A1;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X9Y119_A2;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X9Y119_A3;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X9Y119_A4;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X9Y119_A5;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X9Y119_A6;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X9Y119_AO5;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X9Y119_AO6;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X9Y119_AQ;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X9Y119_A_CY;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X9Y119_A_XOR;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X9Y119_B;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X9Y119_B1;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X9Y119_B2;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X9Y119_B3;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X9Y119_B4;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X9Y119_B5;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X9Y119_B6;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X9Y119_BO5;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X9Y119_BO6;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X9Y119_BQ;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X9Y119_B_CY;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X9Y119_B_XOR;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X9Y119_C;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X9Y119_C1;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X9Y119_C2;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X9Y119_C3;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X9Y119_C4;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X9Y119_C5;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X9Y119_C6;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X9Y119_CLK;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X9Y119_CO5;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X9Y119_CO6;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X9Y119_CQ;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X9Y119_C_CY;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X9Y119_C_XOR;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X9Y119_D;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X9Y119_D1;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X9Y119_D2;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X9Y119_D3;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X9Y119_D4;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X9Y119_D5;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X9Y119_D6;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X9Y119_DMUX;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X9Y119_DO5;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X9Y119_DO6;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X9Y119_D_CY;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X9Y119_D_XOR;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X8Y120_A;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X8Y120_A1;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X8Y120_A2;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X8Y120_A3;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X8Y120_A4;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X8Y120_A5;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X8Y120_A6;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X8Y120_AO5;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X8Y120_AO6;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X8Y120_AQ;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X8Y120_A_CY;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X8Y120_A_XOR;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X8Y120_B;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X8Y120_B1;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X8Y120_B2;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X8Y120_B3;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X8Y120_B4;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X8Y120_B5;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X8Y120_B6;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X8Y120_BO5;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X8Y120_BO6;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X8Y120_BQ;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X8Y120_B_CY;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X8Y120_B_XOR;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X8Y120_C;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X8Y120_C1;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X8Y120_C2;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X8Y120_C3;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X8Y120_C4;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X8Y120_C5;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X8Y120_C6;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X8Y120_CLK;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X8Y120_CO5;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X8Y120_CO6;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X8Y120_CQ;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X8Y120_C_CY;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X8Y120_C_XOR;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X8Y120_D;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X8Y120_D1;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X8Y120_D2;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X8Y120_D3;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X8Y120_D4;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X8Y120_D5;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X8Y120_D6;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X8Y120_DO5;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X8Y120_DO6;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X8Y120_DQ;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X8Y120_D_CY;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X8Y120_D_XOR;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X9Y120_A;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X9Y120_A1;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X9Y120_A2;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X9Y120_A3;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X9Y120_A4;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X9Y120_A5;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X9Y120_A5Q;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X9Y120_A6;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X9Y120_AMUX;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X9Y120_AO5;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X9Y120_AO6;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X9Y120_AQ;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X9Y120_A_CY;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X9Y120_A_XOR;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X9Y120_B;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X9Y120_B1;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X9Y120_B2;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X9Y120_B3;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X9Y120_B4;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X9Y120_B5;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X9Y120_B6;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X9Y120_BO5;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X9Y120_BO6;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X9Y120_BQ;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X9Y120_B_CY;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X9Y120_B_XOR;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X9Y120_C;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X9Y120_C1;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X9Y120_C2;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X9Y120_C3;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X9Y120_C4;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X9Y120_C5;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X9Y120_C6;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X9Y120_CLK;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X9Y120_CO5;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X9Y120_CO6;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X9Y120_CQ;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X9Y120_C_CY;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X9Y120_C_XOR;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X9Y120_D;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X9Y120_D1;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X9Y120_D2;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X9Y120_D3;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X9Y120_D4;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X9Y120_D5;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X9Y120_D5Q;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X9Y120_D6;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X9Y120_DMUX;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X9Y120_DO5;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X9Y120_DO6;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X9Y120_DQ;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X9Y120_D_CY;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X9Y120_D_XOR;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X8Y121_A;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X8Y121_A1;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X8Y121_A2;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X8Y121_A3;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X8Y121_A4;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X8Y121_A5;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X8Y121_A6;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X8Y121_AO5;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X8Y121_AO6;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X8Y121_AQ;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X8Y121_A_CY;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X8Y121_A_XOR;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X8Y121_B;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X8Y121_B1;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X8Y121_B2;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X8Y121_B3;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X8Y121_B4;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X8Y121_B5;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X8Y121_B6;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X8Y121_BO5;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X8Y121_BO6;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X8Y121_BQ;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X8Y121_B_CY;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X8Y121_B_XOR;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X8Y121_C;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X8Y121_C1;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X8Y121_C2;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X8Y121_C3;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X8Y121_C4;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X8Y121_C5;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X8Y121_C5Q;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X8Y121_C6;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X8Y121_CLK;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X8Y121_CMUX;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X8Y121_CO5;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X8Y121_CO6;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X8Y121_CQ;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X8Y121_C_CY;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X8Y121_C_XOR;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X8Y121_D;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X8Y121_D1;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X8Y121_D2;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X8Y121_D3;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X8Y121_D4;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X8Y121_D5;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X8Y121_D6;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X8Y121_DO5;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X8Y121_DO6;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X8Y121_D_CY;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X8Y121_D_XOR;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X9Y121_A;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X9Y121_A1;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X9Y121_A2;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X9Y121_A3;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X9Y121_A4;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X9Y121_A5;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X9Y121_A5Q;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X9Y121_A6;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X9Y121_AMUX;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X9Y121_AO5;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X9Y121_AO6;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X9Y121_AQ;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X9Y121_AX;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X9Y121_A_CY;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X9Y121_A_XOR;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X9Y121_B;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X9Y121_B1;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X9Y121_B2;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X9Y121_B3;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X9Y121_B4;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X9Y121_B5;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X9Y121_B6;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X9Y121_BO5;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X9Y121_BO6;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X9Y121_BQ;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X9Y121_B_CY;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X9Y121_B_XOR;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X9Y121_C;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X9Y121_C1;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X9Y121_C2;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X9Y121_C3;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X9Y121_C4;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X9Y121_C5;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X9Y121_C6;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X9Y121_CLK;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X9Y121_CMUX;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X9Y121_CO5;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X9Y121_CO6;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X9Y121_C_CY;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X9Y121_C_XOR;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X9Y121_D;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X9Y121_D1;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X9Y121_D2;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X9Y121_D3;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X9Y121_D4;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X9Y121_D5;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X9Y121_D6;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X9Y121_DMUX;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X9Y121_DO5;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X9Y121_DO6;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X9Y121_D_CY;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X9Y121_D_XOR;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X8Y122_A;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X8Y122_A1;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X8Y122_A2;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X8Y122_A3;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X8Y122_A4;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X8Y122_A5;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X8Y122_A6;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X8Y122_AO5;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X8Y122_AO6;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X8Y122_AQ;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X8Y122_A_CY;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X8Y122_A_XOR;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X8Y122_B;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X8Y122_B1;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X8Y122_B2;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X8Y122_B3;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X8Y122_B4;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X8Y122_B5;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X8Y122_B6;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X8Y122_BO5;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X8Y122_BO6;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X8Y122_BQ;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X8Y122_B_CY;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X8Y122_B_XOR;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X8Y122_C;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X8Y122_C1;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X8Y122_C2;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X8Y122_C3;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X8Y122_C4;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X8Y122_C5;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X8Y122_C6;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X8Y122_CLK;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X8Y122_CO5;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X8Y122_CO6;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X8Y122_CQ;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X8Y122_C_CY;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X8Y122_C_XOR;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X8Y122_D;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X8Y122_D1;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X8Y122_D2;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X8Y122_D3;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X8Y122_D4;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X8Y122_D5;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X8Y122_D6;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X8Y122_DO5;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X8Y122_DO6;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X8Y122_DQ;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X8Y122_D_CY;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X8Y122_D_XOR;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X9Y122_A;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X9Y122_A1;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X9Y122_A2;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X9Y122_A3;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X9Y122_A4;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X9Y122_A5;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X9Y122_A5Q;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X9Y122_A6;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X9Y122_AMUX;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X9Y122_AO5;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X9Y122_AO6;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X9Y122_AQ;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X9Y122_A_CY;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X9Y122_A_XOR;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X9Y122_B;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X9Y122_B1;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X9Y122_B2;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X9Y122_B3;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X9Y122_B4;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X9Y122_B5;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X9Y122_B6;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X9Y122_BO5;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X9Y122_BO6;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X9Y122_BQ;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X9Y122_B_CY;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X9Y122_B_XOR;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X9Y122_C;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X9Y122_C1;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X9Y122_C2;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X9Y122_C3;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X9Y122_C4;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X9Y122_C5;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X9Y122_C6;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X9Y122_CLK;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X9Y122_CO5;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X9Y122_CO6;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X9Y122_C_CY;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X9Y122_C_XOR;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X9Y122_D;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X9Y122_D1;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X9Y122_D2;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X9Y122_D3;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X9Y122_D4;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X9Y122_D5;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X9Y122_D6;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X9Y122_DO5;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X9Y122_DO6;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X9Y122_D_CY;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X9Y122_D_XOR;
  wire [0:0] CLBLM_R_X7Y123_SLICE_X8Y123_A;
  wire [0:0] CLBLM_R_X7Y123_SLICE_X8Y123_A1;
  wire [0:0] CLBLM_R_X7Y123_SLICE_X8Y123_A2;
  wire [0:0] CLBLM_R_X7Y123_SLICE_X8Y123_A3;
  wire [0:0] CLBLM_R_X7Y123_SLICE_X8Y123_A4;
  wire [0:0] CLBLM_R_X7Y123_SLICE_X8Y123_A5;
  wire [0:0] CLBLM_R_X7Y123_SLICE_X8Y123_A6;
  wire [0:0] CLBLM_R_X7Y123_SLICE_X8Y123_AO5;
  wire [0:0] CLBLM_R_X7Y123_SLICE_X8Y123_AO6;
  wire [0:0] CLBLM_R_X7Y123_SLICE_X8Y123_AQ;
  wire [0:0] CLBLM_R_X7Y123_SLICE_X8Y123_A_CY;
  wire [0:0] CLBLM_R_X7Y123_SLICE_X8Y123_A_XOR;
  wire [0:0] CLBLM_R_X7Y123_SLICE_X8Y123_B;
  wire [0:0] CLBLM_R_X7Y123_SLICE_X8Y123_B1;
  wire [0:0] CLBLM_R_X7Y123_SLICE_X8Y123_B2;
  wire [0:0] CLBLM_R_X7Y123_SLICE_X8Y123_B3;
  wire [0:0] CLBLM_R_X7Y123_SLICE_X8Y123_B4;
  wire [0:0] CLBLM_R_X7Y123_SLICE_X8Y123_B5;
  wire [0:0] CLBLM_R_X7Y123_SLICE_X8Y123_B6;
  wire [0:0] CLBLM_R_X7Y123_SLICE_X8Y123_BO5;
  wire [0:0] CLBLM_R_X7Y123_SLICE_X8Y123_BO6;
  wire [0:0] CLBLM_R_X7Y123_SLICE_X8Y123_BQ;
  wire [0:0] CLBLM_R_X7Y123_SLICE_X8Y123_B_CY;
  wire [0:0] CLBLM_R_X7Y123_SLICE_X8Y123_B_XOR;
  wire [0:0] CLBLM_R_X7Y123_SLICE_X8Y123_C;
  wire [0:0] CLBLM_R_X7Y123_SLICE_X8Y123_C1;
  wire [0:0] CLBLM_R_X7Y123_SLICE_X8Y123_C2;
  wire [0:0] CLBLM_R_X7Y123_SLICE_X8Y123_C3;
  wire [0:0] CLBLM_R_X7Y123_SLICE_X8Y123_C4;
  wire [0:0] CLBLM_R_X7Y123_SLICE_X8Y123_C5;
  wire [0:0] CLBLM_R_X7Y123_SLICE_X8Y123_C6;
  wire [0:0] CLBLM_R_X7Y123_SLICE_X8Y123_CLK;
  wire [0:0] CLBLM_R_X7Y123_SLICE_X8Y123_CO5;
  wire [0:0] CLBLM_R_X7Y123_SLICE_X8Y123_CO6;
  wire [0:0] CLBLM_R_X7Y123_SLICE_X8Y123_CQ;
  wire [0:0] CLBLM_R_X7Y123_SLICE_X8Y123_C_CY;
  wire [0:0] CLBLM_R_X7Y123_SLICE_X8Y123_C_XOR;
  wire [0:0] CLBLM_R_X7Y123_SLICE_X8Y123_D;
  wire [0:0] CLBLM_R_X7Y123_SLICE_X8Y123_D1;
  wire [0:0] CLBLM_R_X7Y123_SLICE_X8Y123_D2;
  wire [0:0] CLBLM_R_X7Y123_SLICE_X8Y123_D3;
  wire [0:0] CLBLM_R_X7Y123_SLICE_X8Y123_D4;
  wire [0:0] CLBLM_R_X7Y123_SLICE_X8Y123_D5;
  wire [0:0] CLBLM_R_X7Y123_SLICE_X8Y123_D6;
  wire [0:0] CLBLM_R_X7Y123_SLICE_X8Y123_DO5;
  wire [0:0] CLBLM_R_X7Y123_SLICE_X8Y123_DO6;
  wire [0:0] CLBLM_R_X7Y123_SLICE_X8Y123_D_CY;
  wire [0:0] CLBLM_R_X7Y123_SLICE_X8Y123_D_XOR;
  wire [0:0] CLBLM_R_X7Y123_SLICE_X9Y123_A;
  wire [0:0] CLBLM_R_X7Y123_SLICE_X9Y123_A1;
  wire [0:0] CLBLM_R_X7Y123_SLICE_X9Y123_A2;
  wire [0:0] CLBLM_R_X7Y123_SLICE_X9Y123_A3;
  wire [0:0] CLBLM_R_X7Y123_SLICE_X9Y123_A4;
  wire [0:0] CLBLM_R_X7Y123_SLICE_X9Y123_A5;
  wire [0:0] CLBLM_R_X7Y123_SLICE_X9Y123_A6;
  wire [0:0] CLBLM_R_X7Y123_SLICE_X9Y123_AO5;
  wire [0:0] CLBLM_R_X7Y123_SLICE_X9Y123_AO6;
  wire [0:0] CLBLM_R_X7Y123_SLICE_X9Y123_AQ;
  wire [0:0] CLBLM_R_X7Y123_SLICE_X9Y123_A_CY;
  wire [0:0] CLBLM_R_X7Y123_SLICE_X9Y123_A_XOR;
  wire [0:0] CLBLM_R_X7Y123_SLICE_X9Y123_B;
  wire [0:0] CLBLM_R_X7Y123_SLICE_X9Y123_B1;
  wire [0:0] CLBLM_R_X7Y123_SLICE_X9Y123_B2;
  wire [0:0] CLBLM_R_X7Y123_SLICE_X9Y123_B3;
  wire [0:0] CLBLM_R_X7Y123_SLICE_X9Y123_B4;
  wire [0:0] CLBLM_R_X7Y123_SLICE_X9Y123_B5;
  wire [0:0] CLBLM_R_X7Y123_SLICE_X9Y123_B6;
  wire [0:0] CLBLM_R_X7Y123_SLICE_X9Y123_BMUX;
  wire [0:0] CLBLM_R_X7Y123_SLICE_X9Y123_BO5;
  wire [0:0] CLBLM_R_X7Y123_SLICE_X9Y123_BO6;
  wire [0:0] CLBLM_R_X7Y123_SLICE_X9Y123_B_CY;
  wire [0:0] CLBLM_R_X7Y123_SLICE_X9Y123_B_XOR;
  wire [0:0] CLBLM_R_X7Y123_SLICE_X9Y123_C;
  wire [0:0] CLBLM_R_X7Y123_SLICE_X9Y123_C1;
  wire [0:0] CLBLM_R_X7Y123_SLICE_X9Y123_C2;
  wire [0:0] CLBLM_R_X7Y123_SLICE_X9Y123_C3;
  wire [0:0] CLBLM_R_X7Y123_SLICE_X9Y123_C4;
  wire [0:0] CLBLM_R_X7Y123_SLICE_X9Y123_C5;
  wire [0:0] CLBLM_R_X7Y123_SLICE_X9Y123_C6;
  wire [0:0] CLBLM_R_X7Y123_SLICE_X9Y123_CLK;
  wire [0:0] CLBLM_R_X7Y123_SLICE_X9Y123_CO5;
  wire [0:0] CLBLM_R_X7Y123_SLICE_X9Y123_CO6;
  wire [0:0] CLBLM_R_X7Y123_SLICE_X9Y123_C_CY;
  wire [0:0] CLBLM_R_X7Y123_SLICE_X9Y123_C_XOR;
  wire [0:0] CLBLM_R_X7Y123_SLICE_X9Y123_D;
  wire [0:0] CLBLM_R_X7Y123_SLICE_X9Y123_D1;
  wire [0:0] CLBLM_R_X7Y123_SLICE_X9Y123_D2;
  wire [0:0] CLBLM_R_X7Y123_SLICE_X9Y123_D3;
  wire [0:0] CLBLM_R_X7Y123_SLICE_X9Y123_D4;
  wire [0:0] CLBLM_R_X7Y123_SLICE_X9Y123_D5;
  wire [0:0] CLBLM_R_X7Y123_SLICE_X9Y123_D6;
  wire [0:0] CLBLM_R_X7Y123_SLICE_X9Y123_DO5;
  wire [0:0] CLBLM_R_X7Y123_SLICE_X9Y123_DO6;
  wire [0:0] CLBLM_R_X7Y123_SLICE_X9Y123_D_CY;
  wire [0:0] CLBLM_R_X7Y123_SLICE_X9Y123_D_XOR;
  wire [0:0] CLBLM_R_X7Y124_SLICE_X8Y124_A;
  wire [0:0] CLBLM_R_X7Y124_SLICE_X8Y124_A1;
  wire [0:0] CLBLM_R_X7Y124_SLICE_X8Y124_A2;
  wire [0:0] CLBLM_R_X7Y124_SLICE_X8Y124_A3;
  wire [0:0] CLBLM_R_X7Y124_SLICE_X8Y124_A4;
  wire [0:0] CLBLM_R_X7Y124_SLICE_X8Y124_A5;
  wire [0:0] CLBLM_R_X7Y124_SLICE_X8Y124_A5Q;
  wire [0:0] CLBLM_R_X7Y124_SLICE_X8Y124_A6;
  wire [0:0] CLBLM_R_X7Y124_SLICE_X8Y124_AMUX;
  wire [0:0] CLBLM_R_X7Y124_SLICE_X8Y124_AO5;
  wire [0:0] CLBLM_R_X7Y124_SLICE_X8Y124_AO6;
  wire [0:0] CLBLM_R_X7Y124_SLICE_X8Y124_AQ;
  wire [0:0] CLBLM_R_X7Y124_SLICE_X8Y124_AX;
  wire [0:0] CLBLM_R_X7Y124_SLICE_X8Y124_A_CY;
  wire [0:0] CLBLM_R_X7Y124_SLICE_X8Y124_A_XOR;
  wire [0:0] CLBLM_R_X7Y124_SLICE_X8Y124_B;
  wire [0:0] CLBLM_R_X7Y124_SLICE_X8Y124_B1;
  wire [0:0] CLBLM_R_X7Y124_SLICE_X8Y124_B2;
  wire [0:0] CLBLM_R_X7Y124_SLICE_X8Y124_B3;
  wire [0:0] CLBLM_R_X7Y124_SLICE_X8Y124_B4;
  wire [0:0] CLBLM_R_X7Y124_SLICE_X8Y124_B5;
  wire [0:0] CLBLM_R_X7Y124_SLICE_X8Y124_B6;
  wire [0:0] CLBLM_R_X7Y124_SLICE_X8Y124_BO5;
  wire [0:0] CLBLM_R_X7Y124_SLICE_X8Y124_BO6;
  wire [0:0] CLBLM_R_X7Y124_SLICE_X8Y124_BQ;
  wire [0:0] CLBLM_R_X7Y124_SLICE_X8Y124_B_CY;
  wire [0:0] CLBLM_R_X7Y124_SLICE_X8Y124_B_XOR;
  wire [0:0] CLBLM_R_X7Y124_SLICE_X8Y124_C;
  wire [0:0] CLBLM_R_X7Y124_SLICE_X8Y124_C1;
  wire [0:0] CLBLM_R_X7Y124_SLICE_X8Y124_C2;
  wire [0:0] CLBLM_R_X7Y124_SLICE_X8Y124_C3;
  wire [0:0] CLBLM_R_X7Y124_SLICE_X8Y124_C4;
  wire [0:0] CLBLM_R_X7Y124_SLICE_X8Y124_C5;
  wire [0:0] CLBLM_R_X7Y124_SLICE_X8Y124_C6;
  wire [0:0] CLBLM_R_X7Y124_SLICE_X8Y124_CLK;
  wire [0:0] CLBLM_R_X7Y124_SLICE_X8Y124_CO5;
  wire [0:0] CLBLM_R_X7Y124_SLICE_X8Y124_CO6;
  wire [0:0] CLBLM_R_X7Y124_SLICE_X8Y124_CQ;
  wire [0:0] CLBLM_R_X7Y124_SLICE_X8Y124_C_CY;
  wire [0:0] CLBLM_R_X7Y124_SLICE_X8Y124_C_XOR;
  wire [0:0] CLBLM_R_X7Y124_SLICE_X8Y124_D;
  wire [0:0] CLBLM_R_X7Y124_SLICE_X8Y124_D1;
  wire [0:0] CLBLM_R_X7Y124_SLICE_X8Y124_D2;
  wire [0:0] CLBLM_R_X7Y124_SLICE_X8Y124_D3;
  wire [0:0] CLBLM_R_X7Y124_SLICE_X8Y124_D4;
  wire [0:0] CLBLM_R_X7Y124_SLICE_X8Y124_D5;
  wire [0:0] CLBLM_R_X7Y124_SLICE_X8Y124_D6;
  wire [0:0] CLBLM_R_X7Y124_SLICE_X8Y124_DMUX;
  wire [0:0] CLBLM_R_X7Y124_SLICE_X8Y124_DO5;
  wire [0:0] CLBLM_R_X7Y124_SLICE_X8Y124_DO6;
  wire [0:0] CLBLM_R_X7Y124_SLICE_X8Y124_D_CY;
  wire [0:0] CLBLM_R_X7Y124_SLICE_X8Y124_D_XOR;
  wire [0:0] CLBLM_R_X7Y124_SLICE_X9Y124_A;
  wire [0:0] CLBLM_R_X7Y124_SLICE_X9Y124_A1;
  wire [0:0] CLBLM_R_X7Y124_SLICE_X9Y124_A2;
  wire [0:0] CLBLM_R_X7Y124_SLICE_X9Y124_A3;
  wire [0:0] CLBLM_R_X7Y124_SLICE_X9Y124_A4;
  wire [0:0] CLBLM_R_X7Y124_SLICE_X9Y124_A5;
  wire [0:0] CLBLM_R_X7Y124_SLICE_X9Y124_A6;
  wire [0:0] CLBLM_R_X7Y124_SLICE_X9Y124_AO5;
  wire [0:0] CLBLM_R_X7Y124_SLICE_X9Y124_AO6;
  wire [0:0] CLBLM_R_X7Y124_SLICE_X9Y124_AQ;
  wire [0:0] CLBLM_R_X7Y124_SLICE_X9Y124_A_CY;
  wire [0:0] CLBLM_R_X7Y124_SLICE_X9Y124_A_XOR;
  wire [0:0] CLBLM_R_X7Y124_SLICE_X9Y124_B;
  wire [0:0] CLBLM_R_X7Y124_SLICE_X9Y124_B1;
  wire [0:0] CLBLM_R_X7Y124_SLICE_X9Y124_B2;
  wire [0:0] CLBLM_R_X7Y124_SLICE_X9Y124_B3;
  wire [0:0] CLBLM_R_X7Y124_SLICE_X9Y124_B4;
  wire [0:0] CLBLM_R_X7Y124_SLICE_X9Y124_B5;
  wire [0:0] CLBLM_R_X7Y124_SLICE_X9Y124_B6;
  wire [0:0] CLBLM_R_X7Y124_SLICE_X9Y124_BO5;
  wire [0:0] CLBLM_R_X7Y124_SLICE_X9Y124_BO6;
  wire [0:0] CLBLM_R_X7Y124_SLICE_X9Y124_B_CY;
  wire [0:0] CLBLM_R_X7Y124_SLICE_X9Y124_B_XOR;
  wire [0:0] CLBLM_R_X7Y124_SLICE_X9Y124_C;
  wire [0:0] CLBLM_R_X7Y124_SLICE_X9Y124_C1;
  wire [0:0] CLBLM_R_X7Y124_SLICE_X9Y124_C2;
  wire [0:0] CLBLM_R_X7Y124_SLICE_X9Y124_C3;
  wire [0:0] CLBLM_R_X7Y124_SLICE_X9Y124_C4;
  wire [0:0] CLBLM_R_X7Y124_SLICE_X9Y124_C5;
  wire [0:0] CLBLM_R_X7Y124_SLICE_X9Y124_C6;
  wire [0:0] CLBLM_R_X7Y124_SLICE_X9Y124_CLK;
  wire [0:0] CLBLM_R_X7Y124_SLICE_X9Y124_CO5;
  wire [0:0] CLBLM_R_X7Y124_SLICE_X9Y124_CO6;
  wire [0:0] CLBLM_R_X7Y124_SLICE_X9Y124_C_CY;
  wire [0:0] CLBLM_R_X7Y124_SLICE_X9Y124_C_XOR;
  wire [0:0] CLBLM_R_X7Y124_SLICE_X9Y124_D;
  wire [0:0] CLBLM_R_X7Y124_SLICE_X9Y124_D1;
  wire [0:0] CLBLM_R_X7Y124_SLICE_X9Y124_D2;
  wire [0:0] CLBLM_R_X7Y124_SLICE_X9Y124_D3;
  wire [0:0] CLBLM_R_X7Y124_SLICE_X9Y124_D4;
  wire [0:0] CLBLM_R_X7Y124_SLICE_X9Y124_D5;
  wire [0:0] CLBLM_R_X7Y124_SLICE_X9Y124_D6;
  wire [0:0] CLBLM_R_X7Y124_SLICE_X9Y124_DO5;
  wire [0:0] CLBLM_R_X7Y124_SLICE_X9Y124_DO6;
  wire [0:0] CLBLM_R_X7Y124_SLICE_X9Y124_D_CY;
  wire [0:0] CLBLM_R_X7Y124_SLICE_X9Y124_D_XOR;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X8Y125_A;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X8Y125_A1;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X8Y125_A2;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X8Y125_A3;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X8Y125_A4;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X8Y125_A5;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X8Y125_A6;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X8Y125_AO5;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X8Y125_AO6;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X8Y125_A_CY;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X8Y125_A_XOR;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X8Y125_B;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X8Y125_B1;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X8Y125_B2;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X8Y125_B3;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X8Y125_B4;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X8Y125_B5;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X8Y125_B6;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X8Y125_BO5;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X8Y125_BO6;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X8Y125_B_CY;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X8Y125_B_XOR;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X8Y125_C;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X8Y125_C1;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X8Y125_C2;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X8Y125_C3;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X8Y125_C4;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X8Y125_C5;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X8Y125_C6;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X8Y125_CO5;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X8Y125_CO6;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X8Y125_C_CY;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X8Y125_C_XOR;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X8Y125_D;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X8Y125_D1;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X8Y125_D2;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X8Y125_D3;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X8Y125_D4;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X8Y125_D5;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X8Y125_D6;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X8Y125_DO5;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X8Y125_DO6;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X8Y125_D_CY;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X8Y125_D_XOR;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X9Y125_A;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X9Y125_A1;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X9Y125_A2;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X9Y125_A3;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X9Y125_A4;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X9Y125_A5;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X9Y125_A6;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X9Y125_AO5;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X9Y125_AO6;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X9Y125_A_CY;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X9Y125_A_XOR;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X9Y125_B;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X9Y125_B1;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X9Y125_B2;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X9Y125_B3;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X9Y125_B4;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X9Y125_B5;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X9Y125_B6;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X9Y125_BO5;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X9Y125_BO6;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X9Y125_B_CY;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X9Y125_B_XOR;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X9Y125_C;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X9Y125_C1;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X9Y125_C2;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X9Y125_C3;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X9Y125_C4;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X9Y125_C5;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X9Y125_C6;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X9Y125_CO5;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X9Y125_CO6;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X9Y125_C_CY;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X9Y125_C_XOR;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X9Y125_D;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X9Y125_D1;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X9Y125_D2;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X9Y125_D3;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X9Y125_D4;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X9Y125_D5;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X9Y125_D6;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X9Y125_DO5;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X9Y125_DO6;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X9Y125_D_CY;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X9Y125_D_XOR;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X8Y127_A;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X8Y127_A1;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X8Y127_A2;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X8Y127_A3;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X8Y127_A4;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X8Y127_A5;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X8Y127_A6;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X8Y127_AO5;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X8Y127_AO6;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X8Y127_AQ;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X8Y127_AX;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X8Y127_A_CY;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X8Y127_A_XOR;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X8Y127_B;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X8Y127_B1;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X8Y127_B2;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X8Y127_B3;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X8Y127_B4;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X8Y127_B5;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X8Y127_B6;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X8Y127_BO5;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X8Y127_BO6;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X8Y127_B_CY;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X8Y127_B_XOR;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X8Y127_C;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X8Y127_C1;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X8Y127_C2;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X8Y127_C3;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X8Y127_C4;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X8Y127_C5;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X8Y127_C6;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X8Y127_CLK;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X8Y127_CO5;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X8Y127_CO6;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X8Y127_C_CY;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X8Y127_C_XOR;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X8Y127_D;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X8Y127_D1;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X8Y127_D2;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X8Y127_D3;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X8Y127_D4;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X8Y127_D5;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X8Y127_D6;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X8Y127_DO5;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X8Y127_DO6;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X8Y127_D_CY;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X8Y127_D_XOR;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X9Y127_A;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X9Y127_A1;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X9Y127_A2;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X9Y127_A3;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X9Y127_A4;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X9Y127_A5;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X9Y127_A6;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X9Y127_AO5;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X9Y127_AO6;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X9Y127_A_CY;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X9Y127_A_XOR;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X9Y127_B;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X9Y127_B1;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X9Y127_B2;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X9Y127_B3;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X9Y127_B4;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X9Y127_B5;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X9Y127_B6;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X9Y127_BO5;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X9Y127_BO6;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X9Y127_B_CY;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X9Y127_B_XOR;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X9Y127_C;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X9Y127_C1;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X9Y127_C2;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X9Y127_C3;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X9Y127_C4;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X9Y127_C5;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X9Y127_C6;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X9Y127_CO5;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X9Y127_CO6;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X9Y127_C_CY;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X9Y127_C_XOR;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X9Y127_D;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X9Y127_D1;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X9Y127_D2;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X9Y127_D3;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X9Y127_D4;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X9Y127_D5;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X9Y127_D6;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X9Y127_DO5;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X9Y127_DO6;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X9Y127_D_CY;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X9Y127_D_XOR;
  wire [0:0] CLBLM_R_X7Y128_SLICE_X8Y128_A;
  wire [0:0] CLBLM_R_X7Y128_SLICE_X8Y128_A1;
  wire [0:0] CLBLM_R_X7Y128_SLICE_X8Y128_A2;
  wire [0:0] CLBLM_R_X7Y128_SLICE_X8Y128_A3;
  wire [0:0] CLBLM_R_X7Y128_SLICE_X8Y128_A4;
  wire [0:0] CLBLM_R_X7Y128_SLICE_X8Y128_A5;
  wire [0:0] CLBLM_R_X7Y128_SLICE_X8Y128_A6;
  wire [0:0] CLBLM_R_X7Y128_SLICE_X8Y128_AMUX;
  wire [0:0] CLBLM_R_X7Y128_SLICE_X8Y128_AO5;
  wire [0:0] CLBLM_R_X7Y128_SLICE_X8Y128_AO6;
  wire [0:0] CLBLM_R_X7Y128_SLICE_X8Y128_AQ;
  wire [0:0] CLBLM_R_X7Y128_SLICE_X8Y128_A_CY;
  wire [0:0] CLBLM_R_X7Y128_SLICE_X8Y128_A_XOR;
  wire [0:0] CLBLM_R_X7Y128_SLICE_X8Y128_B;
  wire [0:0] CLBLM_R_X7Y128_SLICE_X8Y128_B1;
  wire [0:0] CLBLM_R_X7Y128_SLICE_X8Y128_B2;
  wire [0:0] CLBLM_R_X7Y128_SLICE_X8Y128_B3;
  wire [0:0] CLBLM_R_X7Y128_SLICE_X8Y128_B4;
  wire [0:0] CLBLM_R_X7Y128_SLICE_X8Y128_B5;
  wire [0:0] CLBLM_R_X7Y128_SLICE_X8Y128_B6;
  wire [0:0] CLBLM_R_X7Y128_SLICE_X8Y128_BO5;
  wire [0:0] CLBLM_R_X7Y128_SLICE_X8Y128_BO6;
  wire [0:0] CLBLM_R_X7Y128_SLICE_X8Y128_B_CY;
  wire [0:0] CLBLM_R_X7Y128_SLICE_X8Y128_B_XOR;
  wire [0:0] CLBLM_R_X7Y128_SLICE_X8Y128_C;
  wire [0:0] CLBLM_R_X7Y128_SLICE_X8Y128_C1;
  wire [0:0] CLBLM_R_X7Y128_SLICE_X8Y128_C2;
  wire [0:0] CLBLM_R_X7Y128_SLICE_X8Y128_C3;
  wire [0:0] CLBLM_R_X7Y128_SLICE_X8Y128_C4;
  wire [0:0] CLBLM_R_X7Y128_SLICE_X8Y128_C5;
  wire [0:0] CLBLM_R_X7Y128_SLICE_X8Y128_C6;
  wire [0:0] CLBLM_R_X7Y128_SLICE_X8Y128_CLK;
  wire [0:0] CLBLM_R_X7Y128_SLICE_X8Y128_CO5;
  wire [0:0] CLBLM_R_X7Y128_SLICE_X8Y128_CO6;
  wire [0:0] CLBLM_R_X7Y128_SLICE_X8Y128_C_CY;
  wire [0:0] CLBLM_R_X7Y128_SLICE_X8Y128_C_XOR;
  wire [0:0] CLBLM_R_X7Y128_SLICE_X8Y128_D;
  wire [0:0] CLBLM_R_X7Y128_SLICE_X8Y128_D1;
  wire [0:0] CLBLM_R_X7Y128_SLICE_X8Y128_D2;
  wire [0:0] CLBLM_R_X7Y128_SLICE_X8Y128_D3;
  wire [0:0] CLBLM_R_X7Y128_SLICE_X8Y128_D4;
  wire [0:0] CLBLM_R_X7Y128_SLICE_X8Y128_D5;
  wire [0:0] CLBLM_R_X7Y128_SLICE_X8Y128_D6;
  wire [0:0] CLBLM_R_X7Y128_SLICE_X8Y128_DO5;
  wire [0:0] CLBLM_R_X7Y128_SLICE_X8Y128_DO6;
  wire [0:0] CLBLM_R_X7Y128_SLICE_X8Y128_D_CY;
  wire [0:0] CLBLM_R_X7Y128_SLICE_X8Y128_D_XOR;
  wire [0:0] CLBLM_R_X7Y128_SLICE_X9Y128_A;
  wire [0:0] CLBLM_R_X7Y128_SLICE_X9Y128_A1;
  wire [0:0] CLBLM_R_X7Y128_SLICE_X9Y128_A2;
  wire [0:0] CLBLM_R_X7Y128_SLICE_X9Y128_A3;
  wire [0:0] CLBLM_R_X7Y128_SLICE_X9Y128_A4;
  wire [0:0] CLBLM_R_X7Y128_SLICE_X9Y128_A5;
  wire [0:0] CLBLM_R_X7Y128_SLICE_X9Y128_A6;
  wire [0:0] CLBLM_R_X7Y128_SLICE_X9Y128_AO5;
  wire [0:0] CLBLM_R_X7Y128_SLICE_X9Y128_AO6;
  wire [0:0] CLBLM_R_X7Y128_SLICE_X9Y128_A_CY;
  wire [0:0] CLBLM_R_X7Y128_SLICE_X9Y128_A_XOR;
  wire [0:0] CLBLM_R_X7Y128_SLICE_X9Y128_B;
  wire [0:0] CLBLM_R_X7Y128_SLICE_X9Y128_B1;
  wire [0:0] CLBLM_R_X7Y128_SLICE_X9Y128_B2;
  wire [0:0] CLBLM_R_X7Y128_SLICE_X9Y128_B3;
  wire [0:0] CLBLM_R_X7Y128_SLICE_X9Y128_B4;
  wire [0:0] CLBLM_R_X7Y128_SLICE_X9Y128_B5;
  wire [0:0] CLBLM_R_X7Y128_SLICE_X9Y128_B6;
  wire [0:0] CLBLM_R_X7Y128_SLICE_X9Y128_BO5;
  wire [0:0] CLBLM_R_X7Y128_SLICE_X9Y128_BO6;
  wire [0:0] CLBLM_R_X7Y128_SLICE_X9Y128_B_CY;
  wire [0:0] CLBLM_R_X7Y128_SLICE_X9Y128_B_XOR;
  wire [0:0] CLBLM_R_X7Y128_SLICE_X9Y128_C;
  wire [0:0] CLBLM_R_X7Y128_SLICE_X9Y128_C1;
  wire [0:0] CLBLM_R_X7Y128_SLICE_X9Y128_C2;
  wire [0:0] CLBLM_R_X7Y128_SLICE_X9Y128_C3;
  wire [0:0] CLBLM_R_X7Y128_SLICE_X9Y128_C4;
  wire [0:0] CLBLM_R_X7Y128_SLICE_X9Y128_C5;
  wire [0:0] CLBLM_R_X7Y128_SLICE_X9Y128_C6;
  wire [0:0] CLBLM_R_X7Y128_SLICE_X9Y128_CO5;
  wire [0:0] CLBLM_R_X7Y128_SLICE_X9Y128_CO6;
  wire [0:0] CLBLM_R_X7Y128_SLICE_X9Y128_C_CY;
  wire [0:0] CLBLM_R_X7Y128_SLICE_X9Y128_C_XOR;
  wire [0:0] CLBLM_R_X7Y128_SLICE_X9Y128_D;
  wire [0:0] CLBLM_R_X7Y128_SLICE_X9Y128_D1;
  wire [0:0] CLBLM_R_X7Y128_SLICE_X9Y128_D2;
  wire [0:0] CLBLM_R_X7Y128_SLICE_X9Y128_D3;
  wire [0:0] CLBLM_R_X7Y128_SLICE_X9Y128_D4;
  wire [0:0] CLBLM_R_X7Y128_SLICE_X9Y128_D5;
  wire [0:0] CLBLM_R_X7Y128_SLICE_X9Y128_D6;
  wire [0:0] CLBLM_R_X7Y128_SLICE_X9Y128_DO5;
  wire [0:0] CLBLM_R_X7Y128_SLICE_X9Y128_DO6;
  wire [0:0] CLBLM_R_X7Y128_SLICE_X9Y128_D_CY;
  wire [0:0] CLBLM_R_X7Y128_SLICE_X9Y128_D_XOR;
  wire [0:0] CLBLM_R_X7Y151_SLICE_X8Y151_A;
  wire [0:0] CLBLM_R_X7Y151_SLICE_X8Y151_A1;
  wire [0:0] CLBLM_R_X7Y151_SLICE_X8Y151_A2;
  wire [0:0] CLBLM_R_X7Y151_SLICE_X8Y151_A3;
  wire [0:0] CLBLM_R_X7Y151_SLICE_X8Y151_A4;
  wire [0:0] CLBLM_R_X7Y151_SLICE_X8Y151_A5;
  wire [0:0] CLBLM_R_X7Y151_SLICE_X8Y151_A6;
  wire [0:0] CLBLM_R_X7Y151_SLICE_X8Y151_AO5;
  wire [0:0] CLBLM_R_X7Y151_SLICE_X8Y151_AO6;
  wire [0:0] CLBLM_R_X7Y151_SLICE_X8Y151_A_CY;
  wire [0:0] CLBLM_R_X7Y151_SLICE_X8Y151_A_XOR;
  wire [0:0] CLBLM_R_X7Y151_SLICE_X8Y151_B;
  wire [0:0] CLBLM_R_X7Y151_SLICE_X8Y151_B1;
  wire [0:0] CLBLM_R_X7Y151_SLICE_X8Y151_B2;
  wire [0:0] CLBLM_R_X7Y151_SLICE_X8Y151_B3;
  wire [0:0] CLBLM_R_X7Y151_SLICE_X8Y151_B4;
  wire [0:0] CLBLM_R_X7Y151_SLICE_X8Y151_B5;
  wire [0:0] CLBLM_R_X7Y151_SLICE_X8Y151_B6;
  wire [0:0] CLBLM_R_X7Y151_SLICE_X8Y151_BO5;
  wire [0:0] CLBLM_R_X7Y151_SLICE_X8Y151_BO6;
  wire [0:0] CLBLM_R_X7Y151_SLICE_X8Y151_B_CY;
  wire [0:0] CLBLM_R_X7Y151_SLICE_X8Y151_B_XOR;
  wire [0:0] CLBLM_R_X7Y151_SLICE_X8Y151_C;
  wire [0:0] CLBLM_R_X7Y151_SLICE_X8Y151_C1;
  wire [0:0] CLBLM_R_X7Y151_SLICE_X8Y151_C2;
  wire [0:0] CLBLM_R_X7Y151_SLICE_X8Y151_C3;
  wire [0:0] CLBLM_R_X7Y151_SLICE_X8Y151_C4;
  wire [0:0] CLBLM_R_X7Y151_SLICE_X8Y151_C5;
  wire [0:0] CLBLM_R_X7Y151_SLICE_X8Y151_C6;
  wire [0:0] CLBLM_R_X7Y151_SLICE_X8Y151_CO5;
  wire [0:0] CLBLM_R_X7Y151_SLICE_X8Y151_CO6;
  wire [0:0] CLBLM_R_X7Y151_SLICE_X8Y151_C_CY;
  wire [0:0] CLBLM_R_X7Y151_SLICE_X8Y151_C_XOR;
  wire [0:0] CLBLM_R_X7Y151_SLICE_X8Y151_D;
  wire [0:0] CLBLM_R_X7Y151_SLICE_X8Y151_D1;
  wire [0:0] CLBLM_R_X7Y151_SLICE_X8Y151_D2;
  wire [0:0] CLBLM_R_X7Y151_SLICE_X8Y151_D3;
  wire [0:0] CLBLM_R_X7Y151_SLICE_X8Y151_D4;
  wire [0:0] CLBLM_R_X7Y151_SLICE_X8Y151_D5;
  wire [0:0] CLBLM_R_X7Y151_SLICE_X8Y151_D6;
  wire [0:0] CLBLM_R_X7Y151_SLICE_X8Y151_DO5;
  wire [0:0] CLBLM_R_X7Y151_SLICE_X8Y151_DO6;
  wire [0:0] CLBLM_R_X7Y151_SLICE_X8Y151_D_CY;
  wire [0:0] CLBLM_R_X7Y151_SLICE_X8Y151_D_XOR;
  wire [0:0] CLBLM_R_X7Y151_SLICE_X9Y151_A;
  wire [0:0] CLBLM_R_X7Y151_SLICE_X9Y151_A1;
  wire [0:0] CLBLM_R_X7Y151_SLICE_X9Y151_A2;
  wire [0:0] CLBLM_R_X7Y151_SLICE_X9Y151_A3;
  wire [0:0] CLBLM_R_X7Y151_SLICE_X9Y151_A4;
  wire [0:0] CLBLM_R_X7Y151_SLICE_X9Y151_A5;
  wire [0:0] CLBLM_R_X7Y151_SLICE_X9Y151_A6;
  wire [0:0] CLBLM_R_X7Y151_SLICE_X9Y151_AO5;
  wire [0:0] CLBLM_R_X7Y151_SLICE_X9Y151_AO6;
  wire [0:0] CLBLM_R_X7Y151_SLICE_X9Y151_A_CY;
  wire [0:0] CLBLM_R_X7Y151_SLICE_X9Y151_A_XOR;
  wire [0:0] CLBLM_R_X7Y151_SLICE_X9Y151_B;
  wire [0:0] CLBLM_R_X7Y151_SLICE_X9Y151_B1;
  wire [0:0] CLBLM_R_X7Y151_SLICE_X9Y151_B2;
  wire [0:0] CLBLM_R_X7Y151_SLICE_X9Y151_B3;
  wire [0:0] CLBLM_R_X7Y151_SLICE_X9Y151_B4;
  wire [0:0] CLBLM_R_X7Y151_SLICE_X9Y151_B5;
  wire [0:0] CLBLM_R_X7Y151_SLICE_X9Y151_B6;
  wire [0:0] CLBLM_R_X7Y151_SLICE_X9Y151_BO5;
  wire [0:0] CLBLM_R_X7Y151_SLICE_X9Y151_BO6;
  wire [0:0] CLBLM_R_X7Y151_SLICE_X9Y151_B_CY;
  wire [0:0] CLBLM_R_X7Y151_SLICE_X9Y151_B_XOR;
  wire [0:0] CLBLM_R_X7Y151_SLICE_X9Y151_C;
  wire [0:0] CLBLM_R_X7Y151_SLICE_X9Y151_C1;
  wire [0:0] CLBLM_R_X7Y151_SLICE_X9Y151_C2;
  wire [0:0] CLBLM_R_X7Y151_SLICE_X9Y151_C3;
  wire [0:0] CLBLM_R_X7Y151_SLICE_X9Y151_C4;
  wire [0:0] CLBLM_R_X7Y151_SLICE_X9Y151_C5;
  wire [0:0] CLBLM_R_X7Y151_SLICE_X9Y151_C6;
  wire [0:0] CLBLM_R_X7Y151_SLICE_X9Y151_CO5;
  wire [0:0] CLBLM_R_X7Y151_SLICE_X9Y151_CO6;
  wire [0:0] CLBLM_R_X7Y151_SLICE_X9Y151_C_CY;
  wire [0:0] CLBLM_R_X7Y151_SLICE_X9Y151_C_XOR;
  wire [0:0] CLBLM_R_X7Y151_SLICE_X9Y151_D;
  wire [0:0] CLBLM_R_X7Y151_SLICE_X9Y151_D1;
  wire [0:0] CLBLM_R_X7Y151_SLICE_X9Y151_D2;
  wire [0:0] CLBLM_R_X7Y151_SLICE_X9Y151_D3;
  wire [0:0] CLBLM_R_X7Y151_SLICE_X9Y151_D4;
  wire [0:0] CLBLM_R_X7Y151_SLICE_X9Y151_D5;
  wire [0:0] CLBLM_R_X7Y151_SLICE_X9Y151_D6;
  wire [0:0] CLBLM_R_X7Y151_SLICE_X9Y151_DO5;
  wire [0:0] CLBLM_R_X7Y151_SLICE_X9Y151_DO6;
  wire [0:0] CLBLM_R_X7Y151_SLICE_X9Y151_D_CY;
  wire [0:0] CLBLM_R_X7Y151_SLICE_X9Y151_D_XOR;
  wire [0:0] CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_CE0;
  wire [0:0] CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_CE1;
  wire [0:0] CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_I0;
  wire [0:0] CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_I1;
  wire [0:0] CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_IGNORE0;
  wire [0:0] CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_IGNORE1;
  wire [0:0] CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_O;
  wire [0:0] CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_S0;
  wire [0:0] CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_S1;
  wire [0:0] CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_CE;
  wire [0:0] CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_I;
  wire [0:0] CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  wire [0:0] LIOB33_SING_X0Y100_IOB_X0Y100_O;
  wire [0:0] LIOB33_SING_X0Y149_IOB_X0Y149_O;
  wire [0:0] LIOB33_SING_X0Y150_IOB_X0Y150_O;
  wire [0:0] LIOB33_SING_X0Y199_IOB_X0Y199_O;
  wire [0:0] LIOB33_SING_X0Y50_IOB_X0Y50_I;
  wire [0:0] LIOB33_X0Y101_IOB_X0Y101_O;
  wire [0:0] LIOB33_X0Y101_IOB_X0Y102_O;
  wire [0:0] LIOB33_X0Y103_IOB_X0Y103_O;
  wire [0:0] LIOB33_X0Y103_IOB_X0Y104_O;
  wire [0:0] LIOB33_X0Y105_IOB_X0Y105_O;
  wire [0:0] LIOB33_X0Y105_IOB_X0Y106_O;
  wire [0:0] LIOB33_X0Y107_IOB_X0Y107_O;
  wire [0:0] LIOB33_X0Y107_IOB_X0Y108_O;
  wire [0:0] LIOB33_X0Y109_IOB_X0Y109_O;
  wire [0:0] LIOB33_X0Y109_IOB_X0Y110_O;
  wire [0:0] LIOB33_X0Y111_IOB_X0Y111_O;
  wire [0:0] LIOB33_X0Y111_IOB_X0Y112_O;
  wire [0:0] LIOB33_X0Y113_IOB_X0Y113_O;
  wire [0:0] LIOB33_X0Y113_IOB_X0Y114_O;
  wire [0:0] LIOB33_X0Y115_IOB_X0Y115_O;
  wire [0:0] LIOB33_X0Y115_IOB_X0Y116_O;
  wire [0:0] LIOB33_X0Y117_IOB_X0Y117_O;
  wire [0:0] LIOB33_X0Y117_IOB_X0Y118_O;
  wire [0:0] LIOB33_X0Y119_IOB_X0Y119_O;
  wire [0:0] LIOB33_X0Y119_IOB_X0Y120_O;
  wire [0:0] LIOB33_X0Y121_IOB_X0Y121_O;
  wire [0:0] LIOB33_X0Y121_IOB_X0Y122_O;
  wire [0:0] LIOB33_X0Y123_IOB_X0Y123_O;
  wire [0:0] LIOB33_X0Y123_IOB_X0Y124_O;
  wire [0:0] LIOB33_X0Y125_IOB_X0Y125_O;
  wire [0:0] LIOB33_X0Y125_IOB_X0Y126_O;
  wire [0:0] LIOB33_X0Y127_IOB_X0Y127_O;
  wire [0:0] LIOB33_X0Y127_IOB_X0Y128_O;
  wire [0:0] LIOB33_X0Y129_IOB_X0Y129_O;
  wire [0:0] LIOB33_X0Y129_IOB_X0Y130_O;
  wire [0:0] LIOB33_X0Y131_IOB_X0Y131_O;
  wire [0:0] LIOB33_X0Y131_IOB_X0Y132_O;
  wire [0:0] LIOB33_X0Y133_IOB_X0Y133_O;
  wire [0:0] LIOB33_X0Y133_IOB_X0Y134_O;
  wire [0:0] LIOB33_X0Y135_IOB_X0Y135_O;
  wire [0:0] LIOB33_X0Y135_IOB_X0Y136_O;
  wire [0:0] LIOB33_X0Y137_IOB_X0Y137_O;
  wire [0:0] LIOB33_X0Y137_IOB_X0Y138_O;
  wire [0:0] LIOB33_X0Y139_IOB_X0Y139_O;
  wire [0:0] LIOB33_X0Y139_IOB_X0Y140_O;
  wire [0:0] LIOB33_X0Y141_IOB_X0Y141_O;
  wire [0:0] LIOB33_X0Y141_IOB_X0Y142_O;
  wire [0:0] LIOB33_X0Y143_IOB_X0Y143_O;
  wire [0:0] LIOB33_X0Y145_IOB_X0Y145_O;
  wire [0:0] LIOB33_X0Y145_IOB_X0Y146_O;
  wire [0:0] LIOB33_X0Y147_IOB_X0Y147_O;
  wire [0:0] LIOB33_X0Y147_IOB_X0Y148_O;
  wire [0:0] LIOB33_X0Y151_IOB_X0Y151_O;
  wire [0:0] LIOB33_X0Y151_IOB_X0Y152_O;
  wire [0:0] LIOB33_X0Y153_IOB_X0Y153_O;
  wire [0:0] LIOB33_X0Y153_IOB_X0Y154_O;
  wire [0:0] LIOB33_X0Y155_IOB_X0Y155_O;
  wire [0:0] LIOB33_X0Y155_IOB_X0Y156_O;
  wire [0:0] LIOB33_X0Y157_IOB_X0Y157_O;
  wire [0:0] LIOB33_X0Y157_IOB_X0Y158_O;
  wire [0:0] LIOB33_X0Y159_IOB_X0Y159_O;
  wire [0:0] LIOB33_X0Y159_IOB_X0Y160_O;
  wire [0:0] LIOB33_X0Y161_IOB_X0Y161_O;
  wire [0:0] LIOB33_X0Y161_IOB_X0Y162_O;
  wire [0:0] LIOB33_X0Y163_IOB_X0Y163_O;
  wire [0:0] LIOB33_X0Y163_IOB_X0Y164_O;
  wire [0:0] LIOB33_X0Y165_IOB_X0Y165_O;
  wire [0:0] LIOB33_X0Y165_IOB_X0Y166_O;
  wire [0:0] LIOB33_X0Y167_IOB_X0Y167_O;
  wire [0:0] LIOB33_X0Y167_IOB_X0Y168_O;
  wire [0:0] LIOB33_X0Y169_IOB_X0Y169_O;
  wire [0:0] LIOB33_X0Y169_IOB_X0Y170_O;
  wire [0:0] LIOB33_X0Y171_IOB_X0Y171_O;
  wire [0:0] LIOB33_X0Y171_IOB_X0Y172_O;
  wire [0:0] LIOB33_X0Y173_IOB_X0Y173_O;
  wire [0:0] LIOB33_X0Y173_IOB_X0Y174_O;
  wire [0:0] LIOB33_X0Y175_IOB_X0Y175_O;
  wire [0:0] LIOB33_X0Y175_IOB_X0Y176_O;
  wire [0:0] LIOB33_X0Y177_IOB_X0Y177_O;
  wire [0:0] LIOB33_X0Y177_IOB_X0Y178_O;
  wire [0:0] LIOB33_X0Y179_IOB_X0Y179_O;
  wire [0:0] LIOB33_X0Y179_IOB_X0Y180_O;
  wire [0:0] LIOB33_X0Y181_IOB_X0Y181_O;
  wire [0:0] LIOB33_X0Y181_IOB_X0Y182_O;
  wire [0:0] LIOB33_X0Y183_IOB_X0Y183_O;
  wire [0:0] LIOB33_X0Y183_IOB_X0Y184_O;
  wire [0:0] LIOB33_X0Y185_IOB_X0Y185_O;
  wire [0:0] LIOB33_X0Y185_IOB_X0Y186_O;
  wire [0:0] LIOB33_X0Y187_IOB_X0Y187_O;
  wire [0:0] LIOB33_X0Y187_IOB_X0Y188_O;
  wire [0:0] LIOB33_X0Y189_IOB_X0Y189_O;
  wire [0:0] LIOB33_X0Y189_IOB_X0Y190_O;
  wire [0:0] LIOB33_X0Y191_IOB_X0Y191_O;
  wire [0:0] LIOB33_X0Y191_IOB_X0Y192_O;
  wire [0:0] LIOB33_X0Y193_IOB_X0Y193_O;
  wire [0:0] LIOB33_X0Y193_IOB_X0Y194_O;
  wire [0:0] LIOB33_X0Y195_IOB_X0Y195_O;
  wire [0:0] LIOB33_X0Y195_IOB_X0Y196_O;
  wire [0:0] LIOB33_X0Y197_IOB_X0Y197_O;
  wire [0:0] LIOB33_X0Y197_IOB_X0Y198_O;
  wire [0:0] LIOB33_X0Y51_IOB_X0Y51_I;
  wire [0:0] LIOB33_X0Y51_IOB_X0Y52_I;
  wire [0:0] LIOB33_X0Y53_IOB_X0Y53_I;
  wire [0:0] LIOB33_X0Y53_IOB_X0Y54_I;
  wire [0:0] LIOB33_X0Y55_IOB_X0Y55_I;
  wire [0:0] LIOB33_X0Y55_IOB_X0Y56_I;
  wire [0:0] LIOB33_X0Y57_IOB_X0Y57_I;
  wire [0:0] LIOB33_X0Y57_IOB_X0Y58_I;
  wire [0:0] LIOB33_X0Y59_IOB_X0Y59_I;
  wire [0:0] LIOB33_X0Y59_IOB_X0Y60_I;
  wire [0:0] LIOB33_X0Y61_IOB_X0Y61_I;
  wire [0:0] LIOB33_X0Y61_IOB_X0Y62_I;
  wire [0:0] LIOB33_X0Y63_IOB_X0Y63_I;
  wire [0:0] LIOB33_X0Y63_IOB_X0Y64_I;
  wire [0:0] LIOB33_X0Y65_IOB_X0Y65_I;
  wire [0:0] LIOB33_X0Y65_IOB_X0Y66_I;
  wire [0:0] LIOB33_X0Y67_IOB_X0Y67_I;
  wire [0:0] LIOB33_X0Y67_IOB_X0Y68_I;
  wire [0:0] LIOB33_X0Y69_IOB_X0Y69_I;
  wire [0:0] LIOB33_X0Y69_IOB_X0Y70_I;
  wire [0:0] LIOB33_X0Y71_IOB_X0Y71_I;
  wire [0:0] LIOB33_X0Y71_IOB_X0Y72_I;
  wire [0:0] LIOB33_X0Y73_IOB_X0Y73_I;
  wire [0:0] LIOB33_X0Y73_IOB_X0Y74_I;
  wire [0:0] LIOB33_X0Y75_IOB_X0Y75_I;
  wire [0:0] LIOB33_X0Y75_IOB_X0Y76_I;
  wire [0:0] LIOB33_X0Y77_IOB_X0Y77_I;
  wire [0:0] LIOB33_X0Y77_IOB_X0Y78_I;
  wire [0:0] LIOB33_X0Y79_IOB_X0Y79_I;
  wire [0:0] LIOB33_X0Y79_IOB_X0Y80_O;
  wire [0:0] LIOI3_SING_X0Y100_OLOGIC_X0Y100_D1;
  wire [0:0] LIOI3_SING_X0Y100_OLOGIC_X0Y100_OQ;
  wire [0:0] LIOI3_SING_X0Y100_OLOGIC_X0Y100_T1;
  wire [0:0] LIOI3_SING_X0Y100_OLOGIC_X0Y100_TQ;
  wire [0:0] LIOI3_SING_X0Y149_OLOGIC_X0Y149_D1;
  wire [0:0] LIOI3_SING_X0Y149_OLOGIC_X0Y149_OQ;
  wire [0:0] LIOI3_SING_X0Y149_OLOGIC_X0Y149_T1;
  wire [0:0] LIOI3_SING_X0Y149_OLOGIC_X0Y149_TQ;
  wire [0:0] LIOI3_SING_X0Y150_OLOGIC_X0Y150_D1;
  wire [0:0] LIOI3_SING_X0Y150_OLOGIC_X0Y150_OQ;
  wire [0:0] LIOI3_SING_X0Y150_OLOGIC_X0Y150_T1;
  wire [0:0] LIOI3_SING_X0Y150_OLOGIC_X0Y150_TQ;
  wire [0:0] LIOI3_SING_X0Y199_OLOGIC_X0Y199_D1;
  wire [0:0] LIOI3_SING_X0Y199_OLOGIC_X0Y199_OQ;
  wire [0:0] LIOI3_SING_X0Y199_OLOGIC_X0Y199_T1;
  wire [0:0] LIOI3_SING_X0Y199_OLOGIC_X0Y199_TQ;
  wire [0:0] LIOI3_SING_X0Y50_ILOGIC_X0Y50_D;
  wire [0:0] LIOI3_SING_X0Y50_ILOGIC_X0Y50_O;
  wire [0:0] LIOI3_TBYTESRC_X0Y107_OLOGIC_X0Y107_D1;
  wire [0:0] LIOI3_TBYTESRC_X0Y107_OLOGIC_X0Y107_OQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y107_OLOGIC_X0Y107_T1;
  wire [0:0] LIOI3_TBYTESRC_X0Y107_OLOGIC_X0Y107_TQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y107_OLOGIC_X0Y108_D1;
  wire [0:0] LIOI3_TBYTESRC_X0Y107_OLOGIC_X0Y108_OQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y107_OLOGIC_X0Y108_T1;
  wire [0:0] LIOI3_TBYTESRC_X0Y107_OLOGIC_X0Y108_TQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y119_OLOGIC_X0Y119_D1;
  wire [0:0] LIOI3_TBYTESRC_X0Y119_OLOGIC_X0Y119_OQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y119_OLOGIC_X0Y119_T1;
  wire [0:0] LIOI3_TBYTESRC_X0Y119_OLOGIC_X0Y119_TQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y119_OLOGIC_X0Y120_D1;
  wire [0:0] LIOI3_TBYTESRC_X0Y119_OLOGIC_X0Y120_OQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y119_OLOGIC_X0Y120_T1;
  wire [0:0] LIOI3_TBYTESRC_X0Y119_OLOGIC_X0Y120_TQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y131_OLOGIC_X0Y131_D1;
  wire [0:0] LIOI3_TBYTESRC_X0Y131_OLOGIC_X0Y131_OQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y131_OLOGIC_X0Y131_T1;
  wire [0:0] LIOI3_TBYTESRC_X0Y131_OLOGIC_X0Y131_TQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y131_OLOGIC_X0Y132_D1;
  wire [0:0] LIOI3_TBYTESRC_X0Y131_OLOGIC_X0Y132_OQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y131_OLOGIC_X0Y132_T1;
  wire [0:0] LIOI3_TBYTESRC_X0Y131_OLOGIC_X0Y132_TQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y143_OLOGIC_X0Y143_D1;
  wire [0:0] LIOI3_TBYTESRC_X0Y143_OLOGIC_X0Y143_OQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y143_OLOGIC_X0Y143_T1;
  wire [0:0] LIOI3_TBYTESRC_X0Y143_OLOGIC_X0Y143_TQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y143_OLOGIC_X0Y144_D1;
  wire [0:0] LIOI3_TBYTESRC_X0Y143_OLOGIC_X0Y144_OQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y143_OLOGIC_X0Y144_T1;
  wire [0:0] LIOI3_TBYTESRC_X0Y143_OLOGIC_X0Y144_TQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y157_OLOGIC_X0Y157_D1;
  wire [0:0] LIOI3_TBYTESRC_X0Y157_OLOGIC_X0Y157_OQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y157_OLOGIC_X0Y157_T1;
  wire [0:0] LIOI3_TBYTESRC_X0Y157_OLOGIC_X0Y157_TQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y157_OLOGIC_X0Y158_D1;
  wire [0:0] LIOI3_TBYTESRC_X0Y157_OLOGIC_X0Y158_OQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y157_OLOGIC_X0Y158_T1;
  wire [0:0] LIOI3_TBYTESRC_X0Y157_OLOGIC_X0Y158_TQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y169_OLOGIC_X0Y169_D1;
  wire [0:0] LIOI3_TBYTESRC_X0Y169_OLOGIC_X0Y169_OQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y169_OLOGIC_X0Y169_T1;
  wire [0:0] LIOI3_TBYTESRC_X0Y169_OLOGIC_X0Y169_TQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y169_OLOGIC_X0Y170_D1;
  wire [0:0] LIOI3_TBYTESRC_X0Y169_OLOGIC_X0Y170_OQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y169_OLOGIC_X0Y170_T1;
  wire [0:0] LIOI3_TBYTESRC_X0Y169_OLOGIC_X0Y170_TQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y181_OLOGIC_X0Y181_D1;
  wire [0:0] LIOI3_TBYTESRC_X0Y181_OLOGIC_X0Y181_OQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y181_OLOGIC_X0Y181_T1;
  wire [0:0] LIOI3_TBYTESRC_X0Y181_OLOGIC_X0Y181_TQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y181_OLOGIC_X0Y182_D1;
  wire [0:0] LIOI3_TBYTESRC_X0Y181_OLOGIC_X0Y182_OQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y181_OLOGIC_X0Y182_T1;
  wire [0:0] LIOI3_TBYTESRC_X0Y181_OLOGIC_X0Y182_TQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y193_OLOGIC_X0Y193_D1;
  wire [0:0] LIOI3_TBYTESRC_X0Y193_OLOGIC_X0Y193_OQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y193_OLOGIC_X0Y193_T1;
  wire [0:0] LIOI3_TBYTESRC_X0Y193_OLOGIC_X0Y193_TQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y193_OLOGIC_X0Y194_D1;
  wire [0:0] LIOI3_TBYTESRC_X0Y193_OLOGIC_X0Y194_OQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y193_OLOGIC_X0Y194_T1;
  wire [0:0] LIOI3_TBYTESRC_X0Y193_OLOGIC_X0Y194_TQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y57_ILOGIC_X0Y57_D;
  wire [0:0] LIOI3_TBYTESRC_X0Y57_ILOGIC_X0Y57_O;
  wire [0:0] LIOI3_TBYTESRC_X0Y57_ILOGIC_X0Y58_D;
  wire [0:0] LIOI3_TBYTESRC_X0Y57_ILOGIC_X0Y58_O;
  wire [0:0] LIOI3_TBYTESRC_X0Y69_ILOGIC_X0Y69_D;
  wire [0:0] LIOI3_TBYTESRC_X0Y69_ILOGIC_X0Y69_O;
  wire [0:0] LIOI3_TBYTESRC_X0Y69_ILOGIC_X0Y70_D;
  wire [0:0] LIOI3_TBYTESRC_X0Y69_ILOGIC_X0Y70_O;
  wire [0:0] LIOI3_TBYTETERM_X0Y113_OLOGIC_X0Y113_D1;
  wire [0:0] LIOI3_TBYTETERM_X0Y113_OLOGIC_X0Y113_OQ;
  wire [0:0] LIOI3_TBYTETERM_X0Y113_OLOGIC_X0Y113_T1;
  wire [0:0] LIOI3_TBYTETERM_X0Y113_OLOGIC_X0Y113_TQ;
  wire [0:0] LIOI3_TBYTETERM_X0Y113_OLOGIC_X0Y114_D1;
  wire [0:0] LIOI3_TBYTETERM_X0Y113_OLOGIC_X0Y114_OQ;
  wire [0:0] LIOI3_TBYTETERM_X0Y113_OLOGIC_X0Y114_T1;
  wire [0:0] LIOI3_TBYTETERM_X0Y113_OLOGIC_X0Y114_TQ;
  wire [0:0] LIOI3_TBYTETERM_X0Y137_OLOGIC_X0Y137_D1;
  wire [0:0] LIOI3_TBYTETERM_X0Y137_OLOGIC_X0Y137_OQ;
  wire [0:0] LIOI3_TBYTETERM_X0Y137_OLOGIC_X0Y137_T1;
  wire [0:0] LIOI3_TBYTETERM_X0Y137_OLOGIC_X0Y137_TQ;
  wire [0:0] LIOI3_TBYTETERM_X0Y137_OLOGIC_X0Y138_D1;
  wire [0:0] LIOI3_TBYTETERM_X0Y137_OLOGIC_X0Y138_OQ;
  wire [0:0] LIOI3_TBYTETERM_X0Y137_OLOGIC_X0Y138_T1;
  wire [0:0] LIOI3_TBYTETERM_X0Y137_OLOGIC_X0Y138_TQ;
  wire [0:0] LIOI3_TBYTETERM_X0Y163_OLOGIC_X0Y163_D1;
  wire [0:0] LIOI3_TBYTETERM_X0Y163_OLOGIC_X0Y163_OQ;
  wire [0:0] LIOI3_TBYTETERM_X0Y163_OLOGIC_X0Y163_T1;
  wire [0:0] LIOI3_TBYTETERM_X0Y163_OLOGIC_X0Y163_TQ;
  wire [0:0] LIOI3_TBYTETERM_X0Y163_OLOGIC_X0Y164_D1;
  wire [0:0] LIOI3_TBYTETERM_X0Y163_OLOGIC_X0Y164_OQ;
  wire [0:0] LIOI3_TBYTETERM_X0Y163_OLOGIC_X0Y164_T1;
  wire [0:0] LIOI3_TBYTETERM_X0Y163_OLOGIC_X0Y164_TQ;
  wire [0:0] LIOI3_TBYTETERM_X0Y187_OLOGIC_X0Y187_D1;
  wire [0:0] LIOI3_TBYTETERM_X0Y187_OLOGIC_X0Y187_OQ;
  wire [0:0] LIOI3_TBYTETERM_X0Y187_OLOGIC_X0Y187_T1;
  wire [0:0] LIOI3_TBYTETERM_X0Y187_OLOGIC_X0Y187_TQ;
  wire [0:0] LIOI3_TBYTETERM_X0Y187_OLOGIC_X0Y188_D1;
  wire [0:0] LIOI3_TBYTETERM_X0Y187_OLOGIC_X0Y188_OQ;
  wire [0:0] LIOI3_TBYTETERM_X0Y187_OLOGIC_X0Y188_T1;
  wire [0:0] LIOI3_TBYTETERM_X0Y187_OLOGIC_X0Y188_TQ;
  wire [0:0] LIOI3_TBYTETERM_X0Y63_ILOGIC_X0Y63_D;
  wire [0:0] LIOI3_TBYTETERM_X0Y63_ILOGIC_X0Y63_O;
  wire [0:0] LIOI3_TBYTETERM_X0Y63_ILOGIC_X0Y64_D;
  wire [0:0] LIOI3_TBYTETERM_X0Y63_ILOGIC_X0Y64_O;
  wire [0:0] LIOI3_X0Y101_OLOGIC_X0Y101_D1;
  wire [0:0] LIOI3_X0Y101_OLOGIC_X0Y101_OQ;
  wire [0:0] LIOI3_X0Y101_OLOGIC_X0Y101_T1;
  wire [0:0] LIOI3_X0Y101_OLOGIC_X0Y101_TQ;
  wire [0:0] LIOI3_X0Y101_OLOGIC_X0Y102_D1;
  wire [0:0] LIOI3_X0Y101_OLOGIC_X0Y102_OQ;
  wire [0:0] LIOI3_X0Y101_OLOGIC_X0Y102_T1;
  wire [0:0] LIOI3_X0Y101_OLOGIC_X0Y102_TQ;
  wire [0:0] LIOI3_X0Y103_OLOGIC_X0Y103_D1;
  wire [0:0] LIOI3_X0Y103_OLOGIC_X0Y103_OQ;
  wire [0:0] LIOI3_X0Y103_OLOGIC_X0Y103_T1;
  wire [0:0] LIOI3_X0Y103_OLOGIC_X0Y103_TQ;
  wire [0:0] LIOI3_X0Y103_OLOGIC_X0Y104_D1;
  wire [0:0] LIOI3_X0Y103_OLOGIC_X0Y104_OQ;
  wire [0:0] LIOI3_X0Y103_OLOGIC_X0Y104_T1;
  wire [0:0] LIOI3_X0Y103_OLOGIC_X0Y104_TQ;
  wire [0:0] LIOI3_X0Y105_OLOGIC_X0Y105_D1;
  wire [0:0] LIOI3_X0Y105_OLOGIC_X0Y105_OQ;
  wire [0:0] LIOI3_X0Y105_OLOGIC_X0Y105_T1;
  wire [0:0] LIOI3_X0Y105_OLOGIC_X0Y105_TQ;
  wire [0:0] LIOI3_X0Y105_OLOGIC_X0Y106_D1;
  wire [0:0] LIOI3_X0Y105_OLOGIC_X0Y106_OQ;
  wire [0:0] LIOI3_X0Y105_OLOGIC_X0Y106_T1;
  wire [0:0] LIOI3_X0Y105_OLOGIC_X0Y106_TQ;
  wire [0:0] LIOI3_X0Y109_OLOGIC_X0Y109_D1;
  wire [0:0] LIOI3_X0Y109_OLOGIC_X0Y109_OQ;
  wire [0:0] LIOI3_X0Y109_OLOGIC_X0Y109_T1;
  wire [0:0] LIOI3_X0Y109_OLOGIC_X0Y109_TQ;
  wire [0:0] LIOI3_X0Y109_OLOGIC_X0Y110_D1;
  wire [0:0] LIOI3_X0Y109_OLOGIC_X0Y110_OQ;
  wire [0:0] LIOI3_X0Y109_OLOGIC_X0Y110_T1;
  wire [0:0] LIOI3_X0Y109_OLOGIC_X0Y110_TQ;
  wire [0:0] LIOI3_X0Y111_OLOGIC_X0Y111_D1;
  wire [0:0] LIOI3_X0Y111_OLOGIC_X0Y111_OQ;
  wire [0:0] LIOI3_X0Y111_OLOGIC_X0Y111_T1;
  wire [0:0] LIOI3_X0Y111_OLOGIC_X0Y111_TQ;
  wire [0:0] LIOI3_X0Y111_OLOGIC_X0Y112_D1;
  wire [0:0] LIOI3_X0Y111_OLOGIC_X0Y112_OQ;
  wire [0:0] LIOI3_X0Y111_OLOGIC_X0Y112_T1;
  wire [0:0] LIOI3_X0Y111_OLOGIC_X0Y112_TQ;
  wire [0:0] LIOI3_X0Y115_OLOGIC_X0Y115_D1;
  wire [0:0] LIOI3_X0Y115_OLOGIC_X0Y115_OQ;
  wire [0:0] LIOI3_X0Y115_OLOGIC_X0Y115_T1;
  wire [0:0] LIOI3_X0Y115_OLOGIC_X0Y115_TQ;
  wire [0:0] LIOI3_X0Y115_OLOGIC_X0Y116_D1;
  wire [0:0] LIOI3_X0Y115_OLOGIC_X0Y116_OQ;
  wire [0:0] LIOI3_X0Y115_OLOGIC_X0Y116_T1;
  wire [0:0] LIOI3_X0Y115_OLOGIC_X0Y116_TQ;
  wire [0:0] LIOI3_X0Y117_OLOGIC_X0Y117_D1;
  wire [0:0] LIOI3_X0Y117_OLOGIC_X0Y117_OQ;
  wire [0:0] LIOI3_X0Y117_OLOGIC_X0Y117_T1;
  wire [0:0] LIOI3_X0Y117_OLOGIC_X0Y117_TQ;
  wire [0:0] LIOI3_X0Y117_OLOGIC_X0Y118_D1;
  wire [0:0] LIOI3_X0Y117_OLOGIC_X0Y118_OQ;
  wire [0:0] LIOI3_X0Y117_OLOGIC_X0Y118_T1;
  wire [0:0] LIOI3_X0Y117_OLOGIC_X0Y118_TQ;
  wire [0:0] LIOI3_X0Y121_OLOGIC_X0Y121_D1;
  wire [0:0] LIOI3_X0Y121_OLOGIC_X0Y121_OQ;
  wire [0:0] LIOI3_X0Y121_OLOGIC_X0Y121_T1;
  wire [0:0] LIOI3_X0Y121_OLOGIC_X0Y121_TQ;
  wire [0:0] LIOI3_X0Y121_OLOGIC_X0Y122_D1;
  wire [0:0] LIOI3_X0Y121_OLOGIC_X0Y122_OQ;
  wire [0:0] LIOI3_X0Y121_OLOGIC_X0Y122_T1;
  wire [0:0] LIOI3_X0Y121_OLOGIC_X0Y122_TQ;
  wire [0:0] LIOI3_X0Y123_OLOGIC_X0Y123_D1;
  wire [0:0] LIOI3_X0Y123_OLOGIC_X0Y123_OQ;
  wire [0:0] LIOI3_X0Y123_OLOGIC_X0Y123_T1;
  wire [0:0] LIOI3_X0Y123_OLOGIC_X0Y123_TQ;
  wire [0:0] LIOI3_X0Y123_OLOGIC_X0Y124_D1;
  wire [0:0] LIOI3_X0Y123_OLOGIC_X0Y124_OQ;
  wire [0:0] LIOI3_X0Y123_OLOGIC_X0Y124_T1;
  wire [0:0] LIOI3_X0Y123_OLOGIC_X0Y124_TQ;
  wire [0:0] LIOI3_X0Y125_OLOGIC_X0Y125_D1;
  wire [0:0] LIOI3_X0Y125_OLOGIC_X0Y125_OQ;
  wire [0:0] LIOI3_X0Y125_OLOGIC_X0Y125_T1;
  wire [0:0] LIOI3_X0Y125_OLOGIC_X0Y125_TQ;
  wire [0:0] LIOI3_X0Y125_OLOGIC_X0Y126_D1;
  wire [0:0] LIOI3_X0Y125_OLOGIC_X0Y126_OQ;
  wire [0:0] LIOI3_X0Y125_OLOGIC_X0Y126_T1;
  wire [0:0] LIOI3_X0Y125_OLOGIC_X0Y126_TQ;
  wire [0:0] LIOI3_X0Y127_OLOGIC_X0Y127_D1;
  wire [0:0] LIOI3_X0Y127_OLOGIC_X0Y127_OQ;
  wire [0:0] LIOI3_X0Y127_OLOGIC_X0Y127_T1;
  wire [0:0] LIOI3_X0Y127_OLOGIC_X0Y127_TQ;
  wire [0:0] LIOI3_X0Y127_OLOGIC_X0Y128_D1;
  wire [0:0] LIOI3_X0Y127_OLOGIC_X0Y128_OQ;
  wire [0:0] LIOI3_X0Y127_OLOGIC_X0Y128_T1;
  wire [0:0] LIOI3_X0Y127_OLOGIC_X0Y128_TQ;
  wire [0:0] LIOI3_X0Y129_OLOGIC_X0Y129_D1;
  wire [0:0] LIOI3_X0Y129_OLOGIC_X0Y129_OQ;
  wire [0:0] LIOI3_X0Y129_OLOGIC_X0Y129_T1;
  wire [0:0] LIOI3_X0Y129_OLOGIC_X0Y129_TQ;
  wire [0:0] LIOI3_X0Y129_OLOGIC_X0Y130_D1;
  wire [0:0] LIOI3_X0Y129_OLOGIC_X0Y130_OQ;
  wire [0:0] LIOI3_X0Y129_OLOGIC_X0Y130_T1;
  wire [0:0] LIOI3_X0Y129_OLOGIC_X0Y130_TQ;
  wire [0:0] LIOI3_X0Y133_OLOGIC_X0Y133_D1;
  wire [0:0] LIOI3_X0Y133_OLOGIC_X0Y133_OQ;
  wire [0:0] LIOI3_X0Y133_OLOGIC_X0Y133_T1;
  wire [0:0] LIOI3_X0Y133_OLOGIC_X0Y133_TQ;
  wire [0:0] LIOI3_X0Y133_OLOGIC_X0Y134_D1;
  wire [0:0] LIOI3_X0Y133_OLOGIC_X0Y134_OQ;
  wire [0:0] LIOI3_X0Y133_OLOGIC_X0Y134_T1;
  wire [0:0] LIOI3_X0Y133_OLOGIC_X0Y134_TQ;
  wire [0:0] LIOI3_X0Y135_OLOGIC_X0Y135_D1;
  wire [0:0] LIOI3_X0Y135_OLOGIC_X0Y135_OQ;
  wire [0:0] LIOI3_X0Y135_OLOGIC_X0Y135_T1;
  wire [0:0] LIOI3_X0Y135_OLOGIC_X0Y135_TQ;
  wire [0:0] LIOI3_X0Y135_OLOGIC_X0Y136_D1;
  wire [0:0] LIOI3_X0Y135_OLOGIC_X0Y136_OQ;
  wire [0:0] LIOI3_X0Y135_OLOGIC_X0Y136_T1;
  wire [0:0] LIOI3_X0Y135_OLOGIC_X0Y136_TQ;
  wire [0:0] LIOI3_X0Y139_OLOGIC_X0Y139_D1;
  wire [0:0] LIOI3_X0Y139_OLOGIC_X0Y139_OQ;
  wire [0:0] LIOI3_X0Y139_OLOGIC_X0Y139_T1;
  wire [0:0] LIOI3_X0Y139_OLOGIC_X0Y139_TQ;
  wire [0:0] LIOI3_X0Y139_OLOGIC_X0Y140_D1;
  wire [0:0] LIOI3_X0Y139_OLOGIC_X0Y140_OQ;
  wire [0:0] LIOI3_X0Y139_OLOGIC_X0Y140_T1;
  wire [0:0] LIOI3_X0Y139_OLOGIC_X0Y140_TQ;
  wire [0:0] LIOI3_X0Y141_OLOGIC_X0Y141_D1;
  wire [0:0] LIOI3_X0Y141_OLOGIC_X0Y141_OQ;
  wire [0:0] LIOI3_X0Y141_OLOGIC_X0Y141_T1;
  wire [0:0] LIOI3_X0Y141_OLOGIC_X0Y141_TQ;
  wire [0:0] LIOI3_X0Y141_OLOGIC_X0Y142_D1;
  wire [0:0] LIOI3_X0Y141_OLOGIC_X0Y142_OQ;
  wire [0:0] LIOI3_X0Y141_OLOGIC_X0Y142_T1;
  wire [0:0] LIOI3_X0Y141_OLOGIC_X0Y142_TQ;
  wire [0:0] LIOI3_X0Y145_OLOGIC_X0Y145_D1;
  wire [0:0] LIOI3_X0Y145_OLOGIC_X0Y145_OQ;
  wire [0:0] LIOI3_X0Y145_OLOGIC_X0Y145_T1;
  wire [0:0] LIOI3_X0Y145_OLOGIC_X0Y145_TQ;
  wire [0:0] LIOI3_X0Y145_OLOGIC_X0Y146_D1;
  wire [0:0] LIOI3_X0Y145_OLOGIC_X0Y146_OQ;
  wire [0:0] LIOI3_X0Y145_OLOGIC_X0Y146_T1;
  wire [0:0] LIOI3_X0Y145_OLOGIC_X0Y146_TQ;
  wire [0:0] LIOI3_X0Y147_OLOGIC_X0Y147_D1;
  wire [0:0] LIOI3_X0Y147_OLOGIC_X0Y147_OQ;
  wire [0:0] LIOI3_X0Y147_OLOGIC_X0Y147_T1;
  wire [0:0] LIOI3_X0Y147_OLOGIC_X0Y147_TQ;
  wire [0:0] LIOI3_X0Y147_OLOGIC_X0Y148_D1;
  wire [0:0] LIOI3_X0Y147_OLOGIC_X0Y148_OQ;
  wire [0:0] LIOI3_X0Y147_OLOGIC_X0Y148_T1;
  wire [0:0] LIOI3_X0Y147_OLOGIC_X0Y148_TQ;
  wire [0:0] LIOI3_X0Y151_OLOGIC_X0Y151_D1;
  wire [0:0] LIOI3_X0Y151_OLOGIC_X0Y151_OQ;
  wire [0:0] LIOI3_X0Y151_OLOGIC_X0Y151_T1;
  wire [0:0] LIOI3_X0Y151_OLOGIC_X0Y151_TQ;
  wire [0:0] LIOI3_X0Y151_OLOGIC_X0Y152_D1;
  wire [0:0] LIOI3_X0Y151_OLOGIC_X0Y152_OQ;
  wire [0:0] LIOI3_X0Y151_OLOGIC_X0Y152_T1;
  wire [0:0] LIOI3_X0Y151_OLOGIC_X0Y152_TQ;
  wire [0:0] LIOI3_X0Y153_OLOGIC_X0Y153_D1;
  wire [0:0] LIOI3_X0Y153_OLOGIC_X0Y153_OQ;
  wire [0:0] LIOI3_X0Y153_OLOGIC_X0Y153_T1;
  wire [0:0] LIOI3_X0Y153_OLOGIC_X0Y153_TQ;
  wire [0:0] LIOI3_X0Y153_OLOGIC_X0Y154_D1;
  wire [0:0] LIOI3_X0Y153_OLOGIC_X0Y154_OQ;
  wire [0:0] LIOI3_X0Y153_OLOGIC_X0Y154_T1;
  wire [0:0] LIOI3_X0Y153_OLOGIC_X0Y154_TQ;
  wire [0:0] LIOI3_X0Y155_OLOGIC_X0Y155_D1;
  wire [0:0] LIOI3_X0Y155_OLOGIC_X0Y155_OQ;
  wire [0:0] LIOI3_X0Y155_OLOGIC_X0Y155_T1;
  wire [0:0] LIOI3_X0Y155_OLOGIC_X0Y155_TQ;
  wire [0:0] LIOI3_X0Y155_OLOGIC_X0Y156_D1;
  wire [0:0] LIOI3_X0Y155_OLOGIC_X0Y156_OQ;
  wire [0:0] LIOI3_X0Y155_OLOGIC_X0Y156_T1;
  wire [0:0] LIOI3_X0Y155_OLOGIC_X0Y156_TQ;
  wire [0:0] LIOI3_X0Y159_OLOGIC_X0Y159_D1;
  wire [0:0] LIOI3_X0Y159_OLOGIC_X0Y159_OQ;
  wire [0:0] LIOI3_X0Y159_OLOGIC_X0Y159_T1;
  wire [0:0] LIOI3_X0Y159_OLOGIC_X0Y159_TQ;
  wire [0:0] LIOI3_X0Y159_OLOGIC_X0Y160_D1;
  wire [0:0] LIOI3_X0Y159_OLOGIC_X0Y160_OQ;
  wire [0:0] LIOI3_X0Y159_OLOGIC_X0Y160_T1;
  wire [0:0] LIOI3_X0Y159_OLOGIC_X0Y160_TQ;
  wire [0:0] LIOI3_X0Y161_OLOGIC_X0Y161_D1;
  wire [0:0] LIOI3_X0Y161_OLOGIC_X0Y161_OQ;
  wire [0:0] LIOI3_X0Y161_OLOGIC_X0Y161_T1;
  wire [0:0] LIOI3_X0Y161_OLOGIC_X0Y161_TQ;
  wire [0:0] LIOI3_X0Y161_OLOGIC_X0Y162_D1;
  wire [0:0] LIOI3_X0Y161_OLOGIC_X0Y162_OQ;
  wire [0:0] LIOI3_X0Y161_OLOGIC_X0Y162_T1;
  wire [0:0] LIOI3_X0Y161_OLOGIC_X0Y162_TQ;
  wire [0:0] LIOI3_X0Y165_OLOGIC_X0Y165_D1;
  wire [0:0] LIOI3_X0Y165_OLOGIC_X0Y165_OQ;
  wire [0:0] LIOI3_X0Y165_OLOGIC_X0Y165_T1;
  wire [0:0] LIOI3_X0Y165_OLOGIC_X0Y165_TQ;
  wire [0:0] LIOI3_X0Y165_OLOGIC_X0Y166_D1;
  wire [0:0] LIOI3_X0Y165_OLOGIC_X0Y166_OQ;
  wire [0:0] LIOI3_X0Y165_OLOGIC_X0Y166_T1;
  wire [0:0] LIOI3_X0Y165_OLOGIC_X0Y166_TQ;
  wire [0:0] LIOI3_X0Y167_OLOGIC_X0Y167_D1;
  wire [0:0] LIOI3_X0Y167_OLOGIC_X0Y167_OQ;
  wire [0:0] LIOI3_X0Y167_OLOGIC_X0Y167_T1;
  wire [0:0] LIOI3_X0Y167_OLOGIC_X0Y167_TQ;
  wire [0:0] LIOI3_X0Y167_OLOGIC_X0Y168_D1;
  wire [0:0] LIOI3_X0Y167_OLOGIC_X0Y168_OQ;
  wire [0:0] LIOI3_X0Y167_OLOGIC_X0Y168_T1;
  wire [0:0] LIOI3_X0Y167_OLOGIC_X0Y168_TQ;
  wire [0:0] LIOI3_X0Y171_OLOGIC_X0Y171_D1;
  wire [0:0] LIOI3_X0Y171_OLOGIC_X0Y171_OQ;
  wire [0:0] LIOI3_X0Y171_OLOGIC_X0Y171_T1;
  wire [0:0] LIOI3_X0Y171_OLOGIC_X0Y171_TQ;
  wire [0:0] LIOI3_X0Y171_OLOGIC_X0Y172_D1;
  wire [0:0] LIOI3_X0Y171_OLOGIC_X0Y172_OQ;
  wire [0:0] LIOI3_X0Y171_OLOGIC_X0Y172_T1;
  wire [0:0] LIOI3_X0Y171_OLOGIC_X0Y172_TQ;
  wire [0:0] LIOI3_X0Y173_OLOGIC_X0Y173_D1;
  wire [0:0] LIOI3_X0Y173_OLOGIC_X0Y173_OQ;
  wire [0:0] LIOI3_X0Y173_OLOGIC_X0Y173_T1;
  wire [0:0] LIOI3_X0Y173_OLOGIC_X0Y173_TQ;
  wire [0:0] LIOI3_X0Y173_OLOGIC_X0Y174_D1;
  wire [0:0] LIOI3_X0Y173_OLOGIC_X0Y174_OQ;
  wire [0:0] LIOI3_X0Y173_OLOGIC_X0Y174_T1;
  wire [0:0] LIOI3_X0Y173_OLOGIC_X0Y174_TQ;
  wire [0:0] LIOI3_X0Y175_OLOGIC_X0Y175_D1;
  wire [0:0] LIOI3_X0Y175_OLOGIC_X0Y175_OQ;
  wire [0:0] LIOI3_X0Y175_OLOGIC_X0Y175_T1;
  wire [0:0] LIOI3_X0Y175_OLOGIC_X0Y175_TQ;
  wire [0:0] LIOI3_X0Y175_OLOGIC_X0Y176_D1;
  wire [0:0] LIOI3_X0Y175_OLOGIC_X0Y176_OQ;
  wire [0:0] LIOI3_X0Y175_OLOGIC_X0Y176_T1;
  wire [0:0] LIOI3_X0Y175_OLOGIC_X0Y176_TQ;
  wire [0:0] LIOI3_X0Y177_OLOGIC_X0Y177_D1;
  wire [0:0] LIOI3_X0Y177_OLOGIC_X0Y177_OQ;
  wire [0:0] LIOI3_X0Y177_OLOGIC_X0Y177_T1;
  wire [0:0] LIOI3_X0Y177_OLOGIC_X0Y177_TQ;
  wire [0:0] LIOI3_X0Y177_OLOGIC_X0Y178_D1;
  wire [0:0] LIOI3_X0Y177_OLOGIC_X0Y178_OQ;
  wire [0:0] LIOI3_X0Y177_OLOGIC_X0Y178_T1;
  wire [0:0] LIOI3_X0Y177_OLOGIC_X0Y178_TQ;
  wire [0:0] LIOI3_X0Y179_OLOGIC_X0Y179_D1;
  wire [0:0] LIOI3_X0Y179_OLOGIC_X0Y179_OQ;
  wire [0:0] LIOI3_X0Y179_OLOGIC_X0Y179_T1;
  wire [0:0] LIOI3_X0Y179_OLOGIC_X0Y179_TQ;
  wire [0:0] LIOI3_X0Y179_OLOGIC_X0Y180_D1;
  wire [0:0] LIOI3_X0Y179_OLOGIC_X0Y180_OQ;
  wire [0:0] LIOI3_X0Y179_OLOGIC_X0Y180_T1;
  wire [0:0] LIOI3_X0Y179_OLOGIC_X0Y180_TQ;
  wire [0:0] LIOI3_X0Y183_OLOGIC_X0Y183_D1;
  wire [0:0] LIOI3_X0Y183_OLOGIC_X0Y183_OQ;
  wire [0:0] LIOI3_X0Y183_OLOGIC_X0Y183_T1;
  wire [0:0] LIOI3_X0Y183_OLOGIC_X0Y183_TQ;
  wire [0:0] LIOI3_X0Y183_OLOGIC_X0Y184_D1;
  wire [0:0] LIOI3_X0Y183_OLOGIC_X0Y184_OQ;
  wire [0:0] LIOI3_X0Y183_OLOGIC_X0Y184_T1;
  wire [0:0] LIOI3_X0Y183_OLOGIC_X0Y184_TQ;
  wire [0:0] LIOI3_X0Y185_OLOGIC_X0Y185_D1;
  wire [0:0] LIOI3_X0Y185_OLOGIC_X0Y185_OQ;
  wire [0:0] LIOI3_X0Y185_OLOGIC_X0Y185_T1;
  wire [0:0] LIOI3_X0Y185_OLOGIC_X0Y185_TQ;
  wire [0:0] LIOI3_X0Y185_OLOGIC_X0Y186_D1;
  wire [0:0] LIOI3_X0Y185_OLOGIC_X0Y186_OQ;
  wire [0:0] LIOI3_X0Y185_OLOGIC_X0Y186_T1;
  wire [0:0] LIOI3_X0Y185_OLOGIC_X0Y186_TQ;
  wire [0:0] LIOI3_X0Y189_OLOGIC_X0Y189_D1;
  wire [0:0] LIOI3_X0Y189_OLOGIC_X0Y189_OQ;
  wire [0:0] LIOI3_X0Y189_OLOGIC_X0Y189_T1;
  wire [0:0] LIOI3_X0Y189_OLOGIC_X0Y189_TQ;
  wire [0:0] LIOI3_X0Y189_OLOGIC_X0Y190_D1;
  wire [0:0] LIOI3_X0Y189_OLOGIC_X0Y190_OQ;
  wire [0:0] LIOI3_X0Y189_OLOGIC_X0Y190_T1;
  wire [0:0] LIOI3_X0Y189_OLOGIC_X0Y190_TQ;
  wire [0:0] LIOI3_X0Y191_OLOGIC_X0Y191_D1;
  wire [0:0] LIOI3_X0Y191_OLOGIC_X0Y191_OQ;
  wire [0:0] LIOI3_X0Y191_OLOGIC_X0Y191_T1;
  wire [0:0] LIOI3_X0Y191_OLOGIC_X0Y191_TQ;
  wire [0:0] LIOI3_X0Y191_OLOGIC_X0Y192_D1;
  wire [0:0] LIOI3_X0Y191_OLOGIC_X0Y192_OQ;
  wire [0:0] LIOI3_X0Y191_OLOGIC_X0Y192_T1;
  wire [0:0] LIOI3_X0Y191_OLOGIC_X0Y192_TQ;
  wire [0:0] LIOI3_X0Y195_OLOGIC_X0Y195_D1;
  wire [0:0] LIOI3_X0Y195_OLOGIC_X0Y195_OQ;
  wire [0:0] LIOI3_X0Y195_OLOGIC_X0Y195_T1;
  wire [0:0] LIOI3_X0Y195_OLOGIC_X0Y195_TQ;
  wire [0:0] LIOI3_X0Y195_OLOGIC_X0Y196_D1;
  wire [0:0] LIOI3_X0Y195_OLOGIC_X0Y196_OQ;
  wire [0:0] LIOI3_X0Y195_OLOGIC_X0Y196_T1;
  wire [0:0] LIOI3_X0Y195_OLOGIC_X0Y196_TQ;
  wire [0:0] LIOI3_X0Y197_OLOGIC_X0Y197_D1;
  wire [0:0] LIOI3_X0Y197_OLOGIC_X0Y197_OQ;
  wire [0:0] LIOI3_X0Y197_OLOGIC_X0Y197_T1;
  wire [0:0] LIOI3_X0Y197_OLOGIC_X0Y197_TQ;
  wire [0:0] LIOI3_X0Y197_OLOGIC_X0Y198_D1;
  wire [0:0] LIOI3_X0Y197_OLOGIC_X0Y198_OQ;
  wire [0:0] LIOI3_X0Y197_OLOGIC_X0Y198_T1;
  wire [0:0] LIOI3_X0Y197_OLOGIC_X0Y198_TQ;
  wire [0:0] LIOI3_X0Y51_ILOGIC_X0Y51_D;
  wire [0:0] LIOI3_X0Y51_ILOGIC_X0Y51_O;
  wire [0:0] LIOI3_X0Y51_ILOGIC_X0Y52_D;
  wire [0:0] LIOI3_X0Y51_ILOGIC_X0Y52_O;
  wire [0:0] LIOI3_X0Y53_ILOGIC_X0Y53_D;
  wire [0:0] LIOI3_X0Y53_ILOGIC_X0Y53_O;
  wire [0:0] LIOI3_X0Y53_ILOGIC_X0Y54_D;
  wire [0:0] LIOI3_X0Y53_ILOGIC_X0Y54_O;
  wire [0:0] LIOI3_X0Y55_ILOGIC_X0Y55_D;
  wire [0:0] LIOI3_X0Y55_ILOGIC_X0Y55_O;
  wire [0:0] LIOI3_X0Y55_ILOGIC_X0Y56_D;
  wire [0:0] LIOI3_X0Y55_ILOGIC_X0Y56_O;
  wire [0:0] LIOI3_X0Y59_ILOGIC_X0Y59_D;
  wire [0:0] LIOI3_X0Y59_ILOGIC_X0Y59_O;
  wire [0:0] LIOI3_X0Y59_ILOGIC_X0Y60_D;
  wire [0:0] LIOI3_X0Y59_ILOGIC_X0Y60_O;
  wire [0:0] LIOI3_X0Y61_ILOGIC_X0Y61_D;
  wire [0:0] LIOI3_X0Y61_ILOGIC_X0Y61_O;
  wire [0:0] LIOI3_X0Y61_ILOGIC_X0Y62_D;
  wire [0:0] LIOI3_X0Y61_ILOGIC_X0Y62_O;
  wire [0:0] LIOI3_X0Y65_ILOGIC_X0Y65_D;
  wire [0:0] LIOI3_X0Y65_ILOGIC_X0Y65_O;
  wire [0:0] LIOI3_X0Y65_ILOGIC_X0Y66_D;
  wire [0:0] LIOI3_X0Y65_ILOGIC_X0Y66_O;
  wire [0:0] LIOI3_X0Y67_ILOGIC_X0Y67_D;
  wire [0:0] LIOI3_X0Y67_ILOGIC_X0Y67_O;
  wire [0:0] LIOI3_X0Y67_ILOGIC_X0Y68_D;
  wire [0:0] LIOI3_X0Y67_ILOGIC_X0Y68_O;
  wire [0:0] LIOI3_X0Y71_ILOGIC_X0Y71_D;
  wire [0:0] LIOI3_X0Y71_ILOGIC_X0Y71_O;
  wire [0:0] LIOI3_X0Y71_ILOGIC_X0Y72_D;
  wire [0:0] LIOI3_X0Y71_ILOGIC_X0Y72_O;
  wire [0:0] LIOI3_X0Y73_ILOGIC_X0Y73_D;
  wire [0:0] LIOI3_X0Y73_ILOGIC_X0Y73_O;
  wire [0:0] LIOI3_X0Y73_ILOGIC_X0Y74_D;
  wire [0:0] LIOI3_X0Y73_ILOGIC_X0Y74_O;
  wire [0:0] LIOI3_X0Y75_ILOGIC_X0Y75_D;
  wire [0:0] LIOI3_X0Y75_ILOGIC_X0Y75_O;
  wire [0:0] LIOI3_X0Y75_ILOGIC_X0Y76_D;
  wire [0:0] LIOI3_X0Y75_ILOGIC_X0Y76_O;
  wire [0:0] LIOI3_X0Y77_ILOGIC_X0Y77_D;
  wire [0:0] LIOI3_X0Y77_ILOGIC_X0Y77_O;
  wire [0:0] LIOI3_X0Y77_ILOGIC_X0Y78_D;
  wire [0:0] LIOI3_X0Y77_ILOGIC_X0Y78_O;
  wire [0:0] LIOI3_X0Y79_ILOGIC_X0Y79_D;
  wire [0:0] LIOI3_X0Y79_ILOGIC_X0Y79_O;
  wire [0:0] LIOI3_X0Y79_OLOGIC_X0Y80_D1;
  wire [0:0] LIOI3_X0Y79_OLOGIC_X0Y80_OQ;
  wire [0:0] LIOI3_X0Y79_OLOGIC_X0Y80_T1;
  wire [0:0] LIOI3_X0Y79_OLOGIC_X0Y80_TQ;
  wire [0:0] RIOB33_SING_X105Y100_IOB_X1Y100_I;
  wire [0:0] RIOB33_SING_X105Y149_IOB_X1Y149_I;
  wire [0:0] RIOB33_SING_X105Y150_IOB_X1Y150_O;
  wire [0:0] RIOB33_SING_X105Y199_IOB_X1Y199_O;
  wire [0:0] RIOB33_X105Y101_IOB_X1Y101_I;
  wire [0:0] RIOB33_X105Y101_IOB_X1Y102_I;
  wire [0:0] RIOB33_X105Y103_IOB_X1Y103_I;
  wire [0:0] RIOB33_X105Y103_IOB_X1Y104_I;
  wire [0:0] RIOB33_X105Y105_IOB_X1Y105_I;
  wire [0:0] RIOB33_X105Y105_IOB_X1Y106_I;
  wire [0:0] RIOB33_X105Y107_IOB_X1Y107_I;
  wire [0:0] RIOB33_X105Y107_IOB_X1Y108_I;
  wire [0:0] RIOB33_X105Y109_IOB_X1Y109_I;
  wire [0:0] RIOB33_X105Y109_IOB_X1Y110_I;
  wire [0:0] RIOB33_X105Y111_IOB_X1Y111_I;
  wire [0:0] RIOB33_X105Y111_IOB_X1Y112_I;
  wire [0:0] RIOB33_X105Y113_IOB_X1Y113_I;
  wire [0:0] RIOB33_X105Y113_IOB_X1Y114_I;
  wire [0:0] RIOB33_X105Y115_IOB_X1Y115_I;
  wire [0:0] RIOB33_X105Y115_IOB_X1Y116_I;
  wire [0:0] RIOB33_X105Y117_IOB_X1Y117_I;
  wire [0:0] RIOB33_X105Y117_IOB_X1Y118_I;
  wire [0:0] RIOB33_X105Y119_IOB_X1Y119_I;
  wire [0:0] RIOB33_X105Y119_IOB_X1Y120_I;
  wire [0:0] RIOB33_X105Y121_IOB_X1Y121_I;
  wire [0:0] RIOB33_X105Y121_IOB_X1Y122_I;
  wire [0:0] RIOB33_X105Y123_IOB_X1Y123_I;
  wire [0:0] RIOB33_X105Y123_IOB_X1Y124_I;
  wire [0:0] RIOB33_X105Y125_IOB_X1Y125_I;
  wire [0:0] RIOB33_X105Y125_IOB_X1Y126_I;
  wire [0:0] RIOB33_X105Y127_IOB_X1Y127_I;
  wire [0:0] RIOB33_X105Y127_IOB_X1Y128_I;
  wire [0:0] RIOB33_X105Y129_IOB_X1Y129_I;
  wire [0:0] RIOB33_X105Y129_IOB_X1Y130_I;
  wire [0:0] RIOB33_X105Y131_IOB_X1Y131_I;
  wire [0:0] RIOB33_X105Y131_IOB_X1Y132_I;
  wire [0:0] RIOB33_X105Y133_IOB_X1Y133_I;
  wire [0:0] RIOB33_X105Y133_IOB_X1Y134_I;
  wire [0:0] RIOB33_X105Y135_IOB_X1Y135_I;
  wire [0:0] RIOB33_X105Y135_IOB_X1Y136_I;
  wire [0:0] RIOB33_X105Y137_IOB_X1Y137_I;
  wire [0:0] RIOB33_X105Y137_IOB_X1Y138_I;
  wire [0:0] RIOB33_X105Y139_IOB_X1Y139_I;
  wire [0:0] RIOB33_X105Y139_IOB_X1Y140_I;
  wire [0:0] RIOB33_X105Y141_IOB_X1Y141_I;
  wire [0:0] RIOB33_X105Y141_IOB_X1Y142_I;
  wire [0:0] RIOB33_X105Y143_IOB_X1Y143_I;
  wire [0:0] RIOB33_X105Y143_IOB_X1Y144_I;
  wire [0:0] RIOB33_X105Y145_IOB_X1Y145_I;
  wire [0:0] RIOB33_X105Y145_IOB_X1Y146_I;
  wire [0:0] RIOB33_X105Y147_IOB_X1Y147_I;
  wire [0:0] RIOB33_X105Y147_IOB_X1Y148_I;
  wire [0:0] RIOB33_X105Y151_IOB_X1Y151_O;
  wire [0:0] RIOB33_X105Y151_IOB_X1Y152_O;
  wire [0:0] RIOB33_X105Y153_IOB_X1Y153_O;
  wire [0:0] RIOB33_X105Y153_IOB_X1Y154_O;
  wire [0:0] RIOB33_X105Y155_IOB_X1Y155_O;
  wire [0:0] RIOB33_X105Y155_IOB_X1Y156_O;
  wire [0:0] RIOB33_X105Y157_IOB_X1Y157_O;
  wire [0:0] RIOB33_X105Y157_IOB_X1Y158_O;
  wire [0:0] RIOB33_X105Y159_IOB_X1Y159_O;
  wire [0:0] RIOB33_X105Y159_IOB_X1Y160_O;
  wire [0:0] RIOB33_X105Y161_IOB_X1Y161_O;
  wire [0:0] RIOB33_X105Y161_IOB_X1Y162_O;
  wire [0:0] RIOB33_X105Y163_IOB_X1Y163_O;
  wire [0:0] RIOB33_X105Y163_IOB_X1Y164_O;
  wire [0:0] RIOB33_X105Y165_IOB_X1Y165_O;
  wire [0:0] RIOB33_X105Y165_IOB_X1Y166_O;
  wire [0:0] RIOB33_X105Y167_IOB_X1Y167_O;
  wire [0:0] RIOB33_X105Y167_IOB_X1Y168_O;
  wire [0:0] RIOB33_X105Y169_IOB_X1Y169_O;
  wire [0:0] RIOB33_X105Y169_IOB_X1Y170_O;
  wire [0:0] RIOB33_X105Y171_IOB_X1Y171_O;
  wire [0:0] RIOB33_X105Y171_IOB_X1Y172_O;
  wire [0:0] RIOB33_X105Y173_IOB_X1Y173_O;
  wire [0:0] RIOB33_X105Y173_IOB_X1Y174_O;
  wire [0:0] RIOB33_X105Y175_IOB_X1Y175_O;
  wire [0:0] RIOB33_X105Y175_IOB_X1Y176_O;
  wire [0:0] RIOB33_X105Y177_IOB_X1Y177_O;
  wire [0:0] RIOB33_X105Y177_IOB_X1Y178_O;
  wire [0:0] RIOB33_X105Y179_IOB_X1Y179_O;
  wire [0:0] RIOB33_X105Y179_IOB_X1Y180_O;
  wire [0:0] RIOB33_X105Y181_IOB_X1Y181_O;
  wire [0:0] RIOB33_X105Y181_IOB_X1Y182_O;
  wire [0:0] RIOB33_X105Y183_IOB_X1Y183_O;
  wire [0:0] RIOB33_X105Y183_IOB_X1Y184_O;
  wire [0:0] RIOB33_X105Y185_IOB_X1Y185_O;
  wire [0:0] RIOB33_X105Y185_IOB_X1Y186_O;
  wire [0:0] RIOB33_X105Y187_IOB_X1Y187_O;
  wire [0:0] RIOB33_X105Y187_IOB_X1Y188_O;
  wire [0:0] RIOB33_X105Y189_IOB_X1Y189_O;
  wire [0:0] RIOB33_X105Y189_IOB_X1Y190_O;
  wire [0:0] RIOB33_X105Y191_IOB_X1Y191_O;
  wire [0:0] RIOB33_X105Y191_IOB_X1Y192_O;
  wire [0:0] RIOB33_X105Y193_IOB_X1Y193_O;
  wire [0:0] RIOB33_X105Y193_IOB_X1Y194_O;
  wire [0:0] RIOB33_X105Y195_IOB_X1Y195_O;
  wire [0:0] RIOB33_X105Y195_IOB_X1Y196_O;
  wire [0:0] RIOB33_X105Y197_IOB_X1Y197_O;
  wire [0:0] RIOB33_X105Y197_IOB_X1Y198_O;
  wire [0:0] RIOI3_SING_X105Y100_ILOGIC_X1Y100_D;
  wire [0:0] RIOI3_SING_X105Y100_ILOGIC_X1Y100_O;
  wire [0:0] RIOI3_SING_X105Y149_ILOGIC_X1Y149_D;
  wire [0:0] RIOI3_SING_X105Y149_ILOGIC_X1Y149_O;
  wire [0:0] RIOI3_SING_X105Y150_OLOGIC_X1Y150_D1;
  wire [0:0] RIOI3_SING_X105Y150_OLOGIC_X1Y150_OQ;
  wire [0:0] RIOI3_SING_X105Y150_OLOGIC_X1Y150_T1;
  wire [0:0] RIOI3_SING_X105Y150_OLOGIC_X1Y150_TQ;
  wire [0:0] RIOI3_SING_X105Y199_OLOGIC_X1Y199_D1;
  wire [0:0] RIOI3_SING_X105Y199_OLOGIC_X1Y199_OQ;
  wire [0:0] RIOI3_SING_X105Y199_OLOGIC_X1Y199_T1;
  wire [0:0] RIOI3_SING_X105Y199_OLOGIC_X1Y199_TQ;
  wire [0:0] RIOI3_TBYTESRC_X105Y107_ILOGIC_X1Y107_D;
  wire [0:0] RIOI3_TBYTESRC_X105Y107_ILOGIC_X1Y107_O;
  wire [0:0] RIOI3_TBYTESRC_X105Y107_ILOGIC_X1Y108_D;
  wire [0:0] RIOI3_TBYTESRC_X105Y107_ILOGIC_X1Y108_O;
  wire [0:0] RIOI3_TBYTESRC_X105Y119_ILOGIC_X1Y119_D;
  wire [0:0] RIOI3_TBYTESRC_X105Y119_ILOGIC_X1Y119_O;
  wire [0:0] RIOI3_TBYTESRC_X105Y131_ILOGIC_X1Y131_D;
  wire [0:0] RIOI3_TBYTESRC_X105Y131_ILOGIC_X1Y131_O;
  wire [0:0] RIOI3_TBYTESRC_X105Y131_ILOGIC_X1Y132_D;
  wire [0:0] RIOI3_TBYTESRC_X105Y131_ILOGIC_X1Y132_O;
  wire [0:0] RIOI3_TBYTESRC_X105Y143_ILOGIC_X1Y143_D;
  wire [0:0] RIOI3_TBYTESRC_X105Y143_ILOGIC_X1Y143_O;
  wire [0:0] RIOI3_TBYTESRC_X105Y143_ILOGIC_X1Y144_D;
  wire [0:0] RIOI3_TBYTESRC_X105Y143_ILOGIC_X1Y144_O;
  wire [0:0] RIOI3_TBYTESRC_X105Y157_OLOGIC_X1Y157_D1;
  wire [0:0] RIOI3_TBYTESRC_X105Y157_OLOGIC_X1Y157_OQ;
  wire [0:0] RIOI3_TBYTESRC_X105Y157_OLOGIC_X1Y157_T1;
  wire [0:0] RIOI3_TBYTESRC_X105Y157_OLOGIC_X1Y157_TQ;
  wire [0:0] RIOI3_TBYTESRC_X105Y157_OLOGIC_X1Y158_D1;
  wire [0:0] RIOI3_TBYTESRC_X105Y157_OLOGIC_X1Y158_OQ;
  wire [0:0] RIOI3_TBYTESRC_X105Y157_OLOGIC_X1Y158_T1;
  wire [0:0] RIOI3_TBYTESRC_X105Y157_OLOGIC_X1Y158_TQ;
  wire [0:0] RIOI3_TBYTESRC_X105Y169_OLOGIC_X1Y169_D1;
  wire [0:0] RIOI3_TBYTESRC_X105Y169_OLOGIC_X1Y169_OQ;
  wire [0:0] RIOI3_TBYTESRC_X105Y169_OLOGIC_X1Y169_T1;
  wire [0:0] RIOI3_TBYTESRC_X105Y169_OLOGIC_X1Y169_TQ;
  wire [0:0] RIOI3_TBYTESRC_X105Y169_OLOGIC_X1Y170_D1;
  wire [0:0] RIOI3_TBYTESRC_X105Y169_OLOGIC_X1Y170_OQ;
  wire [0:0] RIOI3_TBYTESRC_X105Y169_OLOGIC_X1Y170_T1;
  wire [0:0] RIOI3_TBYTESRC_X105Y169_OLOGIC_X1Y170_TQ;
  wire [0:0] RIOI3_TBYTESRC_X105Y181_OLOGIC_X1Y181_D1;
  wire [0:0] RIOI3_TBYTESRC_X105Y181_OLOGIC_X1Y181_OQ;
  wire [0:0] RIOI3_TBYTESRC_X105Y181_OLOGIC_X1Y181_T1;
  wire [0:0] RIOI3_TBYTESRC_X105Y181_OLOGIC_X1Y181_TQ;
  wire [0:0] RIOI3_TBYTESRC_X105Y181_OLOGIC_X1Y182_D1;
  wire [0:0] RIOI3_TBYTESRC_X105Y181_OLOGIC_X1Y182_OQ;
  wire [0:0] RIOI3_TBYTESRC_X105Y181_OLOGIC_X1Y182_T1;
  wire [0:0] RIOI3_TBYTESRC_X105Y181_OLOGIC_X1Y182_TQ;
  wire [0:0] RIOI3_TBYTESRC_X105Y193_OLOGIC_X1Y193_D1;
  wire [0:0] RIOI3_TBYTESRC_X105Y193_OLOGIC_X1Y193_OQ;
  wire [0:0] RIOI3_TBYTESRC_X105Y193_OLOGIC_X1Y193_T1;
  wire [0:0] RIOI3_TBYTESRC_X105Y193_OLOGIC_X1Y193_TQ;
  wire [0:0] RIOI3_TBYTESRC_X105Y193_OLOGIC_X1Y194_D1;
  wire [0:0] RIOI3_TBYTESRC_X105Y193_OLOGIC_X1Y194_OQ;
  wire [0:0] RIOI3_TBYTESRC_X105Y193_OLOGIC_X1Y194_T1;
  wire [0:0] RIOI3_TBYTESRC_X105Y193_OLOGIC_X1Y194_TQ;
  wire [0:0] RIOI3_TBYTETERM_X105Y113_ILOGIC_X1Y113_D;
  wire [0:0] RIOI3_TBYTETERM_X105Y113_ILOGIC_X1Y113_O;
  wire [0:0] RIOI3_TBYTETERM_X105Y113_ILOGIC_X1Y114_D;
  wire [0:0] RIOI3_TBYTETERM_X105Y113_ILOGIC_X1Y114_O;
  wire [0:0] RIOI3_TBYTETERM_X105Y137_ILOGIC_X1Y137_D;
  wire [0:0] RIOI3_TBYTETERM_X105Y137_ILOGIC_X1Y137_O;
  wire [0:0] RIOI3_TBYTETERM_X105Y137_ILOGIC_X1Y138_D;
  wire [0:0] RIOI3_TBYTETERM_X105Y137_ILOGIC_X1Y138_O;
  wire [0:0] RIOI3_TBYTETERM_X105Y163_OLOGIC_X1Y163_D1;
  wire [0:0] RIOI3_TBYTETERM_X105Y163_OLOGIC_X1Y163_OQ;
  wire [0:0] RIOI3_TBYTETERM_X105Y163_OLOGIC_X1Y163_T1;
  wire [0:0] RIOI3_TBYTETERM_X105Y163_OLOGIC_X1Y163_TQ;
  wire [0:0] RIOI3_TBYTETERM_X105Y163_OLOGIC_X1Y164_D1;
  wire [0:0] RIOI3_TBYTETERM_X105Y163_OLOGIC_X1Y164_OQ;
  wire [0:0] RIOI3_TBYTETERM_X105Y163_OLOGIC_X1Y164_T1;
  wire [0:0] RIOI3_TBYTETERM_X105Y163_OLOGIC_X1Y164_TQ;
  wire [0:0] RIOI3_TBYTETERM_X105Y187_OLOGIC_X1Y187_D1;
  wire [0:0] RIOI3_TBYTETERM_X105Y187_OLOGIC_X1Y187_OQ;
  wire [0:0] RIOI3_TBYTETERM_X105Y187_OLOGIC_X1Y187_T1;
  wire [0:0] RIOI3_TBYTETERM_X105Y187_OLOGIC_X1Y187_TQ;
  wire [0:0] RIOI3_TBYTETERM_X105Y187_OLOGIC_X1Y188_D1;
  wire [0:0] RIOI3_TBYTETERM_X105Y187_OLOGIC_X1Y188_OQ;
  wire [0:0] RIOI3_TBYTETERM_X105Y187_OLOGIC_X1Y188_T1;
  wire [0:0] RIOI3_TBYTETERM_X105Y187_OLOGIC_X1Y188_TQ;
  wire [0:0] RIOI3_X105Y101_ILOGIC_X1Y101_D;
  wire [0:0] RIOI3_X105Y101_ILOGIC_X1Y101_O;
  wire [0:0] RIOI3_X105Y101_ILOGIC_X1Y102_D;
  wire [0:0] RIOI3_X105Y101_ILOGIC_X1Y102_O;
  wire [0:0] RIOI3_X105Y103_ILOGIC_X1Y103_D;
  wire [0:0] RIOI3_X105Y103_ILOGIC_X1Y103_O;
  wire [0:0] RIOI3_X105Y103_ILOGIC_X1Y104_D;
  wire [0:0] RIOI3_X105Y103_ILOGIC_X1Y104_O;
  wire [0:0] RIOI3_X105Y105_ILOGIC_X1Y105_D;
  wire [0:0] RIOI3_X105Y105_ILOGIC_X1Y105_O;
  wire [0:0] RIOI3_X105Y105_ILOGIC_X1Y106_D;
  wire [0:0] RIOI3_X105Y105_ILOGIC_X1Y106_O;
  wire [0:0] RIOI3_X105Y109_ILOGIC_X1Y109_D;
  wire [0:0] RIOI3_X105Y109_ILOGIC_X1Y109_O;
  wire [0:0] RIOI3_X105Y109_ILOGIC_X1Y110_D;
  wire [0:0] RIOI3_X105Y109_ILOGIC_X1Y110_O;
  wire [0:0] RIOI3_X105Y111_ILOGIC_X1Y111_D;
  wire [0:0] RIOI3_X105Y111_ILOGIC_X1Y111_O;
  wire [0:0] RIOI3_X105Y111_ILOGIC_X1Y112_D;
  wire [0:0] RIOI3_X105Y111_ILOGIC_X1Y112_O;
  wire [0:0] RIOI3_X105Y115_ILOGIC_X1Y115_D;
  wire [0:0] RIOI3_X105Y115_ILOGIC_X1Y115_O;
  wire [0:0] RIOI3_X105Y115_ILOGIC_X1Y116_D;
  wire [0:0] RIOI3_X105Y115_ILOGIC_X1Y116_O;
  wire [0:0] RIOI3_X105Y117_ILOGIC_X1Y117_D;
  wire [0:0] RIOI3_X105Y117_ILOGIC_X1Y117_O;
  wire [0:0] RIOI3_X105Y117_ILOGIC_X1Y118_D;
  wire [0:0] RIOI3_X105Y117_ILOGIC_X1Y118_O;
  wire [0:0] RIOI3_X105Y121_ILOGIC_X1Y121_D;
  wire [0:0] RIOI3_X105Y121_ILOGIC_X1Y121_O;
  wire [0:0] RIOI3_X105Y121_ILOGIC_X1Y122_D;
  wire [0:0] RIOI3_X105Y121_ILOGIC_X1Y122_O;
  wire [0:0] RIOI3_X105Y123_ILOGIC_X1Y123_D;
  wire [0:0] RIOI3_X105Y123_ILOGIC_X1Y123_O;
  wire [0:0] RIOI3_X105Y123_ILOGIC_X1Y124_D;
  wire [0:0] RIOI3_X105Y123_ILOGIC_X1Y124_O;
  wire [0:0] RIOI3_X105Y125_ILOGIC_X1Y125_D;
  wire [0:0] RIOI3_X105Y125_ILOGIC_X1Y125_O;
  wire [0:0] RIOI3_X105Y125_ILOGIC_X1Y126_D;
  wire [0:0] RIOI3_X105Y125_ILOGIC_X1Y126_O;
  wire [0:0] RIOI3_X105Y127_ILOGIC_X1Y127_D;
  wire [0:0] RIOI3_X105Y127_ILOGIC_X1Y127_O;
  wire [0:0] RIOI3_X105Y127_ILOGIC_X1Y128_D;
  wire [0:0] RIOI3_X105Y127_ILOGIC_X1Y128_O;
  wire [0:0] RIOI3_X105Y129_ILOGIC_X1Y129_D;
  wire [0:0] RIOI3_X105Y129_ILOGIC_X1Y129_O;
  wire [0:0] RIOI3_X105Y129_ILOGIC_X1Y130_D;
  wire [0:0] RIOI3_X105Y129_ILOGIC_X1Y130_O;
  wire [0:0] RIOI3_X105Y133_ILOGIC_X1Y133_D;
  wire [0:0] RIOI3_X105Y133_ILOGIC_X1Y133_O;
  wire [0:0] RIOI3_X105Y133_ILOGIC_X1Y134_D;
  wire [0:0] RIOI3_X105Y133_ILOGIC_X1Y134_O;
  wire [0:0] RIOI3_X105Y135_ILOGIC_X1Y135_D;
  wire [0:0] RIOI3_X105Y135_ILOGIC_X1Y135_O;
  wire [0:0] RIOI3_X105Y135_ILOGIC_X1Y136_D;
  wire [0:0] RIOI3_X105Y135_ILOGIC_X1Y136_O;
  wire [0:0] RIOI3_X105Y139_ILOGIC_X1Y139_D;
  wire [0:0] RIOI3_X105Y139_ILOGIC_X1Y139_O;
  wire [0:0] RIOI3_X105Y139_ILOGIC_X1Y140_D;
  wire [0:0] RIOI3_X105Y139_ILOGIC_X1Y140_O;
  wire [0:0] RIOI3_X105Y141_ILOGIC_X1Y141_D;
  wire [0:0] RIOI3_X105Y141_ILOGIC_X1Y141_O;
  wire [0:0] RIOI3_X105Y141_ILOGIC_X1Y142_D;
  wire [0:0] RIOI3_X105Y141_ILOGIC_X1Y142_O;
  wire [0:0] RIOI3_X105Y145_ILOGIC_X1Y145_D;
  wire [0:0] RIOI3_X105Y145_ILOGIC_X1Y145_O;
  wire [0:0] RIOI3_X105Y145_ILOGIC_X1Y146_D;
  wire [0:0] RIOI3_X105Y145_ILOGIC_X1Y146_O;
  wire [0:0] RIOI3_X105Y147_ILOGIC_X1Y147_D;
  wire [0:0] RIOI3_X105Y147_ILOGIC_X1Y147_O;
  wire [0:0] RIOI3_X105Y147_ILOGIC_X1Y148_D;
  wire [0:0] RIOI3_X105Y147_ILOGIC_X1Y148_O;
  wire [0:0] RIOI3_X105Y151_OLOGIC_X1Y151_D1;
  wire [0:0] RIOI3_X105Y151_OLOGIC_X1Y151_OQ;
  wire [0:0] RIOI3_X105Y151_OLOGIC_X1Y151_T1;
  wire [0:0] RIOI3_X105Y151_OLOGIC_X1Y151_TQ;
  wire [0:0] RIOI3_X105Y151_OLOGIC_X1Y152_D1;
  wire [0:0] RIOI3_X105Y151_OLOGIC_X1Y152_OQ;
  wire [0:0] RIOI3_X105Y151_OLOGIC_X1Y152_T1;
  wire [0:0] RIOI3_X105Y151_OLOGIC_X1Y152_TQ;
  wire [0:0] RIOI3_X105Y153_OLOGIC_X1Y153_D1;
  wire [0:0] RIOI3_X105Y153_OLOGIC_X1Y153_OQ;
  wire [0:0] RIOI3_X105Y153_OLOGIC_X1Y153_T1;
  wire [0:0] RIOI3_X105Y153_OLOGIC_X1Y153_TQ;
  wire [0:0] RIOI3_X105Y153_OLOGIC_X1Y154_D1;
  wire [0:0] RIOI3_X105Y153_OLOGIC_X1Y154_OQ;
  wire [0:0] RIOI3_X105Y153_OLOGIC_X1Y154_T1;
  wire [0:0] RIOI3_X105Y153_OLOGIC_X1Y154_TQ;
  wire [0:0] RIOI3_X105Y155_OLOGIC_X1Y155_D1;
  wire [0:0] RIOI3_X105Y155_OLOGIC_X1Y155_OQ;
  wire [0:0] RIOI3_X105Y155_OLOGIC_X1Y155_T1;
  wire [0:0] RIOI3_X105Y155_OLOGIC_X1Y155_TQ;
  wire [0:0] RIOI3_X105Y155_OLOGIC_X1Y156_D1;
  wire [0:0] RIOI3_X105Y155_OLOGIC_X1Y156_OQ;
  wire [0:0] RIOI3_X105Y155_OLOGIC_X1Y156_T1;
  wire [0:0] RIOI3_X105Y155_OLOGIC_X1Y156_TQ;
  wire [0:0] RIOI3_X105Y159_OLOGIC_X1Y159_D1;
  wire [0:0] RIOI3_X105Y159_OLOGIC_X1Y159_OQ;
  wire [0:0] RIOI3_X105Y159_OLOGIC_X1Y159_T1;
  wire [0:0] RIOI3_X105Y159_OLOGIC_X1Y159_TQ;
  wire [0:0] RIOI3_X105Y159_OLOGIC_X1Y160_D1;
  wire [0:0] RIOI3_X105Y159_OLOGIC_X1Y160_OQ;
  wire [0:0] RIOI3_X105Y159_OLOGIC_X1Y160_T1;
  wire [0:0] RIOI3_X105Y159_OLOGIC_X1Y160_TQ;
  wire [0:0] RIOI3_X105Y161_OLOGIC_X1Y161_D1;
  wire [0:0] RIOI3_X105Y161_OLOGIC_X1Y161_OQ;
  wire [0:0] RIOI3_X105Y161_OLOGIC_X1Y161_T1;
  wire [0:0] RIOI3_X105Y161_OLOGIC_X1Y161_TQ;
  wire [0:0] RIOI3_X105Y161_OLOGIC_X1Y162_D1;
  wire [0:0] RIOI3_X105Y161_OLOGIC_X1Y162_OQ;
  wire [0:0] RIOI3_X105Y161_OLOGIC_X1Y162_T1;
  wire [0:0] RIOI3_X105Y161_OLOGIC_X1Y162_TQ;
  wire [0:0] RIOI3_X105Y165_OLOGIC_X1Y165_D1;
  wire [0:0] RIOI3_X105Y165_OLOGIC_X1Y165_OQ;
  wire [0:0] RIOI3_X105Y165_OLOGIC_X1Y165_T1;
  wire [0:0] RIOI3_X105Y165_OLOGIC_X1Y165_TQ;
  wire [0:0] RIOI3_X105Y165_OLOGIC_X1Y166_D1;
  wire [0:0] RIOI3_X105Y165_OLOGIC_X1Y166_OQ;
  wire [0:0] RIOI3_X105Y165_OLOGIC_X1Y166_T1;
  wire [0:0] RIOI3_X105Y165_OLOGIC_X1Y166_TQ;
  wire [0:0] RIOI3_X105Y167_OLOGIC_X1Y167_D1;
  wire [0:0] RIOI3_X105Y167_OLOGIC_X1Y167_OQ;
  wire [0:0] RIOI3_X105Y167_OLOGIC_X1Y167_T1;
  wire [0:0] RIOI3_X105Y167_OLOGIC_X1Y167_TQ;
  wire [0:0] RIOI3_X105Y167_OLOGIC_X1Y168_D1;
  wire [0:0] RIOI3_X105Y167_OLOGIC_X1Y168_OQ;
  wire [0:0] RIOI3_X105Y167_OLOGIC_X1Y168_T1;
  wire [0:0] RIOI3_X105Y167_OLOGIC_X1Y168_TQ;
  wire [0:0] RIOI3_X105Y171_OLOGIC_X1Y171_D1;
  wire [0:0] RIOI3_X105Y171_OLOGIC_X1Y171_OQ;
  wire [0:0] RIOI3_X105Y171_OLOGIC_X1Y171_T1;
  wire [0:0] RIOI3_X105Y171_OLOGIC_X1Y171_TQ;
  wire [0:0] RIOI3_X105Y171_OLOGIC_X1Y172_D1;
  wire [0:0] RIOI3_X105Y171_OLOGIC_X1Y172_OQ;
  wire [0:0] RIOI3_X105Y171_OLOGIC_X1Y172_T1;
  wire [0:0] RIOI3_X105Y171_OLOGIC_X1Y172_TQ;
  wire [0:0] RIOI3_X105Y173_OLOGIC_X1Y173_D1;
  wire [0:0] RIOI3_X105Y173_OLOGIC_X1Y173_OQ;
  wire [0:0] RIOI3_X105Y173_OLOGIC_X1Y173_T1;
  wire [0:0] RIOI3_X105Y173_OLOGIC_X1Y173_TQ;
  wire [0:0] RIOI3_X105Y173_OLOGIC_X1Y174_D1;
  wire [0:0] RIOI3_X105Y173_OLOGIC_X1Y174_OQ;
  wire [0:0] RIOI3_X105Y173_OLOGIC_X1Y174_T1;
  wire [0:0] RIOI3_X105Y173_OLOGIC_X1Y174_TQ;
  wire [0:0] RIOI3_X105Y175_OLOGIC_X1Y175_D1;
  wire [0:0] RIOI3_X105Y175_OLOGIC_X1Y175_OQ;
  wire [0:0] RIOI3_X105Y175_OLOGIC_X1Y175_T1;
  wire [0:0] RIOI3_X105Y175_OLOGIC_X1Y175_TQ;
  wire [0:0] RIOI3_X105Y175_OLOGIC_X1Y176_D1;
  wire [0:0] RIOI3_X105Y175_OLOGIC_X1Y176_OQ;
  wire [0:0] RIOI3_X105Y175_OLOGIC_X1Y176_T1;
  wire [0:0] RIOI3_X105Y175_OLOGIC_X1Y176_TQ;
  wire [0:0] RIOI3_X105Y177_OLOGIC_X1Y177_D1;
  wire [0:0] RIOI3_X105Y177_OLOGIC_X1Y177_OQ;
  wire [0:0] RIOI3_X105Y177_OLOGIC_X1Y177_T1;
  wire [0:0] RIOI3_X105Y177_OLOGIC_X1Y177_TQ;
  wire [0:0] RIOI3_X105Y177_OLOGIC_X1Y178_D1;
  wire [0:0] RIOI3_X105Y177_OLOGIC_X1Y178_OQ;
  wire [0:0] RIOI3_X105Y177_OLOGIC_X1Y178_T1;
  wire [0:0] RIOI3_X105Y177_OLOGIC_X1Y178_TQ;
  wire [0:0] RIOI3_X105Y179_OLOGIC_X1Y179_D1;
  wire [0:0] RIOI3_X105Y179_OLOGIC_X1Y179_OQ;
  wire [0:0] RIOI3_X105Y179_OLOGIC_X1Y179_T1;
  wire [0:0] RIOI3_X105Y179_OLOGIC_X1Y179_TQ;
  wire [0:0] RIOI3_X105Y179_OLOGIC_X1Y180_D1;
  wire [0:0] RIOI3_X105Y179_OLOGIC_X1Y180_OQ;
  wire [0:0] RIOI3_X105Y179_OLOGIC_X1Y180_T1;
  wire [0:0] RIOI3_X105Y179_OLOGIC_X1Y180_TQ;
  wire [0:0] RIOI3_X105Y183_OLOGIC_X1Y183_D1;
  wire [0:0] RIOI3_X105Y183_OLOGIC_X1Y183_OQ;
  wire [0:0] RIOI3_X105Y183_OLOGIC_X1Y183_T1;
  wire [0:0] RIOI3_X105Y183_OLOGIC_X1Y183_TQ;
  wire [0:0] RIOI3_X105Y183_OLOGIC_X1Y184_D1;
  wire [0:0] RIOI3_X105Y183_OLOGIC_X1Y184_OQ;
  wire [0:0] RIOI3_X105Y183_OLOGIC_X1Y184_T1;
  wire [0:0] RIOI3_X105Y183_OLOGIC_X1Y184_TQ;
  wire [0:0] RIOI3_X105Y185_OLOGIC_X1Y185_D1;
  wire [0:0] RIOI3_X105Y185_OLOGIC_X1Y185_OQ;
  wire [0:0] RIOI3_X105Y185_OLOGIC_X1Y185_T1;
  wire [0:0] RIOI3_X105Y185_OLOGIC_X1Y185_TQ;
  wire [0:0] RIOI3_X105Y185_OLOGIC_X1Y186_D1;
  wire [0:0] RIOI3_X105Y185_OLOGIC_X1Y186_OQ;
  wire [0:0] RIOI3_X105Y185_OLOGIC_X1Y186_T1;
  wire [0:0] RIOI3_X105Y185_OLOGIC_X1Y186_TQ;
  wire [0:0] RIOI3_X105Y189_OLOGIC_X1Y189_D1;
  wire [0:0] RIOI3_X105Y189_OLOGIC_X1Y189_OQ;
  wire [0:0] RIOI3_X105Y189_OLOGIC_X1Y189_T1;
  wire [0:0] RIOI3_X105Y189_OLOGIC_X1Y189_TQ;
  wire [0:0] RIOI3_X105Y189_OLOGIC_X1Y190_D1;
  wire [0:0] RIOI3_X105Y189_OLOGIC_X1Y190_OQ;
  wire [0:0] RIOI3_X105Y189_OLOGIC_X1Y190_T1;
  wire [0:0] RIOI3_X105Y189_OLOGIC_X1Y190_TQ;
  wire [0:0] RIOI3_X105Y191_OLOGIC_X1Y191_D1;
  wire [0:0] RIOI3_X105Y191_OLOGIC_X1Y191_OQ;
  wire [0:0] RIOI3_X105Y191_OLOGIC_X1Y191_T1;
  wire [0:0] RIOI3_X105Y191_OLOGIC_X1Y191_TQ;
  wire [0:0] RIOI3_X105Y191_OLOGIC_X1Y192_D1;
  wire [0:0] RIOI3_X105Y191_OLOGIC_X1Y192_OQ;
  wire [0:0] RIOI3_X105Y191_OLOGIC_X1Y192_T1;
  wire [0:0] RIOI3_X105Y191_OLOGIC_X1Y192_TQ;
  wire [0:0] RIOI3_X105Y195_OLOGIC_X1Y195_D1;
  wire [0:0] RIOI3_X105Y195_OLOGIC_X1Y195_OQ;
  wire [0:0] RIOI3_X105Y195_OLOGIC_X1Y195_T1;
  wire [0:0] RIOI3_X105Y195_OLOGIC_X1Y195_TQ;
  wire [0:0] RIOI3_X105Y195_OLOGIC_X1Y196_D1;
  wire [0:0] RIOI3_X105Y195_OLOGIC_X1Y196_OQ;
  wire [0:0] RIOI3_X105Y195_OLOGIC_X1Y196_T1;
  wire [0:0] RIOI3_X105Y195_OLOGIC_X1Y196_TQ;
  wire [0:0] RIOI3_X105Y197_OLOGIC_X1Y197_D1;
  wire [0:0] RIOI3_X105Y197_OLOGIC_X1Y197_OQ;
  wire [0:0] RIOI3_X105Y197_OLOGIC_X1Y197_T1;
  wire [0:0] RIOI3_X105Y197_OLOGIC_X1Y197_TQ;
  wire [0:0] RIOI3_X105Y197_OLOGIC_X1Y198_D1;
  wire [0:0] RIOI3_X105Y197_OLOGIC_X1Y198_OQ;
  wire [0:0] RIOI3_X105Y197_OLOGIC_X1Y198_T1;
  wire [0:0] RIOI3_X105Y197_OLOGIC_X1Y198_TQ;


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y109_SLICE_X0Y109_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y109_SLICE_X0Y109_DO5),
.O6(CLBLL_L_X2Y109_SLICE_X0Y109_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y109_SLICE_X0Y109_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y109_SLICE_X0Y109_CO5),
.O6(CLBLL_L_X2Y109_SLICE_X0Y109_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y109_SLICE_X0Y109_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y109_SLICE_X0Y109_BO5),
.O6(CLBLL_L_X2Y109_SLICE_X0Y109_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h00ff00ff00ff00ff)
  ) CLBLL_L_X2Y109_SLICE_X0Y109_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(CLBLL_L_X2Y110_SLICE_X0Y110_BO6),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y109_SLICE_X0Y109_AO5),
.O6(CLBLL_L_X2Y109_SLICE_X0Y109_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y109_SLICE_X1Y109_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y109_SLICE_X1Y109_DO5),
.O6(CLBLL_L_X2Y109_SLICE_X1Y109_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y109_SLICE_X1Y109_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y109_SLICE_X1Y109_CO5),
.O6(CLBLL_L_X2Y109_SLICE_X1Y109_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y109_SLICE_X1Y109_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y109_SLICE_X1Y109_BO5),
.O6(CLBLL_L_X2Y109_SLICE_X1Y109_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y109_SLICE_X1Y109_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y109_SLICE_X1Y109_AO5),
.O6(CLBLL_L_X2Y109_SLICE_X1Y109_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y110_SLICE_X0Y110_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y110_SLICE_X0Y110_DO5),
.O6(CLBLL_L_X2Y110_SLICE_X0Y110_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y110_SLICE_X0Y110_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y110_SLICE_X0Y110_CO5),
.O6(CLBLL_L_X2Y110_SLICE_X0Y110_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hffec0000ecec0000)
  ) CLBLL_L_X2Y110_SLICE_X0Y110_BLUT (
.I0(LIOB33_X0Y51_IOB_X0Y51_I),
.I1(CLBLM_R_X3Y111_SLICE_X2Y111_CO6),
.I2(CLBLL_L_X2Y120_SLICE_X0Y120_CO6),
.I3(LIOB33_X0Y53_IOB_X0Y53_I),
.I4(RIOB33_X105Y105_IOB_X1Y105_I),
.I5(CLBLL_L_X4Y120_SLICE_X4Y120_AO6),
.O5(CLBLL_L_X2Y110_SLICE_X0Y110_BO5),
.O6(CLBLL_L_X2Y110_SLICE_X0Y110_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0f0ff0f000f000f0)
  ) CLBLL_L_X2Y110_SLICE_X0Y110_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(CLBLM_R_X3Y111_SLICE_X3Y111_CO6),
.I3(CLBLL_L_X2Y110_SLICE_X0Y110_BO6),
.I4(CLBLL_L_X4Y121_SLICE_X5Y121_BO5),
.I5(1'b1),
.O5(CLBLL_L_X2Y110_SLICE_X0Y110_AO5),
.O6(CLBLL_L_X2Y110_SLICE_X0Y110_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y110_SLICE_X1Y110_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y110_SLICE_X1Y110_DO5),
.O6(CLBLL_L_X2Y110_SLICE_X1Y110_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y110_SLICE_X1Y110_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y110_SLICE_X1Y110_CO5),
.O6(CLBLL_L_X2Y110_SLICE_X1Y110_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y110_SLICE_X1Y110_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y110_SLICE_X1Y110_BO5),
.O6(CLBLL_L_X2Y110_SLICE_X1Y110_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y110_SLICE_X1Y110_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y110_SLICE_X1Y110_AO5),
.O6(CLBLL_L_X2Y110_SLICE_X1Y110_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffff5fffffdfd)
  ) CLBLL_L_X2Y111_SLICE_X0Y111_DLUT (
.I0(RIOB33_X105Y137_IOB_X1Y137_I),
.I1(CLBLL_L_X2Y120_SLICE_X1Y120_DO6),
.I2(RIOB33_X105Y127_IOB_X1Y128_I),
.I3(CLBLL_L_X4Y120_SLICE_X5Y120_DO6),
.I4(RIOB33_X105Y129_IOB_X1Y129_I),
.I5(1'b1),
.O5(CLBLL_L_X2Y111_SLICE_X0Y111_DO5),
.O6(CLBLL_L_X2Y111_SLICE_X0Y111_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffafffffffcff)
  ) CLBLL_L_X2Y111_SLICE_X0Y111_CLUT (
.I0(CLBLL_L_X2Y120_SLICE_X0Y120_CO6),
.I1(CLBLM_R_X3Y120_SLICE_X3Y120_BO6),
.I2(RIOB33_X105Y127_IOB_X1Y128_I),
.I3(RIOB33_X105Y137_IOB_X1Y137_I),
.I4(RIOB33_X105Y129_IOB_X1Y129_I),
.I5(1'b1),
.O5(CLBLL_L_X2Y111_SLICE_X0Y111_CO5),
.O6(CLBLL_L_X2Y111_SLICE_X0Y111_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hffddfffffffcffff)
  ) CLBLL_L_X2Y111_SLICE_X0Y111_BLUT (
.I0(CLBLL_L_X2Y119_SLICE_X0Y119_BO6),
.I1(RIOB33_X105Y127_IOB_X1Y128_I),
.I2(CLBLL_L_X4Y121_SLICE_X5Y121_BO5),
.I3(RIOB33_X105Y129_IOB_X1Y129_I),
.I4(RIOB33_X105Y137_IOB_X1Y137_I),
.I5(1'b1),
.O5(CLBLL_L_X2Y111_SLICE_X0Y111_BO5),
.O6(CLBLL_L_X2Y111_SLICE_X0Y111_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffeefffffefeffff)
  ) CLBLL_L_X2Y111_SLICE_X0Y111_ALUT (
.I0(RIOB33_X105Y129_IOB_X1Y129_I),
.I1(RIOB33_X105Y127_IOB_X1Y128_I),
.I2(CLBLL_L_X4Y120_SLICE_X4Y120_AO6),
.I3(CLBLM_R_X3Y119_SLICE_X2Y119_AO6),
.I4(RIOB33_X105Y137_IOB_X1Y137_I),
.I5(1'b1),
.O5(CLBLL_L_X2Y111_SLICE_X0Y111_AO5),
.O6(CLBLL_L_X2Y111_SLICE_X0Y111_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y111_SLICE_X1Y111_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y111_SLICE_X1Y111_DO5),
.O6(CLBLL_L_X2Y111_SLICE_X1Y111_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y111_SLICE_X1Y111_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y111_SLICE_X1Y111_CO5),
.O6(CLBLL_L_X2Y111_SLICE_X1Y111_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y111_SLICE_X1Y111_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y111_SLICE_X1Y111_BO5),
.O6(CLBLL_L_X2Y111_SLICE_X1Y111_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y111_SLICE_X1Y111_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y111_SLICE_X1Y111_AO5),
.O6(CLBLL_L_X2Y111_SLICE_X1Y111_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y112_SLICE_X0Y112_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y112_SLICE_X0Y112_DO5),
.O6(CLBLL_L_X2Y112_SLICE_X0Y112_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y112_SLICE_X0Y112_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y112_SLICE_X0Y112_CO5),
.O6(CLBLL_L_X2Y112_SLICE_X0Y112_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y112_SLICE_X0Y112_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y112_SLICE_X0Y112_BO5),
.O6(CLBLL_L_X2Y112_SLICE_X0Y112_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y112_SLICE_X0Y112_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y112_SLICE_X0Y112_AO5),
.O6(CLBLL_L_X2Y112_SLICE_X0Y112_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X2Y112_SLICE_X1Y112_A5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X2Y112_SLICE_X1Y112_CO6),
.Q(CLBLL_L_X2Y112_SLICE_X1Y112_A5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X2Y112_SLICE_X1Y112_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X2Y112_SLICE_X1Y112_AO6),
.Q(CLBLL_L_X2Y112_SLICE_X1Y112_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X2Y112_SLICE_X1Y112_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X2Y112_SLICE_X1Y112_BO6),
.Q(CLBLL_L_X2Y112_SLICE_X1Y112_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y112_SLICE_X1Y112_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y112_SLICE_X1Y112_DO5),
.O6(CLBLL_L_X2Y112_SLICE_X1Y112_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hcecd0a05aaffaaff)
  ) CLBLL_L_X2Y112_SLICE_X1Y112_CLUT (
.I0(CLBLM_L_X10Y113_SLICE_X13Y113_BO6),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(CLBLM_R_X3Y112_SLICE_X2Y112_CO6),
.I3(CLBLL_L_X2Y112_SLICE_X1Y112_A5Q),
.I4(CLBLM_R_X5Y119_SLICE_X6Y119_B5Q),
.I5(1'b1),
.O5(CLBLL_L_X2Y112_SLICE_X1Y112_CO5),
.O6(CLBLL_L_X2Y112_SLICE_X1Y112_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hcccc0000dddd1111)
  ) CLBLL_L_X2Y112_SLICE_X1Y112_BLUT (
.I0(CLBLM_R_X3Y112_SLICE_X3Y112_B5Q),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(1'b1),
.I3(1'b1),
.I4(CLBLL_L_X2Y113_SLICE_X1Y113_CQ),
.I5(CLBLM_L_X8Y112_SLICE_X10Y112_CQ),
.O5(CLBLL_L_X2Y112_SLICE_X1Y112_BO5),
.O6(CLBLL_L_X2Y112_SLICE_X1Y112_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f8f0f800080008)
  ) CLBLL_L_X2Y112_SLICE_X1Y112_ALUT (
.I0(CLBLM_L_X8Y112_SLICE_X10Y112_CQ),
.I1(CLBLL_L_X2Y112_SLICE_X1Y112_BQ),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(RIOB33_X105Y105_IOB_X1Y105_I),
.I4(1'b1),
.I5(CLBLM_R_X3Y114_SLICE_X2Y114_BQ),
.O5(CLBLL_L_X2Y112_SLICE_X1Y112_AO5),
.O6(CLBLL_L_X2Y112_SLICE_X1Y112_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y113_SLICE_X0Y113_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y113_SLICE_X0Y113_DO5),
.O6(CLBLL_L_X2Y113_SLICE_X0Y113_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y113_SLICE_X0Y113_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y113_SLICE_X0Y113_CO5),
.O6(CLBLL_L_X2Y113_SLICE_X0Y113_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y113_SLICE_X0Y113_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y113_SLICE_X0Y113_BO5),
.O6(CLBLL_L_X2Y113_SLICE_X0Y113_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffaf8c8c8c8c)
  ) CLBLL_L_X2Y113_SLICE_X0Y113_ALUT (
.I0(RIOB33_X105Y129_IOB_X1Y129_I),
.I1(CLBLL_L_X2Y113_SLICE_X1Y113_CQ),
.I2(RIOB33_X105Y137_IOB_X1Y137_I),
.I3(CLBLL_L_X4Y120_SLICE_X4Y120_BO6),
.I4(RIOB33_X105Y127_IOB_X1Y128_I),
.I5(1'b1),
.O5(CLBLL_L_X2Y113_SLICE_X0Y113_AO5),
.O6(CLBLL_L_X2Y113_SLICE_X0Y113_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X2Y113_SLICE_X1Y113_C5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X2Y113_SLICE_X1Y113_CO5),
.Q(CLBLL_L_X2Y113_SLICE_X1Y113_C5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X2Y113_SLICE_X1Y113_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X2Y113_SLICE_X1Y113_AO6),
.Q(CLBLL_L_X2Y113_SLICE_X1Y113_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X2Y113_SLICE_X1Y113_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X2Y113_SLICE_X1Y113_BO6),
.Q(CLBLL_L_X2Y113_SLICE_X1Y113_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X2Y113_SLICE_X1Y113_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X2Y113_SLICE_X1Y113_CO6),
.Q(CLBLL_L_X2Y113_SLICE_X1Y113_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y113_SLICE_X1Y113_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y113_SLICE_X1Y113_DO5),
.O6(CLBLL_L_X2Y113_SLICE_X1Y113_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'haf05af058888dddd)
  ) CLBLL_L_X2Y113_SLICE_X1Y113_CLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLL_L_X4Y113_SLICE_X4Y113_BQ),
.I2(CLBLL_L_X2Y119_SLICE_X0Y119_BO6),
.I3(CLBLM_R_X3Y114_SLICE_X3Y114_BQ),
.I4(CLBLL_L_X2Y114_SLICE_X1Y114_DO6),
.I5(1'b1),
.O5(CLBLL_L_X2Y113_SLICE_X1Y113_CO5),
.O6(CLBLL_L_X2Y113_SLICE_X1Y113_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hff000303ff000c0c)
  ) CLBLL_L_X2Y113_SLICE_X1Y113_BLUT (
.I0(1'b1),
.I1(CLBLL_L_X4Y113_SLICE_X4Y113_BQ),
.I2(RIOB33_X105Y105_IOB_X1Y105_I),
.I3(CLBLL_L_X4Y116_SLICE_X4Y116_C5Q),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(CLBLM_R_X5Y112_SLICE_X6Y112_DO6),
.O5(CLBLL_L_X2Y113_SLICE_X1Y113_BO5),
.O6(CLBLL_L_X2Y113_SLICE_X1Y113_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0fff0fff0aaf0aa)
  ) CLBLL_L_X2Y113_SLICE_X1Y113_ALUT (
.I0(CLBLM_R_X7Y120_SLICE_X9Y120_DQ),
.I1(1'b1),
.I2(LIOB33_X0Y79_IOB_X0Y79_I),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(1'b1),
.I5(CLBLL_L_X2Y113_SLICE_X1Y113_AQ),
.O5(CLBLL_L_X2Y113_SLICE_X1Y113_AO5),
.O6(CLBLL_L_X2Y113_SLICE_X1Y113_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y114_SLICE_X0Y114_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y114_SLICE_X0Y114_DO5),
.O6(CLBLL_L_X2Y114_SLICE_X0Y114_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y114_SLICE_X0Y114_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y114_SLICE_X0Y114_CO5),
.O6(CLBLL_L_X2Y114_SLICE_X0Y114_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y114_SLICE_X0Y114_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y114_SLICE_X0Y114_BO5),
.O6(CLBLL_L_X2Y114_SLICE_X0Y114_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y114_SLICE_X0Y114_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y114_SLICE_X0Y114_AO5),
.O6(CLBLL_L_X2Y114_SLICE_X0Y114_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X2Y114_SLICE_X1Y114_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X2Y114_SLICE_X1Y114_AO6),
.Q(CLBLL_L_X2Y114_SLICE_X1Y114_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hdfffffffffffffff)
  ) CLBLL_L_X2Y114_SLICE_X1Y114_DLUT (
.I0(CLBLM_R_X3Y114_SLICE_X2Y114_CQ),
.I1(CLBLM_L_X8Y116_SLICE_X10Y116_AO6),
.I2(CLBLM_R_X5Y111_SLICE_X7Y111_DO6),
.I3(CLBLL_L_X2Y115_SLICE_X1Y115_BQ),
.I4(CLBLL_L_X2Y114_SLICE_X1Y114_AQ),
.I5(CLBLM_R_X3Y114_SLICE_X2Y114_AQ),
.O5(CLBLL_L_X2Y114_SLICE_X1Y114_DO5),
.O6(CLBLL_L_X2Y114_SLICE_X1Y114_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hfff7f7f700000800)
  ) CLBLL_L_X2Y114_SLICE_X1Y114_CLUT (
.I0(CLBLM_R_X3Y114_SLICE_X2Y114_CQ),
.I1(CLBLM_R_X3Y114_SLICE_X2Y114_AQ),
.I2(CLBLM_R_X5Y111_SLICE_X7Y111_DO6),
.I3(CLBLL_L_X2Y115_SLICE_X1Y115_BQ),
.I4(CLBLL_L_X2Y114_SLICE_X1Y114_AQ),
.I5(1'b1),
.O5(CLBLL_L_X2Y114_SLICE_X1Y114_CO5),
.O6(CLBLL_L_X2Y114_SLICE_X1Y114_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h00ff4c3380008000)
  ) CLBLL_L_X2Y114_SLICE_X1Y114_BLUT (
.I0(CLBLL_L_X2Y115_SLICE_X1Y115_BQ),
.I1(CLBLM_R_X3Y114_SLICE_X2Y114_CQ),
.I2(CLBLL_L_X2Y114_SLICE_X1Y114_AQ),
.I3(CLBLM_R_X3Y114_SLICE_X2Y114_AQ),
.I4(CLBLM_R_X5Y119_SLICE_X7Y119_AO6),
.I5(1'b1),
.O5(CLBLL_L_X2Y114_SLICE_X1Y114_BO5),
.O6(CLBLL_L_X2Y114_SLICE_X1Y114_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hff00ff0022222020)
  ) CLBLL_L_X2Y114_SLICE_X1Y114_ALUT (
.I0(RIOB33_X105Y105_IOB_X1Y105_I),
.I1(CLBLM_R_X5Y115_SLICE_X7Y115_AQ),
.I2(CLBLL_L_X2Y114_SLICE_X1Y114_AQ),
.I3(CLBLM_R_X3Y114_SLICE_X3Y114_AQ),
.I4(CLBLL_L_X2Y114_SLICE_X1Y114_CO5),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLL_L_X2Y114_SLICE_X1Y114_AO5),
.O6(CLBLL_L_X2Y114_SLICE_X1Y114_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y115_SLICE_X0Y115_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y115_SLICE_X0Y115_DO5),
.O6(CLBLL_L_X2Y115_SLICE_X0Y115_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y115_SLICE_X0Y115_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y115_SLICE_X0Y115_CO5),
.O6(CLBLL_L_X2Y115_SLICE_X0Y115_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y115_SLICE_X0Y115_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y115_SLICE_X0Y115_BO5),
.O6(CLBLL_L_X2Y115_SLICE_X0Y115_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y115_SLICE_X0Y115_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y115_SLICE_X0Y115_AO5),
.O6(CLBLL_L_X2Y115_SLICE_X0Y115_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X2Y115_SLICE_X1Y115_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X2Y115_SLICE_X1Y115_AO6),
.Q(CLBLL_L_X2Y115_SLICE_X1Y115_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X2Y115_SLICE_X1Y115_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X2Y115_SLICE_X1Y115_BO6),
.Q(CLBLL_L_X2Y115_SLICE_X1Y115_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y115_SLICE_X1Y115_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y115_SLICE_X1Y115_DO5),
.O6(CLBLL_L_X2Y115_SLICE_X1Y115_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y115_SLICE_X1Y115_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y115_SLICE_X1Y115_CO5),
.O6(CLBLL_L_X2Y115_SLICE_X1Y115_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'ha0e4a0b1a0a0a0a0)
  ) CLBLL_L_X2Y115_SLICE_X1Y115_BLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLL_L_X2Y115_SLICE_X1Y115_BQ),
.I2(CLBLM_R_X3Y123_SLICE_X3Y123_AQ),
.I3(CLBLM_R_X5Y115_SLICE_X7Y115_AQ),
.I4(CLBLL_L_X2Y114_SLICE_X1Y114_CO6),
.I5(RIOB33_X105Y105_IOB_X1Y105_I),
.O5(CLBLL_L_X2Y115_SLICE_X1Y115_BO5),
.O6(CLBLL_L_X2Y115_SLICE_X1Y115_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hff00ff00e2e2aaaa)
  ) CLBLL_L_X2Y115_SLICE_X1Y115_ALUT (
.I0(CLBLM_R_X5Y113_SLICE_X6Y113_BQ),
.I1(CLBLM_L_X8Y112_SLICE_X10Y112_CQ),
.I2(CLBLL_L_X2Y115_SLICE_X1Y115_AQ),
.I3(CLBLM_R_X3Y113_SLICE_X2Y113_AQ),
.I4(CLBLL_L_X2Y112_SLICE_X1Y112_BQ),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLL_L_X2Y115_SLICE_X1Y115_AO5),
.O6(CLBLL_L_X2Y115_SLICE_X1Y115_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y116_SLICE_X0Y116_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y116_SLICE_X0Y116_DO5),
.O6(CLBLL_L_X2Y116_SLICE_X0Y116_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y116_SLICE_X0Y116_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y116_SLICE_X0Y116_CO5),
.O6(CLBLL_L_X2Y116_SLICE_X0Y116_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y116_SLICE_X0Y116_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y116_SLICE_X0Y116_BO5),
.O6(CLBLL_L_X2Y116_SLICE_X0Y116_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y116_SLICE_X0Y116_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y116_SLICE_X0Y116_AO5),
.O6(CLBLL_L_X2Y116_SLICE_X0Y116_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X2Y116_SLICE_X1Y116_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X2Y116_SLICE_X1Y116_AO6),
.Q(CLBLL_L_X2Y116_SLICE_X1Y116_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y116_SLICE_X1Y116_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y116_SLICE_X1Y116_DO5),
.O6(CLBLL_L_X2Y116_SLICE_X1Y116_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y116_SLICE_X1Y116_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y116_SLICE_X1Y116_CO5),
.O6(CLBLL_L_X2Y116_SLICE_X1Y116_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y116_SLICE_X1Y116_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y116_SLICE_X1Y116_BO5),
.O6(CLBLL_L_X2Y116_SLICE_X1Y116_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h8888bbb8bbb8bbb8)
  ) CLBLL_L_X2Y116_SLICE_X1Y116_ALUT (
.I0(CLBLL_L_X2Y115_SLICE_X1Y115_BQ),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(CLBLL_L_X2Y116_SLICE_X1Y116_AQ),
.I3(CLBLM_R_X3Y113_SLICE_X2Y113_BQ),
.I4(CLBLL_L_X2Y112_SLICE_X1Y112_BQ),
.I5(CLBLM_L_X8Y112_SLICE_X10Y112_CQ),
.O5(CLBLL_L_X2Y116_SLICE_X1Y116_AO5),
.O6(CLBLL_L_X2Y116_SLICE_X1Y116_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X2Y117_SLICE_X0Y117_A5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X2Y117_SLICE_X0Y117_DO5),
.Q(CLBLL_L_X2Y117_SLICE_X0Y117_A5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X2Y117_SLICE_X0Y117_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X2Y117_SLICE_X0Y117_AO6),
.Q(CLBLL_L_X2Y117_SLICE_X0Y117_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X2Y117_SLICE_X0Y117_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X2Y117_SLICE_X0Y117_BO6),
.Q(CLBLL_L_X2Y117_SLICE_X0Y117_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X2Y117_SLICE_X0Y117_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X2Y117_SLICE_X0Y117_CO6),
.Q(CLBLL_L_X2Y117_SLICE_X0Y117_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hc0000000eaaa0000)
  ) CLBLL_L_X2Y117_SLICE_X0Y117_DLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLL_L_X2Y117_SLICE_X0Y117_CQ),
.I2(CLBLL_L_X2Y117_SLICE_X0Y117_AQ),
.I3(CLBLL_L_X2Y117_SLICE_X0Y117_BQ),
.I4(CLBLL_L_X2Y117_SLICE_X1Y117_BQ),
.I5(1'b1),
.O5(CLBLL_L_X2Y117_SLICE_X0Y117_DO5),
.O6(CLBLL_L_X2Y117_SLICE_X0Y117_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'he4b1e4b1a0a0a0a0)
  ) CLBLL_L_X2Y117_SLICE_X0Y117_CLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLL_L_X2Y117_SLICE_X0Y117_CQ),
.I2(CLBLL_L_X2Y117_SLICE_X0Y117_BQ),
.I3(CLBLL_L_X2Y114_SLICE_X1Y114_DO6),
.I4(1'b1),
.I5(CLBLM_R_X3Y117_SLICE_X2Y117_BO6),
.O5(CLBLL_L_X2Y117_SLICE_X0Y117_CO5),
.O6(CLBLL_L_X2Y117_SLICE_X0Y117_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hffc400c4ff040004)
  ) CLBLL_L_X2Y117_SLICE_X0Y117_BLUT (
.I0(CLBLL_L_X2Y117_SLICE_X0Y117_DO6),
.I1(CLBLM_R_X3Y117_SLICE_X2Y117_BO6),
.I2(CLBLL_L_X2Y117_SLICE_X1Y117_CO6),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLM_R_X3Y116_SLICE_X3Y116_AQ),
.I5(CLBLL_L_X2Y117_SLICE_X0Y117_BQ),
.O5(CLBLL_L_X2Y117_SLICE_X0Y117_BO5),
.O6(CLBLL_L_X2Y117_SLICE_X0Y117_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hff00c0c0ff004848)
  ) CLBLL_L_X2Y117_SLICE_X0Y117_ALUT (
.I0(CLBLL_L_X2Y117_SLICE_X0Y117_CQ),
.I1(CLBLM_R_X3Y117_SLICE_X2Y117_BO6),
.I2(CLBLL_L_X2Y117_SLICE_X0Y117_AQ),
.I3(CLBLL_L_X4Y117_SLICE_X4Y117_BQ),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(CLBLL_L_X2Y114_SLICE_X1Y114_DO6),
.O5(CLBLL_L_X2Y117_SLICE_X0Y117_AO5),
.O6(CLBLL_L_X2Y117_SLICE_X0Y117_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X2Y117_SLICE_X1Y117_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X2Y117_SLICE_X1Y117_AO6),
.Q(CLBLL_L_X2Y117_SLICE_X1Y117_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X2Y117_SLICE_X1Y117_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X2Y117_SLICE_X1Y117_BO6),
.Q(CLBLL_L_X2Y117_SLICE_X1Y117_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hf5fffffff5ffffff)
  ) CLBLL_L_X2Y117_SLICE_X1Y117_DLUT (
.I0(CLBLM_R_X5Y111_SLICE_X7Y111_DO6),
.I1(1'b1),
.I2(CLBLM_L_X8Y116_SLICE_X10Y116_AO6),
.I3(CLBLL_L_X2Y117_SLICE_X0Y117_CQ),
.I4(CLBLL_L_X2Y114_SLICE_X1Y114_BO5),
.I5(1'b1),
.O5(CLBLL_L_X2Y117_SLICE_X1Y117_DO5),
.O6(CLBLL_L_X2Y117_SLICE_X1Y117_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffff7fffffff)
  ) CLBLL_L_X2Y117_SLICE_X1Y117_CLUT (
.I0(CLBLL_L_X2Y117_SLICE_X0Y117_AQ),
.I1(CLBLM_R_X5Y111_SLICE_X7Y111_DO6),
.I2(CLBLL_L_X2Y117_SLICE_X0Y117_CQ),
.I3(CLBLL_L_X2Y117_SLICE_X1Y117_BQ),
.I4(CLBLL_L_X2Y114_SLICE_X1Y114_BO5),
.I5(CLBLM_L_X8Y116_SLICE_X10Y116_AO6),
.O5(CLBLL_L_X2Y117_SLICE_X1Y117_CO5),
.O6(CLBLL_L_X2Y117_SLICE_X1Y117_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf909f000fc0cf000)
  ) CLBLL_L_X2Y117_SLICE_X1Y117_BLUT (
.I0(CLBLL_L_X2Y117_SLICE_X1Y117_DO6),
.I1(CLBLL_L_X2Y117_SLICE_X1Y117_BQ),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLM_L_X10Y117_SLICE_X12Y117_AQ),
.I4(CLBLM_R_X3Y117_SLICE_X2Y117_BO6),
.I5(CLBLL_L_X2Y117_SLICE_X0Y117_AQ),
.O5(CLBLL_L_X2Y117_SLICE_X1Y117_BO5),
.O6(CLBLL_L_X2Y117_SLICE_X1Y117_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hb8b8bb88bb88bb88)
  ) CLBLL_L_X2Y117_SLICE_X1Y117_ALUT (
.I0(CLBLM_R_X3Y116_SLICE_X2Y116_BQ),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(CLBLL_L_X2Y117_SLICE_X1Y117_AQ),
.I3(CLBLM_R_X5Y116_SLICE_X6Y116_BQ),
.I4(CLBLL_L_X2Y112_SLICE_X1Y112_BQ),
.I5(CLBLM_L_X8Y112_SLICE_X10Y112_CQ),
.O5(CLBLL_L_X2Y117_SLICE_X1Y117_AO5),
.O6(CLBLL_L_X2Y117_SLICE_X1Y117_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffffffffafffe)
  ) CLBLL_L_X2Y118_SLICE_X0Y118_DLUT (
.I0(CLBLL_L_X2Y118_SLICE_X0Y118_AO6),
.I1(CLBLL_L_X2Y117_SLICE_X1Y117_AQ),
.I2(CLBLL_L_X2Y118_SLICE_X0Y118_CO6),
.I3(CLBLM_R_X3Y117_SLICE_X2Y117_CO6),
.I4(CLBLM_R_X3Y121_SLICE_X2Y121_AO6),
.I5(CLBLL_L_X2Y118_SLICE_X0Y118_BO6),
.O5(CLBLL_L_X2Y118_SLICE_X0Y118_DO5),
.O6(CLBLL_L_X2Y118_SLICE_X0Y118_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000004000000000)
  ) CLBLL_L_X2Y118_SLICE_X0Y118_CLUT (
.I0(CLBLM_R_X3Y122_SLICE_X3Y122_AO6),
.I1(RIOB33_X105Y133_IOB_X1Y133_I),
.I2(RIOB33_X105Y131_IOB_X1Y131_I),
.I3(RIOB33_X105Y133_IOB_X1Y134_I),
.I4(RIOB33_X105Y131_IOB_X1Y132_I),
.I5(CLBLM_R_X7Y119_SLICE_X8Y119_AQ),
.O5(CLBLL_L_X2Y118_SLICE_X0Y118_CO5),
.O6(CLBLL_L_X2Y118_SLICE_X0Y118_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffff05450044)
  ) CLBLL_L_X2Y118_SLICE_X0Y118_BLUT (
.I0(CLBLM_R_X3Y124_SLICE_X2Y124_AO5),
.I1(LIOB33_X0Y67_IOB_X0Y68_I),
.I2(CLBLL_L_X2Y120_SLICE_X1Y120_AO6),
.I3(CLBLL_L_X2Y121_SLICE_X1Y121_BO6),
.I4(CLBLM_R_X5Y119_SLICE_X6Y119_CQ),
.I5(CLBLL_L_X2Y113_SLICE_X0Y113_AO5),
.O5(CLBLL_L_X2Y118_SLICE_X0Y118_BO5),
.O6(CLBLL_L_X2Y118_SLICE_X0Y118_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000320010)
  ) CLBLL_L_X2Y118_SLICE_X0Y118_ALUT (
.I0(RIOB33_X105Y135_IOB_X1Y136_I),
.I1(CLBLM_R_X3Y122_SLICE_X3Y122_AO5),
.I2(CLBLL_L_X4Y117_SLICE_X4Y117_AQ),
.I3(CLBLL_L_X2Y121_SLICE_X1Y121_BO6),
.I4(RIOB33_X105Y113_IOB_X1Y113_I),
.I5(RIOB33_X105Y135_IOB_X1Y135_I),
.O5(CLBLL_L_X2Y118_SLICE_X0Y118_AO5),
.O6(CLBLL_L_X2Y118_SLICE_X0Y118_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y118_SLICE_X1Y118_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y118_SLICE_X1Y118_DO5),
.O6(CLBLL_L_X2Y118_SLICE_X1Y118_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0404040455550404)
  ) CLBLL_L_X2Y118_SLICE_X1Y118_CLUT (
.I0(CLBLM_R_X3Y124_SLICE_X2Y124_AO6),
.I1(CLBLL_L_X4Y118_SLICE_X5Y118_BQ),
.I2(CLBLL_L_X2Y121_SLICE_X1Y121_BO5),
.I3(1'b1),
.I4(RIOB33_X105Y105_IOB_X1Y106_I),
.I5(CLBLL_L_X2Y121_SLICE_X1Y121_BO6),
.O5(CLBLL_L_X2Y118_SLICE_X1Y118_CO5),
.O6(CLBLL_L_X2Y118_SLICE_X1Y118_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffffffffddcc)
  ) CLBLL_L_X2Y118_SLICE_X1Y118_BLUT (
.I0(CLBLM_R_X3Y122_SLICE_X2Y122_BO5),
.I1(CLBLM_R_X3Y118_SLICE_X2Y118_CO6),
.I2(1'b1),
.I3(CLBLM_R_X5Y116_SLICE_X7Y116_AQ),
.I4(CLBLL_L_X2Y118_SLICE_X1Y118_AO6),
.I5(CLBLL_L_X2Y118_SLICE_X1Y118_CO6),
.O5(CLBLL_L_X2Y118_SLICE_X1Y118_BO5),
.O6(CLBLL_L_X2Y118_SLICE_X1Y118_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h003000300030aaba)
  ) CLBLL_L_X2Y118_SLICE_X1Y118_ALUT (
.I0(CLBLL_L_X2Y112_SLICE_X1Y112_A5Q),
.I1(CLBLL_L_X2Y121_SLICE_X0Y121_BO6),
.I2(CLBLM_R_X5Y115_SLICE_X6Y115_AQ),
.I3(CLBLM_R_X3Y122_SLICE_X3Y122_AO6),
.I4(CLBLM_R_X3Y124_SLICE_X2Y124_AO6),
.I5(CLBLL_L_X2Y120_SLICE_X1Y120_AO6),
.O5(CLBLL_L_X2Y118_SLICE_X1Y118_AO5),
.O6(CLBLL_L_X2Y118_SLICE_X1Y118_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hcfcccfccefeeefee)
  ) CLBLL_L_X2Y119_SLICE_X0Y119_DLUT (
.I0(CLBLL_L_X4Y117_SLICE_X4Y117_AQ),
.I1(CLBLM_R_X3Y117_SLICE_X2Y117_CO6),
.I2(CLBLL_L_X2Y122_SLICE_X0Y122_AO6),
.I3(RIOB33_X105Y113_IOB_X1Y113_I),
.I4(1'b1),
.I5(CLBLL_L_X2Y120_SLICE_X0Y120_AO6),
.O5(CLBLL_L_X2Y119_SLICE_X0Y119_DO5),
.O6(CLBLL_L_X2Y119_SLICE_X0Y119_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hbbfbbbfbaafaaafa)
  ) CLBLL_L_X2Y119_SLICE_X0Y119_CLUT (
.I0(CLBLL_L_X2Y119_SLICE_X0Y119_AO6),
.I1(CLBLL_L_X2Y121_SLICE_X0Y121_AO6),
.I2(CLBLL_L_X2Y117_SLICE_X1Y117_AQ),
.I3(CLBLM_R_X3Y121_SLICE_X2Y121_AO6),
.I4(1'b1),
.I5(LIOB33_X0Y67_IOB_X0Y68_I),
.O5(CLBLL_L_X2Y119_SLICE_X0Y119_CO5),
.O6(CLBLL_L_X2Y119_SLICE_X0Y119_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000055051101)
  ) CLBLL_L_X2Y119_SLICE_X0Y119_BLUT (
.I0(CLBLL_L_X2Y119_SLICE_X0Y119_DO6),
.I1(CLBLM_R_X7Y119_SLICE_X8Y119_AQ),
.I2(CLBLM_R_X3Y121_SLICE_X2Y121_DO6),
.I3(CLBLL_L_X2Y120_SLICE_X0Y120_BO6),
.I4(CLBLL_L_X2Y120_SLICE_X0Y120_AO5),
.I5(CLBLL_L_X2Y119_SLICE_X0Y119_CO6),
.O5(CLBLL_L_X2Y119_SLICE_X0Y119_BO5),
.O6(CLBLL_L_X2Y119_SLICE_X0Y119_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hcdcd05cdcccc00cc)
  ) CLBLL_L_X2Y119_SLICE_X0Y119_ALUT (
.I0(CLBLM_R_X3Y124_SLICE_X2Y124_AO5),
.I1(CLBLL_L_X2Y113_SLICE_X1Y113_CQ),
.I2(CLBLL_L_X2Y120_SLICE_X1Y120_AO6),
.I3(RIOB33_X105Y137_IOB_X1Y137_I),
.I4(RIOB33_X105Y129_IOB_X1Y129_I),
.I5(CLBLM_R_X5Y119_SLICE_X6Y119_CQ),
.O5(CLBLL_L_X2Y119_SLICE_X0Y119_AO5),
.O6(CLBLL_L_X2Y119_SLICE_X0Y119_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h5f55dfdd0f00cfcc)
  ) CLBLL_L_X2Y119_SLICE_X1Y119_DLUT (
.I0(CLBLL_L_X2Y121_SLICE_X1Y121_AO6),
.I1(RIOB33_X105Y105_IOB_X1Y106_I),
.I2(CLBLM_R_X3Y122_SLICE_X2Y122_BO5),
.I3(CLBLM_R_X5Y116_SLICE_X7Y116_AQ),
.I4(CLBLL_L_X2Y122_SLICE_X0Y122_AO6),
.I5(CLBLL_L_X4Y118_SLICE_X5Y118_BQ),
.O5(CLBLL_L_X2Y119_SLICE_X1Y119_DO5),
.O6(CLBLL_L_X2Y119_SLICE_X1Y119_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000100)
  ) CLBLL_L_X2Y119_SLICE_X1Y119_CLUT (
.I0(CLBLL_L_X2Y118_SLICE_X1Y118_BO6),
.I1(CLBLL_L_X2Y122_SLICE_X0Y122_BO6),
.I2(CLBLL_L_X2Y118_SLICE_X0Y118_DO6),
.I3(CLBLL_L_X2Y120_SLICE_X1Y120_BO6),
.I4(CLBLL_L_X2Y121_SLICE_X1Y121_CO6),
.I5(CLBLL_L_X4Y118_SLICE_X4Y118_CO6),
.O5(CLBLL_L_X2Y119_SLICE_X1Y119_CO5),
.O6(CLBLL_L_X2Y119_SLICE_X1Y119_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000100000000)
  ) CLBLL_L_X2Y119_SLICE_X1Y119_BLUT (
.I0(CLBLL_L_X4Y120_SLICE_X5Y120_DO6),
.I1(CLBLM_R_X3Y120_SLICE_X3Y120_BO6),
.I2(CLBLM_R_X3Y121_SLICE_X2Y121_CO6),
.I3(CLBLL_L_X4Y120_SLICE_X4Y120_AO6),
.I4(CLBLL_L_X4Y120_SLICE_X4Y120_BO6),
.I5(CLBLL_L_X2Y119_SLICE_X1Y119_CO6),
.O5(CLBLL_L_X2Y119_SLICE_X1Y119_BO5),
.O6(CLBLL_L_X2Y119_SLICE_X1Y119_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h41400000feffffff)
  ) CLBLL_L_X2Y119_SLICE_X1Y119_ALUT (
.I0(CLBLM_R_X3Y124_SLICE_X2Y124_AO6),
.I1(RIOB33_X105Y131_IOB_X1Y132_I),
.I2(RIOB33_X105Y133_IOB_X1Y133_I),
.I3(RIOB33_X105Y133_IOB_X1Y134_I),
.I4(RIOB33_X105Y131_IOB_X1Y131_I),
.I5(1'b1),
.O5(CLBLL_L_X2Y119_SLICE_X1Y119_AO5),
.O6(CLBLL_L_X2Y119_SLICE_X1Y119_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y120_SLICE_X0Y120_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y120_SLICE_X0Y120_DO5),
.O6(CLBLL_L_X2Y120_SLICE_X0Y120_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffffffffffffe)
  ) CLBLL_L_X2Y120_SLICE_X0Y120_CLUT (
.I0(CLBLM_R_X5Y122_SLICE_X6Y122_CO6),
.I1(CLBLL_L_X4Y118_SLICE_X4Y118_CO6),
.I2(CLBLL_L_X2Y122_SLICE_X0Y122_CO6),
.I3(CLBLM_R_X3Y118_SLICE_X2Y118_DO6),
.I4(CLBLL_L_X2Y119_SLICE_X1Y119_DO6),
.I5(CLBLL_L_X2Y121_SLICE_X1Y121_CO6),
.O5(CLBLL_L_X2Y120_SLICE_X0Y120_CO5),
.O6(CLBLL_L_X2Y120_SLICE_X0Y120_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hbabaaaaaabaaaaaa)
  ) CLBLL_L_X2Y120_SLICE_X0Y120_BLUT (
.I0(CLBLL_L_X4Y122_SLICE_X5Y122_DO6),
.I1(CLBLM_R_X3Y124_SLICE_X2Y124_AO6),
.I2(RIOB33_X105Y131_IOB_X1Y132_I),
.I3(RIOB33_X105Y133_IOB_X1Y134_I),
.I4(RIOB33_X105Y131_IOB_X1Y131_I),
.I5(RIOB33_X105Y133_IOB_X1Y133_I),
.O5(CLBLL_L_X2Y120_SLICE_X0Y120_BO5),
.O6(CLBLL_L_X2Y120_SLICE_X0Y120_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffdffffffffdffff)
  ) CLBLL_L_X2Y120_SLICE_X0Y120_ALUT (
.I0(RIOB33_X105Y133_IOB_X1Y133_I),
.I1(CLBLM_R_X3Y122_SLICE_X3Y122_AO6),
.I2(RIOB33_X105Y131_IOB_X1Y132_I),
.I3(RIOB33_X105Y133_IOB_X1Y134_I),
.I4(RIOB33_X105Y131_IOB_X1Y131_I),
.I5(1'b1),
.O5(CLBLL_L_X2Y120_SLICE_X0Y120_AO5),
.O6(CLBLL_L_X2Y120_SLICE_X0Y120_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffffffcfcfcfe)
  ) CLBLL_L_X2Y120_SLICE_X1Y120_DLUT (
.I0(CLBLL_L_X2Y120_SLICE_X1Y120_CO6),
.I1(CLBLM_R_X3Y119_SLICE_X3Y119_CO6),
.I2(CLBLM_R_X3Y120_SLICE_X2Y120_DO6),
.I3(CLBLL_L_X2Y120_SLICE_X1Y120_AO5),
.I4(CLBLL_L_X4Y122_SLICE_X5Y122_DO6),
.I5(CLBLM_R_X3Y121_SLICE_X3Y121_DO6),
.O5(CLBLL_L_X2Y120_SLICE_X1Y120_DO5),
.O6(CLBLL_L_X2Y120_SLICE_X1Y120_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000080000000)
  ) CLBLL_L_X2Y120_SLICE_X1Y120_CLUT (
.I0(CLBLL_L_X2Y121_SLICE_X1Y121_AO6),
.I1(CLBLM_R_X3Y122_SLICE_X2Y122_AO6),
.I2(CLBLM_R_X3Y121_SLICE_X2Y121_AO5),
.I3(CLBLL_L_X4Y121_SLICE_X4Y121_CO5),
.I4(CLBLL_L_X2Y120_SLICE_X0Y120_AO6),
.I5(CLBLM_R_X3Y122_SLICE_X2Y122_CO6),
.O5(CLBLL_L_X2Y120_SLICE_X1Y120_CO5),
.O6(CLBLL_L_X2Y120_SLICE_X1Y120_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffffffffff7f)
  ) CLBLL_L_X2Y120_SLICE_X1Y120_BLUT (
.I0(CLBLL_L_X4Y121_SLICE_X4Y121_CO5),
.I1(CLBLM_R_X3Y122_SLICE_X2Y122_AO6),
.I2(CLBLL_L_X2Y120_SLICE_X0Y120_AO6),
.I3(CLBLL_L_X4Y122_SLICE_X5Y122_DO6),
.I4(CLBLL_L_X2Y119_SLICE_X1Y119_AO6),
.I5(CLBLM_R_X3Y122_SLICE_X2Y122_CO6),
.O5(CLBLL_L_X2Y120_SLICE_X1Y120_BO5),
.O6(CLBLL_L_X2Y120_SLICE_X1Y120_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffdfffdf0000c000)
  ) CLBLL_L_X2Y120_SLICE_X1Y120_ALUT (
.I0(RIOB33_X105Y133_IOB_X1Y134_I),
.I1(RIOB33_X105Y133_IOB_X1Y133_I),
.I2(RIOB33_X105Y131_IOB_X1Y131_I),
.I3(RIOB33_X105Y131_IOB_X1Y132_I),
.I4(CLBLM_R_X3Y124_SLICE_X2Y124_AO6),
.I5(1'b1),
.O5(CLBLL_L_X2Y120_SLICE_X1Y120_AO5),
.O6(CLBLL_L_X2Y120_SLICE_X1Y120_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0303070300000500)
  ) CLBLL_L_X2Y121_SLICE_X0Y121_DLUT (
.I0(RIOB33_X105Y131_IOB_X1Y132_I),
.I1(CLBLL_L_X2Y120_SLICE_X1Y120_AO6),
.I2(CLBLM_R_X3Y124_SLICE_X2Y124_AO5),
.I3(CLBLL_L_X4Y117_SLICE_X4Y117_BQ),
.I4(CLBLL_L_X2Y121_SLICE_X0Y121_BO5),
.I5(CLBLL_L_X2Y117_SLICE_X0Y117_BQ),
.O5(CLBLL_L_X2Y121_SLICE_X0Y121_DO5),
.O6(CLBLL_L_X2Y121_SLICE_X0Y121_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h000010ff00001010)
  ) CLBLL_L_X2Y121_SLICE_X0Y121_CLUT (
.I0(RIOB33_X105Y131_IOB_X1Y132_I),
.I1(CLBLL_L_X2Y121_SLICE_X0Y121_BO5),
.I2(CLBLM_R_X5Y121_SLICE_X6Y121_B5Q),
.I3(CLBLL_L_X2Y121_SLICE_X0Y121_AO5),
.I4(CLBLM_R_X3Y124_SLICE_X2Y124_AO5),
.I5(LIOB33_X0Y53_IOB_X0Y54_I),
.O5(CLBLL_L_X2Y121_SLICE_X0Y121_CO5),
.O6(CLBLL_L_X2Y121_SLICE_X0Y121_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfff3ffff3fff3fff)
  ) CLBLL_L_X2Y121_SLICE_X0Y121_BLUT (
.I0(1'b1),
.I1(RIOB33_X105Y133_IOB_X1Y133_I),
.I2(RIOB33_X105Y131_IOB_X1Y131_I),
.I3(RIOB33_X105Y133_IOB_X1Y134_I),
.I4(RIOB33_X105Y131_IOB_X1Y132_I),
.I5(1'b1),
.O5(CLBLL_L_X2Y121_SLICE_X0Y121_BO5),
.O6(CLBLL_L_X2Y121_SLICE_X0Y121_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffbfffffcfffffff)
  ) CLBLL_L_X2Y121_SLICE_X0Y121_ALUT (
.I0(CLBLM_R_X3Y124_SLICE_X2Y124_AO5),
.I1(RIOB33_X105Y133_IOB_X1Y133_I),
.I2(RIOB33_X105Y131_IOB_X1Y131_I),
.I3(RIOB33_X105Y133_IOB_X1Y134_I),
.I4(RIOB33_X105Y131_IOB_X1Y132_I),
.I5(1'b1),
.O5(CLBLL_L_X2Y121_SLICE_X0Y121_AO5),
.O6(CLBLL_L_X2Y121_SLICE_X0Y121_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000200000)
  ) CLBLL_L_X2Y121_SLICE_X1Y121_DLUT (
.I0(CLBLM_R_X3Y122_SLICE_X2Y122_AO6),
.I1(CLBLM_R_X3Y122_SLICE_X2Y122_CO6),
.I2(CLBLL_L_X2Y121_SLICE_X1Y121_AO6),
.I3(CLBLL_L_X4Y121_SLICE_X4Y121_DO6),
.I4(CLBLM_R_X3Y121_SLICE_X2Y121_AO5),
.I5(CLBLL_L_X2Y120_SLICE_X1Y120_AO5),
.O5(CLBLL_L_X2Y121_SLICE_X1Y121_DO5),
.O6(CLBLL_L_X2Y121_SLICE_X1Y121_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000002)
  ) CLBLL_L_X2Y121_SLICE_X1Y121_CLUT (
.I0(CLBLM_R_X3Y122_SLICE_X2Y122_AO6),
.I1(CLBLM_R_X3Y122_SLICE_X2Y122_CO6),
.I2(CLBLL_L_X2Y121_SLICE_X1Y121_AO5),
.I3(CLBLL_L_X4Y121_SLICE_X4Y121_DO6),
.I4(CLBLL_L_X4Y122_SLICE_X5Y122_AO6),
.I5(CLBLL_L_X2Y119_SLICE_X1Y119_AO6),
.O5(CLBLL_L_X2Y121_SLICE_X1Y121_CO5),
.O6(CLBLL_L_X2Y121_SLICE_X1Y121_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hcffffffffffffff3)
  ) CLBLL_L_X2Y121_SLICE_X1Y121_BLUT (
.I0(1'b1),
.I1(RIOB33_X105Y133_IOB_X1Y134_I),
.I2(RIOB33_X105Y131_IOB_X1Y132_I),
.I3(RIOB33_X105Y131_IOB_X1Y131_I),
.I4(RIOB33_X105Y133_IOB_X1Y133_I),
.I5(1'b1),
.O5(CLBLL_L_X2Y121_SLICE_X1Y121_BO5),
.O6(CLBLL_L_X2Y121_SLICE_X1Y121_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffffb00004004)
  ) CLBLL_L_X2Y121_SLICE_X1Y121_ALUT (
.I0(CLBLM_R_X3Y124_SLICE_X2Y124_AO6),
.I1(RIOB33_X105Y133_IOB_X1Y134_I),
.I2(RIOB33_X105Y131_IOB_X1Y132_I),
.I3(RIOB33_X105Y133_IOB_X1Y133_I),
.I4(RIOB33_X105Y131_IOB_X1Y131_I),
.I5(1'b1),
.O5(CLBLL_L_X2Y121_SLICE_X1Y121_AO5),
.O6(CLBLL_L_X2Y121_SLICE_X1Y121_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h004400f4004400f4)
  ) CLBLL_L_X2Y122_SLICE_X0Y122_DLUT (
.I0(CLBLL_L_X2Y121_SLICE_X0Y121_BO6),
.I1(LIOB33_X0Y69_IOB_X0Y70_I),
.I2(CLBLL_L_X2Y117_SLICE_X0Y117_CQ),
.I3(CLBLM_R_X3Y124_SLICE_X2Y124_AO5),
.I4(CLBLL_L_X2Y120_SLICE_X1Y120_AO6),
.I5(1'b1),
.O5(CLBLL_L_X2Y122_SLICE_X0Y122_DO5),
.O6(CLBLL_L_X2Y122_SLICE_X0Y122_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffffffffffcfe)
  ) CLBLL_L_X2Y122_SLICE_X0Y122_CLUT (
.I0(RIOB33_X105Y113_IOB_X1Y114_I),
.I1(CLBLL_L_X2Y121_SLICE_X0Y121_CO6),
.I2(CLBLL_L_X2Y122_SLICE_X1Y122_BO6),
.I3(CLBLL_L_X2Y122_SLICE_X0Y122_AO5),
.I4(CLBLL_L_X2Y122_SLICE_X0Y122_DO6),
.I5(CLBLL_L_X4Y122_SLICE_X5Y122_BO6),
.O5(CLBLL_L_X2Y122_SLICE_X0Y122_CO5),
.O6(CLBLL_L_X2Y122_SLICE_X0Y122_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffffffffffffe)
  ) CLBLL_L_X2Y122_SLICE_X0Y122_BLUT (
.I0(CLBLL_L_X2Y122_SLICE_X0Y122_DO6),
.I1(CLBLL_L_X2Y122_SLICE_X1Y122_BO6),
.I2(CLBLL_L_X2Y123_SLICE_X0Y123_AO6),
.I3(CLBLL_L_X4Y122_SLICE_X5Y122_BO6),
.I4(CLBLM_R_X5Y122_SLICE_X6Y122_CO6),
.I5(CLBLL_L_X2Y121_SLICE_X0Y121_CO6),
.O5(CLBLL_L_X2Y122_SLICE_X0Y122_BO5),
.O6(CLBLL_L_X2Y122_SLICE_X0Y122_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfff7fffffffdffff)
  ) CLBLL_L_X2Y122_SLICE_X0Y122_ALUT (
.I0(RIOB33_X105Y133_IOB_X1Y133_I),
.I1(RIOB33_X105Y131_IOB_X1Y131_I),
.I2(RIOB33_X105Y133_IOB_X1Y134_I),
.I3(CLBLM_R_X3Y124_SLICE_X2Y124_AO6),
.I4(RIOB33_X105Y131_IOB_X1Y132_I),
.I5(1'b1),
.O5(CLBLL_L_X2Y122_SLICE_X0Y122_AO5),
.O6(CLBLL_L_X2Y122_SLICE_X0Y122_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hff33ff33ff33ff33)
  ) CLBLL_L_X2Y122_SLICE_X1Y122_DLUT (
.I0(1'b1),
.I1(RIOB33_X105Y133_IOB_X1Y133_I),
.I2(1'b1),
.I3(RIOB33_X105Y133_IOB_X1Y134_I),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y122_SLICE_X1Y122_DO5),
.O6(CLBLL_L_X2Y122_SLICE_X1Y122_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0033000000f300f0)
  ) CLBLL_L_X2Y122_SLICE_X1Y122_CLUT (
.I0(1'b1),
.I1(CLBLL_L_X2Y121_SLICE_X1Y121_BO5),
.I2(LIOB33_X0Y63_IOB_X0Y63_I),
.I3(CLBLM_R_X3Y124_SLICE_X2Y124_AO5),
.I4(CLBLM_R_X3Y116_SLICE_X3Y116_CQ),
.I5(CLBLL_L_X2Y121_SLICE_X1Y121_BO6),
.O5(CLBLL_L_X2Y122_SLICE_X1Y122_CO5),
.O6(CLBLL_L_X2Y122_SLICE_X1Y122_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h1155005511110000)
  ) CLBLL_L_X2Y122_SLICE_X1Y122_BLUT (
.I0(CLBLM_R_X3Y124_SLICE_X2Y124_AO5),
.I1(CLBLL_L_X2Y121_SLICE_X1Y121_BO5),
.I2(1'b1),
.I3(CLBLL_L_X2Y121_SLICE_X1Y121_BO6),
.I4(CLBLM_R_X5Y122_SLICE_X7Y122_DQ),
.I5(LIOB33_X0Y59_IOB_X0Y59_I),
.O5(CLBLL_L_X2Y122_SLICE_X1Y122_BO5),
.O6(CLBLL_L_X2Y122_SLICE_X1Y122_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000050400040)
  ) CLBLL_L_X2Y122_SLICE_X1Y122_ALUT (
.I0(CLBLL_L_X2Y122_SLICE_X1Y122_DO6),
.I1(LIOB33_X0Y71_IOB_X0Y71_I),
.I2(RIOB33_X105Y131_IOB_X1Y132_I),
.I3(RIOB33_X105Y131_IOB_X1Y131_I),
.I4(LIOB33_X0Y61_IOB_X0Y61_I),
.I5(CLBLM_R_X3Y124_SLICE_X2Y124_AO5),
.O5(CLBLL_L_X2Y122_SLICE_X1Y122_AO5),
.O6(CLBLL_L_X2Y122_SLICE_X1Y122_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y123_SLICE_X0Y123_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y123_SLICE_X0Y123_DO5),
.O6(CLBLL_L_X2Y123_SLICE_X0Y123_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y123_SLICE_X0Y123_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y123_SLICE_X0Y123_CO5),
.O6(CLBLL_L_X2Y123_SLICE_X0Y123_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y123_SLICE_X0Y123_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y123_SLICE_X0Y123_BO5),
.O6(CLBLL_L_X2Y123_SLICE_X0Y123_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000002000000000)
  ) CLBLL_L_X2Y123_SLICE_X0Y123_ALUT (
.I0(RIOB33_X105Y113_IOB_X1Y114_I),
.I1(CLBLM_R_X3Y124_SLICE_X2Y124_AO6),
.I2(RIOB33_X105Y133_IOB_X1Y133_I),
.I3(RIOB33_X105Y133_IOB_X1Y134_I),
.I4(RIOB33_X105Y131_IOB_X1Y131_I),
.I5(RIOB33_X105Y131_IOB_X1Y132_I),
.O5(CLBLL_L_X2Y123_SLICE_X0Y123_AO5),
.O6(CLBLL_L_X2Y123_SLICE_X0Y123_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y123_SLICE_X1Y123_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y123_SLICE_X1Y123_DO5),
.O6(CLBLL_L_X2Y123_SLICE_X1Y123_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y123_SLICE_X1Y123_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y123_SLICE_X1Y123_CO5),
.O6(CLBLL_L_X2Y123_SLICE_X1Y123_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y123_SLICE_X1Y123_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y123_SLICE_X1Y123_BO5),
.O6(CLBLL_L_X2Y123_SLICE_X1Y123_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y123_SLICE_X1Y123_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y123_SLICE_X1Y123_AO5),
.O6(CLBLL_L_X2Y123_SLICE_X1Y123_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y110_SLICE_X4Y110_A5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y110_SLICE_X4Y110_BO6),
.Q(CLBLL_L_X4Y110_SLICE_X4Y110_A5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y110_SLICE_X4Y110_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y110_SLICE_X4Y110_AO6),
.Q(CLBLL_L_X4Y110_SLICE_X4Y110_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y110_SLICE_X4Y110_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y110_SLICE_X4Y110_CO6),
.Q(CLBLL_L_X4Y110_SLICE_X4Y110_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y110_SLICE_X4Y110_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y110_SLICE_X4Y110_DO6),
.Q(CLBLL_L_X4Y110_SLICE_X4Y110_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffc3330eeec2220)
  ) CLBLL_L_X4Y110_SLICE_X4Y110_DLUT (
.I0(CLBLM_R_X3Y118_SLICE_X2Y118_AQ),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(CLBLL_L_X4Y110_SLICE_X4Y110_DQ),
.I3(CLBLM_R_X5Y112_SLICE_X7Y112_AO6),
.I4(CLBLM_R_X3Y111_SLICE_X3Y111_BQ),
.I5(RIOB33_X105Y117_IOB_X1Y118_I),
.O5(CLBLL_L_X4Y110_SLICE_X4Y110_DO5),
.O6(CLBLL_L_X4Y110_SLICE_X4Y110_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hcccccccc05055050)
  ) CLBLL_L_X4Y110_SLICE_X4Y110_CLUT (
.I0(RIOB33_X105Y105_IOB_X1Y105_I),
.I1(CLBLL_L_X4Y110_SLICE_X4Y110_AQ),
.I2(CLBLM_L_X10Y116_SLICE_X12Y116_CQ),
.I3(1'b1),
.I4(CLBLL_L_X4Y110_SLICE_X4Y110_BO5),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLL_L_X4Y110_SLICE_X4Y110_CO5),
.O6(CLBLL_L_X4Y110_SLICE_X4Y110_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf3e2c0c0ffaa0000)
  ) CLBLL_L_X4Y110_SLICE_X4Y110_BLUT (
.I0(CLBLM_L_X8Y120_SLICE_X11Y120_CQ),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(CLBLM_R_X5Y121_SLICE_X6Y121_B5Q),
.I3(CLBLL_L_X4Y110_SLICE_X4Y110_DQ),
.I4(RIOB33_X105Y121_IOB_X1Y121_I),
.I5(1'b1),
.O5(CLBLL_L_X4Y110_SLICE_X4Y110_BO5),
.O6(CLBLL_L_X4Y110_SLICE_X4Y110_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaaaaaac0f0c0f0)
  ) CLBLL_L_X4Y110_SLICE_X4Y110_ALUT (
.I0(CLBLM_R_X3Y112_SLICE_X3Y112_C5Q),
.I1(CLBLM_R_X3Y118_SLICE_X2Y118_AQ),
.I2(CLBLL_L_X4Y110_SLICE_X4Y110_AQ),
.I3(RIOB33_X105Y117_IOB_X1Y118_I),
.I4(1'b1),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLL_L_X4Y110_SLICE_X4Y110_AO5),
.O6(CLBLL_L_X4Y110_SLICE_X4Y110_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y110_SLICE_X5Y110_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y110_SLICE_X5Y110_AO6),
.Q(CLBLL_L_X4Y110_SLICE_X5Y110_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y110_SLICE_X5Y110_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y110_SLICE_X5Y110_BO6),
.Q(CLBLL_L_X4Y110_SLICE_X5Y110_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000001100000011)
  ) CLBLL_L_X4Y110_SLICE_X5Y110_DLUT (
.I0(CLBLM_R_X5Y109_SLICE_X6Y109_BQ),
.I1(CLBLM_R_X3Y110_SLICE_X3Y110_BQ),
.I2(1'b1),
.I3(CLBLM_R_X5Y109_SLICE_X6Y109_AQ),
.I4(CLBLL_L_X4Y110_SLICE_X4Y110_AQ),
.I5(1'b1),
.O5(CLBLL_L_X4Y110_SLICE_X5Y110_DO5),
.O6(CLBLL_L_X4Y110_SLICE_X5Y110_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h00005050ff000c0c)
  ) CLBLL_L_X4Y110_SLICE_X5Y110_CLUT (
.I0(CLBLM_L_X8Y118_SLICE_X10Y118_DQ),
.I1(CLBLM_R_X5Y114_SLICE_X6Y114_BQ),
.I2(RIOB33_X105Y105_IOB_X1Y105_I),
.I3(CLBLM_R_X3Y110_SLICE_X3Y110_BQ),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(1'b1),
.O5(CLBLL_L_X4Y110_SLICE_X5Y110_CO5),
.O6(CLBLL_L_X4Y110_SLICE_X5Y110_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hff540054ff540054)
  ) CLBLL_L_X4Y110_SLICE_X5Y110_BLUT (
.I0(CLBLM_R_X5Y111_SLICE_X7Y111_DO6),
.I1(CLBLL_L_X4Y110_SLICE_X5Y110_BQ),
.I2(CLBLM_R_X5Y114_SLICE_X6Y114_DQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLL_L_X4Y113_SLICE_X5Y113_AQ),
.I5(1'b1),
.O5(CLBLL_L_X4Y110_SLICE_X5Y110_BO5),
.O6(CLBLL_L_X4Y110_SLICE_X5Y110_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h88ff88f888888888)
  ) CLBLL_L_X4Y110_SLICE_X5Y110_ALUT (
.I0(CLBLM_R_X3Y111_SLICE_X2Y111_AQ),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(CLBLL_L_X4Y110_SLICE_X5Y110_AQ),
.I3(CLBLM_L_X10Y111_SLICE_X13Y111_BO6),
.I4(CLBLM_R_X7Y110_SLICE_X8Y110_DO5),
.I5(CLBLL_L_X4Y110_SLICE_X5Y110_CO6),
.O5(CLBLL_L_X4Y110_SLICE_X5Y110_AO5),
.O6(CLBLL_L_X4Y110_SLICE_X5Y110_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y111_SLICE_X4Y111_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y111_SLICE_X4Y111_AO6),
.Q(CLBLL_L_X4Y111_SLICE_X4Y111_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y111_SLICE_X4Y111_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y111_SLICE_X4Y111_BO6),
.Q(CLBLL_L_X4Y111_SLICE_X4Y111_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y111_SLICE_X4Y111_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y111_SLICE_X4Y111_CO6),
.Q(CLBLL_L_X4Y111_SLICE_X4Y111_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y111_SLICE_X4Y111_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y111_SLICE_X4Y111_DO6),
.Q(CLBLL_L_X4Y111_SLICE_X4Y111_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'haa00aa00aaf0aaf0)
  ) CLBLL_L_X4Y111_SLICE_X4Y111_DLUT (
.I0(CLBLL_L_X4Y112_SLICE_X5Y112_AQ),
.I1(1'b1),
.I2(CLBLL_L_X4Y111_SLICE_X4Y111_DQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(1'b1),
.I5(RIOB33_X105Y105_IOB_X1Y105_I),
.O5(CLBLL_L_X4Y111_SLICE_X4Y111_DO5),
.O6(CLBLL_L_X4Y111_SLICE_X4Y111_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hc0c0c0c0d1e2d1e2)
  ) CLBLL_L_X4Y111_SLICE_X4Y111_CLUT (
.I0(CLBLL_L_X4Y112_SLICE_X5Y112_AQ),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(CLBLM_R_X7Y121_SLICE_X9Y121_AQ),
.I3(CLBLM_R_X5Y112_SLICE_X7Y112_CO6),
.I4(1'b1),
.I5(RIOB33_X105Y105_IOB_X1Y105_I),
.O5(CLBLL_L_X4Y111_SLICE_X4Y111_CO5),
.O6(CLBLL_L_X4Y111_SLICE_X4Y111_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hffaaff88aaaa8888)
  ) CLBLL_L_X4Y111_SLICE_X4Y111_BLUT (
.I0(CLBLM_R_X5Y115_SLICE_X6Y115_CO6),
.I1(CLBLL_L_X4Y111_SLICE_X4Y111_BQ),
.I2(1'b1),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLM_R_X5Y111_SLICE_X6Y111_BQ),
.I5(CLBLM_R_X7Y109_SLICE_X8Y109_BQ),
.O5(CLBLL_L_X4Y111_SLICE_X4Y111_BO5),
.O6(CLBLL_L_X4Y111_SLICE_X4Y111_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'haa03aa00f0f00000)
  ) CLBLL_L_X4Y111_SLICE_X4Y111_ALUT (
.I0(CLBLL_L_X2Y113_SLICE_X1Y113_BQ),
.I1(CLBLL_L_X4Y111_SLICE_X5Y111_DO6),
.I2(RIOB33_X105Y117_IOB_X1Y118_I),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLM_R_X3Y118_SLICE_X2Y118_AQ),
.I5(1'b1),
.O5(CLBLL_L_X4Y111_SLICE_X4Y111_AO5),
.O6(CLBLL_L_X4Y111_SLICE_X4Y111_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y111_SLICE_X5Y111_A5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y110_SLICE_X5Y110_CO5),
.Q(CLBLL_L_X4Y111_SLICE_X5Y111_A5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y111_SLICE_X5Y111_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y111_SLICE_X5Y111_AO6),
.Q(CLBLL_L_X4Y111_SLICE_X5Y111_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y111_SLICE_X5Y111_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y111_SLICE_X5Y111_BO6),
.Q(CLBLL_L_X4Y111_SLICE_X5Y111_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0055005500550005)
  ) CLBLL_L_X4Y111_SLICE_X5Y111_DLUT (
.I0(CLBLL_L_X4Y111_SLICE_X4Y111_AQ),
.I1(1'b1),
.I2(CLBLL_L_X4Y120_SLICE_X4Y120_BO6),
.I3(CLBLM_R_X5Y116_SLICE_X7Y116_CQ),
.I4(CLBLM_R_X7Y109_SLICE_X8Y109_AQ),
.I5(RIOB33_X105Y105_IOB_X1Y105_I),
.O5(CLBLL_L_X4Y111_SLICE_X5Y111_DO5),
.O6(CLBLL_L_X4Y111_SLICE_X5Y111_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0040000000000000)
  ) CLBLL_L_X4Y111_SLICE_X5Y111_CLUT (
.I0(CLBLL_L_X4Y114_SLICE_X5Y114_DO6),
.I1(CLBLM_R_X5Y111_SLICE_X6Y111_CQ),
.I2(CLBLM_R_X7Y113_SLICE_X8Y113_AQ),
.I3(CLBLL_L_X4Y114_SLICE_X5Y114_BO6),
.I4(CLBLM_R_X3Y115_SLICE_X3Y115_DQ),
.I5(CLBLL_L_X4Y115_SLICE_X4Y115_BQ),
.O5(CLBLL_L_X4Y111_SLICE_X5Y111_CO5),
.O6(CLBLL_L_X4Y111_SLICE_X5Y111_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hff300030ffc000c0)
  ) CLBLL_L_X4Y111_SLICE_X5Y111_BLUT (
.I0(1'b1),
.I1(CLBLM_R_X5Y110_SLICE_X6Y110_BO6),
.I2(RIOB33_X105Y105_IOB_X1Y105_I),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLM_R_X7Y120_SLICE_X8Y120_DQ),
.I5(CLBLL_L_X4Y112_SLICE_X5Y112_DO6),
.O5(CLBLL_L_X4Y111_SLICE_X5Y111_BO5),
.O6(CLBLL_L_X4Y111_SLICE_X5Y111_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hcc00ccf0cc00ccf0)
  ) CLBLL_L_X4Y111_SLICE_X5Y111_ALUT (
.I0(1'b1),
.I1(CLBLL_L_X4Y111_SLICE_X5Y111_BQ),
.I2(CLBLL_L_X4Y111_SLICE_X5Y111_AQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(RIOB33_X105Y105_IOB_X1Y105_I),
.I5(1'b1),
.O5(CLBLL_L_X4Y111_SLICE_X5Y111_AO5),
.O6(CLBLL_L_X4Y111_SLICE_X5Y111_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y112_SLICE_X4Y112_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y112_SLICE_X4Y112_AO6),
.Q(CLBLL_L_X4Y112_SLICE_X4Y112_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y112_SLICE_X4Y112_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y112_SLICE_X4Y112_BO6),
.Q(CLBLL_L_X4Y112_SLICE_X4Y112_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h00000000ff00ff00)
  ) CLBLL_L_X4Y112_SLICE_X4Y112_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(CLBLM_R_X7Y120_SLICE_X9Y120_CQ),
.I4(1'b1),
.I5(CLBLM_R_X5Y114_SLICE_X7Y114_AQ),
.O5(CLBLL_L_X4Y112_SLICE_X4Y112_DO5),
.O6(CLBLL_L_X4Y112_SLICE_X4Y112_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hc000c00000000000)
  ) CLBLL_L_X4Y112_SLICE_X4Y112_CLUT (
.I0(1'b1),
.I1(CLBLL_L_X4Y111_SLICE_X4Y111_CQ),
.I2(CLBLM_R_X7Y122_SLICE_X9Y122_BQ),
.I3(CLBLL_L_X4Y111_SLICE_X5Y111_A5Q),
.I4(1'b1),
.I5(CLBLL_L_X4Y111_SLICE_X5Y111_BQ),
.O5(CLBLL_L_X4Y112_SLICE_X4Y112_CO5),
.O6(CLBLL_L_X4Y112_SLICE_X4Y112_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hcccccffc00000330)
  ) CLBLL_L_X4Y112_SLICE_X4Y112_BLUT (
.I0(1'b1),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(CLBLM_R_X5Y112_SLICE_X6Y112_BO6),
.I3(CLBLL_L_X4Y113_SLICE_X5Y113_CQ),
.I4(RIOB33_X105Y105_IOB_X1Y105_I),
.I5(CLBLM_R_X3Y115_SLICE_X2Y115_CQ),
.O5(CLBLL_L_X4Y112_SLICE_X4Y112_BO5),
.O6(CLBLL_L_X4Y112_SLICE_X4Y112_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'haaffaafcaa00aa30)
  ) CLBLL_L_X4Y112_SLICE_X4Y112_ALUT (
.I0(CLBLM_R_X5Y114_SLICE_X6Y114_AQ),
.I1(RIOB33_X105Y117_IOB_X1Y118_I),
.I2(CLBLL_L_X4Y112_SLICE_X4Y112_AQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLM_R_X3Y118_SLICE_X2Y118_AQ),
.I5(CLBLM_R_X3Y115_SLICE_X2Y115_CQ),
.O5(CLBLL_L_X4Y112_SLICE_X4Y112_AO5),
.O6(CLBLL_L_X4Y112_SLICE_X4Y112_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y112_SLICE_X5Y112_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y112_SLICE_X5Y112_AO6),
.Q(CLBLL_L_X4Y112_SLICE_X5Y112_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0ff0f00ff00f0ff0)
  ) CLBLL_L_X4Y112_SLICE_X5Y112_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(CLBLM_L_X8Y120_SLICE_X10Y120_BQ),
.I3(CLBLM_L_X10Y116_SLICE_X13Y116_AQ),
.I4(CLBLM_R_X7Y122_SLICE_X9Y122_BQ),
.I5(CLBLL_L_X4Y111_SLICE_X5Y111_BQ),
.O5(CLBLL_L_X4Y112_SLICE_X5Y112_DO5),
.O6(CLBLL_L_X4Y112_SLICE_X5Y112_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hddffffffffffffff)
  ) CLBLL_L_X4Y112_SLICE_X5Y112_CLUT (
.I0(CLBLL_L_X2Y113_SLICE_X1Y113_BQ),
.I1(CLBLM_R_X5Y114_SLICE_X6Y114_BQ),
.I2(1'b1),
.I3(CLBLM_R_X5Y111_SLICE_X6Y111_BQ),
.I4(CLBLL_L_X4Y113_SLICE_X4Y113_BQ),
.I5(CLBLM_R_X7Y117_SLICE_X8Y117_CQ),
.O5(CLBLL_L_X4Y112_SLICE_X5Y112_CO5),
.O6(CLBLL_L_X4Y112_SLICE_X5Y112_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000500)
  ) CLBLL_L_X4Y112_SLICE_X5Y112_BLUT (
.I0(CLBLM_L_X10Y116_SLICE_X13Y116_AQ),
.I1(1'b1),
.I2(CLBLM_R_X3Y112_SLICE_X3Y112_BQ),
.I3(CLBLL_L_X4Y112_SLICE_X4Y112_CO6),
.I4(CLBLL_L_X4Y114_SLICE_X5Y114_CO6),
.I5(CLBLL_L_X4Y112_SLICE_X5Y112_CO6),
.O5(CLBLL_L_X4Y112_SLICE_X5Y112_BO5),
.O6(CLBLL_L_X4Y112_SLICE_X5Y112_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hccde0012ccde0012)
  ) CLBLL_L_X4Y112_SLICE_X5Y112_ALUT (
.I0(CLBLM_R_X5Y114_SLICE_X7Y114_DO6),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(CLBLM_R_X5Y111_SLICE_X6Y111_BQ),
.I3(RIOB33_X105Y105_IOB_X1Y105_I),
.I4(CLBLL_L_X4Y112_SLICE_X4Y112_AQ),
.I5(1'b1),
.O5(CLBLL_L_X4Y112_SLICE_X5Y112_AO5),
.O6(CLBLL_L_X4Y112_SLICE_X5Y112_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y113_SLICE_X4Y113_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y113_SLICE_X4Y113_AO6),
.Q(CLBLL_L_X4Y113_SLICE_X4Y113_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y113_SLICE_X4Y113_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y113_SLICE_X4Y113_BO6),
.Q(CLBLL_L_X4Y113_SLICE_X4Y113_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hacaca3acacacacac)
  ) CLBLL_L_X4Y113_SLICE_X4Y113_DLUT (
.I0(CLBLM_L_X8Y120_SLICE_X11Y120_CQ),
.I1(CLBLL_L_X4Y111_SLICE_X4Y111_DQ),
.I2(RIOB33_X105Y121_IOB_X1Y121_I),
.I3(CLBLL_L_X4Y112_SLICE_X4Y112_DO6),
.I4(CLBLL_L_X4Y121_SLICE_X4Y121_AQ),
.I5(CLBLL_L_X4Y114_SLICE_X4Y114_BQ),
.O5(CLBLL_L_X4Y113_SLICE_X4Y113_DO5),
.O6(CLBLL_L_X4Y113_SLICE_X4Y113_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0080000000000000)
  ) CLBLL_L_X4Y113_SLICE_X4Y113_CLUT (
.I0(CLBLM_R_X3Y111_SLICE_X3Y111_BQ),
.I1(CLBLL_L_X4Y118_SLICE_X5Y118_AQ),
.I2(RIOB33_X105Y117_IOB_X1Y118_I),
.I3(CLBLM_R_X3Y118_SLICE_X2Y118_AQ),
.I4(CLBLM_R_X3Y112_SLICE_X3Y112_AQ),
.I5(CLBLM_R_X5Y116_SLICE_X6Y116_BQ),
.O5(CLBLL_L_X4Y113_SLICE_X4Y113_CO5),
.O6(CLBLL_L_X4Y113_SLICE_X4Y113_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hc0c0c0c0c5cac5ca)
  ) CLBLL_L_X4Y113_SLICE_X4Y113_BLUT (
.I0(CLBLL_L_X4Y113_SLICE_X4Y113_DO6),
.I1(CLBLM_R_X5Y115_SLICE_X6Y115_BQ),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLL_L_X4Y111_SLICE_X5Y111_BQ),
.I4(1'b1),
.I5(RIOB33_X105Y105_IOB_X1Y105_I),
.O5(CLBLL_L_X4Y113_SLICE_X4Y113_BO5),
.O6(CLBLL_L_X4Y113_SLICE_X4Y113_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hab01ab01ba10ba10)
  ) CLBLL_L_X4Y113_SLICE_X4Y113_ALUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_R_X5Y110_SLICE_X7Y110_BQ),
.I2(CLBLL_L_X4Y113_SLICE_X4Y113_AQ),
.I3(CLBLM_R_X11Y113_SLICE_X15Y113_AQ),
.I4(1'b1),
.I5(CLBLL_L_X4Y113_SLICE_X4Y113_CO6),
.O5(CLBLL_L_X4Y113_SLICE_X4Y113_AO5),
.O6(CLBLL_L_X4Y113_SLICE_X4Y113_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y113_SLICE_X5Y113_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y113_SLICE_X5Y113_AO6),
.Q(CLBLL_L_X4Y113_SLICE_X5Y113_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y113_SLICE_X5Y113_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y113_SLICE_X5Y113_BO6),
.Q(CLBLL_L_X4Y113_SLICE_X5Y113_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y113_SLICE_X5Y113_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y113_SLICE_X5Y113_CO6),
.Q(CLBLL_L_X4Y113_SLICE_X5Y113_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hfc00fc00ff00aa00)
  ) CLBLL_L_X4Y113_SLICE_X5Y113_DLUT (
.I0(CLBLM_R_X5Y113_SLICE_X6Y113_AQ),
.I1(CLBLM_L_X8Y115_SLICE_X11Y115_C5Q),
.I2(CLBLM_R_X3Y113_SLICE_X2Y113_AQ),
.I3(RIOB33_X105Y121_IOB_X1Y121_I),
.I4(CLBLM_R_X3Y116_SLICE_X3Y116_BQ),
.I5(1'b1),
.O5(CLBLL_L_X4Y113_SLICE_X5Y113_DO5),
.O6(CLBLL_L_X4Y113_SLICE_X5Y113_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f00033f0f03300)
  ) CLBLL_L_X4Y113_SLICE_X5Y113_CLUT (
.I0(1'b1),
.I1(RIOB33_X105Y105_IOB_X1Y105_I),
.I2(CLBLM_R_X3Y117_SLICE_X3Y117_BQ),
.I3(CLBLM_R_X5Y114_SLICE_X6Y114_CQ),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(CLBLL_L_X4Y113_SLICE_X5Y113_DO5),
.O5(CLBLL_L_X4Y113_SLICE_X5Y113_CO5),
.O6(CLBLL_L_X4Y113_SLICE_X5Y113_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hffeeffccaaaa0000)
  ) CLBLL_L_X4Y113_SLICE_X5Y113_BLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLL_L_X4Y113_SLICE_X5Y113_BQ),
.I2(1'b1),
.I3(CLBLL_L_X4Y113_SLICE_X4Y113_BQ),
.I4(CLBLM_R_X11Y114_SLICE_X14Y114_D5Q),
.I5(CLBLM_R_X5Y115_SLICE_X6Y115_CO6),
.O5(CLBLL_L_X4Y113_SLICE_X5Y113_BO5),
.O6(CLBLL_L_X4Y113_SLICE_X5Y113_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hb8b8b8b8bbb8bbb8)
  ) CLBLL_L_X4Y113_SLICE_X5Y113_ALUT (
.I0(CLBLM_R_X5Y117_SLICE_X6Y117_BQ),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(CLBLL_L_X4Y112_SLICE_X5Y112_BO6),
.I3(CLBLL_L_X4Y113_SLICE_X5Y113_AQ),
.I4(1'b1),
.I5(RIOB33_X105Y105_IOB_X1Y105_I),
.O5(CLBLL_L_X4Y113_SLICE_X5Y113_AO5),
.O6(CLBLL_L_X4Y113_SLICE_X5Y113_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y114_SLICE_X4Y114_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y114_SLICE_X4Y114_AO6),
.Q(CLBLL_L_X4Y114_SLICE_X4Y114_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y114_SLICE_X4Y114_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y114_SLICE_X4Y114_BO6),
.Q(CLBLL_L_X4Y114_SLICE_X4Y114_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y114_SLICE_X4Y114_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y114_SLICE_X4Y114_CO6),
.Q(CLBLL_L_X4Y114_SLICE_X4Y114_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0e0a0a3f0f0a0a0)
  ) CLBLL_L_X4Y114_SLICE_X4Y114_DLUT (
.I0(CLBLL_L_X4Y114_SLICE_X5Y114_AQ),
.I1(CLBLM_R_X5Y114_SLICE_X7Y114_AQ),
.I2(RIOB33_X105Y121_IOB_X1Y121_I),
.I3(CLBLM_R_X5Y114_SLICE_X7Y114_BO5),
.I4(CLBLL_L_X4Y116_SLICE_X4Y116_BQ),
.I5(CLBLM_R_X7Y120_SLICE_X9Y120_CQ),
.O5(CLBLL_L_X4Y114_SLICE_X4Y114_DO5),
.O6(CLBLL_L_X4Y114_SLICE_X4Y114_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hffa8fffc00a800fc)
  ) CLBLL_L_X4Y114_SLICE_X4Y114_CLUT (
.I0(CLBLM_L_X10Y113_SLICE_X13Y113_BO6),
.I1(CLBLL_L_X4Y114_SLICE_X4Y114_CQ),
.I2(CLBLL_L_X4Y113_SLICE_X4Y113_AQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLM_R_X7Y119_SLICE_X8Y119_D5Q),
.I5(CLBLL_L_X4Y116_SLICE_X4Y116_BQ),
.O5(CLBLL_L_X4Y114_SLICE_X4Y114_CO5),
.O6(CLBLL_L_X4Y114_SLICE_X4Y114_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hff40ff4000400040)
  ) CLBLL_L_X4Y114_SLICE_X4Y114_BLUT (
.I0(CLBLL_L_X4Y115_SLICE_X4Y115_CQ),
.I1(CLBLL_L_X4Y114_SLICE_X4Y114_BQ),
.I2(RIOB33_X105Y105_IOB_X1Y105_I),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(1'b1),
.I5(CLBLL_L_X4Y113_SLICE_X5Y113_CQ),
.O5(CLBLL_L_X4Y114_SLICE_X4Y114_BO5),
.O6(CLBLL_L_X4Y114_SLICE_X4Y114_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffc8c8c8ffc8c8c8)
  ) CLBLL_L_X4Y114_SLICE_X4Y114_ALUT (
.I0(CLBLM_R_X3Y115_SLICE_X3Y115_DQ),
.I1(CLBLM_R_X5Y115_SLICE_X6Y115_CO6),
.I2(CLBLL_L_X4Y114_SLICE_X4Y114_AQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLL_L_X4Y111_SLICE_X4Y111_BQ),
.I5(1'b1),
.O5(CLBLL_L_X4Y114_SLICE_X4Y114_AO5),
.O6(CLBLL_L_X4Y114_SLICE_X4Y114_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y114_SLICE_X5Y114_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y114_SLICE_X5Y114_AO6),
.Q(CLBLL_L_X4Y114_SLICE_X5Y114_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffffffefefefe)
  ) CLBLL_L_X4Y114_SLICE_X5Y114_DLUT (
.I0(CLBLL_L_X4Y116_SLICE_X5Y116_DQ),
.I1(CLBLL_L_X4Y113_SLICE_X5Y113_CQ),
.I2(CLBLM_R_X5Y116_SLICE_X6Y116_DQ),
.I3(1'b1),
.I4(1'b1),
.I5(CLBLL_L_X4Y112_SLICE_X4Y112_BQ),
.O5(CLBLL_L_X4Y114_SLICE_X5Y114_DO5),
.O6(CLBLL_L_X4Y114_SLICE_X5Y114_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffffffbfffff)
  ) CLBLL_L_X4Y114_SLICE_X5Y114_CLUT (
.I0(RIOB33_X105Y105_IOB_X1Y105_I),
.I1(CLBLM_R_X7Y119_SLICE_X9Y119_AQ),
.I2(CLBLM_L_X8Y120_SLICE_X10Y120_BQ),
.I3(CLBLM_R_X5Y121_SLICE_X6Y121_AQ),
.I4(CLBLL_L_X4Y114_SLICE_X5Y114_BO5),
.I5(CLBLL_L_X4Y112_SLICE_X5Y112_AQ),
.O5(CLBLL_L_X4Y114_SLICE_X5Y114_CO5),
.O6(CLBLL_L_X4Y114_SLICE_X5Y114_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfefffeff0f000f00)
  ) CLBLL_L_X4Y114_SLICE_X5Y114_BLUT (
.I0(CLBLM_R_X5Y121_SLICE_X6Y121_AQ),
.I1(CLBLM_R_X5Y115_SLICE_X6Y115_BQ),
.I2(RIOB33_X105Y121_IOB_X1Y121_I),
.I3(CLBLM_R_X7Y114_SLICE_X8Y114_BQ),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y114_SLICE_X5Y114_BO5),
.O6(CLBLL_L_X4Y114_SLICE_X5Y114_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hff88ff8800880088)
  ) CLBLL_L_X4Y114_SLICE_X5Y114_ALUT (
.I0(CLBLL_L_X4Y115_SLICE_X5Y115_CQ),
.I1(RIOB33_X105Y105_IOB_X1Y105_I),
.I2(1'b1),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(1'b1),
.I5(CLBLM_R_X3Y114_SLICE_X2Y114_DQ),
.O5(CLBLL_L_X4Y114_SLICE_X5Y114_AO5),
.O6(CLBLL_L_X4Y114_SLICE_X5Y114_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y115_SLICE_X4Y115_C5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y115_SLICE_X4Y115_CO5),
.Q(CLBLL_L_X4Y115_SLICE_X4Y115_C5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y115_SLICE_X4Y115_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y115_SLICE_X4Y115_AO6),
.Q(CLBLL_L_X4Y115_SLICE_X4Y115_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y115_SLICE_X4Y115_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y115_SLICE_X4Y115_BO6),
.Q(CLBLL_L_X4Y115_SLICE_X4Y115_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y115_SLICE_X4Y115_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y115_SLICE_X4Y115_CO6),
.Q(CLBLL_L_X4Y115_SLICE_X4Y115_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y115_SLICE_X4Y115_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y115_SLICE_X4Y115_DO6),
.Q(CLBLL_L_X4Y115_SLICE_X4Y115_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hddccddcc11001100)
  ) CLBLL_L_X4Y115_SLICE_X4Y115_DLUT (
.I0(RIOB33_X105Y105_IOB_X1Y105_I),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(1'b1),
.I3(CLBLM_R_X5Y115_SLICE_X6Y115_BQ),
.I4(1'b1),
.I5(CLBLM_R_X3Y115_SLICE_X3Y115_AQ),
.O5(CLBLL_L_X4Y115_SLICE_X4Y115_DO5),
.O6(CLBLL_L_X4Y115_SLICE_X4Y115_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hfc30fc30ddcc1100)
  ) CLBLL_L_X4Y115_SLICE_X4Y115_CLUT (
.I0(RIOB33_X105Y105_IOB_X1Y105_I),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(CLBLM_R_X5Y117_SLICE_X6Y117_BQ),
.I3(CLBLM_L_X8Y115_SLICE_X10Y115_CQ),
.I4(CLBLM_R_X3Y115_SLICE_X2Y115_AQ),
.I5(1'b1),
.O5(CLBLL_L_X4Y115_SLICE_X4Y115_CO5),
.O6(CLBLL_L_X4Y115_SLICE_X4Y115_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf000f0ccf000f0cc)
  ) CLBLL_L_X4Y115_SLICE_X4Y115_BLUT (
.I0(1'b1),
.I1(CLBLL_L_X4Y115_SLICE_X4Y115_DQ),
.I2(CLBLL_L_X2Y115_SLICE_X1Y115_AQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(RIOB33_X105Y105_IOB_X1Y105_I),
.I5(1'b1),
.O5(CLBLL_L_X4Y115_SLICE_X4Y115_BO5),
.O6(CLBLL_L_X4Y115_SLICE_X4Y115_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hff540054ff540054)
  ) CLBLL_L_X4Y115_SLICE_X4Y115_ALUT (
.I0(CLBLM_R_X5Y115_SLICE_X6Y115_CO5),
.I1(CLBLL_L_X4Y115_SLICE_X4Y115_DQ),
.I2(CLBLL_L_X4Y115_SLICE_X4Y115_AQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLL_L_X4Y111_SLICE_X4Y111_AQ),
.I5(1'b1),
.O5(CLBLL_L_X4Y115_SLICE_X4Y115_AO5),
.O6(CLBLL_L_X4Y115_SLICE_X4Y115_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y115_SLICE_X5Y115_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y115_SLICE_X5Y115_AO6),
.Q(CLBLL_L_X4Y115_SLICE_X5Y115_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y115_SLICE_X5Y115_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y115_SLICE_X5Y115_BO6),
.Q(CLBLL_L_X4Y115_SLICE_X5Y115_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y115_SLICE_X5Y115_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y115_SLICE_X5Y115_CO6),
.Q(CLBLL_L_X4Y115_SLICE_X5Y115_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y115_SLICE_X5Y115_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y115_SLICE_X5Y115_DO6),
.Q(CLBLL_L_X4Y115_SLICE_X5Y115_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'heeea4440fffa5550)
  ) CLBLL_L_X4Y115_SLICE_X5Y115_DLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_L_X10Y113_SLICE_X13Y113_BO6),
.I2(CLBLL_L_X4Y115_SLICE_X5Y115_DQ),
.I3(CLBLM_R_X3Y115_SLICE_X2Y115_BQ),
.I4(CLBLL_L_X4Y111_SLICE_X5Y111_AQ),
.I5(CLBLM_R_X7Y119_SLICE_X8Y119_D5Q),
.O5(CLBLL_L_X4Y115_SLICE_X5Y115_DO5),
.O6(CLBLL_L_X4Y115_SLICE_X5Y115_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'haa00aa00aaccaacc)
  ) CLBLL_L_X4Y115_SLICE_X5Y115_CLUT (
.I0(CLBLM_R_X5Y115_SLICE_X7Y115_AQ),
.I1(CLBLM_R_X7Y118_SLICE_X9Y118_CQ),
.I2(1'b1),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(1'b1),
.I5(RIOB33_X105Y105_IOB_X1Y105_I),
.O5(CLBLL_L_X4Y115_SLICE_X5Y115_CO5),
.O6(CLBLL_L_X4Y115_SLICE_X5Y115_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hcd01cd01ce02ce02)
  ) CLBLL_L_X4Y115_SLICE_X5Y115_BLUT (
.I0(CLBLL_L_X4Y113_SLICE_X5Y113_DO6),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(RIOB33_X105Y105_IOB_X1Y105_I),
.I3(CLBLL_L_X4Y115_SLICE_X4Y115_DQ),
.I4(1'b1),
.I5(CLBLM_R_X5Y116_SLICE_X6Y116_DQ),
.O5(CLBLL_L_X4Y115_SLICE_X5Y115_BO5),
.O6(CLBLL_L_X4Y115_SLICE_X5Y115_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hccccccccfafafa00)
  ) CLBLL_L_X4Y115_SLICE_X5Y115_ALUT (
.I0(CLBLL_L_X4Y113_SLICE_X4Y113_DO6),
.I1(CLBLM_R_X11Y116_SLICE_X14Y116_CQ),
.I2(CLBLL_L_X4Y115_SLICE_X5Y115_AQ),
.I3(RIOB33_X105Y117_IOB_X1Y118_I),
.I4(CLBLM_R_X3Y118_SLICE_X2Y118_AQ),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLL_L_X4Y115_SLICE_X5Y115_AO5),
.O6(CLBLL_L_X4Y115_SLICE_X5Y115_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y116_SLICE_X4Y116_C5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y116_SLICE_X4Y116_CO5),
.Q(CLBLL_L_X4Y116_SLICE_X4Y116_C5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y116_SLICE_X4Y116_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y116_SLICE_X4Y116_AO6),
.Q(CLBLL_L_X4Y116_SLICE_X4Y116_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y116_SLICE_X4Y116_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y116_SLICE_X4Y116_BO6),
.Q(CLBLL_L_X4Y116_SLICE_X4Y116_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y116_SLICE_X4Y116_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y116_SLICE_X4Y116_CO6),
.Q(CLBLL_L_X4Y116_SLICE_X4Y116_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y116_SLICE_X4Y116_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y116_SLICE_X4Y116_DO6),
.Q(CLBLL_L_X4Y116_SLICE_X4Y116_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hccffcc55ccf0cc50)
  ) CLBLL_L_X4Y116_SLICE_X4Y116_DLUT (
.I0(CLBLM_R_X7Y119_SLICE_X8Y119_D5Q),
.I1(CLBLM_R_X7Y115_SLICE_X9Y115_C5Q),
.I2(CLBLL_L_X4Y116_SLICE_X4Y116_DQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLM_L_X10Y113_SLICE_X13Y113_BO6),
.I5(CLBLM_R_X3Y113_SLICE_X2Y113_BQ),
.O5(CLBLL_L_X4Y116_SLICE_X4Y116_DO5),
.O6(CLBLL_L_X4Y116_SLICE_X4Y116_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0aaf0aaccaaccaa)
  ) CLBLL_L_X4Y116_SLICE_X4Y116_CLUT (
.I0(RIOB33_X105Y101_IOB_X1Y102_I),
.I1(CLBLL_L_X4Y116_SLICE_X4Y116_AQ),
.I2(CLBLL_L_X4Y111_SLICE_X4Y111_CQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y116_SLICE_X4Y116_CO5),
.O6(CLBLL_L_X4Y116_SLICE_X4Y116_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf000f000f0ccf0cc)
  ) CLBLL_L_X4Y116_SLICE_X4Y116_BLUT (
.I0(1'b1),
.I1(CLBLL_L_X4Y116_SLICE_X4Y116_BQ),
.I2(CLBLL_L_X4Y119_SLICE_X5Y119_AQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(1'b1),
.I5(RIOB33_X105Y105_IOB_X1Y105_I),
.O5(CLBLL_L_X4Y116_SLICE_X4Y116_BO5),
.O6(CLBLL_L_X4Y116_SLICE_X4Y116_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfc30ee22ee22ee22)
  ) CLBLL_L_X4Y116_SLICE_X4Y116_ALUT (
.I0(CLBLL_L_X4Y113_SLICE_X4Y113_AQ),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(CLBLL_L_X4Y116_SLICE_X4Y116_AQ),
.I3(CLBLL_L_X4Y116_SLICE_X5Y116_A5Q),
.I4(CLBLL_L_X2Y112_SLICE_X1Y112_BQ),
.I5(CLBLM_L_X8Y112_SLICE_X10Y112_CQ),
.O5(CLBLL_L_X4Y116_SLICE_X4Y116_AO5),
.O6(CLBLL_L_X4Y116_SLICE_X4Y116_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y116_SLICE_X5Y116_A5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y116_SLICE_X5Y116_CO6),
.Q(CLBLL_L_X4Y116_SLICE_X5Y116_A5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y116_SLICE_X5Y116_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y116_SLICE_X5Y116_AO6),
.Q(CLBLL_L_X4Y116_SLICE_X5Y116_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y116_SLICE_X5Y116_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y116_SLICE_X5Y116_BO6),
.Q(CLBLL_L_X4Y116_SLICE_X5Y116_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y116_SLICE_X5Y116_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y116_SLICE_X5Y116_DO6),
.Q(CLBLL_L_X4Y116_SLICE_X5Y116_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaaaaaa0c0c0c0c)
  ) CLBLL_L_X4Y116_SLICE_X5Y116_DLUT (
.I0(CLBLL_L_X4Y116_SLICE_X5Y116_AQ),
.I1(CLBLM_R_X5Y111_SLICE_X6Y111_CQ),
.I2(RIOB33_X105Y105_IOB_X1Y105_I),
.I3(1'b1),
.I4(1'b1),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLL_L_X4Y116_SLICE_X5Y116_DO5),
.O6(CLBLL_L_X4Y116_SLICE_X5Y116_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'heeec2220aaa0aaa0)
  ) CLBLL_L_X4Y116_SLICE_X5Y116_CLUT (
.I0(RIOB33_X105Y121_IOB_X1Y121_I),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(CLBLM_R_X11Y116_SLICE_X15Y116_AQ),
.I3(CLBLM_R_X7Y118_SLICE_X9Y118_CQ),
.I4(CLBLM_R_X11Y113_SLICE_X14Y113_BQ),
.I5(1'b1),
.O5(CLBLL_L_X4Y116_SLICE_X5Y116_CO5),
.O6(CLBLL_L_X4Y116_SLICE_X5Y116_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaaaaaacfc0cfc0)
  ) CLBLL_L_X4Y116_SLICE_X5Y116_BLUT (
.I0(CLBLL_L_X4Y110_SLICE_X5Y110_AQ),
.I1(CLBLL_L_X4Y116_SLICE_X5Y116_BQ),
.I2(CLBLM_R_X5Y115_SLICE_X6Y115_CO5),
.I3(CLBLL_L_X4Y116_SLICE_X5Y116_DQ),
.I4(1'b1),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLL_L_X4Y116_SLICE_X5Y116_BO5),
.O6(CLBLL_L_X4Y116_SLICE_X5Y116_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfedc3210fedc3210)
  ) CLBLL_L_X4Y116_SLICE_X5Y116_ALUT (
.I0(CLBLM_R_X5Y115_SLICE_X6Y115_CO5),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(CLBLL_L_X4Y116_SLICE_X5Y116_AQ),
.I3(CLBLM_R_X5Y115_SLICE_X6Y115_BQ),
.I4(CLBLM_R_X5Y115_SLICE_X7Y115_BQ),
.I5(1'b1),
.O5(CLBLL_L_X4Y116_SLICE_X5Y116_AO5),
.O6(CLBLL_L_X4Y116_SLICE_X5Y116_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y117_SLICE_X4Y117_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y117_SLICE_X4Y117_AO6),
.Q(CLBLL_L_X4Y117_SLICE_X4Y117_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y117_SLICE_X4Y117_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y117_SLICE_X4Y117_BO6),
.Q(CLBLL_L_X4Y117_SLICE_X4Y117_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hff0aff0affffff0a)
  ) CLBLL_L_X4Y117_SLICE_X4Y117_DLUT (
.I0(CLBLL_L_X4Y116_SLICE_X5Y116_BQ),
.I1(1'b1),
.I2(CLBLL_L_X4Y120_SLICE_X5Y120_BO6),
.I3(CLBLM_R_X3Y117_SLICE_X2Y117_DO6),
.I4(CLBLL_L_X4Y116_SLICE_X4Y116_DQ),
.I5(CLBLL_L_X2Y121_SLICE_X1Y121_AO6),
.O5(CLBLL_L_X4Y117_SLICE_X4Y117_DO5),
.O6(CLBLL_L_X4Y117_SLICE_X4Y117_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h000033bb000000aa)
  ) CLBLL_L_X4Y117_SLICE_X4Y117_CLUT (
.I0(CLBLL_L_X4Y115_SLICE_X4Y115_AQ),
.I1(CLBLL_L_X2Y121_SLICE_X1Y121_BO5),
.I2(1'b1),
.I3(CLBLL_L_X2Y121_SLICE_X1Y121_BO6),
.I4(CLBLM_R_X3Y122_SLICE_X3Y122_AO6),
.I5(CLBLL_L_X4Y111_SLICE_X4Y111_BQ),
.O5(CLBLL_L_X4Y117_SLICE_X4Y117_CO5),
.O6(CLBLL_L_X4Y117_SLICE_X4Y117_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0fcf0fc00cc00cc)
  ) CLBLL_L_X4Y117_SLICE_X4Y117_BLUT (
.I0(1'b1),
.I1(CLBLL_L_X4Y117_SLICE_X4Y117_BQ),
.I2(CLBLM_L_X10Y112_SLICE_X13Y112_CQ),
.I3(CLBLM_R_X3Y116_SLICE_X2Y116_CO6),
.I4(1'b1),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLL_L_X4Y117_SLICE_X4Y117_BO5),
.O6(CLBLL_L_X4Y117_SLICE_X4Y117_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffcc00ccfff000f0)
  ) CLBLL_L_X4Y117_SLICE_X4Y117_ALUT (
.I0(1'b1),
.I1(CLBLM_R_X5Y114_SLICE_X6Y114_CQ),
.I2(CLBLL_L_X4Y117_SLICE_X4Y117_AQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLL_L_X4Y116_SLICE_X5Y116_BQ),
.I5(CLBLM_R_X5Y115_SLICE_X6Y115_CO5),
.O5(CLBLL_L_X4Y117_SLICE_X4Y117_AO5),
.O6(CLBLL_L_X4Y117_SLICE_X4Y117_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y117_SLICE_X5Y117_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y117_SLICE_X5Y117_AO6),
.Q(CLBLL_L_X4Y117_SLICE_X5Y117_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y117_SLICE_X5Y117_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y117_SLICE_X5Y117_BO6),
.Q(CLBLL_L_X4Y117_SLICE_X5Y117_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y117_SLICE_X5Y117_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y117_SLICE_X5Y117_CO6),
.Q(CLBLL_L_X4Y117_SLICE_X5Y117_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y117_SLICE_X5Y117_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y117_SLICE_X5Y117_DO6),
.Q(CLBLL_L_X4Y117_SLICE_X5Y117_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hcc00cc00dd11ee22)
  ) CLBLL_L_X4Y117_SLICE_X5Y117_DLUT (
.I0(CLBLL_L_X4Y116_SLICE_X5Y116_CO5),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(1'b1),
.I3(CLBLL_L_X4Y115_SLICE_X5Y115_DQ),
.I4(CLBLM_L_X8Y115_SLICE_X10Y115_AQ),
.I5(RIOB33_X105Y105_IOB_X1Y105_I),
.O5(CLBLL_L_X4Y117_SLICE_X5Y117_DO5),
.O6(CLBLL_L_X4Y117_SLICE_X5Y117_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaaf0f0aaaacccc)
  ) CLBLL_L_X4Y117_SLICE_X5Y117_CLUT (
.I0(CLBLM_R_X3Y116_SLICE_X3Y116_BQ),
.I1(CLBLL_L_X4Y117_SLICE_X5Y117_CQ),
.I2(CLBLM_R_X7Y119_SLICE_X9Y119_BQ),
.I3(1'b1),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(CLBLM_R_X11Y121_SLICE_X14Y121_CO6),
.O5(CLBLL_L_X4Y117_SLICE_X5Y117_CO5),
.O6(CLBLL_L_X4Y117_SLICE_X5Y117_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0ff000ff0fc000c)
  ) CLBLL_L_X4Y117_SLICE_X5Y117_BLUT (
.I0(1'b1),
.I1(CLBLL_L_X4Y117_SLICE_X5Y117_BQ),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLM_R_X11Y121_SLICE_X14Y121_CO6),
.I4(CLBLL_L_X4Y117_SLICE_X4Y117_AQ),
.I5(CLBLL_L_X4Y110_SLICE_X4Y110_CQ),
.O5(CLBLL_L_X4Y117_SLICE_X5Y117_BO5),
.O6(CLBLL_L_X4Y117_SLICE_X5Y117_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfedcfcfc32103030)
  ) CLBLL_L_X4Y117_SLICE_X5Y117_ALUT (
.I0(CLBLM_L_X8Y112_SLICE_X10Y112_CQ),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(CLBLM_R_X3Y111_SLICE_X3Y111_BQ),
.I3(CLBLL_L_X4Y117_SLICE_X5Y117_AQ),
.I4(CLBLL_L_X2Y112_SLICE_X1Y112_BQ),
.I5(CLBLM_R_X5Y117_SLICE_X7Y117_BQ),
.O5(CLBLL_L_X4Y117_SLICE_X5Y117_AO5),
.O6(CLBLL_L_X4Y117_SLICE_X5Y117_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y118_SLICE_X4Y118_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y118_SLICE_X4Y118_AO6),
.Q(CLBLL_L_X4Y118_SLICE_X4Y118_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0fafffff0faf0fa)
  ) CLBLL_L_X4Y118_SLICE_X4Y118_DLUT (
.I0(CLBLL_L_X4Y116_SLICE_X4Y116_AQ),
.I1(1'b1),
.I2(CLBLL_L_X4Y118_SLICE_X5Y118_DO6),
.I3(CLBLM_R_X3Y121_SLICE_X2Y121_AO5),
.I4(CLBLM_R_X3Y121_SLICE_X2Y121_AO6),
.I5(CLBLM_R_X5Y118_SLICE_X6Y118_AQ),
.O5(CLBLL_L_X4Y118_SLICE_X4Y118_DO5),
.O6(CLBLL_L_X4Y118_SLICE_X4Y118_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hcfccefeecfccefee)
  ) CLBLL_L_X4Y118_SLICE_X4Y118_CLUT (
.I0(CLBLL_L_X4Y117_SLICE_X5Y117_BQ),
.I1(CLBLM_R_X3Y118_SLICE_X3Y118_BO6),
.I2(CLBLL_L_X4Y121_SLICE_X4Y121_CO6),
.I3(CLBLM_R_X7Y118_SLICE_X9Y118_BQ),
.I4(CLBLL_L_X4Y120_SLICE_X5Y120_BO5),
.I5(1'b1),
.O5(CLBLL_L_X4Y118_SLICE_X4Y118_CO5),
.O6(CLBLL_L_X4Y118_SLICE_X4Y118_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h77f733f355f500f0)
  ) CLBLL_L_X4Y118_SLICE_X4Y118_BLUT (
.I0(CLBLL_L_X2Y119_SLICE_X1Y119_AO5),
.I1(CLBLL_L_X4Y120_SLICE_X5Y120_BO6),
.I2(CLBLM_L_X10Y117_SLICE_X13Y117_CQ),
.I3(CLBLL_L_X2Y121_SLICE_X1Y121_AO6),
.I4(CLBLM_R_X3Y112_SLICE_X2Y112_AQ),
.I5(CLBLM_R_X5Y121_SLICE_X6Y121_BQ),
.O5(CLBLL_L_X4Y118_SLICE_X4Y118_BO5),
.O6(CLBLL_L_X4Y118_SLICE_X4Y118_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h5554005455540054)
  ) CLBLL_L_X4Y118_SLICE_X4Y118_ALUT (
.I0(CLBLM_R_X5Y115_SLICE_X6Y115_CO6),
.I1(CLBLL_L_X4Y112_SLICE_X5Y112_AQ),
.I2(CLBLL_L_X4Y118_SLICE_X4Y118_AQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLM_R_X5Y118_SLICE_X6Y118_AQ),
.I5(1'b1),
.O5(CLBLL_L_X4Y118_SLICE_X4Y118_AO5),
.O6(CLBLL_L_X4Y118_SLICE_X4Y118_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y118_SLICE_X5Y118_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y118_SLICE_X5Y118_AO6),
.Q(CLBLL_L_X4Y118_SLICE_X5Y118_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y118_SLICE_X5Y118_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y118_SLICE_X5Y118_BO6),
.Q(CLBLL_L_X4Y118_SLICE_X5Y118_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y118_SLICE_X5Y118_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y118_SLICE_X5Y118_CO6),
.Q(CLBLL_L_X4Y118_SLICE_X5Y118_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000a0c)
  ) CLBLL_L_X4Y118_SLICE_X5Y118_DLUT (
.I0(CLBLM_L_X8Y118_SLICE_X11Y118_AQ),
.I1(CLBLM_R_X11Y116_SLICE_X14Y116_AQ),
.I2(CLBLL_L_X2Y122_SLICE_X1Y122_DO6),
.I3(RIOB33_X105Y131_IOB_X1Y131_I),
.I4(RIOB33_X105Y131_IOB_X1Y132_I),
.I5(CLBLM_R_X3Y122_SLICE_X3Y122_AO6),
.O5(CLBLL_L_X4Y118_SLICE_X5Y118_DO5),
.O6(CLBLL_L_X4Y118_SLICE_X5Y118_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hff55af05ee44ae04)
  ) CLBLL_L_X4Y118_SLICE_X5Y118_CLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLL_L_X4Y118_SLICE_X5Y118_CQ),
.I2(CLBLM_R_X7Y119_SLICE_X8Y119_D5Q),
.I3(CLBLL_L_X4Y117_SLICE_X5Y117_CQ),
.I4(CLBLM_L_X10Y113_SLICE_X13Y113_BO6),
.I5(CLBLL_L_X4Y118_SLICE_X5Y118_AQ),
.O5(CLBLL_L_X4Y118_SLICE_X5Y118_CO5),
.O6(CLBLL_L_X4Y118_SLICE_X5Y118_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hff00e4e4ff00f0f0)
  ) CLBLL_L_X4Y118_SLICE_X5Y118_BLUT (
.I0(CLBLM_L_X10Y113_SLICE_X13Y113_BO6),
.I1(CLBLL_L_X4Y118_SLICE_X5Y118_BQ),
.I2(CLBLM_R_X3Y111_SLICE_X3Y111_BQ),
.I3(CLBLM_R_X5Y122_SLICE_X6Y122_AQ),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(CLBLM_R_X7Y119_SLICE_X8Y119_D5Q),
.O5(CLBLL_L_X4Y118_SLICE_X5Y118_BO5),
.O6(CLBLL_L_X4Y118_SLICE_X5Y118_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'haaffaaffaaf0aa3c)
  ) CLBLL_L_X4Y118_SLICE_X5Y118_ALUT (
.I0(CLBLM_R_X7Y119_SLICE_X9Y119_BQ),
.I1(RIOB33_X105Y117_IOB_X1Y118_I),
.I2(CLBLL_L_X4Y118_SLICE_X5Y118_AQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLM_R_X3Y118_SLICE_X2Y118_AQ),
.I5(CLBLM_R_X5Y110_SLICE_X7Y110_BQ),
.O5(CLBLL_L_X4Y118_SLICE_X5Y118_AO5),
.O6(CLBLL_L_X4Y118_SLICE_X5Y118_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y119_SLICE_X4Y119_B5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y119_SLICE_X4Y119_BO5),
.Q(CLBLL_L_X4Y119_SLICE_X4Y119_B5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "C5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y119_SLICE_X4Y119_C5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y119_SLICE_X4Y119_CO5),
.Q(CLBLL_L_X4Y119_SLICE_X4Y119_C5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y119_SLICE_X4Y119_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y119_SLICE_X4Y119_AO6),
.Q(CLBLL_L_X4Y119_SLICE_X4Y119_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y119_SLICE_X4Y119_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y119_SLICE_X4Y119_BO6),
.Q(CLBLL_L_X4Y119_SLICE_X4Y119_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y119_SLICE_X4Y119_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y119_SLICE_X4Y119_CO6),
.Q(CLBLL_L_X4Y119_SLICE_X4Y119_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y119_SLICE_X4Y119_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y119_SLICE_X4Y119_DO6),
.Q(CLBLL_L_X4Y119_SLICE_X4Y119_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hfbfbeaea51514040)
  ) CLBLL_L_X4Y119_SLICE_X4Y119_DLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_R_X3Y116_SLICE_X2Y116_DO6),
.I2(CLBLL_L_X4Y119_SLICE_X4Y119_DQ),
.I3(1'b1),
.I4(CLBLL_L_X4Y119_SLICE_X4Y119_B5Q),
.I5(CLBLM_R_X11Y119_SLICE_X15Y119_AQ),
.O5(CLBLL_L_X4Y119_SLICE_X4Y119_DO5),
.O6(CLBLL_L_X4Y119_SLICE_X4Y119_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hf5a0f5a0eeee4444)
  ) CLBLL_L_X4Y119_SLICE_X4Y119_CLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_R_X5Y110_SLICE_X7Y110_BQ),
.I2(CLBLM_R_X3Y119_SLICE_X3Y119_AQ),
.I3(CLBLL_L_X4Y116_SLICE_X5Y116_A5Q),
.I4(CLBLL_L_X2Y117_SLICE_X0Y117_A5Q),
.I5(1'b1),
.O5(CLBLL_L_X4Y119_SLICE_X4Y119_CO5),
.O6(CLBLL_L_X4Y119_SLICE_X4Y119_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f0ff00ccccaaaa)
  ) CLBLL_L_X4Y119_SLICE_X4Y119_BLUT (
.I0(CLBLM_R_X7Y121_SLICE_X9Y121_AQ),
.I1(CLBLL_L_X4Y119_SLICE_X4Y119_BQ),
.I2(CLBLL_L_X2Y116_SLICE_X1Y116_AQ),
.I3(RIOB33_X105Y127_IOB_X1Y127_I),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(1'b1),
.O5(CLBLL_L_X4Y119_SLICE_X4Y119_BO5),
.O6(CLBLL_L_X4Y119_SLICE_X4Y119_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hccccff00ccccf0f0)
  ) CLBLL_L_X4Y119_SLICE_X4Y119_ALUT (
.I0(1'b1),
.I1(CLBLM_R_X5Y120_SLICE_X7Y120_AQ),
.I2(CLBLL_L_X4Y119_SLICE_X4Y119_AQ),
.I3(CLBLL_L_X4Y115_SLICE_X4Y115_BQ),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(CLBLM_R_X5Y115_SLICE_X6Y115_CO5),
.O5(CLBLL_L_X4Y119_SLICE_X4Y119_AO5),
.O6(CLBLL_L_X4Y119_SLICE_X4Y119_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y119_SLICE_X5Y119_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y119_SLICE_X5Y119_AO6),
.Q(CLBLL_L_X4Y119_SLICE_X5Y119_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hffcfffefffccffee)
  ) CLBLL_L_X4Y119_SLICE_X5Y119_DLUT (
.I0(CLBLL_L_X2Y116_SLICE_X1Y116_AQ),
.I1(CLBLM_R_X5Y119_SLICE_X6Y119_DO6),
.I2(CLBLL_L_X4Y120_SLICE_X5Y120_BO5),
.I3(CLBLL_L_X4Y119_SLICE_X5Y119_CO6),
.I4(CLBLM_R_X3Y121_SLICE_X2Y121_AO5),
.I5(CLBLM_L_X8Y116_SLICE_X11Y116_AQ),
.O5(CLBLL_L_X4Y119_SLICE_X5Y119_DO5),
.O6(CLBLL_L_X4Y119_SLICE_X5Y119_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000001000)
  ) CLBLL_L_X4Y119_SLICE_X5Y119_CLUT (
.I0(CLBLM_R_X3Y122_SLICE_X3Y122_AO6),
.I1(RIOB33_X105Y133_IOB_X1Y133_I),
.I2(RIOB33_X105Y131_IOB_X1Y132_I),
.I3(CLBLM_R_X7Y120_SLICE_X8Y120_AQ),
.I4(RIOB33_X105Y133_IOB_X1Y134_I),
.I5(RIOB33_X105Y131_IOB_X1Y131_I),
.O5(CLBLL_L_X4Y119_SLICE_X5Y119_CO5),
.O6(CLBLL_L_X4Y119_SLICE_X5Y119_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h73ff737350ff5050)
  ) CLBLL_L_X4Y119_SLICE_X5Y119_BLUT (
.I0(CLBLL_L_X4Y121_SLICE_X4Y121_DO5),
.I1(CLBLL_L_X4Y120_SLICE_X5Y120_BO6),
.I2(CLBLL_L_X4Y119_SLICE_X5Y119_AQ),
.I3(CLBLL_L_X2Y120_SLICE_X0Y120_AO6),
.I4(CLBLL_L_X4Y116_SLICE_X5Y116_AQ),
.I5(CLBLM_R_X7Y118_SLICE_X8Y118_CQ),
.O5(CLBLL_L_X4Y119_SLICE_X5Y119_BO5),
.O6(CLBLL_L_X4Y119_SLICE_X5Y119_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaafcfcaaaa3030)
  ) CLBLL_L_X4Y119_SLICE_X5Y119_ALUT (
.I0(CLBLM_R_X5Y120_SLICE_X6Y120_A5Q),
.I1(CLBLM_R_X5Y115_SLICE_X6Y115_CO5),
.I2(CLBLL_L_X4Y119_SLICE_X5Y119_AQ),
.I3(1'b1),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(CLBLM_R_X7Y117_SLICE_X8Y117_CQ),
.O5(CLBLL_L_X4Y119_SLICE_X5Y119_AO5),
.O6(CLBLL_L_X4Y119_SLICE_X5Y119_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hf2f2f2f2fff2fff2)
  ) CLBLL_L_X4Y120_SLICE_X4Y120_DLUT (
.I0(RIOB33_X105Y107_IOB_X1Y108_I),
.I1(CLBLL_L_X2Y122_SLICE_X0Y122_AO6),
.I2(CLBLM_R_X3Y120_SLICE_X3Y120_CO6),
.I3(CLBLM_R_X7Y120_SLICE_X8Y120_BQ),
.I4(1'b1),
.I5(CLBLM_R_X3Y122_SLICE_X2Y122_BO5),
.O5(CLBLL_L_X4Y120_SLICE_X4Y120_DO5),
.O6(CLBLL_L_X4Y120_SLICE_X4Y120_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hcecececeffceffce)
  ) CLBLL_L_X4Y120_SLICE_X4Y120_CLUT (
.I0(RIOB33_X105Y107_IOB_X1Y107_I),
.I1(CLBLL_L_X4Y117_SLICE_X4Y117_CO6),
.I2(CLBLL_L_X2Y122_SLICE_X0Y122_AO6),
.I3(CLBLM_R_X7Y118_SLICE_X8Y118_BQ),
.I4(1'b1),
.I5(CLBLM_R_X3Y122_SLICE_X2Y122_BO5),
.O5(CLBLL_L_X4Y120_SLICE_X4Y120_CO5),
.O6(CLBLL_L_X4Y120_SLICE_X4Y120_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffffffffffffe)
  ) CLBLL_L_X4Y120_SLICE_X4Y120_BLUT (
.I0(CLBLL_L_X4Y118_SLICE_X4Y118_DO6),
.I1(CLBLL_L_X2Y121_SLICE_X1Y121_CO6),
.I2(CLBLM_R_X3Y123_SLICE_X3Y123_DO6),
.I3(CLBLL_L_X4Y120_SLICE_X4Y120_DO6),
.I4(CLBLL_L_X4Y119_SLICE_X5Y119_BO6),
.I5(CLBLL_L_X4Y121_SLICE_X5Y121_CO5),
.O5(CLBLL_L_X4Y120_SLICE_X4Y120_BO5),
.O6(CLBLL_L_X4Y120_SLICE_X4Y120_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffffffffffffe)
  ) CLBLL_L_X4Y120_SLICE_X4Y120_ALUT (
.I0(CLBLM_R_X5Y121_SLICE_X6Y121_DO6),
.I1(CLBLL_L_X4Y118_SLICE_X4Y118_BO6),
.I2(CLBLM_R_X3Y123_SLICE_X2Y123_BO6),
.I3(CLBLL_L_X2Y121_SLICE_X1Y121_CO6),
.I4(CLBLM_R_X5Y120_SLICE_X6Y120_CO6),
.I5(CLBLL_L_X4Y120_SLICE_X4Y120_CO6),
.O5(CLBLL_L_X4Y120_SLICE_X4Y120_AO5),
.O6(CLBLL_L_X4Y120_SLICE_X4Y120_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffffffffffdfc)
  ) CLBLL_L_X4Y120_SLICE_X5Y120_DLUT (
.I0(CLBLL_L_X4Y122_SLICE_X5Y122_CO6),
.I1(CLBLM_R_X5Y120_SLICE_X6Y120_DO6),
.I2(CLBLL_L_X4Y119_SLICE_X5Y119_DO6),
.I3(CLBLL_L_X2Y121_SLICE_X1Y121_DO6),
.I4(CLBLL_L_X4Y122_SLICE_X4Y122_CO6),
.I5(CLBLL_L_X4Y117_SLICE_X4Y117_DO6),
.O5(CLBLL_L_X4Y120_SLICE_X5Y120_DO5),
.O6(CLBLL_L_X4Y120_SLICE_X5Y120_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h3f330f00bfbbafaa)
  ) CLBLL_L_X4Y120_SLICE_X5Y120_CLUT (
.I0(CLBLM_R_X5Y120_SLICE_X6Y120_BQ),
.I1(CLBLM_R_X3Y122_SLICE_X2Y122_BO5),
.I2(CLBLL_L_X4Y121_SLICE_X4Y121_DO5),
.I3(CLBLM_R_X7Y117_SLICE_X9Y117_DQ),
.I4(CLBLL_L_X4Y121_SLICE_X5Y121_AQ),
.I5(CLBLL_L_X4Y120_SLICE_X5Y120_BO6),
.O5(CLBLL_L_X4Y120_SLICE_X5Y120_CO5),
.O6(CLBLL_L_X4Y120_SLICE_X5Y120_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffdfffffffeffff)
  ) CLBLL_L_X4Y120_SLICE_X5Y120_BLUT (
.I0(RIOB33_X105Y131_IOB_X1Y132_I),
.I1(CLBLM_R_X3Y122_SLICE_X3Y122_AO6),
.I2(RIOB33_X105Y133_IOB_X1Y134_I),
.I3(RIOB33_X105Y131_IOB_X1Y131_I),
.I4(RIOB33_X105Y133_IOB_X1Y133_I),
.I5(1'b1),
.O5(CLBLL_L_X4Y120_SLICE_X5Y120_BO5),
.O6(CLBLL_L_X4Y120_SLICE_X5Y120_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfcfcfcfc69699696)
  ) CLBLL_L_X4Y120_SLICE_X5Y120_ALUT (
.I0(CLBLL_L_X2Y120_SLICE_X0Y120_CO6),
.I1(CLBLL_L_X4Y120_SLICE_X4Y120_BO6),
.I2(CLBLL_L_X4Y120_SLICE_X4Y120_AO6),
.I3(1'b1),
.I4(CLBLL_L_X2Y119_SLICE_X0Y119_BO6),
.I5(1'b1),
.O5(CLBLL_L_X4Y120_SLICE_X5Y120_AO5),
.O6(CLBLL_L_X4Y120_SLICE_X5Y120_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y121_SLICE_X4Y121_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y121_SLICE_X4Y121_AO6),
.Q(CLBLL_L_X4Y121_SLICE_X4Y121_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y121_SLICE_X4Y121_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y121_SLICE_X4Y121_BO6),
.Q(CLBLL_L_X4Y121_SLICE_X4Y121_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h00002022fffeffff)
  ) CLBLL_L_X4Y121_SLICE_X4Y121_DLUT (
.I0(RIOB33_X105Y133_IOB_X1Y133_I),
.I1(CLBLM_R_X3Y122_SLICE_X3Y122_AO6),
.I2(RIOB33_X105Y131_IOB_X1Y131_I),
.I3(RIOB33_X105Y131_IOB_X1Y132_I),
.I4(RIOB33_X105Y133_IOB_X1Y134_I),
.I5(1'b1),
.O5(CLBLL_L_X4Y121_SLICE_X4Y121_DO5),
.O6(CLBLL_L_X4Y121_SLICE_X4Y121_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffefffffffffdd)
  ) CLBLL_L_X4Y121_SLICE_X4Y121_CLUT (
.I0(RIOB33_X105Y133_IOB_X1Y133_I),
.I1(CLBLM_R_X3Y122_SLICE_X3Y122_AO6),
.I2(RIOB33_X105Y131_IOB_X1Y131_I),
.I3(RIOB33_X105Y131_IOB_X1Y132_I),
.I4(RIOB33_X105Y133_IOB_X1Y134_I),
.I5(1'b1),
.O5(CLBLL_L_X4Y121_SLICE_X4Y121_CO5),
.O6(CLBLL_L_X4Y121_SLICE_X4Y121_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'he2c0c0c0c0c0c0c0)
  ) CLBLL_L_X4Y121_SLICE_X4Y121_BLUT (
.I0(CLBLM_R_X5Y122_SLICE_X6Y122_AQ),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(CLBLM_L_X8Y115_SLICE_X11Y115_BQ),
.I3(CLBLM_R_X7Y120_SLICE_X8Y120_CQ),
.I4(CLBLM_R_X5Y121_SLICE_X6Y121_B5Q),
.I5(CLBLL_L_X4Y117_SLICE_X4Y117_BQ),
.O5(CLBLL_L_X4Y121_SLICE_X4Y121_BO5),
.O6(CLBLL_L_X4Y121_SLICE_X4Y121_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hcc00cc00fc30cc00)
  ) CLBLL_L_X4Y121_SLICE_X4Y121_ALUT (
.I0(1'b1),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(CLBLL_L_X4Y121_SLICE_X4Y121_AQ),
.I3(CLBLM_R_X5Y124_SLICE_X6Y124_BQ),
.I4(RIOB33_X105Y105_IOB_X1Y105_I),
.I5(CLBLL_L_X4Y115_SLICE_X4Y115_CQ),
.O5(CLBLL_L_X4Y121_SLICE_X4Y121_AO5),
.O6(CLBLL_L_X4Y121_SLICE_X4Y121_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y121_SLICE_X5Y121_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y121_SLICE_X5Y121_AO6),
.Q(CLBLL_L_X4Y121_SLICE_X5Y121_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000001000000000)
  ) CLBLL_L_X4Y121_SLICE_X5Y121_DLUT (
.I0(RIOB33_X105Y133_IOB_X1Y133_I),
.I1(RIOB33_X105Y131_IOB_X1Y132_I),
.I2(RIOB33_X105Y133_IOB_X1Y134_I),
.I3(CLBLM_R_X3Y122_SLICE_X3Y122_AO6),
.I4(RIOB33_X105Y131_IOB_X1Y131_I),
.I5(CLBLL_L_X4Y113_SLICE_X5Y113_BQ),
.O5(CLBLL_L_X4Y121_SLICE_X5Y121_DO5),
.O6(CLBLL_L_X4Y121_SLICE_X5Y121_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff00ff30302222)
  ) CLBLL_L_X4Y121_SLICE_X5Y121_CLUT (
.I0(CLBLM_L_X8Y121_SLICE_X10Y121_BQ),
.I1(CLBLL_L_X4Y122_SLICE_X4Y122_AO5),
.I2(CLBLL_L_X4Y113_SLICE_X5Y113_AQ),
.I3(RIOB33_X105Y135_IOB_X1Y136_I),
.I4(RIOB33_X105Y131_IOB_X1Y131_I),
.I5(1'b1),
.O5(CLBLL_L_X4Y121_SLICE_X5Y121_CO5),
.O6(CLBLL_L_X4Y121_SLICE_X5Y121_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hafafafaf23dcdc23)
  ) CLBLL_L_X4Y121_SLICE_X5Y121_BLUT (
.I0(RIOB33_X105Y129_IOB_X1Y129_I),
.I1(CLBLM_R_X7Y127_SLICE_X8Y127_AQ),
.I2(RIOB33_X105Y137_IOB_X1Y137_I),
.I3(CLBLL_L_X4Y120_SLICE_X5Y120_AO5),
.I4(CLBLM_R_X5Y120_SLICE_X7Y120_DO5),
.I5(1'b1),
.O5(CLBLL_L_X4Y121_SLICE_X5Y121_BO5),
.O6(CLBLL_L_X4Y121_SLICE_X5Y121_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffcc00ccfff000f0)
  ) CLBLL_L_X4Y121_SLICE_X5Y121_ALUT (
.I0(1'b1),
.I1(CLBLM_R_X7Y122_SLICE_X9Y122_BQ),
.I2(CLBLL_L_X4Y121_SLICE_X5Y121_AQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLL_L_X4Y119_SLICE_X4Y119_AQ),
.I5(CLBLM_R_X5Y115_SLICE_X6Y115_CO5),
.O5(CLBLL_L_X4Y121_SLICE_X5Y121_AO5),
.O6(CLBLL_L_X4Y121_SLICE_X5Y121_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000454500004040)
  ) CLBLL_L_X4Y122_SLICE_X4Y122_DLUT (
.I0(CLBLL_L_X4Y122_SLICE_X4Y122_AO6),
.I1(CLBLM_R_X5Y122_SLICE_X7Y122_CQ),
.I2(RIOB33_X105Y131_IOB_X1Y131_I),
.I3(1'b1),
.I4(CLBLM_R_X3Y124_SLICE_X2Y124_AO5),
.I5(CLBLM_R_X5Y122_SLICE_X6Y122_BQ),
.O5(CLBLL_L_X4Y122_SLICE_X4Y122_DO5),
.O6(CLBLL_L_X4Y122_SLICE_X4Y122_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffffff0affce)
  ) CLBLL_L_X4Y122_SLICE_X4Y122_CLUT (
.I0(RIOB33_X105Y109_IOB_X1Y110_I),
.I1(CLBLL_L_X4Y123_SLICE_X4Y123_CQ),
.I2(CLBLL_L_X2Y122_SLICE_X0Y122_AO6),
.I3(CLBLL_L_X4Y121_SLICE_X5Y121_DO6),
.I4(CLBLM_R_X3Y123_SLICE_X3Y123_BO5),
.I5(CLBLL_L_X4Y122_SLICE_X4Y122_BO6),
.O5(CLBLL_L_X4Y122_SLICE_X4Y122_CO5),
.O6(CLBLL_L_X4Y122_SLICE_X4Y122_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf000f222f0f0f2f2)
  ) CLBLL_L_X4Y122_SLICE_X4Y122_BLUT (
.I0(LIOB33_X0Y65_IOB_X0Y65_I),
.I1(CLBLL_L_X2Y121_SLICE_X1Y121_BO6),
.I2(CLBLM_L_X8Y120_SLICE_X10Y120_D5Q),
.I3(RIOB33_X105Y129_IOB_X1Y129_I),
.I4(CLBLM_R_X3Y124_SLICE_X2Y124_AO5),
.I5(RIOB33_X105Y137_IOB_X1Y137_I),
.O5(CLBLL_L_X4Y122_SLICE_X4Y122_BO5),
.O6(CLBLL_L_X4Y122_SLICE_X4Y122_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfcfcfffffffffff3)
  ) CLBLL_L_X4Y122_SLICE_X4Y122_ALUT (
.I0(1'b1),
.I1(RIOB33_X105Y131_IOB_X1Y132_I),
.I2(RIOB33_X105Y133_IOB_X1Y133_I),
.I3(CLBLM_R_X3Y122_SLICE_X3Y122_AO6),
.I4(RIOB33_X105Y133_IOB_X1Y134_I),
.I5(1'b1),
.O5(CLBLL_L_X4Y122_SLICE_X4Y122_AO5),
.O6(CLBLL_L_X4Y122_SLICE_X4Y122_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000004000000000)
  ) CLBLL_L_X4Y122_SLICE_X5Y122_DLUT (
.I0(RIOB33_X105Y129_IOB_X1Y130_I),
.I1(RIOB33_X105Y135_IOB_X1Y135_I),
.I2(CLBLL_L_X4Y123_SLICE_X5Y123_AO5),
.I3(RIOB33_X105Y131_IOB_X1Y131_I),
.I4(CLBLL_L_X4Y121_SLICE_X5Y121_BO6),
.I5(RIOB33_X105Y135_IOB_X1Y136_I),
.O5(CLBLL_L_X4Y122_SLICE_X5Y122_DO5),
.O6(CLBLL_L_X4Y122_SLICE_X5Y122_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h000000c000001111)
  ) CLBLL_L_X4Y122_SLICE_X5Y122_CLUT (
.I0(CLBLM_R_X3Y124_SLICE_X2Y124_BO6),
.I1(RIOB33_X105Y135_IOB_X1Y135_I),
.I2(CLBLL_L_X4Y123_SLICE_X5Y123_AO5),
.I3(RIOB33_X105Y131_IOB_X1Y131_I),
.I4(CLBLM_R_X3Y122_SLICE_X3Y122_AO5),
.I5(RIOB33_X105Y135_IOB_X1Y136_I),
.O5(CLBLL_L_X4Y122_SLICE_X5Y122_CO5),
.O6(CLBLL_L_X4Y122_SLICE_X5Y122_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hc0c0c0c0c0c0e2c0)
  ) CLBLL_L_X4Y122_SLICE_X5Y122_BLUT (
.I0(RIOB33_X105Y135_IOB_X1Y135_I),
.I1(CLBLL_L_X4Y121_SLICE_X5Y121_BO6),
.I2(CLBLM_R_X7Y113_SLICE_X9Y113_AQ),
.I3(CLBLL_L_X4Y123_SLICE_X5Y123_AO5),
.I4(RIOB33_X105Y129_IOB_X1Y130_I),
.I5(CLBLL_L_X4Y121_SLICE_X5Y121_CO6),
.O5(CLBLL_L_X4Y122_SLICE_X5Y122_BO5),
.O6(CLBLL_L_X4Y122_SLICE_X5Y122_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h000000000c001d11)
  ) CLBLL_L_X4Y122_SLICE_X5Y122_ALUT (
.I0(RIOB33_X105Y135_IOB_X1Y135_I),
.I1(RIOB33_X105Y135_IOB_X1Y136_I),
.I2(RIOB33_X105Y131_IOB_X1Y131_I),
.I3(CLBLL_L_X4Y123_SLICE_X5Y123_AO5),
.I4(CLBLM_R_X3Y124_SLICE_X2Y124_BO6),
.I5(CLBLM_R_X3Y122_SLICE_X3Y122_AO5),
.O5(CLBLL_L_X4Y122_SLICE_X5Y122_AO5),
.O6(CLBLL_L_X4Y122_SLICE_X5Y122_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y123_SLICE_X4Y123_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y123_SLICE_X4Y123_AO6),
.Q(CLBLL_L_X4Y123_SLICE_X4Y123_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y123_SLICE_X4Y123_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y123_SLICE_X4Y123_BO6),
.Q(CLBLL_L_X4Y123_SLICE_X4Y123_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y123_SLICE_X4Y123_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y123_SLICE_X4Y123_CO6),
.Q(CLBLL_L_X4Y123_SLICE_X4Y123_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0400000000000000)
  ) CLBLL_L_X4Y123_SLICE_X4Y123_DLUT (
.I0(RIOB33_X105Y131_IOB_X1Y132_I),
.I1(RIOB33_X105Y131_IOB_X1Y131_I),
.I2(CLBLM_R_X3Y124_SLICE_X2Y124_AO5),
.I3(RIOB33_X105Y133_IOB_X1Y134_I),
.I4(CLBLM_R_X5Y122_SLICE_X6Y122_AQ),
.I5(RIOB33_X105Y133_IOB_X1Y133_I),
.O5(CLBLL_L_X4Y123_SLICE_X4Y123_DO5),
.O6(CLBLL_L_X4Y123_SLICE_X4Y123_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h8d8d8d888d8d8d88)
  ) CLBLL_L_X4Y123_SLICE_X4Y123_CLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLL_L_X4Y117_SLICE_X5Y117_DQ),
.I2(CLBLM_R_X3Y116_SLICE_X2Y116_DO6),
.I3(CLBLM_R_X5Y116_SLICE_X6Y116_A5Q),
.I4(CLBLL_L_X4Y123_SLICE_X4Y123_CQ),
.I5(1'b1),
.O5(CLBLL_L_X4Y123_SLICE_X4Y123_CO5),
.O6(CLBLL_L_X4Y123_SLICE_X4Y123_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f00066f0f00000)
  ) CLBLL_L_X4Y123_SLICE_X4Y123_BLUT (
.I0(CLBLM_R_X5Y125_SLICE_X6Y125_BO5),
.I1(CLBLL_L_X4Y123_SLICE_X4Y123_BQ),
.I2(CLBLL_L_X2Y113_SLICE_X1Y113_C5Q),
.I3(CLBLL_L_X4Y119_SLICE_X4Y119_C5Q),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(RIOB33_X105Y105_IOB_X1Y105_I),
.O5(CLBLL_L_X4Y123_SLICE_X4Y123_BO5),
.O6(CLBLL_L_X4Y123_SLICE_X4Y123_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hbe3caa00faf0aa00)
  ) CLBLL_L_X4Y123_SLICE_X4Y123_ALUT (
.I0(CLBLL_L_X4Y123_SLICE_X4Y123_CQ),
.I1(CLBLM_R_X7Y124_SLICE_X8Y124_BQ),
.I2(CLBLL_L_X4Y123_SLICE_X4Y123_AQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLM_R_X7Y124_SLICE_X8Y124_DO5),
.I5(CLBLM_R_X7Y124_SLICE_X8Y124_A5Q),
.O5(CLBLL_L_X4Y123_SLICE_X4Y123_AO5),
.O6(CLBLL_L_X4Y123_SLICE_X4Y123_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X4Y123_SLICE_X5Y123_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y123_SLICE_X5Y123_DO5),
.O6(CLBLL_L_X4Y123_SLICE_X5Y123_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X4Y123_SLICE_X5Y123_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y123_SLICE_X5Y123_CO5),
.O6(CLBLL_L_X4Y123_SLICE_X5Y123_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X4Y123_SLICE_X5Y123_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y123_SLICE_X5Y123_BO5),
.O6(CLBLL_L_X4Y123_SLICE_X5Y123_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffff0ff0000f000)
  ) CLBLL_L_X4Y123_SLICE_X5Y123_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(RIOB33_X105Y131_IOB_X1Y132_I),
.I3(RIOB33_X105Y133_IOB_X1Y133_I),
.I4(RIOB33_X105Y133_IOB_X1Y134_I),
.I5(1'b1),
.O5(CLBLL_L_X4Y123_SLICE_X5Y123_AO5),
.O6(CLBLL_L_X4Y123_SLICE_X5Y123_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X52Y126_SLICE_X78Y126_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X52Y126_SLICE_X78Y126_DO5),
.O6(CLBLL_L_X52Y126_SLICE_X78Y126_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X52Y126_SLICE_X78Y126_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X52Y126_SLICE_X78Y126_CO5),
.O6(CLBLL_L_X52Y126_SLICE_X78Y126_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X52Y126_SLICE_X78Y126_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X52Y126_SLICE_X78Y126_BO5),
.O6(CLBLL_L_X52Y126_SLICE_X78Y126_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h00ff00ff00ff00ff)
  ) CLBLL_L_X52Y126_SLICE_X78Y126_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(RIOB33_X105Y123_IOB_X1Y124_I),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X52Y126_SLICE_X78Y126_AO5),
.O6(CLBLL_L_X52Y126_SLICE_X78Y126_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X52Y126_SLICE_X79Y126_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X52Y126_SLICE_X79Y126_DO5),
.O6(CLBLL_L_X52Y126_SLICE_X79Y126_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X52Y126_SLICE_X79Y126_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X52Y126_SLICE_X79Y126_CO5),
.O6(CLBLL_L_X52Y126_SLICE_X79Y126_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X52Y126_SLICE_X79Y126_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X52Y126_SLICE_X79Y126_BO5),
.O6(CLBLL_L_X52Y126_SLICE_X79Y126_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X52Y126_SLICE_X79Y126_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X52Y126_SLICE_X79Y126_AO5),
.O6(CLBLL_L_X52Y126_SLICE_X79Y126_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y110_SLICE_X10Y110_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y110_SLICE_X10Y110_AO6),
.Q(CLBLM_L_X8Y110_SLICE_X10Y110_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y110_SLICE_X10Y110_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y110_SLICE_X10Y110_BO6),
.Q(CLBLM_L_X8Y110_SLICE_X10Y110_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h5faf5faff5faf5fa)
  ) CLBLM_L_X8Y110_SLICE_X10Y110_DLUT (
.I0(CLBLM_R_X7Y115_SLICE_X9Y115_BQ),
.I1(1'b1),
.I2(CLBLM_L_X8Y116_SLICE_X11Y116_BQ),
.I3(CLBLM_R_X7Y110_SLICE_X9Y110_BQ),
.I4(1'b1),
.I5(CLBLM_L_X10Y116_SLICE_X13Y116_CQ),
.O5(CLBLM_L_X8Y110_SLICE_X10Y110_DO5),
.O6(CLBLM_L_X8Y110_SLICE_X10Y110_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff7dbeffff7dbe)
  ) CLBLM_L_X8Y110_SLICE_X10Y110_CLUT (
.I0(CLBLM_R_X5Y111_SLICE_X6Y111_C5Q),
.I1(CLBLM_L_X10Y118_SLICE_X12Y118_BQ),
.I2(CLBLM_L_X10Y115_SLICE_X12Y115_DQ),
.I3(CLBLM_L_X10Y110_SLICE_X12Y110_BQ),
.I4(CLBLM_L_X8Y110_SLICE_X10Y110_DO6),
.I5(1'b1),
.O5(CLBLM_L_X8Y110_SLICE_X10Y110_CO5),
.O6(CLBLM_L_X8Y110_SLICE_X10Y110_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff0e0000000e00)
  ) CLBLM_L_X8Y110_SLICE_X10Y110_BLUT (
.I0(CLBLM_L_X10Y111_SLICE_X13Y111_BO6),
.I1(CLBLM_L_X8Y110_SLICE_X10Y110_BQ),
.I2(CLBLM_L_X8Y118_SLICE_X10Y118_DQ),
.I3(RIOB33_X105Y105_IOB_X1Y105_I),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(CLBLM_L_X10Y115_SLICE_X12Y115_AQ),
.O5(CLBLM_L_X8Y110_SLICE_X10Y110_BO5),
.O6(CLBLM_L_X8Y110_SLICE_X10Y110_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hff54ff5400540054)
  ) CLBLM_L_X8Y110_SLICE_X10Y110_ALUT (
.I0(CLBLM_R_X5Y111_SLICE_X7Y111_DO6),
.I1(CLBLL_L_X4Y110_SLICE_X5Y110_BQ),
.I2(CLBLM_L_X8Y110_SLICE_X10Y110_AQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(1'b1),
.I5(CLBLL_L_X4Y110_SLICE_X4Y110_A5Q),
.O5(CLBLM_L_X8Y110_SLICE_X10Y110_AO5),
.O6(CLBLM_L_X8Y110_SLICE_X10Y110_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X8Y110_SLICE_X11Y110_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X8Y110_SLICE_X11Y110_DO5),
.O6(CLBLM_L_X8Y110_SLICE_X11Y110_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X8Y110_SLICE_X11Y110_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X8Y110_SLICE_X11Y110_CO5),
.O6(CLBLM_L_X8Y110_SLICE_X11Y110_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X8Y110_SLICE_X11Y110_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X8Y110_SLICE_X11Y110_BO5),
.O6(CLBLM_L_X8Y110_SLICE_X11Y110_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X8Y110_SLICE_X11Y110_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X8Y110_SLICE_X11Y110_AO5),
.O6(CLBLM_L_X8Y110_SLICE_X11Y110_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y111_SLICE_X10Y111_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y111_SLICE_X10Y111_AO6),
.Q(CLBLM_L_X8Y111_SLICE_X10Y111_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h7d7d7d7dbebebebe)
  ) CLBLM_L_X8Y111_SLICE_X10Y111_DLUT (
.I0(CLBLM_R_X7Y110_SLICE_X8Y110_AQ),
.I1(CLBLM_L_X8Y118_SLICE_X10Y118_CQ),
.I2(CLBLM_R_X11Y114_SLICE_X14Y114_BQ),
.I3(1'b1),
.I4(1'b1),
.I5(CLBLM_R_X11Y113_SLICE_X15Y113_BQ),
.O5(CLBLM_L_X8Y111_SLICE_X10Y111_DO5),
.O6(CLBLM_L_X8Y111_SLICE_X10Y111_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h6699996666999966)
  ) CLBLM_L_X8Y111_SLICE_X10Y111_CLUT (
.I0(CLBLM_R_X7Y110_SLICE_X8Y110_AQ),
.I1(CLBLM_L_X8Y118_SLICE_X10Y118_CQ),
.I2(1'b1),
.I3(CLBLM_R_X5Y114_SLICE_X6Y114_AQ),
.I4(CLBLM_L_X8Y117_SLICE_X10Y117_BQ),
.I5(1'b1),
.O5(CLBLM_L_X8Y111_SLICE_X10Y111_CO5),
.O6(CLBLM_L_X8Y111_SLICE_X10Y111_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0d00fff2000df2ff)
  ) CLBLM_L_X8Y111_SLICE_X10Y111_BLUT (
.I0(CLBLM_R_X5Y111_SLICE_X7Y111_CO6),
.I1(CLBLM_R_X7Y111_SLICE_X9Y111_AO5),
.I2(CLBLM_R_X5Y119_SLICE_X7Y119_CO6),
.I3(CLBLM_R_X7Y111_SLICE_X9Y111_BO5),
.I4(CLBLM_R_X5Y111_SLICE_X6Y111_C5Q),
.I5(CLBLM_R_X5Y114_SLICE_X6Y114_DQ),
.O5(CLBLM_L_X8Y111_SLICE_X10Y111_BO5),
.O6(CLBLM_L_X8Y111_SLICE_X10Y111_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hb8bb88bbb8888888)
  ) CLBLM_L_X8Y111_SLICE_X10Y111_ALUT (
.I0(CLBLM_R_X5Y111_SLICE_X7Y111_BQ),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(CLBLM_L_X8Y111_SLICE_X10Y111_AQ),
.I3(CLBLM_L_X10Y113_SLICE_X12Y113_DO6),
.I4(RIOB33_X105Y105_IOB_X1Y105_I),
.I5(CLBLM_R_X11Y113_SLICE_X15Y113_BQ),
.O5(CLBLM_L_X8Y111_SLICE_X10Y111_AO5),
.O6(CLBLM_L_X8Y111_SLICE_X10Y111_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h3b3b3f3f31313030)
  ) CLBLM_L_X8Y111_SLICE_X11Y111_DLUT (
.I0(CLBLM_R_X7Y111_SLICE_X9Y111_AO5),
.I1(CLBLM_L_X10Y127_SLICE_X12Y127_AQ),
.I2(CLBLM_R_X5Y119_SLICE_X7Y119_CO6),
.I3(1'b1),
.I4(CLBLM_R_X5Y111_SLICE_X7Y111_CO6),
.I5(CLBLM_L_X10Y111_SLICE_X12Y111_AO6),
.O5(CLBLM_L_X8Y111_SLICE_X11Y111_DO5),
.O6(CLBLM_L_X8Y111_SLICE_X11Y111_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h02020303f7f7f3f3)
  ) CLBLM_L_X8Y111_SLICE_X11Y111_CLUT (
.I0(CLBLM_R_X7Y111_SLICE_X9Y111_AO5),
.I1(CLBLM_L_X10Y111_SLICE_X13Y111_CO5),
.I2(CLBLM_R_X5Y119_SLICE_X7Y119_CO6),
.I3(1'b1),
.I4(CLBLM_R_X5Y111_SLICE_X7Y111_CO6),
.I5(CLBLM_R_X7Y115_SLICE_X9Y115_BQ),
.O5(CLBLM_L_X8Y111_SLICE_X11Y111_CO5),
.O6(CLBLM_L_X8Y111_SLICE_X11Y111_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hffde00120012ffde)
  ) CLBLM_L_X8Y111_SLICE_X11Y111_BLUT (
.I0(CLBLM_L_X8Y112_SLICE_X11Y112_BO5),
.I1(CLBLL_L_X2Y119_SLICE_X1Y119_BO6),
.I2(CLBLM_R_X7Y111_SLICE_X9Y111_BO6),
.I3(CLBLM_R_X5Y119_SLICE_X7Y119_CO6),
.I4(CLBLM_L_X10Y118_SLICE_X12Y118_BQ),
.I5(CLBLL_L_X4Y119_SLICE_X4Y119_CQ),
.O5(CLBLM_L_X8Y111_SLICE_X11Y111_BO5),
.O6(CLBLM_L_X8Y111_SLICE_X11Y111_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h6996966996696996)
  ) CLBLM_L_X8Y111_SLICE_X11Y111_ALUT (
.I0(CLBLM_L_X8Y111_SLICE_X11Y111_DO6),
.I1(CLBLM_L_X8Y111_SLICE_X10Y111_BO6),
.I2(CLBLM_L_X10Y111_SLICE_X12Y111_DO6),
.I3(CLBLM_L_X8Y111_SLICE_X11Y111_BO6),
.I4(CLBLM_L_X8Y113_SLICE_X11Y113_DO6),
.I5(CLBLM_L_X8Y111_SLICE_X11Y111_CO6),
.O5(CLBLM_L_X8Y111_SLICE_X11Y111_AO5),
.O6(CLBLM_L_X8Y111_SLICE_X11Y111_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y112_SLICE_X10Y112_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y112_SLICE_X10Y112_AO6),
.Q(CLBLM_L_X8Y112_SLICE_X10Y112_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y112_SLICE_X10Y112_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y112_SLICE_X10Y112_BO6),
.Q(CLBLM_L_X8Y112_SLICE_X10Y112_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y112_SLICE_X10Y112_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y112_SLICE_X10Y112_CO6),
.Q(CLBLM_L_X8Y112_SLICE_X10Y112_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y112_SLICE_X10Y112_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y112_SLICE_X10Y112_DO6),
.Q(CLBLM_L_X8Y112_SLICE_X10Y112_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hf505f505f000f000)
  ) CLBLM_L_X8Y112_SLICE_X10Y112_DLUT (
.I0(RIOB33_X105Y105_IOB_X1Y105_I),
.I1(1'b1),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLM_L_X10Y116_SLICE_X13Y116_CQ),
.I4(1'b1),
.I5(CLBLM_R_X7Y109_SLICE_X8Y109_BQ),
.O5(CLBLM_L_X8Y112_SLICE_X10Y112_DO5),
.O6(CLBLM_L_X8Y112_SLICE_X10Y112_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hee44ee44aa00ee44)
  ) CLBLM_L_X8Y112_SLICE_X10Y112_CLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_L_X8Y112_SLICE_X10Y112_CQ),
.I2(1'b1),
.I3(CLBLM_L_X8Y112_SLICE_X10Y112_BQ),
.I4(RIOB33_X105Y117_IOB_X1Y118_I),
.I5(CLBLM_R_X3Y118_SLICE_X2Y118_AQ),
.O5(CLBLM_L_X8Y112_SLICE_X10Y112_CO5),
.O6(CLBLM_L_X8Y112_SLICE_X10Y112_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'haac0aaffaac0aa00)
  ) CLBLM_L_X8Y112_SLICE_X10Y112_BLUT (
.I0(CLBLM_R_X7Y112_SLICE_X8Y112_CQ),
.I1(CLBLM_L_X8Y112_SLICE_X10Y112_BQ),
.I2(RIOB33_X105Y105_IOB_X1Y105_I),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLM_L_X10Y113_SLICE_X12Y113_DO6),
.I5(CLBLM_R_X11Y113_SLICE_X15Y113_AQ),
.O5(CLBLM_L_X8Y112_SLICE_X10Y112_BO5),
.O6(CLBLM_L_X8Y112_SLICE_X10Y112_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfc30cc00ee22ee22)
  ) CLBLM_L_X8Y112_SLICE_X10Y112_ALUT (
.I0(CLBLM_R_X11Y114_SLICE_X14Y114_BQ),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(CLBLM_L_X8Y112_SLICE_X10Y112_AQ),
.I3(CLBLM_R_X7Y112_SLICE_X9Y112_BQ),
.I4(RIOB33_X105Y105_IOB_X1Y105_I),
.I5(CLBLM_L_X10Y113_SLICE_X12Y113_DO6),
.O5(CLBLM_L_X8Y112_SLICE_X10Y112_AO5),
.O6(CLBLM_L_X8Y112_SLICE_X10Y112_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y112_SLICE_X11Y112_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y112_SLICE_X11Y112_AO6),
.Q(CLBLM_L_X8Y112_SLICE_X11Y112_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h00000000c33c3cc3)
  ) CLBLM_L_X8Y112_SLICE_X11Y112_DLUT (
.I0(1'b1),
.I1(CLBLM_L_X12Y115_SLICE_X16Y115_CQ),
.I2(CLBLM_L_X10Y120_SLICE_X12Y120_BQ),
.I3(CLBLM_L_X8Y111_SLICE_X10Y111_CO6),
.I4(CLBLM_L_X8Y113_SLICE_X10Y113_BO6),
.I5(CLBLM_L_X8Y112_SLICE_X11Y112_AQ),
.O5(CLBLM_L_X8Y112_SLICE_X11Y112_DO5),
.O6(CLBLM_L_X8Y112_SLICE_X11Y112_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h001d002e000c003f)
  ) CLBLM_L_X8Y112_SLICE_X11Y112_CLUT (
.I0(CLBLM_L_X10Y111_SLICE_X12Y111_AO5),
.I1(CLBLM_R_X5Y111_SLICE_X7Y111_DO6),
.I2(CLBLM_L_X8Y115_SLICE_X11Y115_CQ),
.I3(CLBLM_R_X7Y112_SLICE_X9Y112_BQ),
.I4(CLBLM_L_X8Y110_SLICE_X10Y110_AQ),
.I5(CLBLM_L_X8Y112_SLICE_X11Y112_BO6),
.O5(CLBLM_L_X8Y112_SLICE_X11Y112_CO5),
.O6(CLBLM_L_X8Y112_SLICE_X11Y112_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h5050505033333363)
  ) CLBLM_L_X8Y112_SLICE_X11Y112_BLUT (
.I0(CLBLL_L_X4Y110_SLICE_X5Y110_AQ),
.I1(CLBLL_L_X4Y110_SLICE_X5Y110_BQ),
.I2(CLBLM_L_X8Y110_SLICE_X10Y110_BQ),
.I3(CLBLM_L_X10Y112_SLICE_X13Y112_CQ),
.I4(CLBLM_R_X7Y110_SLICE_X8Y110_CQ),
.I5(1'b1),
.O5(CLBLM_L_X8Y112_SLICE_X11Y112_BO5),
.O6(CLBLM_L_X8Y112_SLICE_X11Y112_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfff5ffc400f500c4)
  ) CLBLM_L_X8Y112_SLICE_X11Y112_ALUT (
.I0(CLBLM_L_X8Y112_SLICE_X11Y112_DO6),
.I1(CLBLM_R_X3Y118_SLICE_X2Y118_AQ),
.I2(CLBLM_R_X7Y111_SLICE_X9Y111_AO6),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(RIOB33_X105Y117_IOB_X1Y118_I),
.I5(CLBLM_L_X8Y117_SLICE_X11Y117_CQ),
.O5(CLBLM_L_X8Y112_SLICE_X11Y112_AO5),
.O6(CLBLM_L_X8Y112_SLICE_X11Y112_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h66ff66ffff66ff66)
  ) CLBLM_L_X8Y113_SLICE_X10Y113_DLUT (
.I0(CLBLM_L_X8Y112_SLICE_X10Y112_BQ),
.I1(CLBLM_L_X8Y117_SLICE_X10Y117_BQ),
.I2(1'b1),
.I3(CLBLM_R_X11Y113_SLICE_X14Y113_AQ),
.I4(1'b1),
.I5(CLBLM_R_X5Y118_SLICE_X6Y118_BQ),
.O5(CLBLM_L_X8Y113_SLICE_X10Y113_DO5),
.O6(CLBLM_L_X8Y113_SLICE_X10Y113_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h77bb77bbddeeddee)
  ) CLBLM_L_X8Y113_SLICE_X10Y113_CLUT (
.I0(CLBLM_L_X8Y114_SLICE_X10Y114_AQ),
.I1(CLBLM_R_X7Y112_SLICE_X9Y112_AQ),
.I2(1'b1),
.I3(CLBLM_L_X8Y112_SLICE_X10Y112_AQ),
.I4(1'b1),
.I5(CLBLM_R_X11Y113_SLICE_X15Y113_AQ),
.O5(CLBLM_L_X8Y113_SLICE_X10Y113_CO5),
.O6(CLBLM_L_X8Y113_SLICE_X10Y113_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h3cc3c33c3cc3c33c)
  ) CLBLM_L_X8Y113_SLICE_X10Y113_BLUT (
.I0(1'b1),
.I1(CLBLL_L_X4Y112_SLICE_X4Y112_AQ),
.I2(CLBLM_R_X7Y112_SLICE_X9Y112_AQ),
.I3(CLBLM_R_X5Y118_SLICE_X6Y118_BQ),
.I4(CLBLM_L_X8Y114_SLICE_X10Y114_AQ),
.I5(1'b1),
.O5(CLBLM_L_X8Y113_SLICE_X10Y113_BO5),
.O6(CLBLM_L_X8Y113_SLICE_X10Y113_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffffbbeebbee)
  ) CLBLM_L_X8Y113_SLICE_X10Y113_ALUT (
.I0(CLBLM_L_X8Y113_SLICE_X10Y113_DO6),
.I1(CLBLL_L_X4Y112_SLICE_X4Y112_AQ),
.I2(1'b1),
.I3(CLBLM_L_X8Y113_SLICE_X11Y113_BQ),
.I4(1'b1),
.I5(CLBLM_L_X8Y113_SLICE_X10Y113_CO6),
.O5(CLBLM_L_X8Y113_SLICE_X10Y113_AO5),
.O6(CLBLM_L_X8Y113_SLICE_X10Y113_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y113_SLICE_X11Y113_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y113_SLICE_X11Y113_AO6),
.Q(CLBLM_L_X8Y113_SLICE_X11Y113_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y113_SLICE_X11Y113_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y113_SLICE_X11Y113_BO6),
.Q(CLBLM_L_X8Y113_SLICE_X11Y113_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y113_SLICE_X11Y113_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y113_SLICE_X11Y113_CO6),
.Q(CLBLM_L_X8Y113_SLICE_X11Y113_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hf00ff00ff00f6666)
  ) CLBLM_L_X8Y113_SLICE_X11Y113_DLUT (
.I0(CLBLM_L_X10Y113_SLICE_X12Y113_AO6),
.I1(CLBLM_L_X10Y114_SLICE_X12Y114_AO6),
.I2(CLBLM_R_X7Y115_SLICE_X9Y115_B5Q),
.I3(CLBLM_L_X8Y115_SLICE_X11Y115_CQ),
.I4(CLBLM_R_X5Y119_SLICE_X7Y119_CO6),
.I5(CLBLL_L_X2Y119_SLICE_X1Y119_BO6),
.O5(CLBLM_L_X8Y113_SLICE_X11Y113_DO5),
.O6(CLBLM_L_X8Y113_SLICE_X11Y113_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffffcd00ef00)
  ) CLBLM_L_X8Y113_SLICE_X11Y113_CLUT (
.I0(CLBLM_R_X7Y111_SLICE_X9Y111_AO6),
.I1(CLBLM_L_X8Y113_SLICE_X11Y113_CQ),
.I2(CLBLM_L_X8Y111_SLICE_X11Y111_AO6),
.I3(CLBLM_R_X11Y123_SLICE_X14Y123_CO6),
.I4(CLBLM_L_X10Y113_SLICE_X12Y113_CO6),
.I5(CLBLM_R_X5Y121_SLICE_X6Y121_CO5),
.O5(CLBLM_L_X8Y113_SLICE_X11Y113_CO5),
.O6(CLBLM_L_X8Y113_SLICE_X11Y113_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'heefaaafa44500050)
  ) CLBLM_L_X8Y113_SLICE_X11Y113_BLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_L_X8Y113_SLICE_X11Y113_BQ),
.I2(CLBLM_L_X8Y111_SLICE_X10Y111_AQ),
.I3(CLBLM_L_X10Y113_SLICE_X12Y113_DO6),
.I4(RIOB33_X105Y105_IOB_X1Y105_I),
.I5(CLBLL_L_X4Y115_SLICE_X4Y115_BQ),
.O5(CLBLM_L_X8Y113_SLICE_X11Y113_BO5),
.O6(CLBLM_L_X8Y113_SLICE_X11Y113_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfaee5044aaee0044)
  ) CLBLM_L_X8Y113_SLICE_X11Y113_ALUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_L_X8Y112_SLICE_X10Y112_BQ),
.I2(CLBLM_L_X8Y113_SLICE_X11Y113_AQ),
.I3(CLBLM_L_X10Y113_SLICE_X12Y113_DO6),
.I4(CLBLL_L_X4Y121_SLICE_X4Y121_AQ),
.I5(RIOB33_X105Y105_IOB_X1Y105_I),
.O5(CLBLM_L_X8Y113_SLICE_X11Y113_AO5),
.O6(CLBLM_L_X8Y113_SLICE_X11Y113_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y114_SLICE_X10Y114_B5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y114_SLICE_X10Y114_BO5),
.Q(CLBLM_L_X8Y114_SLICE_X10Y114_B5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "C5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y114_SLICE_X10Y114_C5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y114_SLICE_X10Y114_CO5),
.Q(CLBLM_L_X8Y114_SLICE_X10Y114_C5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y114_SLICE_X10Y114_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y114_SLICE_X10Y114_AO6),
.Q(CLBLM_L_X8Y114_SLICE_X10Y114_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y114_SLICE_X10Y114_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y114_SLICE_X10Y114_BO6),
.Q(CLBLM_L_X8Y114_SLICE_X10Y114_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y114_SLICE_X10Y114_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y114_SLICE_X10Y114_CO6),
.Q(CLBLM_L_X8Y114_SLICE_X10Y114_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y114_SLICE_X10Y114_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y114_SLICE_X10Y114_DO6),
.Q(CLBLM_L_X8Y114_SLICE_X10Y114_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hff00ff00fcfca8a8)
  ) CLBLM_L_X8Y114_SLICE_X10Y114_DLUT (
.I0(CLBLM_R_X3Y118_SLICE_X2Y118_AQ),
.I1(CLBLM_R_X5Y115_SLICE_X7Y115_CO6),
.I2(CLBLM_L_X8Y114_SLICE_X10Y114_DQ),
.I3(CLBLL_L_X4Y116_SLICE_X5Y116_DQ),
.I4(RIOB33_X105Y117_IOB_X1Y118_I),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLM_L_X8Y114_SLICE_X10Y114_DO5),
.O6(CLBLM_L_X8Y114_SLICE_X10Y114_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hff00aaaacccc0f00)
  ) CLBLM_L_X8Y114_SLICE_X10Y114_CLUT (
.I0(RIOB33_X105Y103_IOB_X1Y103_I),
.I1(CLBLM_R_X5Y113_SLICE_X6Y113_BQ),
.I2(RIOB33_X105Y105_IOB_X1Y105_I),
.I3(CLBLM_L_X8Y114_SLICE_X11Y114_CQ),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(1'b1),
.O5(CLBLM_L_X8Y114_SLICE_X10Y114_CO5),
.O6(CLBLM_L_X8Y114_SLICE_X10Y114_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'ha0a0acacc0c0cfc0)
  ) CLBLM_L_X8Y114_SLICE_X10Y114_BLUT (
.I0(CLBLM_R_X11Y115_SLICE_X14Y115_CQ),
.I1(CLBLM_L_X8Y112_SLICE_X10Y112_DQ),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLM_R_X3Y116_SLICE_X3Y116_BQ),
.I4(RIOB33_X105Y105_IOB_X1Y105_I),
.I5(1'b1),
.O5(CLBLM_L_X8Y114_SLICE_X10Y114_BO5),
.O6(CLBLM_L_X8Y114_SLICE_X10Y114_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hccaaccaaccaaccf0)
  ) CLBLM_L_X8Y114_SLICE_X10Y114_ALUT (
.I0(CLBLM_L_X8Y117_SLICE_X10Y117_CQ),
.I1(CLBLM_L_X8Y114_SLICE_X10Y114_DQ),
.I2(CLBLM_L_X8Y114_SLICE_X10Y114_AQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLM_R_X3Y118_SLICE_X2Y118_AQ),
.I5(RIOB33_X105Y117_IOB_X1Y118_I),
.O5(CLBLM_L_X8Y114_SLICE_X10Y114_AO5),
.O6(CLBLM_L_X8Y114_SLICE_X10Y114_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y114_SLICE_X11Y114_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y114_SLICE_X11Y114_AO6),
.Q(CLBLM_L_X8Y114_SLICE_X11Y114_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y114_SLICE_X11Y114_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y114_SLICE_X11Y114_BO6),
.Q(CLBLM_L_X8Y114_SLICE_X11Y114_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y114_SLICE_X11Y114_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y114_SLICE_X11Y114_CO6),
.Q(CLBLM_L_X8Y114_SLICE_X11Y114_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffefffefffefffe)
  ) CLBLM_L_X8Y114_SLICE_X11Y114_DLUT (
.I0(CLBLM_L_X8Y115_SLICE_X11Y115_C5Q),
.I1(CLBLM_L_X8Y114_SLICE_X11Y114_CQ),
.I2(CLBLM_L_X8Y115_SLICE_X11Y115_DQ),
.I3(CLBLM_L_X8Y120_SLICE_X11Y120_CQ),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X8Y114_SLICE_X11Y114_DO5),
.O6(CLBLM_L_X8Y114_SLICE_X11Y114_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h88bb88bb88888888)
  ) CLBLM_L_X8Y114_SLICE_X11Y114_CLUT (
.I0(CLBLM_L_X8Y110_SLICE_X10Y110_BQ),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(1'b1),
.I3(RIOB33_X105Y105_IOB_X1Y105_I),
.I4(1'b1),
.I5(CLBLM_L_X8Y114_SLICE_X10Y114_BQ),
.O5(CLBLM_L_X8Y114_SLICE_X11Y114_CO5),
.O6(CLBLM_L_X8Y114_SLICE_X11Y114_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hc0c0c0c0e2e2e2e2)
  ) CLBLM_L_X8Y114_SLICE_X11Y114_BLUT (
.I0(CLBLM_R_X7Y115_SLICE_X8Y115_CQ),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(CLBLM_L_X8Y114_SLICE_X11Y114_AQ),
.I3(1'b1),
.I4(1'b1),
.I5(RIOB33_X105Y105_IOB_X1Y105_I),
.O5(CLBLM_L_X8Y114_SLICE_X11Y114_BO5),
.O6(CLBLM_L_X8Y114_SLICE_X11Y114_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfdec3120ddcc1100)
  ) CLBLM_L_X8Y114_SLICE_X11Y114_ALUT (
.I0(CLBLM_L_X10Y113_SLICE_X12Y113_DO6),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(CLBLM_L_X8Y114_SLICE_X11Y114_AQ),
.I3(CLBLM_L_X10Y112_SLICE_X12Y112_CQ),
.I4(CLBLM_L_X8Y118_SLICE_X10Y118_AQ),
.I5(RIOB33_X105Y105_IOB_X1Y105_I),
.O5(CLBLM_L_X8Y114_SLICE_X11Y114_AO5),
.O6(CLBLM_L_X8Y114_SLICE_X11Y114_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y115_SLICE_X10Y115_C5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y115_SLICE_X10Y115_CO5),
.Q(CLBLM_L_X8Y115_SLICE_X10Y115_C5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y115_SLICE_X10Y115_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y115_SLICE_X10Y115_AO6),
.Q(CLBLM_L_X8Y115_SLICE_X10Y115_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y115_SLICE_X10Y115_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y115_SLICE_X10Y115_CO6),
.Q(CLBLM_L_X8Y115_SLICE_X10Y115_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y115_SLICE_X10Y115_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y115_SLICE_X10Y115_DO6),
.Q(CLBLM_L_X8Y115_SLICE_X10Y115_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffffaaaaf0c0)
  ) CLBLM_L_X8Y115_SLICE_X10Y115_DLUT (
.I0(CLBLM_R_X3Y114_SLICE_X2Y114_AQ),
.I1(RIOB33_X105Y117_IOB_X1Y118_I),
.I2(CLBLM_L_X8Y115_SLICE_X10Y115_DQ),
.I3(CLBLM_R_X3Y118_SLICE_X2Y118_AQ),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(CLBLM_R_X7Y113_SLICE_X9Y113_CO6),
.O5(CLBLM_L_X8Y115_SLICE_X10Y115_DO5),
.O6(CLBLM_L_X8Y115_SLICE_X10Y115_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hcfc0c0c0fafa0a0a)
  ) CLBLM_L_X8Y115_SLICE_X10Y115_CLUT (
.I0(CLBLM_R_X7Y122_SLICE_X9Y122_AQ),
.I1(CLBLM_R_X7Y116_SLICE_X9Y116_AQ),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(RIOB33_X105Y105_IOB_X1Y105_I),
.I4(CLBLM_L_X8Y114_SLICE_X10Y114_B5Q),
.I5(1'b1),
.O5(CLBLM_L_X8Y115_SLICE_X10Y115_CO5),
.O6(CLBLM_L_X8Y115_SLICE_X10Y115_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfcec3020f0a0f0a0)
  ) CLBLM_L_X8Y115_SLICE_X10Y115_BLUT (
.I0(CLBLM_R_X7Y115_SLICE_X8Y115_CQ),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(RIOB33_X105Y121_IOB_X1Y121_I),
.I3(CLBLM_R_X7Y115_SLICE_X8Y115_AQ),
.I4(CLBLM_R_X11Y113_SLICE_X14Y113_AQ),
.I5(1'b1),
.O5(CLBLM_L_X8Y115_SLICE_X10Y115_BO5),
.O6(CLBLM_L_X8Y115_SLICE_X10Y115_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hff050005ff0a000a)
  ) CLBLM_L_X8Y115_SLICE_X10Y115_ALUT (
.I0(CLBLM_L_X8Y115_SLICE_X10Y115_BO5),
.I1(1'b1),
.I2(RIOB33_X105Y105_IOB_X1Y105_I),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLL_L_X4Y115_SLICE_X5Y115_CQ),
.I5(CLBLM_R_X7Y119_SLICE_X8Y119_BQ),
.O5(CLBLM_L_X8Y115_SLICE_X10Y115_AO5),
.O6(CLBLM_L_X8Y115_SLICE_X10Y115_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y115_SLICE_X11Y115_C5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y115_SLICE_X11Y115_CO5),
.Q(CLBLM_L_X8Y115_SLICE_X11Y115_C5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y115_SLICE_X11Y115_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y115_SLICE_X11Y115_AO6),
.Q(CLBLM_L_X8Y115_SLICE_X11Y115_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y115_SLICE_X11Y115_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y115_SLICE_X11Y115_BO6),
.Q(CLBLM_L_X8Y115_SLICE_X11Y115_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y115_SLICE_X11Y115_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y115_SLICE_X11Y115_CO6),
.Q(CLBLM_L_X8Y115_SLICE_X11Y115_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y115_SLICE_X11Y115_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y115_SLICE_X11Y115_DO6),
.Q(CLBLM_L_X8Y115_SLICE_X11Y115_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hff00ff0022222222)
  ) CLBLM_L_X8Y115_SLICE_X11Y115_DLUT (
.I0(CLBLM_L_X8Y115_SLICE_X11Y115_C5Q),
.I1(RIOB33_X105Y105_IOB_X1Y105_I),
.I2(1'b1),
.I3(CLBLM_L_X10Y120_SLICE_X12Y120_BQ),
.I4(1'b1),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLM_L_X8Y115_SLICE_X11Y115_DO5),
.O6(CLBLM_L_X8Y115_SLICE_X11Y115_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hcfc0cfc0f8f80808)
  ) CLBLM_L_X8Y115_SLICE_X11Y115_CLUT (
.I0(RIOB33_X105Y105_IOB_X1Y105_I),
.I1(CLBLM_R_X7Y119_SLICE_X9Y119_CQ),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLM_L_X8Y119_SLICE_X10Y119_A5Q),
.I4(CLBLM_L_X8Y113_SLICE_X11Y113_AQ),
.I5(1'b1),
.O5(CLBLM_L_X8Y115_SLICE_X11Y115_CO5),
.O6(CLBLM_L_X8Y115_SLICE_X11Y115_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff00e0000000e0)
  ) CLBLM_L_X8Y115_SLICE_X11Y115_BLUT (
.I0(CLBLM_L_X10Y111_SLICE_X13Y111_AQ),
.I1(CLBLM_L_X8Y115_SLICE_X11Y115_BQ),
.I2(CLBLM_R_X3Y118_SLICE_X2Y118_AQ),
.I3(RIOB33_X105Y117_IOB_X1Y118_I),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(CLBLM_L_X10Y115_SLICE_X12Y115_CQ),
.O5(CLBLM_L_X8Y115_SLICE_X11Y115_BO5),
.O6(CLBLM_L_X8Y115_SLICE_X11Y115_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'haa33aa33aa30aa30)
  ) CLBLM_L_X8Y115_SLICE_X11Y115_ALUT (
.I0(CLBLM_L_X10Y111_SLICE_X13Y111_AQ),
.I1(CLBLM_R_X5Y119_SLICE_X7Y119_AO6),
.I2(CLBLM_L_X8Y115_SLICE_X11Y115_AQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(1'b1),
.I5(CLBLM_R_X7Y116_SLICE_X9Y116_AQ),
.O5(CLBLM_L_X8Y115_SLICE_X11Y115_AO5),
.O6(CLBLM_L_X8Y115_SLICE_X11Y115_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y116_SLICE_X10Y116_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(LIOB33_X0Y77_IOB_X0Y77_I),
.D(CLBLM_R_X7Y116_SLICE_X8Y116_AQ),
.Q(CLBLM_L_X8Y116_SLICE_X10Y116_AQ),
.R(CLBLM_R_X11Y123_SLICE_X14Y123_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h6f6ff6f66f6ff6f6)
  ) CLBLM_L_X8Y116_SLICE_X10Y116_DLUT (
.I0(CLBLM_R_X11Y115_SLICE_X15Y115_CQ),
.I1(CLBLM_L_X8Y115_SLICE_X11Y115_CQ),
.I2(CLBLM_L_X10Y122_SLICE_X13Y122_A5Q),
.I3(1'b1),
.I4(CLBLM_R_X7Y116_SLICE_X8Y116_CQ),
.I5(1'b1),
.O5(CLBLM_L_X8Y116_SLICE_X10Y116_DO5),
.O6(CLBLM_L_X8Y116_SLICE_X10Y116_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000a00a00005005)
  ) CLBLM_L_X8Y116_SLICE_X10Y116_CLUT (
.I0(CLBLM_L_X8Y115_SLICE_X11Y115_AQ),
.I1(1'b1),
.I2(CLBLL_L_X4Y119_SLICE_X4Y119_CQ),
.I3(CLBLM_R_X7Y116_SLICE_X9Y116_AQ),
.I4(CLBLM_L_X8Y116_SLICE_X10Y116_DO6),
.I5(CLBLM_L_X10Y127_SLICE_X12Y127_AQ),
.O5(CLBLM_L_X8Y116_SLICE_X10Y116_CO5),
.O6(CLBLM_L_X8Y116_SLICE_X10Y116_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000001)
  ) CLBLM_L_X8Y116_SLICE_X10Y116_BLUT (
.I0(CLBLM_R_X11Y115_SLICE_X15Y115_CQ),
.I1(CLBLM_L_X10Y110_SLICE_X12Y110_BQ),
.I2(CLBLM_L_X8Y117_SLICE_X10Y117_AQ),
.I3(CLBLM_R_X7Y110_SLICE_X9Y110_BQ),
.I4(CLBLM_L_X8Y115_SLICE_X11Y115_AQ),
.I5(CLBLM_L_X10Y115_SLICE_X12Y115_DQ),
.O5(CLBLM_L_X8Y116_SLICE_X10Y116_BO5),
.O6(CLBLM_L_X8Y116_SLICE_X10Y116_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0041008200000000)
  ) CLBLM_L_X8Y116_SLICE_X10Y116_ALUT (
.I0(CLBLM_R_X7Y116_SLICE_X9Y116_CO6),
.I1(CLBLM_R_X7Y115_SLICE_X9Y115_B5Q),
.I2(CLBLM_L_X8Y117_SLICE_X10Y117_AQ),
.I3(CLBLM_L_X8Y110_SLICE_X10Y110_CO6),
.I4(CLBLM_L_X10Y114_SLICE_X13Y114_DQ),
.I5(CLBLM_L_X8Y116_SLICE_X10Y116_CO6),
.O5(CLBLM_L_X8Y116_SLICE_X10Y116_AO5),
.O6(CLBLM_L_X8Y116_SLICE_X10Y116_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y116_SLICE_X11Y116_A5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y116_SLICE_X11Y116_CO6),
.Q(CLBLM_L_X8Y116_SLICE_X11Y116_A5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y116_SLICE_X11Y116_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y116_SLICE_X11Y116_AO6),
.Q(CLBLM_L_X8Y116_SLICE_X11Y116_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y116_SLICE_X11Y116_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y116_SLICE_X11Y116_BO6),
.Q(CLBLM_L_X8Y116_SLICE_X11Y116_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y116_SLICE_X11Y116_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y116_SLICE_X11Y116_DO6),
.Q(CLBLM_L_X8Y116_SLICE_X11Y116_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff00fa000000fa)
  ) CLBLM_L_X8Y116_SLICE_X11Y116_DLUT (
.I0(CLBLM_R_X7Y116_SLICE_X8Y116_AQ),
.I1(1'b1),
.I2(CLBLM_L_X8Y116_SLICE_X11Y116_DQ),
.I3(CLBLM_R_X5Y111_SLICE_X7Y111_DO6),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(CLBLM_L_X10Y115_SLICE_X12Y115_DQ),
.O5(CLBLM_L_X8Y116_SLICE_X11Y116_DO5),
.O6(CLBLM_L_X8Y116_SLICE_X11Y116_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'he2f3f3e200ff0000)
  ) CLBLM_L_X8Y116_SLICE_X11Y116_CLUT (
.I0(CLBLM_R_X11Y119_SLICE_X14Y119_AO6),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(CLBLM_R_X7Y111_SLICE_X8Y111_AQ),
.I3(CLBLM_L_X8Y116_SLICE_X11Y116_A5Q),
.I4(CLBLM_L_X8Y119_SLICE_X10Y119_BQ),
.I5(1'b1),
.O5(CLBLM_L_X8Y116_SLICE_X11Y116_CO5),
.O6(CLBLM_L_X8Y116_SLICE_X11Y116_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hff000000fffc00fc)
  ) CLBLM_L_X8Y116_SLICE_X11Y116_BLUT (
.I0(1'b1),
.I1(CLBLM_L_X8Y116_SLICE_X11Y116_BQ),
.I2(CLBLM_R_X7Y110_SLICE_X9Y110_BQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLM_L_X8Y118_SLICE_X11Y118_AQ),
.I5(CLBLM_R_X5Y111_SLICE_X7Y111_DO6),
.O5(CLBLM_L_X8Y116_SLICE_X11Y116_BO5),
.O6(CLBLM_L_X8Y116_SLICE_X11Y116_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffb8ffb800b800b8)
  ) CLBLM_L_X8Y116_SLICE_X11Y116_ALUT (
.I0(CLBLM_L_X8Y121_SLICE_X10Y121_CQ),
.I1(CLBLM_R_X11Y121_SLICE_X14Y121_CO6),
.I2(CLBLM_L_X8Y116_SLICE_X11Y116_AQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(1'b1),
.I5(CLBLM_L_X8Y111_SLICE_X10Y111_AQ),
.O5(CLBLM_L_X8Y116_SLICE_X11Y116_AO5),
.O6(CLBLM_L_X8Y116_SLICE_X11Y116_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y117_SLICE_X10Y117_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y117_SLICE_X10Y117_AO6),
.Q(CLBLM_L_X8Y117_SLICE_X10Y117_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y117_SLICE_X10Y117_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y117_SLICE_X10Y117_BO6),
.Q(CLBLM_L_X8Y117_SLICE_X10Y117_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y117_SLICE_X10Y117_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y117_SLICE_X10Y117_CO6),
.Q(CLBLM_L_X8Y117_SLICE_X10Y117_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaafc00fc00fc00)
  ) CLBLM_L_X8Y117_SLICE_X10Y117_DLUT (
.I0(CLBLM_L_X8Y117_SLICE_X10Y117_BQ),
.I1(CLBLM_R_X3Y116_SLICE_X3Y116_BQ),
.I2(CLBLM_L_X8Y115_SLICE_X10Y115_DQ),
.I3(RIOB33_X105Y121_IOB_X1Y121_I),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(1'b1),
.O5(CLBLM_L_X8Y117_SLICE_X10Y117_DO5),
.O6(CLBLM_L_X8Y117_SLICE_X10Y117_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hff300030ff200020)
  ) CLBLM_L_X8Y117_SLICE_X10Y117_CLUT (
.I0(CLBLM_L_X8Y117_SLICE_X10Y117_CQ),
.I1(RIOB33_X105Y117_IOB_X1Y118_I),
.I2(CLBLM_R_X3Y118_SLICE_X2Y118_AQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLM_L_X10Y117_SLICE_X12Y117_BQ),
.I5(CLBLM_R_X11Y115_SLICE_X14Y115_CQ),
.O5(CLBLM_L_X8Y117_SLICE_X10Y117_CO5),
.O6(CLBLM_L_X8Y117_SLICE_X10Y117_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hff00ff00f1f1e0e0)
  ) CLBLM_L_X8Y117_SLICE_X10Y117_BLUT (
.I0(CLBLM_R_X3Y118_SLICE_X2Y118_AQ),
.I1(RIOB33_X105Y117_IOB_X1Y118_I),
.I2(CLBLM_R_X3Y116_SLICE_X3Y116_AQ),
.I3(CLBLM_L_X8Y119_SLICE_X10Y119_BQ),
.I4(CLBLM_L_X8Y117_SLICE_X10Y117_BQ),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLM_L_X8Y117_SLICE_X10Y117_BO5),
.O6(CLBLM_L_X8Y117_SLICE_X10Y117_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hcc00cc00ccffccf0)
  ) CLBLM_L_X8Y117_SLICE_X10Y117_ALUT (
.I0(1'b1),
.I1(CLBLM_R_X7Y121_SLICE_X8Y121_AQ),
.I2(CLBLM_L_X8Y117_SLICE_X10Y117_AQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLM_L_X8Y115_SLICE_X11Y115_AQ),
.I5(CLBLM_R_X5Y119_SLICE_X7Y119_AO6),
.O5(CLBLM_L_X8Y117_SLICE_X10Y117_AO5),
.O6(CLBLM_L_X8Y117_SLICE_X10Y117_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y117_SLICE_X11Y117_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y117_SLICE_X11Y117_AO6),
.Q(CLBLM_L_X8Y117_SLICE_X11Y117_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y117_SLICE_X11Y117_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y117_SLICE_X11Y117_BO6),
.Q(CLBLM_L_X8Y117_SLICE_X11Y117_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y117_SLICE_X11Y117_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y117_SLICE_X11Y117_CO6),
.Q(CLBLM_L_X8Y117_SLICE_X11Y117_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y117_SLICE_X11Y117_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y117_SLICE_X11Y117_DO6),
.Q(CLBLM_L_X8Y117_SLICE_X11Y117_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hcccc0000fecc3200)
  ) CLBLM_L_X8Y117_SLICE_X11Y117_DLUT (
.I0(CLBLM_R_X7Y116_SLICE_X8Y116_DO6),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(CLBLM_L_X8Y117_SLICE_X11Y117_DQ),
.I3(CLBLM_R_X3Y118_SLICE_X2Y118_AQ),
.I4(CLBLM_R_X7Y118_SLICE_X8Y118_AQ),
.I5(RIOB33_X105Y117_IOB_X1Y118_I),
.O5(CLBLM_L_X8Y117_SLICE_X11Y117_DO5),
.O6(CLBLM_L_X8Y117_SLICE_X11Y117_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hff00ff00eeeee0e0)
  ) CLBLM_L_X8Y117_SLICE_X11Y117_CLUT (
.I0(CLBLM_R_X7Y116_SLICE_X8Y116_DO6),
.I1(CLBLM_L_X8Y117_SLICE_X11Y117_CQ),
.I2(CLBLM_R_X3Y118_SLICE_X2Y118_AQ),
.I3(CLBLM_R_X7Y120_SLICE_X9Y120_CQ),
.I4(RIOB33_X105Y117_IOB_X1Y118_I),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLM_L_X8Y117_SLICE_X11Y117_CO5),
.O6(CLBLM_L_X8Y117_SLICE_X11Y117_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hff0fff0c000f000c)
  ) CLBLM_L_X8Y117_SLICE_X11Y117_BLUT (
.I0(1'b1),
.I1(CLBLM_L_X8Y117_SLICE_X11Y117_BQ),
.I2(CLBLM_R_X5Y111_SLICE_X7Y111_DO6),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLM_L_X10Y116_SLICE_X13Y116_AO5),
.I5(CLBLM_R_X7Y121_SLICE_X9Y121_A5Q),
.O5(CLBLM_L_X8Y117_SLICE_X11Y117_BO5),
.O6(CLBLM_L_X8Y117_SLICE_X11Y117_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffefff33332333)
  ) CLBLM_L_X8Y117_SLICE_X11Y117_ALUT (
.I0(CLBLM_L_X8Y121_SLICE_X10Y121_DO6),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(RIOB33_X105Y135_IOB_X1Y135_I),
.I3(RIOB33_X105Y131_IOB_X1Y131_I),
.I4(RIOB33_X105Y135_IOB_X1Y136_I),
.I5(CLBLM_L_X10Y114_SLICE_X13Y114_A5Q),
.O5(CLBLM_L_X8Y117_SLICE_X11Y117_AO5),
.O6(CLBLM_L_X8Y117_SLICE_X11Y117_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y118_SLICE_X10Y118_D5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y118_SLICE_X10Y118_DO5),
.Q(CLBLM_L_X8Y118_SLICE_X10Y118_D5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y118_SLICE_X10Y118_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y118_SLICE_X10Y118_AO6),
.Q(CLBLM_L_X8Y118_SLICE_X10Y118_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y118_SLICE_X10Y118_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y118_SLICE_X10Y118_BO6),
.Q(CLBLM_L_X8Y118_SLICE_X10Y118_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y118_SLICE_X10Y118_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y118_SLICE_X10Y118_CO6),
.Q(CLBLM_L_X8Y118_SLICE_X10Y118_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y118_SLICE_X10Y118_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y118_SLICE_X10Y118_DO6),
.Q(CLBLM_L_X8Y118_SLICE_X10Y118_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hfa0afa0afcfc0c0c)
  ) CLBLM_L_X8Y118_SLICE_X10Y118_DLUT (
.I0(CLBLM_L_X8Y120_SLICE_X11Y120_AQ),
.I1(CLBLM_L_X10Y122_SLICE_X12Y122_BQ),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLM_R_X7Y111_SLICE_X8Y111_CQ),
.I4(CLBLM_L_X10Y116_SLICE_X12Y116_CQ),
.I5(1'b1),
.O5(CLBLM_L_X8Y118_SLICE_X10Y118_DO5),
.O6(CLBLM_L_X8Y118_SLICE_X10Y118_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f0aaaaf0f0aacc)
  ) CLBLM_L_X8Y118_SLICE_X10Y118_CLUT (
.I0(CLBLM_L_X8Y115_SLICE_X11Y115_BQ),
.I1(CLBLM_L_X8Y118_SLICE_X10Y118_CQ),
.I2(CLBLM_R_X11Y118_SLICE_X15Y118_CQ),
.I3(RIOB33_X105Y117_IOB_X1Y118_I),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(CLBLM_R_X3Y118_SLICE_X2Y118_AQ),
.O5(CLBLM_L_X8Y118_SLICE_X10Y118_CO5),
.O6(CLBLM_L_X8Y118_SLICE_X10Y118_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hff000f0fff000c0c)
  ) CLBLM_L_X8Y118_SLICE_X10Y118_BLUT (
.I0(1'b1),
.I1(CLBLM_L_X8Y118_SLICE_X10Y118_BQ),
.I2(CLBLM_R_X11Y121_SLICE_X14Y121_CO6),
.I3(CLBLM_L_X10Y112_SLICE_X12Y112_CQ),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(CLBLM_L_X10Y116_SLICE_X12Y116_CQ),
.O5(CLBLM_L_X8Y118_SLICE_X10Y118_BO5),
.O6(CLBLM_L_X8Y118_SLICE_X10Y118_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hcccc00ffcccc00f0)
  ) CLBLM_L_X8Y118_SLICE_X10Y118_ALUT (
.I0(1'b1),
.I1(CLBLM_R_X5Y110_SLICE_X7Y110_CQ),
.I2(CLBLM_L_X8Y118_SLICE_X10Y118_AQ),
.I3(CLBLM_R_X11Y121_SLICE_X14Y121_CO6),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(CLBLM_L_X8Y119_SLICE_X11Y119_CQ),
.O5(CLBLM_L_X8Y118_SLICE_X10Y118_AO5),
.O6(CLBLM_L_X8Y118_SLICE_X10Y118_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y118_SLICE_X11Y118_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y118_SLICE_X11Y118_AO6),
.Q(CLBLM_L_X8Y118_SLICE_X11Y118_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X8Y118_SLICE_X11Y118_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X8Y118_SLICE_X11Y118_DO5),
.O6(CLBLM_L_X8Y118_SLICE_X11Y118_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X8Y118_SLICE_X11Y118_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X8Y118_SLICE_X11Y118_CO5),
.O6(CLBLM_L_X8Y118_SLICE_X11Y118_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hafa0aca0ff00cc00)
  ) CLBLM_L_X8Y118_SLICE_X11Y118_BLUT (
.I0(CLBLM_R_X5Y124_SLICE_X6Y124_CQ),
.I1(CLBLM_L_X8Y114_SLICE_X10Y114_BQ),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(RIOB33_X105Y121_IOB_X1Y121_I),
.I4(CLBLM_L_X8Y117_SLICE_X11Y117_CQ),
.I5(1'b1),
.O5(CLBLM_L_X8Y118_SLICE_X11Y118_BO5),
.O6(CLBLM_L_X8Y118_SLICE_X11Y118_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hcccc00facccc00fa)
  ) CLBLM_L_X8Y118_SLICE_X11Y118_ALUT (
.I0(CLBLM_L_X10Y119_SLICE_X13Y119_DQ),
.I1(CLBLM_L_X10Y118_SLICE_X12Y118_BQ),
.I2(CLBLM_L_X8Y118_SLICE_X11Y118_AQ),
.I3(CLBLM_R_X11Y121_SLICE_X14Y121_CO6),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(1'b1),
.O5(CLBLM_L_X8Y118_SLICE_X11Y118_AO5),
.O6(CLBLM_L_X8Y118_SLICE_X11Y118_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y119_SLICE_X10Y119_A5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y119_SLICE_X10Y119_DO6),
.Q(CLBLM_L_X8Y119_SLICE_X10Y119_A5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y119_SLICE_X10Y119_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y119_SLICE_X10Y119_AO6),
.Q(CLBLM_L_X8Y119_SLICE_X10Y119_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y119_SLICE_X10Y119_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y119_SLICE_X10Y119_BO6),
.Q(CLBLM_L_X8Y119_SLICE_X10Y119_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y119_SLICE_X10Y119_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y119_SLICE_X10Y119_CO6),
.Q(CLBLM_L_X8Y119_SLICE_X10Y119_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hfa50ea40f0f0c0c0)
  ) CLBLM_L_X8Y119_SLICE_X10Y119_DLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_L_X8Y114_SLICE_X10Y114_C5Q),
.I2(RIOB33_X105Y121_IOB_X1Y121_I),
.I3(CLBLM_L_X8Y110_SLICE_X10Y110_AQ),
.I4(CLBLM_L_X10Y119_SLICE_X12Y119_AQ),
.I5(1'b1),
.O5(CLBLM_L_X8Y119_SLICE_X10Y119_DO5),
.O6(CLBLM_L_X8Y119_SLICE_X10Y119_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'ha0a0e4e4a0a0e4e4)
  ) CLBLM_L_X8Y119_SLICE_X10Y119_CLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_L_X10Y119_SLICE_X13Y119_CQ),
.I2(CLBLM_L_X8Y120_SLICE_X10Y120_DQ),
.I3(1'b1),
.I4(CLBLM_L_X12Y120_SLICE_X17Y120_CO6),
.I5(1'b1),
.O5(CLBLM_L_X8Y119_SLICE_X10Y119_CO5),
.O6(CLBLM_L_X8Y119_SLICE_X10Y119_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf505f000f505f000)
  ) CLBLM_L_X8Y119_SLICE_X10Y119_BLUT (
.I0(CLBLM_L_X12Y120_SLICE_X17Y120_CO6),
.I1(1'b1),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLM_L_X8Y115_SLICE_X10Y115_AQ),
.I4(CLBLM_L_X8Y120_SLICE_X10Y120_AQ),
.I5(1'b1),
.O5(CLBLM_L_X8Y119_SLICE_X10Y119_BO5),
.O6(CLBLM_L_X8Y119_SLICE_X10Y119_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffdff33333133)
  ) CLBLM_L_X8Y119_SLICE_X10Y119_ALUT (
.I0(RIOB33_X105Y131_IOB_X1Y131_I),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(RIOB33_X105Y135_IOB_X1Y135_I),
.I3(RIOB33_X105Y135_IOB_X1Y136_I),
.I4(CLBLM_L_X8Y121_SLICE_X10Y121_DO6),
.I5(CLBLM_L_X10Y119_SLICE_X13Y119_CQ),
.O5(CLBLM_L_X8Y119_SLICE_X10Y119_AO5),
.O6(CLBLM_L_X8Y119_SLICE_X10Y119_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y119_SLICE_X11Y119_C5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y119_SLICE_X11Y119_CO5),
.Q(CLBLM_L_X8Y119_SLICE_X11Y119_C5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y119_SLICE_X11Y119_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y119_SLICE_X11Y119_AO6),
.Q(CLBLM_L_X8Y119_SLICE_X11Y119_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y119_SLICE_X11Y119_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y119_SLICE_X11Y119_BO6),
.Q(CLBLM_L_X8Y119_SLICE_X11Y119_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y119_SLICE_X11Y119_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y119_SLICE_X11Y119_CO6),
.Q(CLBLM_L_X8Y119_SLICE_X11Y119_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y119_SLICE_X11Y119_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y119_SLICE_X11Y119_DO6),
.Q(CLBLM_L_X8Y119_SLICE_X11Y119_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaafcfcaaaafcf0)
  ) CLBLM_L_X8Y119_SLICE_X11Y119_DLUT (
.I0(CLBLM_L_X8Y116_SLICE_X11Y116_BQ),
.I1(CLBLM_L_X10Y123_SLICE_X12Y123_AO6),
.I2(CLBLM_L_X8Y122_SLICE_X11Y122_CO6),
.I3(CLBLM_R_X5Y118_SLICE_X7Y118_CO6),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(CLBLM_R_X3Y117_SLICE_X3Y117_BQ),
.O5(CLBLM_L_X8Y119_SLICE_X11Y119_DO5),
.O6(CLBLM_L_X8Y119_SLICE_X11Y119_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaa00ccccccf0f0)
  ) CLBLM_L_X8Y119_SLICE_X11Y119_CLUT (
.I0(CLBLM_R_X7Y116_SLICE_X8Y116_BQ),
.I1(CLBLM_L_X10Y119_SLICE_X13Y119_DQ),
.I2(CLBLM_R_X7Y121_SLICE_X9Y121_A5Q),
.I3(RIOB33_X105Y105_IOB_X1Y105_I),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(1'b1),
.O5(CLBLM_L_X8Y119_SLICE_X11Y119_CO5),
.O6(CLBLM_L_X8Y119_SLICE_X11Y119_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f00055f0f000aa)
  ) CLBLM_L_X8Y119_SLICE_X11Y119_BLUT (
.I0(CLBLM_L_X8Y118_SLICE_X11Y118_BO5),
.I1(1'b1),
.I2(CLBLM_L_X12Y120_SLICE_X17Y120_AQ),
.I3(RIOB33_X105Y105_IOB_X1Y105_I),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(CLBLM_L_X8Y121_SLICE_X10Y121_CQ),
.O5(CLBLM_L_X8Y119_SLICE_X11Y119_BO5),
.O6(CLBLM_L_X8Y119_SLICE_X11Y119_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfb51ea40fb51ea40)
  ) CLBLM_L_X8Y119_SLICE_X11Y119_ALUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_R_X11Y121_SLICE_X14Y121_CO6),
.I2(CLBLM_L_X8Y119_SLICE_X11Y119_AQ),
.I3(CLBLM_L_X10Y120_SLICE_X12Y120_AQ),
.I4(CLBLM_R_X7Y119_SLICE_X8Y119_BQ),
.I5(1'b1),
.O5(CLBLM_L_X8Y119_SLICE_X11Y119_AO5),
.O6(CLBLM_L_X8Y119_SLICE_X11Y119_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y120_SLICE_X10Y120_A5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y120_SLICE_X10Y120_AO5),
.Q(CLBLM_L_X8Y120_SLICE_X10Y120_A5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y120_SLICE_X10Y120_D5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y120_SLICE_X10Y120_DO5),
.Q(CLBLM_L_X8Y120_SLICE_X10Y120_D5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y120_SLICE_X10Y120_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y120_SLICE_X10Y120_AO6),
.Q(CLBLM_L_X8Y120_SLICE_X10Y120_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y120_SLICE_X10Y120_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y120_SLICE_X10Y120_BO6),
.Q(CLBLM_L_X8Y120_SLICE_X10Y120_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y120_SLICE_X10Y120_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y120_SLICE_X10Y120_CO6),
.Q(CLBLM_L_X8Y120_SLICE_X10Y120_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y120_SLICE_X10Y120_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y120_SLICE_X10Y120_DO6),
.Q(CLBLM_L_X8Y120_SLICE_X10Y120_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hee44ee44f5f5a0a0)
  ) CLBLM_L_X8Y120_SLICE_X10Y120_DLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLL_L_X2Y120_SLICE_X1Y120_DO6),
.I2(CLBLM_L_X8Y122_SLICE_X11Y122_BQ),
.I3(CLBLM_R_X7Y112_SLICE_X9Y112_AQ),
.I4(CLBLL_L_X4Y120_SLICE_X5Y120_DO6),
.I5(1'b1),
.O5(CLBLM_L_X8Y120_SLICE_X10Y120_DO5),
.O6(CLBLM_L_X8Y120_SLICE_X10Y120_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hb1f5f5f5f5f5f5f5)
  ) CLBLM_L_X8Y120_SLICE_X10Y120_CLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_L_X8Y120_SLICE_X10Y120_CQ),
.I2(CLBLM_R_X7Y118_SLICE_X9Y118_AQ),
.I3(CLBLM_L_X8Y120_SLICE_X10Y120_A5Q),
.I4(RIOB33_X105Y105_IOB_X1Y105_I),
.I5(CLBLM_L_X8Y120_SLICE_X11Y120_C5Q),
.O5(CLBLM_L_X8Y120_SLICE_X10Y120_CO5),
.O6(CLBLM_L_X8Y120_SLICE_X10Y120_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'ha0a0a0a0afa0afa0)
  ) CLBLM_L_X8Y120_SLICE_X10Y120_BLUT (
.I0(CLBLM_L_X10Y121_SLICE_X12Y121_BQ),
.I1(1'b1),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLM_R_X7Y122_SLICE_X9Y122_BQ),
.I4(1'b1),
.I5(RIOB33_X105Y105_IOB_X1Y105_I),
.O5(CLBLM_L_X8Y120_SLICE_X10Y120_BO5),
.O6(CLBLM_L_X8Y120_SLICE_X10Y120_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hff005050ccccff00)
  ) CLBLM_L_X8Y120_SLICE_X10Y120_ALUT (
.I0(CLBLM_L_X12Y120_SLICE_X17Y120_CO6),
.I1(CLBLM_L_X8Y120_SLICE_X11Y120_CQ),
.I2(CLBLM_L_X8Y119_SLICE_X10Y119_CQ),
.I3(CLBLM_R_X7Y121_SLICE_X8Y121_CQ),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(1'b1),
.O5(CLBLM_L_X8Y120_SLICE_X10Y120_AO5),
.O6(CLBLM_L_X8Y120_SLICE_X10Y120_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y120_SLICE_X11Y120_C5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y120_SLICE_X11Y120_CO5),
.Q(CLBLM_L_X8Y120_SLICE_X11Y120_C5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y120_SLICE_X11Y120_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y120_SLICE_X11Y120_AO6),
.Q(CLBLM_L_X8Y120_SLICE_X11Y120_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y120_SLICE_X11Y120_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y120_SLICE_X11Y120_BO6),
.Q(CLBLM_L_X8Y120_SLICE_X11Y120_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y120_SLICE_X11Y120_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y120_SLICE_X11Y120_CO6),
.Q(CLBLM_L_X8Y120_SLICE_X11Y120_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h5a5a5a5a5a5a5a5a)
  ) CLBLM_L_X8Y120_SLICE_X11Y120_DLUT (
.I0(CLBLM_L_X10Y126_SLICE_X12Y126_AQ),
.I1(1'b1),
.I2(CLBLL_L_X4Y117_SLICE_X5Y117_DQ),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X8Y120_SLICE_X11Y120_DO5),
.O6(CLBLM_L_X8Y120_SLICE_X11Y120_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'haafa0050e4e4e4e4)
  ) CLBLM_L_X8Y120_SLICE_X11Y120_CLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_L_X8Y120_SLICE_X10Y120_A5Q),
.I2(CLBLM_L_X8Y115_SLICE_X11Y115_DQ),
.I3(RIOB33_X105Y105_IOB_X1Y105_I),
.I4(CLBLM_R_X7Y124_SLICE_X8Y124_AQ),
.I5(1'b1),
.O5(CLBLM_L_X8Y120_SLICE_X11Y120_CO5),
.O6(CLBLM_L_X8Y120_SLICE_X11Y120_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'ha0acafafa0aca0a0)
  ) CLBLM_L_X8Y120_SLICE_X11Y120_BLUT (
.I0(CLBLM_L_X8Y115_SLICE_X10Y115_DQ),
.I1(CLBLM_L_X8Y120_SLICE_X11Y120_BQ),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLM_L_X10Y123_SLICE_X12Y123_AO6),
.I4(CLBLM_R_X7Y123_SLICE_X9Y123_CO6),
.I5(CLBLM_L_X10Y121_SLICE_X12Y121_BQ),
.O5(CLBLM_L_X8Y120_SLICE_X11Y120_BO5),
.O6(CLBLM_L_X8Y120_SLICE_X11Y120_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffffb0000fffb)
  ) CLBLM_L_X8Y120_SLICE_X11Y120_ALUT (
.I0(CLBLM_L_X8Y121_SLICE_X10Y121_DO6),
.I1(RIOB33_X105Y135_IOB_X1Y135_I),
.I2(RIOB33_X105Y131_IOB_X1Y131_I),
.I3(RIOB33_X105Y135_IOB_X1Y136_I),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(CLBLM_L_X8Y122_SLICE_X11Y122_A5Q),
.O5(CLBLM_L_X8Y120_SLICE_X11Y120_AO5),
.O6(CLBLM_L_X8Y120_SLICE_X11Y120_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y121_SLICE_X10Y121_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y121_SLICE_X10Y121_AO6),
.Q(CLBLM_L_X8Y121_SLICE_X10Y121_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y121_SLICE_X10Y121_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y121_SLICE_X10Y121_BO6),
.Q(CLBLM_L_X8Y121_SLICE_X10Y121_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y121_SLICE_X10Y121_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y121_SLICE_X10Y121_CO6),
.Q(CLBLM_L_X8Y121_SLICE_X10Y121_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffffffffffffe)
  ) CLBLM_L_X8Y121_SLICE_X10Y121_DLUT (
.I0(RIOB33_X105Y137_IOB_X1Y137_I),
.I1(RIOB33_X105Y131_IOB_X1Y132_I),
.I2(RIOB33_X105Y133_IOB_X1Y133_I),
.I3(RIOB33_X105Y127_IOB_X1Y128_I),
.I4(RIOB33_X105Y133_IOB_X1Y134_I),
.I5(RIOB33_X105Y129_IOB_X1Y130_I),
.O5(CLBLM_L_X8Y121_SLICE_X10Y121_DO5),
.O6(CLBLM_L_X8Y121_SLICE_X10Y121_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'haaee0044aaee0044)
  ) CLBLM_L_X8Y121_SLICE_X10Y121_CLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_L_X8Y121_SLICE_X11Y121_DQ),
.I2(1'b1),
.I3(RIOB33_X105Y105_IOB_X1Y105_I),
.I4(CLBLM_R_X7Y117_SLICE_X9Y117_DQ),
.I5(1'b1),
.O5(CLBLM_L_X8Y121_SLICE_X10Y121_CO5),
.O6(CLBLM_L_X8Y121_SLICE_X10Y121_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'haaccaafcaa00aa00)
  ) CLBLM_L_X8Y121_SLICE_X10Y121_BLUT (
.I0(CLBLM_L_X8Y119_SLICE_X11Y119_DQ),
.I1(CLBLM_L_X8Y121_SLICE_X10Y121_BQ),
.I2(CLBLM_R_X7Y114_SLICE_X8Y114_BQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(RIOB33_X105Y121_IOB_X1Y121_I),
.I5(RIOB33_X105Y105_IOB_X1Y105_I),
.O5(CLBLM_L_X8Y121_SLICE_X10Y121_BO5),
.O6(CLBLM_L_X8Y121_SLICE_X10Y121_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h88d888d8dddd8888)
  ) CLBLM_L_X8Y121_SLICE_X10Y121_ALUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_L_X8Y114_SLICE_X10Y114_CQ),
.I2(CLBLM_L_X8Y121_SLICE_X10Y121_AQ),
.I3(CLBLM_L_X10Y123_SLICE_X12Y123_AO6),
.I4(CLBLM_L_X8Y122_SLICE_X11Y122_AQ),
.I5(CLBLM_R_X7Y123_SLICE_X9Y123_CO6),
.O5(CLBLM_L_X8Y121_SLICE_X10Y121_AO5),
.O6(CLBLM_L_X8Y121_SLICE_X10Y121_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y121_SLICE_X11Y121_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y121_SLICE_X11Y121_AO6),
.Q(CLBLM_L_X8Y121_SLICE_X11Y121_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y121_SLICE_X11Y121_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y121_SLICE_X11Y121_BO6),
.Q(CLBLM_L_X8Y121_SLICE_X11Y121_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y121_SLICE_X11Y121_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y121_SLICE_X11Y121_CO6),
.Q(CLBLM_L_X8Y121_SLICE_X11Y121_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y121_SLICE_X11Y121_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y121_SLICE_X11Y121_DO6),
.Q(CLBLM_L_X8Y121_SLICE_X11Y121_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hab01aa00ea40be14)
  ) CLBLM_L_X8Y121_SLICE_X11Y121_DLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_L_X10Y119_SLICE_X13Y119_DQ),
.I2(CLBLM_L_X8Y121_SLICE_X11Y121_DQ),
.I3(CLBLM_R_X7Y122_SLICE_X9Y122_AQ),
.I4(CLBLM_L_X8Y120_SLICE_X11Y120_DO6),
.I5(RIOB33_X105Y105_IOB_X1Y105_I),
.O5(CLBLM_L_X8Y121_SLICE_X11Y121_DO5),
.O6(CLBLM_L_X8Y121_SLICE_X11Y121_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffff0fe0f0f000e)
  ) CLBLM_L_X8Y121_SLICE_X11Y121_CLUT (
.I0(CLBLM_L_X8Y121_SLICE_X10Y121_AQ),
.I1(CLBLM_L_X8Y121_SLICE_X11Y121_CQ),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLM_R_X7Y123_SLICE_X9Y123_CO6),
.I4(CLBLM_L_X10Y123_SLICE_X12Y123_AO6),
.I5(CLBLM_R_X5Y121_SLICE_X6Y121_AQ),
.O5(CLBLM_L_X8Y121_SLICE_X11Y121_CO5),
.O6(CLBLM_L_X8Y121_SLICE_X11Y121_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hff440044fff000f0)
  ) CLBLM_L_X8Y121_SLICE_X11Y121_BLUT (
.I0(CLBLM_L_X10Y123_SLICE_X12Y123_AO6),
.I1(CLBLM_L_X8Y121_SLICE_X11Y121_BQ),
.I2(CLBLM_L_X8Y121_SLICE_X11Y121_AQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLM_R_X3Y118_SLICE_X2Y118_AQ),
.I5(CLBLM_R_X7Y123_SLICE_X9Y123_CO6),
.O5(CLBLM_L_X8Y121_SLICE_X11Y121_BO5),
.O6(CLBLM_L_X8Y121_SLICE_X11Y121_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hff300030ffaa00aa)
  ) CLBLM_L_X8Y121_SLICE_X11Y121_ALUT (
.I0(CLBLM_L_X8Y120_SLICE_X11Y120_BQ),
.I1(CLBLM_L_X10Y123_SLICE_X12Y123_AO6),
.I2(CLBLM_L_X8Y121_SLICE_X11Y121_AQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLM_L_X8Y119_SLICE_X11Y119_C5Q),
.I5(CLBLM_R_X7Y123_SLICE_X9Y123_CO6),
.O5(CLBLM_L_X8Y121_SLICE_X11Y121_AO5),
.O6(CLBLM_L_X8Y121_SLICE_X11Y121_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y122_SLICE_X10Y122_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(LIOB33_X0Y77_IOB_X0Y77_I),
.D(CLBLM_R_X7Y122_SLICE_X9Y122_BQ),
.Q(CLBLM_L_X8Y122_SLICE_X10Y122_AQ),
.R(CLBLM_R_X11Y123_SLICE_X14Y123_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hc3c63636c3c6c6c6)
  ) CLBLM_L_X8Y122_SLICE_X10Y122_DLUT (
.I0(CLBLM_R_X5Y120_SLICE_X6Y120_A5Q),
.I1(CLBLM_R_X5Y111_SLICE_X7Y111_CO5),
.I2(CLBLM_L_X8Y119_SLICE_X11Y119_DQ),
.I3(CLBLM_R_X7Y120_SLICE_X9Y120_A5Q),
.I4(CLBLM_L_X10Y124_SLICE_X12Y124_AQ),
.I5(CLBLM_R_X7Y124_SLICE_X8Y124_AQ),
.O5(CLBLM_L_X8Y122_SLICE_X10Y122_DO5),
.O6(CLBLM_L_X8Y122_SLICE_X10Y122_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000008cffffffff)
  ) CLBLM_L_X8Y122_SLICE_X10Y122_CLUT (
.I0(CLBLM_L_X8Y122_SLICE_X10Y122_AO6),
.I1(CLBLM_R_X7Y122_SLICE_X8Y122_CQ),
.I2(CLBLM_L_X10Y118_SLICE_X12Y118_B5Q),
.I3(CLBLM_L_X10Y124_SLICE_X13Y124_BO6),
.I4(CLBLM_L_X8Y122_SLICE_X10Y122_DO6),
.I5(CLBLM_L_X10Y122_SLICE_X12Y122_BQ),
.O5(CLBLM_L_X8Y122_SLICE_X10Y122_CO5),
.O6(CLBLM_L_X8Y122_SLICE_X10Y122_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'haa00aaaafffcfffc)
  ) CLBLM_L_X8Y122_SLICE_X10Y122_BLUT (
.I0(CLBLM_L_X8Y120_SLICE_X10Y120_DQ),
.I1(RIOB33_X105Y127_IOB_X1Y128_I),
.I2(RIOB33_X105Y129_IOB_X1Y130_I),
.I3(RIOB33_X105Y129_IOB_X1Y129_I),
.I4(RIOB33_X105Y137_IOB_X1Y137_I),
.I5(1'b1),
.O5(CLBLM_L_X8Y122_SLICE_X10Y122_BO5),
.O6(CLBLM_L_X8Y122_SLICE_X10Y122_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffcc50500000)
  ) CLBLM_L_X8Y122_SLICE_X10Y122_ALUT (
.I0(CLBLM_L_X10Y118_SLICE_X12Y118_B5Q),
.I1(CLBLM_R_X7Y120_SLICE_X9Y120_A5Q),
.I2(CLBLM_L_X10Y124_SLICE_X12Y124_AQ),
.I3(CLBLM_R_X7Y124_SLICE_X8Y124_AQ),
.I4(CLBLM_R_X5Y120_SLICE_X6Y120_A5Q),
.I5(1'b1),
.O5(CLBLM_L_X8Y122_SLICE_X10Y122_AO5),
.O6(CLBLM_L_X8Y122_SLICE_X10Y122_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y122_SLICE_X11Y122_A5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y115_SLICE_X10Y115_BO6),
.Q(CLBLM_L_X8Y122_SLICE_X11Y122_A5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y122_SLICE_X11Y122_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y122_SLICE_X11Y122_AO6),
.Q(CLBLM_L_X8Y122_SLICE_X11Y122_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y122_SLICE_X11Y122_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y122_SLICE_X11Y122_BO6),
.Q(CLBLM_L_X8Y122_SLICE_X11Y122_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h00ff33ff11ff33ff)
  ) CLBLM_L_X8Y122_SLICE_X11Y122_DLUT (
.I0(CLBLM_R_X7Y120_SLICE_X9Y120_A5Q),
.I1(CLBLM_L_X8Y122_SLICE_X10Y122_AO5),
.I2(1'b1),
.I3(CLBLM_R_X7Y123_SLICE_X9Y123_BO5),
.I4(CLBLM_L_X8Y119_SLICE_X11Y119_DQ),
.I5(CLBLM_R_X7Y124_SLICE_X8Y124_AQ),
.O5(CLBLM_L_X8Y122_SLICE_X11Y122_DO5),
.O6(CLBLM_L_X8Y122_SLICE_X11Y122_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h00ffff0000fecc00)
  ) CLBLM_L_X8Y122_SLICE_X11Y122_CLUT (
.I0(CLBLM_R_X5Y120_SLICE_X6Y120_A5Q),
.I1(CLBLM_R_X7Y124_SLICE_X8Y124_AQ),
.I2(CLBLM_L_X10Y124_SLICE_X12Y124_AQ),
.I3(CLBLM_R_X7Y123_SLICE_X9Y123_BO5),
.I4(CLBLM_L_X8Y119_SLICE_X11Y119_DQ),
.I5(CLBLM_R_X7Y120_SLICE_X9Y120_A5Q),
.O5(CLBLM_L_X8Y122_SLICE_X11Y122_CO5),
.O6(CLBLM_L_X8Y122_SLICE_X11Y122_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf055f0ddf000f088)
  ) CLBLM_L_X8Y122_SLICE_X11Y122_BLUT (
.I0(CLBLM_R_X7Y123_SLICE_X9Y123_CO6),
.I1(CLBLM_L_X8Y122_SLICE_X11Y122_BQ),
.I2(CLBLM_R_X5Y123_SLICE_X6Y123_CQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLM_L_X10Y123_SLICE_X12Y123_AO6),
.I5(CLBLM_L_X8Y121_SLICE_X11Y121_CQ),
.O5(CLBLM_L_X8Y122_SLICE_X11Y122_BO5),
.O6(CLBLM_L_X8Y122_SLICE_X11Y122_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h8888b8b8bb88bb88)
  ) CLBLM_L_X8Y122_SLICE_X11Y122_ALUT (
.I0(CLBLM_R_X5Y122_SLICE_X7Y122_CQ),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(CLBLM_L_X8Y122_SLICE_X11Y122_AQ),
.I3(CLBLM_L_X8Y121_SLICE_X11Y121_BQ),
.I4(CLBLM_L_X10Y123_SLICE_X12Y123_AO6),
.I5(CLBLM_R_X7Y123_SLICE_X9Y123_CO6),
.O5(CLBLM_L_X8Y122_SLICE_X11Y122_AO5),
.O6(CLBLM_L_X8Y122_SLICE_X11Y122_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y123_SLICE_X10Y123_A5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y123_SLICE_X10Y123_AO5),
.Q(CLBLM_L_X8Y123_SLICE_X10Y123_A5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y123_SLICE_X10Y123_B5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y123_SLICE_X10Y123_BO5),
.Q(CLBLM_L_X8Y123_SLICE_X10Y123_B5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y123_SLICE_X10Y123_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y123_SLICE_X10Y123_AO6),
.Q(CLBLM_L_X8Y123_SLICE_X10Y123_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y123_SLICE_X10Y123_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y123_SLICE_X10Y123_BO6),
.Q(CLBLM_L_X8Y123_SLICE_X10Y123_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X8Y123_SLICE_X10Y123_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X8Y123_SLICE_X10Y123_DO5),
.O6(CLBLM_L_X8Y123_SLICE_X10Y123_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X8Y123_SLICE_X10Y123_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X8Y123_SLICE_X10Y123_CO5),
.O6(CLBLM_L_X8Y123_SLICE_X10Y123_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hccccc3c3a9a9aaaa)
  ) CLBLM_L_X8Y123_SLICE_X10Y123_BLUT (
.I0(CLBLM_L_X8Y123_SLICE_X10Y123_B5Q),
.I1(CLBLM_L_X8Y123_SLICE_X10Y123_BQ),
.I2(CLBLM_R_X7Y118_SLICE_X9Y118_DO6),
.I3(1'b1),
.I4(CLBLM_L_X8Y123_SLICE_X10Y123_A5Q),
.I5(1'b1),
.O5(CLBLM_L_X8Y123_SLICE_X10Y123_BO5),
.O6(CLBLM_L_X8Y123_SLICE_X10Y123_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h111100000f0ff0f0)
  ) CLBLM_L_X8Y123_SLICE_X10Y123_ALUT (
.I0(CLBLM_L_X8Y123_SLICE_X10Y123_B5Q),
.I1(CLBLM_L_X8Y123_SLICE_X10Y123_BQ),
.I2(CLBLM_R_X7Y118_SLICE_X9Y118_DO6),
.I3(1'b1),
.I4(CLBLM_L_X8Y123_SLICE_X10Y123_A5Q),
.I5(1'b1),
.O5(CLBLM_L_X8Y123_SLICE_X10Y123_AO5),
.O6(CLBLM_L_X8Y123_SLICE_X10Y123_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y123_SLICE_X11Y123_A5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y123_SLICE_X11Y123_AO5),
.Q(CLBLM_L_X8Y123_SLICE_X11Y123_A5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y123_SLICE_X11Y123_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y123_SLICE_X11Y123_AO6),
.Q(CLBLM_L_X8Y123_SLICE_X11Y123_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X8Y123_SLICE_X11Y123_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X8Y123_SLICE_X11Y123_DO5),
.O6(CLBLM_L_X8Y123_SLICE_X11Y123_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X8Y123_SLICE_X11Y123_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X8Y123_SLICE_X11Y123_CO5),
.O6(CLBLM_L_X8Y123_SLICE_X11Y123_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X8Y123_SLICE_X11Y123_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X8Y123_SLICE_X11Y123_BO5),
.O6(CLBLM_L_X8Y123_SLICE_X11Y123_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hff0ff000afafa0a0)
  ) CLBLM_L_X8Y123_SLICE_X11Y123_ALUT (
.I0(CLBLM_R_X11Y120_SLICE_X15Y120_AQ),
.I1(1'b1),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLL_L_X4Y123_SLICE_X4Y123_AQ),
.I4(RIOB33_X105Y125_IOB_X1Y126_I),
.I5(1'b1),
.O5(CLBLM_L_X8Y123_SLICE_X11Y123_AO5),
.O6(CLBLM_L_X8Y123_SLICE_X11Y123_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X8Y128_SLICE_X10Y128_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X8Y128_SLICE_X10Y128_DO5),
.O6(CLBLM_L_X8Y128_SLICE_X10Y128_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X8Y128_SLICE_X10Y128_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X8Y128_SLICE_X10Y128_CO5),
.O6(CLBLM_L_X8Y128_SLICE_X10Y128_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X8Y128_SLICE_X10Y128_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X8Y128_SLICE_X10Y128_BO5),
.O6(CLBLM_L_X8Y128_SLICE_X10Y128_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffaa5500ffff3333)
  ) CLBLM_L_X8Y128_SLICE_X10Y128_ALUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(RIOB33_X105Y143_IOB_X1Y143_I),
.I2(1'b1),
.I3(CLBLL_L_X4Y121_SLICE_X5Y121_BO5),
.I4(CLBLM_L_X8Y122_SLICE_X10Y122_AQ),
.I5(1'b1),
.O5(CLBLM_L_X8Y128_SLICE_X10Y128_AO5),
.O6(CLBLM_L_X8Y128_SLICE_X10Y128_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X8Y128_SLICE_X11Y128_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X8Y128_SLICE_X11Y128_DO5),
.O6(CLBLM_L_X8Y128_SLICE_X11Y128_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X8Y128_SLICE_X11Y128_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X8Y128_SLICE_X11Y128_CO5),
.O6(CLBLM_L_X8Y128_SLICE_X11Y128_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X8Y128_SLICE_X11Y128_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X8Y128_SLICE_X11Y128_BO5),
.O6(CLBLM_L_X8Y128_SLICE_X11Y128_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X8Y128_SLICE_X11Y128_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X8Y128_SLICE_X11Y128_AO5),
.O6(CLBLM_L_X8Y128_SLICE_X11Y128_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X8Y133_SLICE_X10Y133_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X8Y133_SLICE_X10Y133_DO5),
.O6(CLBLM_L_X8Y133_SLICE_X10Y133_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X8Y133_SLICE_X10Y133_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X8Y133_SLICE_X10Y133_CO5),
.O6(CLBLM_L_X8Y133_SLICE_X10Y133_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X8Y133_SLICE_X10Y133_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X8Y133_SLICE_X10Y133_BO5),
.O6(CLBLM_L_X8Y133_SLICE_X10Y133_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X8Y133_SLICE_X10Y133_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X8Y133_SLICE_X10Y133_AO5),
.O6(CLBLM_L_X8Y133_SLICE_X10Y133_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X8Y133_SLICE_X11Y133_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X8Y133_SLICE_X11Y133_DO5),
.O6(CLBLM_L_X8Y133_SLICE_X11Y133_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X8Y133_SLICE_X11Y133_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X8Y133_SLICE_X11Y133_CO5),
.O6(CLBLM_L_X8Y133_SLICE_X11Y133_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X8Y133_SLICE_X11Y133_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X8Y133_SLICE_X11Y133_BO5),
.O6(CLBLM_L_X8Y133_SLICE_X11Y133_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h7777ffffc000c000)
  ) CLBLM_L_X8Y133_SLICE_X11Y133_ALUT (
.I0(CLBLM_L_X8Y120_SLICE_X10Y120_A5Q),
.I1(RIOB33_X105Y105_IOB_X1Y105_I),
.I2(RIOB33_X105Y139_IOB_X1Y140_I),
.I3(RIOB33_X105Y141_IOB_X1Y141_I),
.I4(CLBLM_L_X8Y120_SLICE_X11Y120_C5Q),
.I5(1'b1),
.O5(CLBLM_L_X8Y133_SLICE_X11Y133_AO5),
.O6(CLBLM_L_X8Y133_SLICE_X11Y133_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y110_SLICE_X12Y110_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y110_SLICE_X12Y110_AO6),
.Q(CLBLM_L_X10Y110_SLICE_X12Y110_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y110_SLICE_X12Y110_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y110_SLICE_X12Y110_BO6),
.Q(CLBLM_L_X10Y110_SLICE_X12Y110_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X10Y110_SLICE_X12Y110_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X10Y110_SLICE_X12Y110_DO5),
.O6(CLBLM_L_X10Y110_SLICE_X12Y110_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X10Y110_SLICE_X12Y110_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X10Y110_SLICE_X12Y110_CO5),
.O6(CLBLM_L_X10Y110_SLICE_X12Y110_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f0f0f055445544)
  ) CLBLM_L_X10Y110_SLICE_X12Y110_BLUT (
.I0(CLBLM_R_X5Y111_SLICE_X7Y111_DO6),
.I1(CLBLM_L_X10Y110_SLICE_X12Y110_BQ),
.I2(CLBLM_L_X10Y110_SLICE_X12Y110_AQ),
.I3(CLBLM_L_X8Y116_SLICE_X11Y116_BQ),
.I4(1'b1),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLM_L_X10Y110_SLICE_X12Y110_BO5),
.O6(CLBLM_L_X10Y110_SLICE_X12Y110_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'haabeaaaa00140000)
  ) CLBLM_L_X10Y110_SLICE_X12Y110_ALUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_L_X10Y110_SLICE_X13Y110_DO5),
.I2(CLBLM_L_X10Y110_SLICE_X12Y110_AQ),
.I3(CLBLM_R_X7Y120_SLICE_X9Y120_DQ),
.I4(RIOB33_X105Y105_IOB_X1Y105_I),
.I5(CLBLM_R_X5Y114_SLICE_X7Y114_AQ),
.O5(CLBLM_L_X10Y110_SLICE_X12Y110_AO5),
.O6(CLBLM_L_X10Y110_SLICE_X12Y110_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y110_SLICE_X13Y110_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y110_SLICE_X13Y110_AO6),
.Q(CLBLM_L_X10Y110_SLICE_X13Y110_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y110_SLICE_X13Y110_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y110_SLICE_X13Y110_BO6),
.Q(CLBLM_L_X10Y110_SLICE_X13Y110_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000088800004ccc)
  ) CLBLM_L_X10Y110_SLICE_X13Y110_DLUT (
.I0(CLBLM_L_X10Y110_SLICE_X12Y110_AQ),
.I1(CLBLM_R_X11Y115_SLICE_X14Y115_AQ),
.I2(CLBLM_L_X10Y110_SLICE_X13Y110_BQ),
.I3(CLBLM_L_X10Y110_SLICE_X13Y110_AQ),
.I4(CLBLM_L_X10Y113_SLICE_X12Y113_DO6),
.I5(1'b1),
.O5(CLBLM_L_X10Y110_SLICE_X13Y110_DO5),
.O6(CLBLM_L_X10Y110_SLICE_X13Y110_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h00002000a0000000)
  ) CLBLM_L_X10Y110_SLICE_X13Y110_CLUT (
.I0(CLBLM_L_X10Y110_SLICE_X12Y110_AQ),
.I1(CLBLM_L_X10Y113_SLICE_X12Y113_DO6),
.I2(CLBLM_L_X10Y110_SLICE_X13Y110_BQ),
.I3(CLBLM_R_X11Y115_SLICE_X14Y115_AQ),
.I4(CLBLM_L_X10Y110_SLICE_X13Y110_AQ),
.I5(1'b1),
.O5(CLBLM_L_X10Y110_SLICE_X13Y110_CO5),
.O6(CLBLM_L_X10Y110_SLICE_X13Y110_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf000f000f066f000)
  ) CLBLM_L_X10Y110_SLICE_X13Y110_BLUT (
.I0(CLBLM_L_X10Y110_SLICE_X13Y110_DO6),
.I1(CLBLM_L_X10Y110_SLICE_X13Y110_BQ),
.I2(CLBLM_L_X10Y116_SLICE_X13Y116_AQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(RIOB33_X105Y105_IOB_X1Y105_I),
.I5(CLBLM_R_X7Y120_SLICE_X9Y120_DQ),
.O5(CLBLM_L_X10Y110_SLICE_X13Y110_BO5),
.O6(CLBLM_L_X10Y110_SLICE_X13Y110_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hddcc1100dccc1000)
  ) CLBLM_L_X10Y110_SLICE_X13Y110_ALUT (
.I0(CLBLM_R_X7Y120_SLICE_X9Y120_DQ),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(CLBLM_L_X10Y110_SLICE_X13Y110_AQ),
.I3(RIOB33_X105Y105_IOB_X1Y105_I),
.I4(CLBLM_L_X10Y112_SLICE_X12Y112_DQ),
.I5(CLBLM_L_X10Y110_SLICE_X13Y110_CO6),
.O5(CLBLM_L_X10Y110_SLICE_X13Y110_AO5),
.O6(CLBLM_L_X10Y110_SLICE_X13Y110_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h33cc35c533cc3aca)
  ) CLBLM_L_X10Y111_SLICE_X12Y111_DLUT (
.I0(CLBLM_L_X10Y112_SLICE_X12Y112_AO6),
.I1(CLBLM_L_X10Y122_SLICE_X13Y122_A5Q),
.I2(CLBLM_R_X5Y119_SLICE_X7Y119_CO6),
.I3(CLBLM_L_X10Y116_SLICE_X13Y116_CQ),
.I4(CLBLL_L_X2Y119_SLICE_X1Y119_BO6),
.I5(CLBLM_L_X10Y111_SLICE_X12Y111_BO6),
.O5(CLBLM_L_X10Y111_SLICE_X12Y111_DO5),
.O6(CLBLM_L_X10Y111_SLICE_X12Y111_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h1015101015101515)
  ) CLBLM_L_X10Y111_SLICE_X12Y111_CLUT (
.I0(CLBLM_L_X10Y111_SLICE_X13Y111_AQ),
.I1(CLBLM_R_X7Y115_SLICE_X9Y115_BQ),
.I2(CLBLM_R_X5Y111_SLICE_X7Y111_DO6),
.I3(CLBLM_L_X10Y111_SLICE_X12Y111_AO5),
.I4(CLBLM_L_X10Y111_SLICE_X12Y111_BO5),
.I5(CLBLM_L_X10Y117_SLICE_X12Y117_AQ),
.O5(CLBLM_L_X10Y111_SLICE_X12Y111_CO5),
.O6(CLBLM_L_X10Y111_SLICE_X12Y111_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h00ff08f70c0c0c0c)
  ) CLBLM_L_X10Y111_SLICE_X12Y111_BLUT (
.I0(CLBLM_L_X10Y112_SLICE_X13Y112_CQ),
.I1(CLBLL_L_X4Y110_SLICE_X5Y110_AQ),
.I2(CLBLM_L_X8Y110_SLICE_X10Y110_BQ),
.I3(CLBLM_L_X10Y115_SLICE_X12Y115_BQ),
.I4(CLBLM_R_X7Y110_SLICE_X8Y110_CQ),
.I5(1'b1),
.O5(CLBLM_L_X10Y111_SLICE_X12Y111_BO5),
.O6(CLBLM_L_X10Y111_SLICE_X12Y111_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0f0f0f87bbbbbbbb)
  ) CLBLM_L_X10Y111_SLICE_X12Y111_ALUT (
.I0(CLBLM_L_X10Y112_SLICE_X13Y112_CQ),
.I1(CLBLM_R_X7Y110_SLICE_X8Y110_CQ),
.I2(CLBLM_L_X10Y115_SLICE_X12Y115_AQ),
.I3(CLBLL_L_X4Y110_SLICE_X5Y110_AQ),
.I4(CLBLM_L_X8Y110_SLICE_X10Y110_BQ),
.I5(1'b1),
.O5(CLBLM_L_X10Y111_SLICE_X12Y111_AO5),
.O6(CLBLM_L_X10Y111_SLICE_X12Y111_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y111_SLICE_X13Y111_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y111_SLICE_X13Y111_AO6),
.Q(CLBLM_L_X10Y111_SLICE_X13Y111_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X10Y111_SLICE_X13Y111_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X10Y111_SLICE_X13Y111_DO5),
.O6(CLBLM_L_X10Y111_SLICE_X13Y111_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffff0fcccc9ccc)
  ) CLBLM_L_X10Y111_SLICE_X13Y111_CLUT (
.I0(CLBLM_L_X10Y112_SLICE_X13Y112_CQ),
.I1(CLBLM_L_X10Y117_SLICE_X12Y117_AQ),
.I2(CLBLL_L_X4Y110_SLICE_X5Y110_AQ),
.I3(CLBLM_R_X7Y110_SLICE_X8Y110_CQ),
.I4(CLBLM_L_X8Y110_SLICE_X10Y110_BQ),
.I5(1'b1),
.O5(CLBLM_L_X10Y111_SLICE_X13Y111_CO5),
.O6(CLBLM_L_X10Y111_SLICE_X13Y111_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000400010505050)
  ) CLBLM_L_X10Y111_SLICE_X13Y111_BLUT (
.I0(CLBLM_R_X5Y111_SLICE_X7Y111_DO6),
.I1(CLBLM_L_X10Y112_SLICE_X13Y112_CQ),
.I2(CLBLM_R_X7Y110_SLICE_X8Y110_CQ),
.I3(CLBLL_L_X4Y110_SLICE_X5Y110_AQ),
.I4(CLBLM_L_X8Y110_SLICE_X10Y110_BQ),
.I5(1'b1),
.O5(CLBLM_L_X10Y111_SLICE_X13Y111_BO5),
.O6(CLBLM_L_X10Y111_SLICE_X13Y111_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f0f0f044445555)
  ) CLBLM_L_X10Y111_SLICE_X13Y111_ALUT (
.I0(CLBLM_L_X10Y111_SLICE_X12Y111_CO6),
.I1(CLBLM_R_X7Y128_SLICE_X8Y128_AQ),
.I2(CLBLM_R_X7Y119_SLICE_X8Y119_D5Q),
.I3(1'b1),
.I4(RIOB33_X105Y141_IOB_X1Y142_I),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLM_L_X10Y111_SLICE_X13Y111_AO5),
.O6(CLBLM_L_X10Y111_SLICE_X13Y111_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y112_SLICE_X12Y112_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y112_SLICE_X12Y112_BO6),
.Q(CLBLM_L_X10Y112_SLICE_X12Y112_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y112_SLICE_X12Y112_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y112_SLICE_X12Y112_CO6),
.Q(CLBLM_L_X10Y112_SLICE_X12Y112_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y112_SLICE_X12Y112_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y112_SLICE_X12Y112_DO6),
.Q(CLBLM_L_X10Y112_SLICE_X12Y112_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'haa33aa00aa30aa00)
  ) CLBLM_L_X10Y112_SLICE_X12Y112_DLUT (
.I0(CLBLM_L_X10Y112_SLICE_X12Y112_BQ),
.I1(RIOB33_X105Y117_IOB_X1Y118_I),
.I2(CLBLM_L_X10Y112_SLICE_X12Y112_DQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLM_R_X3Y118_SLICE_X2Y118_AQ),
.I5(CLBLM_L_X10Y113_SLICE_X12Y113_BQ),
.O5(CLBLM_L_X10Y112_SLICE_X12Y112_DO5),
.O6(CLBLM_L_X10Y112_SLICE_X12Y112_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hf8fff8f0080f0800)
  ) CLBLM_L_X10Y112_SLICE_X12Y112_CLUT (
.I0(RIOB33_X105Y105_IOB_X1Y105_I),
.I1(CLBLM_L_X10Y112_SLICE_X12Y112_CQ),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLM_L_X10Y113_SLICE_X12Y113_DO6),
.I4(CLBLM_R_X11Y114_SLICE_X14Y114_AQ),
.I5(CLBLM_R_X5Y112_SLICE_X6Y112_AQ),
.O5(CLBLM_L_X10Y112_SLICE_X12Y112_CO5),
.O6(CLBLM_L_X10Y112_SLICE_X12Y112_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfff5faf0fef4faf0)
  ) CLBLM_L_X10Y112_SLICE_X12Y112_BLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_R_X3Y118_SLICE_X2Y118_AQ),
.I2(CLBLM_R_X7Y112_SLICE_X8Y112_DO6),
.I3(CLBLM_R_X3Y112_SLICE_X3Y112_B5Q),
.I4(CLBLM_L_X10Y112_SLICE_X12Y112_BQ),
.I5(RIOB33_X105Y117_IOB_X1Y118_I),
.O5(CLBLM_L_X10Y112_SLICE_X12Y112_BO5),
.O6(CLBLM_L_X10Y112_SLICE_X12Y112_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h10ef00ff05050505)
  ) CLBLM_L_X10Y112_SLICE_X12Y112_ALUT (
.I0(CLBLL_L_X4Y110_SLICE_X5Y110_AQ),
.I1(CLBLM_R_X7Y110_SLICE_X8Y110_CQ),
.I2(CLBLM_L_X8Y110_SLICE_X10Y110_BQ),
.I3(CLBLM_R_X11Y117_SLICE_X14Y117_BQ),
.I4(CLBLM_L_X10Y112_SLICE_X13Y112_CQ),
.I5(1'b1),
.O5(CLBLM_L_X10Y112_SLICE_X12Y112_AO5),
.O6(CLBLM_L_X10Y112_SLICE_X12Y112_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y112_SLICE_X13Y112_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y112_SLICE_X13Y112_AO6),
.Q(CLBLM_L_X10Y112_SLICE_X13Y112_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y112_SLICE_X13Y112_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y112_SLICE_X13Y112_BO6),
.Q(CLBLM_L_X10Y112_SLICE_X13Y112_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y112_SLICE_X13Y112_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y112_SLICE_X13Y112_CO6),
.Q(CLBLM_L_X10Y112_SLICE_X13Y112_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hdffddffdeffeeffe)
  ) CLBLM_L_X10Y112_SLICE_X13Y112_DLUT (
.I0(CLBLM_L_X8Y111_SLICE_X10Y111_AQ),
.I1(CLBLM_L_X8Y111_SLICE_X10Y111_DO6),
.I2(CLBLM_L_X10Y120_SLICE_X12Y120_BQ),
.I3(CLBLM_L_X10Y112_SLICE_X13Y112_BQ),
.I4(1'b1),
.I5(CLBLM_L_X12Y115_SLICE_X16Y115_CQ),
.O5(CLBLM_L_X10Y112_SLICE_X13Y112_DO5),
.O6(CLBLM_L_X10Y112_SLICE_X13Y112_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hab01aa00ae04aa00)
  ) CLBLM_L_X10Y112_SLICE_X13Y112_CLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_L_X10Y111_SLICE_X13Y111_BO5),
.I2(CLBLM_L_X8Y118_SLICE_X10Y118_DQ),
.I3(CLBLM_L_X12Y120_SLICE_X17Y120_BQ),
.I4(RIOB33_X105Y105_IOB_X1Y105_I),
.I5(CLBLM_L_X10Y112_SLICE_X13Y112_CQ),
.O5(CLBLM_L_X10Y112_SLICE_X13Y112_CO5),
.O6(CLBLM_L_X10Y112_SLICE_X13Y112_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hefafeaaa45054000)
  ) CLBLM_L_X10Y112_SLICE_X13Y112_BLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_L_X10Y112_SLICE_X13Y112_BQ),
.I2(CLBLM_L_X10Y113_SLICE_X12Y113_DO6),
.I3(RIOB33_X105Y105_IOB_X1Y105_I),
.I4(CLBLM_R_X11Y113_SLICE_X14Y113_AQ),
.I5(CLBLM_L_X8Y118_SLICE_X10Y118_DQ),
.O5(CLBLM_L_X10Y112_SLICE_X13Y112_BO5),
.O6(CLBLM_L_X10Y112_SLICE_X13Y112_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffa50ffffea40)
  ) CLBLM_L_X10Y112_SLICE_X13Y112_ALUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_R_X3Y118_SLICE_X2Y118_AQ),
.I2(CLBLM_L_X10Y112_SLICE_X13Y112_AQ),
.I3(CLBLM_R_X5Y114_SLICE_X6Y114_DQ),
.I4(CLBLM_R_X7Y112_SLICE_X8Y112_DO6),
.I5(RIOB33_X105Y117_IOB_X1Y118_I),
.O5(CLBLM_L_X10Y112_SLICE_X13Y112_AO5),
.O6(CLBLM_L_X10Y112_SLICE_X13Y112_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y113_SLICE_X12Y113_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y113_SLICE_X12Y113_BO6),
.Q(CLBLM_L_X10Y113_SLICE_X12Y113_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h00000000000000f0)
  ) CLBLM_L_X10Y113_SLICE_X12Y113_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(CLBLL_L_X2Y113_SLICE_X1Y113_AQ),
.I3(CLBLM_R_X3Y118_SLICE_X2Y118_AQ),
.I4(RIOB33_X105Y117_IOB_X1Y118_I),
.I5(CLBLM_R_X5Y110_SLICE_X7Y110_BQ),
.O5(CLBLM_L_X10Y113_SLICE_X12Y113_DO5),
.O6(CLBLM_L_X10Y113_SLICE_X12Y113_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0f0f0a0a0f0e0a0b)
  ) CLBLM_L_X10Y113_SLICE_X12Y113_CLUT (
.I0(CLBLM_L_X10Y114_SLICE_X13Y114_DQ),
.I1(CLBLM_L_X8Y110_SLICE_X10Y110_BQ),
.I2(CLBLM_R_X5Y111_SLICE_X7Y111_DO6),
.I3(CLBLL_L_X4Y110_SLICE_X5Y110_AQ),
.I4(CLBLM_L_X10Y116_SLICE_X13Y116_AO5),
.I5(CLBLM_L_X10Y111_SLICE_X12Y111_AO5),
.O5(CLBLM_L_X10Y113_SLICE_X12Y113_CO5),
.O6(CLBLM_L_X10Y113_SLICE_X12Y113_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'heca0ffa0ffa0eca0)
  ) CLBLM_L_X10Y113_SLICE_X12Y113_BLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_L_X10Y113_SLICE_X12Y113_BQ),
.I2(CLBLM_L_X10Y114_SLICE_X13Y114_DQ),
.I3(CLBLM_R_X11Y123_SLICE_X14Y123_CO6),
.I4(CLBLM_L_X8Y111_SLICE_X11Y111_AO6),
.I5(CLBLM_L_X10Y113_SLICE_X12Y113_CO6),
.O5(CLBLM_L_X10Y113_SLICE_X12Y113_BO5),
.O6(CLBLM_L_X10Y113_SLICE_X12Y113_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfeff0100ffcfffcf)
  ) CLBLM_L_X10Y113_SLICE_X12Y113_ALUT (
.I0(CLBLM_L_X10Y112_SLICE_X13Y112_CQ),
.I1(CLBLM_R_X7Y110_SLICE_X8Y110_CQ),
.I2(CLBLM_L_X8Y110_SLICE_X10Y110_BQ),
.I3(CLBLL_L_X4Y110_SLICE_X5Y110_AQ),
.I4(CLBLM_R_X7Y112_SLICE_X9Y112_CQ),
.I5(1'b1),
.O5(CLBLM_L_X10Y113_SLICE_X12Y113_AO5),
.O6(CLBLM_L_X10Y113_SLICE_X12Y113_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000001)
  ) CLBLM_L_X10Y113_SLICE_X13Y113_DLUT (
.I0(CLBLM_R_X11Y113_SLICE_X14Y113_AQ),
.I1(CLBLM_R_X11Y113_SLICE_X15Y113_BQ),
.I2(CLBLM_R_X11Y114_SLICE_X14Y114_AQ),
.I3(CLBLM_L_X8Y112_SLICE_X10Y112_AQ),
.I4(CLBLM_R_X11Y114_SLICE_X14Y114_BQ),
.I5(CLBLM_L_X10Y112_SLICE_X12Y112_CQ),
.O5(CLBLM_L_X10Y113_SLICE_X13Y113_DO5),
.O6(CLBLM_L_X10Y113_SLICE_X13Y113_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaaaaaaaaabaaaa)
  ) CLBLM_L_X10Y113_SLICE_X13Y113_CLUT (
.I0(CLBLM_L_X8Y114_SLICE_X11Y114_AQ),
.I1(CLBLM_L_X8Y113_SLICE_X11Y113_AQ),
.I2(CLBLM_R_X11Y113_SLICE_X15Y113_AQ),
.I3(CLBLM_R_X11Y113_SLICE_X14Y113_DO6),
.I4(CLBLM_L_X10Y113_SLICE_X13Y113_DO6),
.I5(CLBLM_L_X8Y112_SLICE_X10Y112_BQ),
.O5(CLBLM_L_X10Y113_SLICE_X13Y113_CO5),
.O6(CLBLM_L_X10Y113_SLICE_X13Y113_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0fff4fff0fff1fff)
  ) CLBLM_L_X10Y113_SLICE_X13Y113_BLUT (
.I0(CLBLM_L_X10Y112_SLICE_X13Y112_DO6),
.I1(CLBLM_R_X7Y111_SLICE_X9Y111_DO6),
.I2(CLBLM_L_X10Y110_SLICE_X13Y110_CO5),
.I3(CLBLM_L_X10Y113_SLICE_X12Y113_DO6),
.I4(CLBLM_L_X8Y113_SLICE_X10Y113_AO6),
.I5(CLBLM_L_X10Y113_SLICE_X13Y113_AO5),
.O5(CLBLM_L_X10Y113_SLICE_X13Y113_BO5),
.O6(CLBLM_L_X10Y113_SLICE_X13Y113_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h3faa0caa3f000c00)
  ) CLBLM_L_X10Y113_SLICE_X13Y113_ALUT (
.I0(CLBLM_R_X7Y111_SLICE_X9Y111_DO6),
.I1(CLBLM_L_X10Y114_SLICE_X13Y114_AQ),
.I2(CLBLM_L_X8Y114_SLICE_X11Y114_AQ),
.I3(CLBLM_L_X10Y110_SLICE_X13Y110_CO5),
.I4(CLBLM_L_X10Y113_SLICE_X13Y113_CO6),
.I5(1'b1),
.O5(CLBLM_L_X10Y113_SLICE_X13Y113_AO5),
.O6(CLBLM_L_X10Y113_SLICE_X13Y113_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y114_SLICE_X12Y114_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(LIOB33_X0Y77_IOB_X0Y77_I),
.D(CLBLM_R_X11Y114_SLICE_X14Y114_DQ),
.Q(CLBLM_L_X10Y114_SLICE_X12Y114_AQ),
.R(CLBLM_R_X11Y123_SLICE_X14Y123_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000001)
  ) CLBLM_L_X10Y114_SLICE_X12Y114_DLUT (
.I0(CLBLM_L_X10Y117_SLICE_X12Y117_AQ),
.I1(CLBLM_L_X8Y110_SLICE_X10Y110_AQ),
.I2(CLBLM_R_X11Y117_SLICE_X14Y117_BQ),
.I3(CLBLL_L_X4Y110_SLICE_X5Y110_BQ),
.I4(CLBLM_R_X7Y112_SLICE_X9Y112_CQ),
.I5(CLBLM_R_X5Y114_SLICE_X6Y114_DQ),
.O5(CLBLM_L_X10Y114_SLICE_X12Y114_DO5),
.O6(CLBLM_L_X10Y114_SLICE_X12Y114_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0505114405051111)
  ) CLBLM_L_X10Y114_SLICE_X12Y114_CLUT (
.I0(CLBLM_L_X10Y114_SLICE_X13Y114_CQ),
.I1(CLBLM_L_X10Y115_SLICE_X12Y115_AQ),
.I2(CLBLM_L_X10Y127_SLICE_X12Y127_AQ),
.I3(CLBLM_L_X10Y114_SLICE_X12Y114_AO5),
.I4(CLBLM_R_X5Y111_SLICE_X7Y111_DO6),
.I5(CLBLM_L_X10Y112_SLICE_X12Y112_AO5),
.O5(CLBLM_L_X10Y114_SLICE_X12Y114_CO5),
.O6(CLBLM_L_X10Y114_SLICE_X12Y114_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hccccfa00fa00fa00)
  ) CLBLM_L_X10Y114_SLICE_X12Y114_BLUT (
.I0(CLBLM_L_X8Y114_SLICE_X10Y114_DQ),
.I1(CLBLM_L_X10Y115_SLICE_X12Y115_BQ),
.I2(CLBLM_L_X8Y115_SLICE_X11Y115_C5Q),
.I3(RIOB33_X105Y121_IOB_X1Y121_I),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(1'b1),
.O5(CLBLM_L_X10Y114_SLICE_X12Y114_BO5),
.O6(CLBLM_L_X10Y114_SLICE_X12Y114_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h5559555533ff33ff)
  ) CLBLM_L_X10Y114_SLICE_X12Y114_ALUT (
.I0(CLBLM_L_X8Y110_SLICE_X10Y110_AQ),
.I1(CLBLM_R_X7Y110_SLICE_X8Y110_CQ),
.I2(CLBLL_L_X4Y110_SLICE_X5Y110_AQ),
.I3(CLBLM_L_X10Y112_SLICE_X13Y112_CQ),
.I4(CLBLM_L_X8Y110_SLICE_X10Y110_BQ),
.I5(1'b1),
.O5(CLBLM_L_X10Y114_SLICE_X12Y114_AO5),
.O6(CLBLM_L_X10Y114_SLICE_X12Y114_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y114_SLICE_X13Y114_A5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y114_SLICE_X13Y114_BO6),
.Q(CLBLM_L_X10Y114_SLICE_X13Y114_A5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y114_SLICE_X13Y114_D5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y114_SLICE_X13Y114_DO5),
.Q(CLBLM_L_X10Y114_SLICE_X13Y114_D5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y114_SLICE_X13Y114_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y114_SLICE_X13Y114_AO6),
.Q(CLBLM_L_X10Y114_SLICE_X13Y114_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y114_SLICE_X13Y114_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y114_SLICE_X13Y114_CO6),
.Q(CLBLM_L_X10Y114_SLICE_X13Y114_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y114_SLICE_X13Y114_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y114_SLICE_X13Y114_DO6),
.Q(CLBLM_L_X10Y114_SLICE_X13Y114_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hbb88bb88fcfc3030)
  ) CLBLM_L_X10Y114_SLICE_X13Y114_DLUT (
.I0(CLBLM_R_X7Y110_SLICE_X8Y110_CQ),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(CLBLM_R_X11Y120_SLICE_X15Y120_CQ),
.I3(CLBLM_L_X10Y114_SLICE_X13Y114_A5Q),
.I4(CLBLM_L_X10Y113_SLICE_X12Y113_BQ),
.I5(1'b1),
.O5(CLBLM_L_X10Y114_SLICE_X13Y114_DO5),
.O6(CLBLM_L_X10Y114_SLICE_X13Y114_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'haa33aa00aa33aa33)
  ) CLBLM_L_X10Y114_SLICE_X13Y114_CLUT (
.I0(CLBLM_R_X3Y113_SLICE_X3Y113_AQ),
.I1(CLBLM_L_X10Y114_SLICE_X12Y114_CO6),
.I2(1'b1),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLM_R_X7Y128_SLICE_X8Y128_AQ),
.I5(RIOB33_X105Y141_IOB_X1Y142_I),
.O5(CLBLM_L_X10Y114_SLICE_X13Y114_CO5),
.O6(CLBLM_L_X10Y114_SLICE_X13Y114_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfecc3200fa00fa00)
  ) CLBLM_L_X10Y114_SLICE_X13Y114_BLUT (
.I0(CLBLL_L_X4Y114_SLICE_X5Y114_AQ),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(CLBLM_L_X10Y112_SLICE_X13Y112_AQ),
.I3(RIOB33_X105Y121_IOB_X1Y121_I),
.I4(CLBLM_R_X11Y116_SLICE_X14Y116_DQ),
.I5(1'b1),
.O5(CLBLM_L_X10Y114_SLICE_X13Y114_BO5),
.O6(CLBLM_L_X10Y114_SLICE_X13Y114_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfd31ec20dd11cc00)
  ) CLBLM_L_X10Y114_SLICE_X13Y114_ALUT (
.I0(CLBLM_L_X10Y113_SLICE_X12Y113_DO6),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(CLBLM_L_X10Y114_SLICE_X13Y114_AQ),
.I3(CLBLM_R_X7Y112_SLICE_X8Y112_BQ),
.I4(CLBLM_L_X8Y114_SLICE_X11Y114_AQ),
.I5(RIOB33_X105Y105_IOB_X1Y105_I),
.O5(CLBLM_L_X10Y114_SLICE_X13Y114_AO5),
.O6(CLBLM_L_X10Y114_SLICE_X13Y114_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y115_SLICE_X12Y115_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y115_SLICE_X12Y115_AO6),
.Q(CLBLM_L_X10Y115_SLICE_X12Y115_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y115_SLICE_X12Y115_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y115_SLICE_X12Y115_BO6),
.Q(CLBLM_L_X10Y115_SLICE_X12Y115_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y115_SLICE_X12Y115_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y115_SLICE_X12Y115_CO6),
.Q(CLBLM_L_X10Y115_SLICE_X12Y115_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y115_SLICE_X12Y115_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y115_SLICE_X12Y115_DO6),
.Q(CLBLM_L_X10Y115_SLICE_X12Y115_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff333000003330)
  ) CLBLM_L_X10Y115_SLICE_X12Y115_DLUT (
.I0(1'b1),
.I1(CLBLM_R_X5Y111_SLICE_X7Y111_DO6),
.I2(CLBLM_L_X10Y115_SLICE_X12Y115_DQ),
.I3(CLBLM_L_X10Y110_SLICE_X12Y110_BQ),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(CLBLM_R_X7Y119_SLICE_X8Y119_BQ),
.O5(CLBLM_L_X10Y115_SLICE_X12Y115_DO5),
.O6(CLBLM_L_X10Y115_SLICE_X12Y115_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaa0000faea5040)
  ) CLBLM_L_X10Y115_SLICE_X12Y115_CLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_L_X10Y115_SLICE_X12Y115_CQ),
.I2(RIOB33_X105Y105_IOB_X1Y105_I),
.I3(CLBLM_R_X7Y115_SLICE_X9Y115_DQ),
.I4(CLBLM_L_X10Y117_SLICE_X13Y117_DQ),
.I5(CLBLM_R_X7Y114_SLICE_X8Y114_BQ),
.O5(CLBLM_L_X10Y115_SLICE_X12Y115_CO5),
.O6(CLBLM_L_X10Y115_SLICE_X12Y115_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hff55ff4400550044)
  ) CLBLM_L_X10Y115_SLICE_X12Y115_BLUT (
.I0(CLBLM_R_X5Y111_SLICE_X7Y111_DO6),
.I1(CLBLM_L_X10Y115_SLICE_X12Y115_BQ),
.I2(1'b1),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLM_L_X10Y117_SLICE_X12Y117_AQ),
.I5(CLBLM_L_X8Y121_SLICE_X10Y121_CQ),
.O5(CLBLM_L_X10Y115_SLICE_X12Y115_BO5),
.O6(CLBLM_L_X10Y115_SLICE_X12Y115_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaa0000fefe5454)
  ) CLBLM_L_X10Y115_SLICE_X12Y115_ALUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_L_X10Y115_SLICE_X12Y115_AQ),
.I2(CLBLM_L_X8Y117_SLICE_X11Y117_BQ),
.I3(1'b1),
.I4(CLBLM_L_X8Y123_SLICE_X11Y123_AQ),
.I5(CLBLM_R_X5Y111_SLICE_X7Y111_DO6),
.O5(CLBLM_L_X10Y115_SLICE_X12Y115_AO5),
.O6(CLBLM_L_X10Y115_SLICE_X12Y115_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffffffffeeee)
  ) CLBLM_L_X10Y115_SLICE_X13Y115_DLUT (
.I0(CLBLM_R_X11Y115_SLICE_X15Y115_BQ),
.I1(CLBLM_R_X11Y115_SLICE_X15Y115_DQ),
.I2(1'b1),
.I3(1'b1),
.I4(CLBLM_L_X10Y115_SLICE_X12Y115_AQ),
.I5(CLBLM_L_X10Y119_SLICE_X12Y119_BQ),
.O5(CLBLM_L_X10Y115_SLICE_X13Y115_DO5),
.O6(CLBLM_L_X10Y115_SLICE_X13Y115_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000001010)
  ) CLBLM_L_X10Y115_SLICE_X13Y115_CLUT (
.I0(CLBLM_L_X8Y117_SLICE_X11Y117_BQ),
.I1(CLBLM_L_X10Y117_SLICE_X13Y117_BQ),
.I2(CLBLM_L_X10Y114_SLICE_X12Y114_DO6),
.I3(1'b1),
.I4(CLBLM_L_X10Y115_SLICE_X13Y115_DO6),
.I5(CLBLM_L_X10Y115_SLICE_X12Y115_BQ),
.O5(CLBLM_L_X10Y115_SLICE_X13Y115_CO5),
.O6(CLBLM_L_X10Y115_SLICE_X13Y115_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0001111044455554)
  ) CLBLM_L_X10Y115_SLICE_X13Y115_BLUT (
.I0(CLBLM_R_X11Y115_SLICE_X14Y115_BQ),
.I1(CLBLM_R_X5Y111_SLICE_X7Y111_DO6),
.I2(CLBLM_L_X10Y111_SLICE_X13Y111_CO6),
.I3(CLBLM_L_X10Y112_SLICE_X13Y112_CQ),
.I4(CLBLM_R_X7Y112_SLICE_X9Y112_CQ),
.I5(CLBLM_R_X7Y115_SLICE_X9Y115_B5Q),
.O5(CLBLM_L_X10Y115_SLICE_X13Y115_BO5),
.O6(CLBLM_L_X10Y115_SLICE_X13Y115_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0110001123322233)
  ) CLBLM_L_X10Y115_SLICE_X13Y115_ALUT (
.I0(CLBLM_R_X5Y111_SLICE_X7Y111_DO6),
.I1(CLBLM_R_X11Y115_SLICE_X14Y115_CQ),
.I2(CLBLM_L_X10Y111_SLICE_X13Y111_CO6),
.I3(CLBLM_L_X10Y115_SLICE_X12Y115_BQ),
.I4(CLBLM_L_X10Y112_SLICE_X13Y112_CQ),
.I5(CLBLM_L_X10Y116_SLICE_X13Y116_CQ),
.O5(CLBLM_L_X10Y115_SLICE_X13Y115_AO5),
.O6(CLBLM_L_X10Y115_SLICE_X13Y115_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y116_SLICE_X12Y116_A5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y114_SLICE_X12Y114_BO6),
.Q(CLBLM_L_X10Y116_SLICE_X12Y116_A5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y116_SLICE_X12Y116_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y116_SLICE_X12Y116_AO6),
.Q(CLBLM_L_X10Y116_SLICE_X12Y116_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y116_SLICE_X12Y116_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y116_SLICE_X12Y116_BO6),
.Q(CLBLM_L_X10Y116_SLICE_X12Y116_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y116_SLICE_X12Y116_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y116_SLICE_X12Y116_CO6),
.Q(CLBLM_L_X10Y116_SLICE_X12Y116_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000030000000100)
  ) CLBLM_L_X10Y116_SLICE_X12Y116_DLUT (
.I0(CLBLM_L_X10Y116_SLICE_X12Y116_BQ),
.I1(CLBLM_L_X8Y116_SLICE_X11Y116_A5Q),
.I2(CLBLM_R_X11Y116_SLICE_X14Y116_CQ),
.I3(CLBLM_L_X8Y119_SLICE_X10Y119_BQ),
.I4(CLBLM_L_X10Y116_SLICE_X12Y116_AQ),
.I5(1'b1),
.O5(CLBLM_L_X10Y116_SLICE_X12Y116_DO5),
.O6(CLBLM_L_X10Y116_SLICE_X12Y116_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h888888888d8dd8d8)
  ) CLBLM_L_X10Y116_SLICE_X12Y116_CLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_L_X10Y116_SLICE_X13Y116_BQ),
.I2(CLBLM_L_X10Y114_SLICE_X12Y114_BO5),
.I3(1'b1),
.I4(CLBLM_L_X10Y119_SLICE_X12Y119_CQ),
.I5(RIOB33_X105Y105_IOB_X1Y105_I),
.O5(CLBLM_L_X10Y116_SLICE_X12Y116_CO5),
.O6(CLBLM_L_X10Y116_SLICE_X12Y116_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f0fffff0f06666)
  ) CLBLM_L_X10Y116_SLICE_X12Y116_BLUT (
.I0(CLBLM_L_X10Y116_SLICE_X12Y116_DO6),
.I1(CLBLM_L_X10Y116_SLICE_X12Y116_BQ),
.I2(CLBLL_L_X4Y116_SLICE_X4Y116_DQ),
.I3(1'b1),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(CLBLM_R_X11Y119_SLICE_X14Y119_AO6),
.O5(CLBLM_L_X10Y116_SLICE_X12Y116_BO5),
.O6(CLBLM_L_X10Y116_SLICE_X12Y116_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h88888888888b88b8)
  ) CLBLM_L_X10Y116_SLICE_X12Y116_ALUT (
.I0(CLBLM_L_X10Y114_SLICE_X12Y114_AQ),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(CLBLM_L_X10Y116_SLICE_X12Y116_AQ),
.I3(CLBLM_L_X10Y116_SLICE_X12Y116_DO5),
.I4(CLBLM_L_X8Y116_SLICE_X11Y116_CO5),
.I5(CLBLM_R_X11Y119_SLICE_X14Y119_AO6),
.O5(CLBLM_L_X10Y116_SLICE_X12Y116_AO5),
.O6(CLBLM_L_X10Y116_SLICE_X12Y116_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y116_SLICE_X13Y116_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y116_SLICE_X14Y116_BO6),
.Q(CLBLM_L_X10Y116_SLICE_X13Y116_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y116_SLICE_X13Y116_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y116_SLICE_X13Y116_BO6),
.Q(CLBLM_L_X10Y116_SLICE_X13Y116_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y116_SLICE_X13Y116_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y116_SLICE_X13Y116_CO6),
.Q(CLBLM_L_X10Y116_SLICE_X13Y116_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y116_SLICE_X13Y116_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y116_SLICE_X13Y116_DO6),
.Q(CLBLM_L_X10Y116_SLICE_X13Y116_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'haa00fe54aa00fe54)
  ) CLBLM_L_X10Y116_SLICE_X13Y116_DLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_L_X10Y117_SLICE_X13Y117_AQ),
.I2(CLBLM_L_X10Y116_SLICE_X13Y116_DQ),
.I3(CLBLM_R_X7Y117_SLICE_X8Y117_A5Q),
.I4(CLBLM_R_X5Y111_SLICE_X7Y111_DO6),
.I5(1'b1),
.O5(CLBLM_L_X10Y116_SLICE_X13Y116_DO5),
.O6(CLBLM_L_X10Y116_SLICE_X13Y116_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaaf0f000440044)
  ) CLBLM_L_X10Y116_SLICE_X13Y116_CLUT (
.I0(CLBLM_L_X10Y116_SLICE_X12Y116_AQ),
.I1(CLBLM_L_X8Y119_SLICE_X10Y119_BQ),
.I2(CLBLM_L_X10Y116_SLICE_X13Y116_BQ),
.I3(CLBLM_L_X8Y116_SLICE_X11Y116_A5Q),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(1'b1),
.O5(CLBLM_L_X10Y116_SLICE_X13Y116_CO5),
.O6(CLBLM_L_X10Y116_SLICE_X13Y116_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hccccfa0005ff05ff)
  ) CLBLM_L_X10Y116_SLICE_X13Y116_BLUT (
.I0(CLBLM_L_X10Y117_SLICE_X13Y117_DQ),
.I1(CLBLM_L_X10Y112_SLICE_X13Y112_BQ),
.I2(CLBLM_R_X5Y119_SLICE_X6Y119_BQ),
.I3(RIOB33_X105Y121_IOB_X1Y121_I),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(1'b1),
.O5(CLBLM_L_X10Y116_SLICE_X13Y116_BO5),
.O6(CLBLM_L_X10Y116_SLICE_X13Y116_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hcacacaca3333ffcc)
  ) CLBLM_L_X10Y116_SLICE_X13Y116_ALUT (
.I0(RIOB33_X105Y103_IOB_X1Y104_I),
.I1(CLBLM_L_X10Y117_SLICE_X13Y117_AQ),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLM_L_X10Y115_SLICE_X13Y115_CO6),
.I4(CLBLM_L_X10Y116_SLICE_X13Y116_DQ),
.I5(1'b1),
.O5(CLBLM_L_X10Y116_SLICE_X13Y116_AO5),
.O6(CLBLM_L_X10Y116_SLICE_X13Y116_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y117_SLICE_X12Y117_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y117_SLICE_X12Y117_AO6),
.Q(CLBLM_L_X10Y117_SLICE_X12Y117_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y117_SLICE_X12Y117_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y117_SLICE_X12Y117_BO6),
.Q(CLBLM_L_X10Y117_SLICE_X12Y117_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X10Y117_SLICE_X12Y117_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X10Y117_SLICE_X12Y117_DO5),
.O6(CLBLM_L_X10Y117_SLICE_X12Y117_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000033330f5a)
  ) CLBLM_L_X10Y117_SLICE_X12Y117_CLUT (
.I0(CLBLM_L_X10Y112_SLICE_X13Y112_CQ),
.I1(CLBLM_L_X10Y118_SLICE_X12Y118_BQ),
.I2(CLBLL_L_X4Y110_SLICE_X5Y110_BQ),
.I3(CLBLM_L_X10Y113_SLICE_X12Y113_AO5),
.I4(CLBLM_R_X5Y111_SLICE_X7Y111_DO6),
.I5(CLBLM_L_X10Y118_SLICE_X12Y118_AQ),
.O5(CLBLM_L_X10Y117_SLICE_X12Y117_CO5),
.O6(CLBLM_L_X10Y117_SLICE_X12Y117_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'ha0a0acacafa0afa0)
  ) CLBLM_L_X10Y117_SLICE_X12Y117_BLUT (
.I0(CLBLL_L_X2Y117_SLICE_X0Y117_AQ),
.I1(CLBLM_L_X10Y117_SLICE_X12Y117_BQ),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLM_R_X11Y117_SLICE_X15Y117_AQ),
.I4(CLBLM_R_X11Y119_SLICE_X14Y119_AO6),
.I5(CLBLM_L_X12Y119_SLICE_X17Y119_AO5),
.O5(CLBLM_L_X10Y117_SLICE_X12Y117_BO5),
.O6(CLBLM_L_X10Y117_SLICE_X12Y117_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hcc00cc00ccffccf0)
  ) CLBLM_L_X10Y117_SLICE_X12Y117_ALUT (
.I0(1'b1),
.I1(CLBLM_R_X11Y116_SLICE_X15Y116_AQ),
.I2(CLBLM_L_X10Y117_SLICE_X12Y117_AQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLM_R_X7Y112_SLICE_X9Y112_CQ),
.I5(CLBLM_R_X5Y111_SLICE_X7Y111_DO6),
.O5(CLBLM_L_X10Y117_SLICE_X12Y117_AO5),
.O6(CLBLM_L_X10Y117_SLICE_X12Y117_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y117_SLICE_X13Y117_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y117_SLICE_X13Y117_AO6),
.Q(CLBLM_L_X10Y117_SLICE_X13Y117_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y117_SLICE_X13Y117_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y117_SLICE_X13Y117_BO6),
.Q(CLBLM_L_X10Y117_SLICE_X13Y117_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y117_SLICE_X13Y117_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y117_SLICE_X13Y117_CO6),
.Q(CLBLM_L_X10Y117_SLICE_X13Y117_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y117_SLICE_X13Y117_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y117_SLICE_X13Y117_DO6),
.Q(CLBLM_L_X10Y117_SLICE_X13Y117_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffffffa50ea40)
  ) CLBLM_L_X10Y117_SLICE_X13Y117_DLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(RIOB33_X105Y117_IOB_X1Y118_I),
.I2(CLBLM_L_X10Y117_SLICE_X13Y117_DQ),
.I3(CLBLM_R_X13Y119_SLICE_X18Y119_AQ),
.I4(CLBLM_R_X3Y118_SLICE_X2Y118_AQ),
.I5(CLBLM_R_X7Y113_SLICE_X8Y113_CO6),
.O5(CLBLM_L_X10Y117_SLICE_X13Y117_DO5),
.O6(CLBLM_L_X10Y117_SLICE_X13Y117_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hf5f5e4e4a0f5a0e4)
  ) CLBLM_L_X10Y117_SLICE_X13Y117_CLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_L_X10Y117_SLICE_X13Y117_CQ),
.I2(CLBLM_L_X10Y116_SLICE_X13Y116_DQ),
.I3(CLBLM_R_X7Y119_SLICE_X8Y119_D5Q),
.I4(CLBLM_R_X3Y112_SLICE_X3Y112_AQ),
.I5(CLBLM_L_X10Y113_SLICE_X13Y113_BO6),
.O5(CLBLM_L_X10Y117_SLICE_X13Y117_CO5),
.O6(CLBLM_L_X10Y117_SLICE_X13Y117_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hff000f0fff000c0c)
  ) CLBLM_L_X10Y117_SLICE_X13Y117_BLUT (
.I0(1'b1),
.I1(CLBLM_L_X10Y117_SLICE_X13Y117_BQ),
.I2(CLBLM_R_X5Y119_SLICE_X7Y119_AO6),
.I3(CLBLM_R_X11Y118_SLICE_X15Y118_BQ),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(CLBLM_R_X11Y115_SLICE_X15Y115_BQ),
.O5(CLBLM_L_X10Y117_SLICE_X13Y117_BO5),
.O6(CLBLM_L_X10Y117_SLICE_X13Y117_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'haa00aafcaa00aafc)
  ) CLBLM_L_X10Y117_SLICE_X13Y117_ALUT (
.I0(CLBLM_L_X10Y119_SLICE_X12Y119_CQ),
.I1(CLBLM_L_X10Y119_SLICE_X12Y119_BQ),
.I2(CLBLM_L_X10Y117_SLICE_X13Y117_AQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLM_R_X5Y119_SLICE_X7Y119_AO6),
.I5(1'b1),
.O5(CLBLM_L_X10Y117_SLICE_X13Y117_AO5),
.O6(CLBLM_L_X10Y117_SLICE_X13Y117_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y118_SLICE_X12Y118_B5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y118_SLICE_X12Y118_BO5),
.Q(CLBLM_L_X10Y118_SLICE_X12Y118_B5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y118_SLICE_X12Y118_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y118_SLICE_X12Y118_AO6),
.Q(CLBLM_L_X10Y118_SLICE_X12Y118_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y118_SLICE_X12Y118_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y118_SLICE_X12Y118_BO6),
.Q(CLBLM_L_X10Y118_SLICE_X12Y118_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffffffffff0ff)
  ) CLBLM_L_X10Y118_SLICE_X12Y118_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(CLBLM_L_X8Y119_SLICE_X11Y119_BQ),
.I3(CLBLM_L_X10Y118_SLICE_X13Y118_CQ),
.I4(CLBLM_L_X10Y119_SLICE_X12Y119_CQ),
.I5(CLBLM_L_X10Y116_SLICE_X12Y116_CQ),
.O5(CLBLM_L_X10Y118_SLICE_X12Y118_DO5),
.O6(CLBLM_L_X10Y118_SLICE_X12Y118_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000400000000)
  ) CLBLM_L_X10Y118_SLICE_X12Y118_CLUT (
.I0(CLBLM_R_X7Y119_SLICE_X8Y119_BQ),
.I1(CLBLM_L_X10Y121_SLICE_X12Y121_DO6),
.I2(CLBLM_L_X10Y119_SLICE_X12Y119_DO6),
.I3(CLBLL_L_X4Y110_SLICE_X4Y110_CQ),
.I4(CLBLM_L_X10Y118_SLICE_X12Y118_DO6),
.I5(CLBLM_R_X7Y119_SLICE_X9Y119_BQ),
.O5(CLBLM_L_X10Y118_SLICE_X12Y118_CO5),
.O6(CLBLM_L_X10Y118_SLICE_X12Y118_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf3f3c0c0eeeeaaaa)
  ) CLBLM_L_X10Y118_SLICE_X12Y118_BLUT (
.I0(CLBLM_L_X10Y123_SLICE_X13Y123_BO6),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(CLBLM_R_X5Y110_SLICE_X7Y110_BQ),
.I3(1'b1),
.I4(CLBLM_L_X10Y116_SLICE_X12Y116_A5Q),
.I5(1'b1),
.O5(CLBLM_L_X10Y118_SLICE_X12Y118_BO5),
.O6(CLBLM_L_X10Y118_SLICE_X12Y118_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hf3f3f0f303030003)
  ) CLBLM_L_X10Y118_SLICE_X12Y118_ALUT (
.I0(1'b1),
.I1(CLBLM_L_X10Y117_SLICE_X12Y117_CO6),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(RIOB33_X105Y141_IOB_X1Y142_I),
.I4(CLBLM_R_X7Y128_SLICE_X8Y128_AQ),
.I5(CLBLM_L_X8Y119_SLICE_X11Y119_CQ),
.O5(CLBLM_L_X10Y118_SLICE_X12Y118_AO5),
.O6(CLBLM_L_X10Y118_SLICE_X12Y118_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y118_SLICE_X13Y118_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y118_SLICE_X13Y118_AO6),
.Q(CLBLM_L_X10Y118_SLICE_X13Y118_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y118_SLICE_X13Y118_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y118_SLICE_X13Y118_BO6),
.Q(CLBLM_L_X10Y118_SLICE_X13Y118_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y118_SLICE_X13Y118_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y118_SLICE_X13Y118_CO6),
.Q(CLBLM_L_X10Y118_SLICE_X13Y118_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffffffdffffff)
  ) CLBLM_L_X10Y118_SLICE_X13Y118_DLUT (
.I0(CLBLM_L_X10Y115_SLICE_X13Y115_CO6),
.I1(CLBLM_R_X11Y113_SLICE_X15Y113_CO6),
.I2(CLBLM_R_X7Y118_SLICE_X8Y118_BQ),
.I3(CLBLM_R_X7Y123_SLICE_X9Y123_CO6),
.I4(CLBLM_R_X11Y119_SLICE_X14Y119_BO5),
.I5(CLBLM_L_X10Y113_SLICE_X13Y113_CO6),
.O5(CLBLM_L_X10Y118_SLICE_X13Y118_DO5),
.O6(CLBLM_L_X10Y118_SLICE_X13Y118_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'haaebaaeb00410041)
  ) CLBLM_L_X10Y118_SLICE_X13Y118_CLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLL_L_X4Y110_SLICE_X4Y110_CQ),
.I2(CLBLM_L_X10Y116_SLICE_X13Y116_BO5),
.I3(RIOB33_X105Y105_IOB_X1Y105_I),
.I4(1'b1),
.I5(CLBLM_L_X8Y122_SLICE_X11Y122_AQ),
.O5(CLBLM_L_X10Y118_SLICE_X13Y118_CO5),
.O6(CLBLM_L_X10Y118_SLICE_X13Y118_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf5f0fdf805000d08)
  ) CLBLM_L_X10Y118_SLICE_X13Y118_BLUT (
.I0(CLBLM_L_X12Y119_SLICE_X17Y119_AO5),
.I1(CLBLM_L_X10Y118_SLICE_X13Y118_BQ),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLM_L_X10Y117_SLICE_X12Y117_BQ),
.I4(CLBLM_R_X11Y119_SLICE_X14Y119_AO6),
.I5(CLBLM_R_X7Y117_SLICE_X8Y117_CQ),
.O5(CLBLM_L_X10Y118_SLICE_X13Y118_BO5),
.O6(CLBLM_L_X10Y118_SLICE_X13Y118_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hbb11fb51aa00ea40)
  ) CLBLM_L_X10Y118_SLICE_X13Y118_ALUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_L_X12Y119_SLICE_X17Y119_AO5),
.I2(CLBLM_L_X10Y118_SLICE_X13Y118_AQ),
.I3(CLBLM_L_X8Y114_SLICE_X11Y114_BQ),
.I4(CLBLM_R_X11Y119_SLICE_X14Y119_AO6),
.I5(CLBLM_L_X10Y120_SLICE_X12Y120_CQ),
.O5(CLBLM_L_X10Y118_SLICE_X13Y118_AO5),
.O6(CLBLM_L_X10Y118_SLICE_X13Y118_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y119_SLICE_X12Y119_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y119_SLICE_X12Y119_AO6),
.Q(CLBLM_L_X10Y119_SLICE_X12Y119_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y119_SLICE_X12Y119_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y119_SLICE_X12Y119_BO6),
.Q(CLBLM_L_X10Y119_SLICE_X12Y119_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y119_SLICE_X12Y119_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y119_SLICE_X12Y119_CO6),
.Q(CLBLM_L_X10Y119_SLICE_X12Y119_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffffffeffffff)
  ) CLBLM_L_X10Y119_SLICE_X12Y119_DLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(RIOB33_X105Y105_IOB_X1Y105_I),
.I2(RIOB33_X105Y121_IOB_X1Y121_I),
.I3(CLBLM_L_X8Y119_SLICE_X11Y119_CQ),
.I4(CLBLM_R_X7Y114_SLICE_X8Y114_BQ),
.I5(CLBLM_R_X13Y119_SLICE_X18Y119_BQ),
.O5(CLBLM_L_X10Y119_SLICE_X12Y119_DO5),
.O6(CLBLM_L_X10Y119_SLICE_X12Y119_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hc0d1c0d1c0e2c0e2)
  ) CLBLM_L_X10Y119_SLICE_X12Y119_CLUT (
.I0(CLBLM_L_X8Y119_SLICE_X11Y119_BQ),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(CLBLM_R_X7Y114_SLICE_X8Y114_BQ),
.I3(RIOB33_X105Y105_IOB_X1Y105_I),
.I4(1'b1),
.I5(CLBLM_L_X8Y119_SLICE_X10Y119_DO5),
.O5(CLBLM_L_X10Y119_SLICE_X12Y119_CO5),
.O6(CLBLM_L_X10Y119_SLICE_X12Y119_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'ha0a0afafa0a0acac)
  ) CLBLM_L_X10Y119_SLICE_X12Y119_BLUT (
.I0(CLBLM_L_X8Y120_SLICE_X11Y120_BQ),
.I1(CLBLM_L_X10Y119_SLICE_X12Y119_BQ),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(1'b1),
.I4(CLBLM_R_X5Y119_SLICE_X7Y119_AO6),
.I5(CLBLM_L_X10Y117_SLICE_X13Y117_BQ),
.O5(CLBLM_L_X10Y119_SLICE_X12Y119_BO5),
.O6(CLBLM_L_X10Y119_SLICE_X12Y119_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hdddddd88d8d8d888)
  ) CLBLM_L_X10Y119_SLICE_X12Y119_ALUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_L_X10Y119_SLICE_X12Y119_BQ),
.I2(CLBLM_L_X10Y119_SLICE_X12Y119_AQ),
.I3(CLBLM_R_X3Y118_SLICE_X2Y118_AQ),
.I4(RIOB33_X105Y117_IOB_X1Y118_I),
.I5(CLBLM_R_X5Y115_SLICE_X7Y115_DO6),
.O5(CLBLM_L_X10Y119_SLICE_X12Y119_AO5),
.O6(CLBLM_L_X10Y119_SLICE_X12Y119_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y119_SLICE_X13Y119_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y119_SLICE_X13Y119_AO6),
.Q(CLBLM_L_X10Y119_SLICE_X13Y119_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y119_SLICE_X13Y119_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y119_SLICE_X13Y119_BO6),
.Q(CLBLM_L_X10Y119_SLICE_X13Y119_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y119_SLICE_X13Y119_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y119_SLICE_X13Y119_CO6),
.Q(CLBLM_L_X10Y119_SLICE_X13Y119_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y119_SLICE_X13Y119_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y119_SLICE_X13Y119_DO6),
.Q(CLBLM_L_X10Y119_SLICE_X13Y119_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hab01ba10ab01ba10)
  ) CLBLM_L_X10Y119_SLICE_X13Y119_DLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(RIOB33_X105Y105_IOB_X1Y105_I),
.I2(CLBLM_L_X10Y114_SLICE_X13Y114_BO5),
.I3(CLBLM_L_X10Y119_SLICE_X13Y119_BQ),
.I4(CLBLL_L_X4Y117_SLICE_X5Y117_DQ),
.I5(1'b1),
.O5(CLBLM_L_X10Y119_SLICE_X13Y119_DO5),
.O6(CLBLM_L_X10Y119_SLICE_X13Y119_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaaf0f0aaaa5040)
  ) CLBLM_L_X10Y119_SLICE_X13Y119_CLUT (
.I0(CLBLM_R_X13Y119_SLICE_X18Y119_CQ),
.I1(CLBLM_L_X10Y119_SLICE_X13Y119_AQ),
.I2(CLBLM_L_X10Y119_SLICE_X13Y119_BQ),
.I3(CLBLM_R_X11Y118_SLICE_X14Y118_BQ),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(CLBLM_R_X11Y119_SLICE_X15Y119_CQ),
.O5(CLBLM_L_X10Y119_SLICE_X13Y119_CO5),
.O6(CLBLM_L_X10Y119_SLICE_X13Y119_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffc0f0cfffc0f0c)
  ) CLBLM_L_X10Y119_SLICE_X13Y119_BLUT (
.I0(1'b1),
.I1(CLBLM_L_X8Y119_SLICE_X10Y119_BQ),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLM_L_X12Y120_SLICE_X17Y120_CO6),
.I4(CLBLM_R_X7Y113_SLICE_X9Y113_A5Q),
.I5(1'b1),
.O5(CLBLM_L_X10Y119_SLICE_X13Y119_BO5),
.O6(CLBLM_L_X10Y119_SLICE_X13Y119_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hc5c5c5c0c0c0c5c0)
  ) CLBLM_L_X10Y119_SLICE_X13Y119_ALUT (
.I0(RIOB33_X105Y121_IOB_X1Y121_I),
.I1(CLBLM_R_X7Y120_SLICE_X9Y120_D5Q),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLM_L_X10Y119_SLICE_X13Y119_AQ),
.I4(CLBLM_L_X12Y120_SLICE_X16Y120_AO6),
.I5(CLBLM_R_X11Y118_SLICE_X14Y118_BQ),
.O5(CLBLM_L_X10Y119_SLICE_X13Y119_AO5),
.O6(CLBLM_L_X10Y119_SLICE_X13Y119_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y120_SLICE_X12Y120_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y120_SLICE_X12Y120_AO6),
.Q(CLBLM_L_X10Y120_SLICE_X12Y120_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y120_SLICE_X12Y120_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y120_SLICE_X12Y120_BO6),
.Q(CLBLM_L_X10Y120_SLICE_X12Y120_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y120_SLICE_X12Y120_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y120_SLICE_X12Y120_CO6),
.Q(CLBLM_L_X10Y120_SLICE_X12Y120_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y120_SLICE_X12Y120_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y120_SLICE_X12Y120_DO6),
.Q(CLBLM_L_X10Y120_SLICE_X12Y120_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff50cc000050cc)
  ) CLBLM_L_X10Y120_SLICE_X12Y120_DLUT (
.I0(CLBLM_R_X11Y119_SLICE_X14Y119_AO6),
.I1(CLBLM_R_X11Y118_SLICE_X15Y118_CQ),
.I2(CLBLM_L_X10Y120_SLICE_X12Y120_DQ),
.I3(CLBLM_L_X12Y119_SLICE_X17Y119_AO5),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(CLBLM_L_X10Y121_SLICE_X12Y121_AQ),
.O5(CLBLM_L_X10Y120_SLICE_X12Y120_DO5),
.O6(CLBLM_L_X10Y120_SLICE_X12Y120_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hffaa00aafffe00fe)
  ) CLBLM_L_X10Y120_SLICE_X12Y120_CLUT (
.I0(CLBLM_R_X11Y119_SLICE_X14Y119_AO6),
.I1(CLBLM_L_X10Y120_SLICE_X12Y120_CQ),
.I2(CLBLM_L_X10Y120_SLICE_X12Y120_DQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLM_L_X8Y121_SLICE_X10Y121_BQ),
.I5(CLBLM_L_X12Y119_SLICE_X17Y119_AO5),
.O5(CLBLM_L_X10Y120_SLICE_X12Y120_CO5),
.O6(CLBLM_L_X10Y120_SLICE_X12Y120_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f0f0f0ffee0044)
  ) CLBLM_L_X10Y120_SLICE_X12Y120_BLUT (
.I0(CLBLM_R_X3Y118_SLICE_X2Y118_AQ),
.I1(CLBLM_L_X10Y120_SLICE_X12Y120_BQ),
.I2(CLBLM_L_X10Y120_SLICE_X12Y120_DQ),
.I3(RIOB33_X105Y117_IOB_X1Y118_I),
.I4(CLBLM_R_X7Y120_SLICE_X9Y120_BQ),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLM_L_X10Y120_SLICE_X12Y120_BO5),
.O6(CLBLM_L_X10Y120_SLICE_X12Y120_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hcccc00aacccc00a0)
  ) CLBLM_L_X10Y120_SLICE_X12Y120_ALUT (
.I0(CLBLM_R_X3Y118_SLICE_X2Y118_AQ),
.I1(CLBLM_L_X10Y121_SLICE_X13Y121_BQ),
.I2(CLBLM_L_X10Y120_SLICE_X12Y120_AQ),
.I3(RIOB33_X105Y117_IOB_X1Y118_I),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(CLBLM_R_X5Y115_SLICE_X7Y115_DO6),
.O5(CLBLM_L_X10Y120_SLICE_X12Y120_AO5),
.O6(CLBLM_L_X10Y120_SLICE_X12Y120_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y120_SLICE_X13Y120_A5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y118_SLICE_X11Y118_BO6),
.Q(CLBLM_L_X10Y120_SLICE_X13Y120_A5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y120_SLICE_X13Y120_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y120_SLICE_X13Y120_AO6),
.Q(CLBLM_L_X10Y120_SLICE_X13Y120_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y120_SLICE_X13Y120_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y120_SLICE_X13Y120_BO6),
.Q(CLBLM_L_X10Y120_SLICE_X13Y120_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h99999999aa999999)
  ) CLBLM_L_X10Y120_SLICE_X13Y120_DLUT (
.I0(CLBLM_L_X10Y120_SLICE_X13Y120_BQ),
.I1(CLBLM_L_X10Y123_SLICE_X12Y123_CO6),
.I2(1'b1),
.I3(CLBLM_L_X10Y120_SLICE_X13Y120_CO6),
.I4(CLBLM_L_X10Y121_SLICE_X12Y121_BQ),
.I5(CLBLM_L_X8Y122_SLICE_X11Y122_DO6),
.O5(CLBLM_L_X10Y120_SLICE_X13Y120_DO5),
.O6(CLBLM_L_X10Y120_SLICE_X13Y120_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h00052004a000a000)
  ) CLBLM_L_X10Y120_SLICE_X13Y120_CLUT (
.I0(CLBLM_L_X10Y121_SLICE_X13Y121_AQ),
.I1(CLBLM_L_X10Y124_SLICE_X12Y124_AQ),
.I2(CLBLM_L_X10Y121_SLICE_X13Y121_CQ),
.I3(CLBLM_L_X10Y120_SLICE_X13Y120_AQ),
.I4(CLBLM_R_X7Y120_SLICE_X9Y120_A5Q),
.I5(CLBLM_R_X7Y124_SLICE_X8Y124_AQ),
.O5(CLBLM_L_X10Y120_SLICE_X13Y120_CO5),
.O6(CLBLM_L_X10Y120_SLICE_X13Y120_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h44440044ffff00ff)
  ) CLBLM_L_X10Y120_SLICE_X13Y120_BLUT (
.I0(CLBLM_L_X10Y120_SLICE_X13Y120_DO6),
.I1(CLBLM_L_X10Y124_SLICE_X13Y124_BO5),
.I2(1'b1),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLM_R_X3Y112_SLICE_X3Y112_AQ),
.I5(CLBLM_L_X10Y124_SLICE_X13Y124_AO5),
.O5(CLBLM_L_X10Y120_SLICE_X13Y120_BO5),
.O6(CLBLM_L_X10Y120_SLICE_X13Y120_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h44004444ff00ffff)
  ) CLBLM_L_X10Y120_SLICE_X13Y120_ALUT (
.I0(CLBLM_L_X10Y121_SLICE_X13Y121_DO6),
.I1(CLBLM_L_X10Y124_SLICE_X13Y124_BO5),
.I2(1'b1),
.I3(CLBLL_L_X2Y113_SLICE_X1Y113_AQ),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(CLBLM_L_X10Y124_SLICE_X13Y124_AO5),
.O5(CLBLM_L_X10Y120_SLICE_X13Y120_AO5),
.O6(CLBLM_L_X10Y120_SLICE_X13Y120_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y121_SLICE_X12Y121_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y121_SLICE_X12Y121_AO6),
.Q(CLBLM_L_X10Y121_SLICE_X12Y121_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y121_SLICE_X12Y121_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y121_SLICE_X12Y121_BO6),
.Q(CLBLM_L_X10Y121_SLICE_X12Y121_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000400)
  ) CLBLM_L_X10Y121_SLICE_X12Y121_DLUT (
.I0(CLBLM_L_X8Y115_SLICE_X10Y115_AQ),
.I1(CLBLM_L_X8Y121_SLICE_X10Y121_CQ),
.I2(CLBLM_L_X10Y119_SLICE_X13Y119_DQ),
.I3(CLBLM_L_X10Y126_SLICE_X12Y126_AQ),
.I4(CLBLM_L_X8Y121_SLICE_X11Y121_DQ),
.I5(CLBLL_L_X4Y117_SLICE_X5Y117_DQ),
.O5(CLBLM_L_X10Y121_SLICE_X12Y121_DO5),
.O6(CLBLM_L_X10Y121_SLICE_X12Y121_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0f0f0f0f0f0b070f)
  ) CLBLM_L_X10Y121_SLICE_X12Y121_CLUT (
.I0(CLBLM_L_X10Y121_SLICE_X13Y121_CQ),
.I1(CLBLM_L_X10Y121_SLICE_X12Y121_AQ),
.I2(CLBLM_L_X10Y123_SLICE_X12Y123_CO6),
.I3(CLBLM_L_X10Y120_SLICE_X13Y120_AQ),
.I4(CLBLM_L_X10Y122_SLICE_X12Y122_CO6),
.I5(CLBLM_L_X8Y122_SLICE_X11Y122_DO6),
.O5(CLBLM_L_X10Y121_SLICE_X12Y121_CO5),
.O6(CLBLM_L_X10Y121_SLICE_X12Y121_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaa00ccaaaaf0f0)
  ) CLBLM_L_X10Y121_SLICE_X12Y121_BLUT (
.I0(CLBLM_L_X8Y116_SLICE_X11Y116_DQ),
.I1(CLBLM_L_X10Y121_SLICE_X12Y121_BQ),
.I2(CLBLM_L_X10Y121_SLICE_X12Y121_AQ),
.I3(CLBLM_L_X10Y123_SLICE_X12Y123_AO6),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(CLBLM_R_X7Y123_SLICE_X9Y123_CO6),
.O5(CLBLM_L_X10Y121_SLICE_X12Y121_BO5),
.O6(CLBLM_L_X10Y121_SLICE_X12Y121_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'haaeefaee00445044)
  ) CLBLM_L_X10Y121_SLICE_X12Y121_ALUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_L_X8Y122_SLICE_X11Y122_BQ),
.I2(CLBLM_L_X10Y121_SLICE_X12Y121_AQ),
.I3(CLBLM_R_X7Y123_SLICE_X9Y123_CO6),
.I4(CLBLM_L_X10Y123_SLICE_X12Y123_AO6),
.I5(CLBLM_R_X7Y120_SLICE_X8Y120_CQ),
.O5(CLBLM_L_X10Y121_SLICE_X12Y121_AO5),
.O6(CLBLM_L_X10Y121_SLICE_X12Y121_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y121_SLICE_X13Y121_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y121_SLICE_X13Y121_AO6),
.Q(CLBLM_L_X10Y121_SLICE_X13Y121_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y121_SLICE_X13Y121_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y121_SLICE_X13Y121_BO6),
.Q(CLBLM_L_X10Y121_SLICE_X13Y121_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y121_SLICE_X13Y121_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y121_SLICE_X13Y121_CO6),
.Q(CLBLM_L_X10Y121_SLICE_X13Y121_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hcc33cc33cc39cc93)
  ) CLBLM_L_X10Y121_SLICE_X13Y121_DLUT (
.I0(CLBLM_L_X8Y122_SLICE_X11Y122_BQ),
.I1(CLBLM_L_X10Y120_SLICE_X13Y120_AQ),
.I2(CLBLM_L_X10Y122_SLICE_X12Y122_CO6),
.I3(CLBLM_L_X10Y123_SLICE_X12Y123_CO6),
.I4(CLBLM_L_X10Y121_SLICE_X13Y121_CQ),
.I5(CLBLM_L_X8Y122_SLICE_X11Y122_DO6),
.O5(CLBLM_L_X10Y121_SLICE_X13Y121_DO5),
.O6(CLBLM_L_X10Y121_SLICE_X13Y121_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h33f333f311511151)
  ) CLBLM_L_X10Y121_SLICE_X13Y121_CLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_L_X10Y124_SLICE_X13Y124_AO5),
.I2(CLBLM_L_X10Y124_SLICE_X13Y124_BO5),
.I3(CLBLM_R_X11Y121_SLICE_X14Y121_DO6),
.I4(1'b1),
.I5(CLBLM_L_X10Y117_SLICE_X13Y117_CQ),
.O5(CLBLM_L_X10Y121_SLICE_X13Y121_CO5),
.O6(CLBLM_L_X10Y121_SLICE_X13Y121_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h00aa000affff0f0f)
  ) CLBLM_L_X10Y121_SLICE_X13Y121_BLUT (
.I0(CLBLM_L_X10Y124_SLICE_X13Y124_BO5),
.I1(1'b1),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLM_L_X10Y123_SLICE_X12Y123_DO6),
.I4(CLBLM_R_X11Y120_SLICE_X15Y120_BQ),
.I5(CLBLM_L_X10Y124_SLICE_X13Y124_AO5),
.O5(CLBLM_L_X10Y121_SLICE_X13Y121_BO5),
.O6(CLBLM_L_X10Y121_SLICE_X13Y121_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'ha00a2002ffff3333)
  ) CLBLM_L_X10Y121_SLICE_X13Y121_ALUT (
.I0(CLBLM_L_X10Y124_SLICE_X13Y124_BO5),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(CLBLM_L_X10Y121_SLICE_X13Y121_AQ),
.I3(CLBLM_L_X10Y121_SLICE_X12Y121_CO6),
.I4(CLBLM_R_X7Y122_SLICE_X8Y122_DQ),
.I5(CLBLM_L_X10Y124_SLICE_X13Y124_AO5),
.O5(CLBLM_L_X10Y121_SLICE_X13Y121_AO5),
.O6(CLBLM_L_X10Y121_SLICE_X13Y121_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y122_SLICE_X12Y122_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y122_SLICE_X12Y122_AO6),
.Q(CLBLM_L_X10Y122_SLICE_X12Y122_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y122_SLICE_X12Y122_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y122_SLICE_X12Y122_BO6),
.Q(CLBLM_L_X10Y122_SLICE_X12Y122_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'haa5aaa59aa55aa55)
  ) CLBLM_L_X10Y122_SLICE_X12Y122_DLUT (
.I0(CLBLM_L_X10Y122_SLICE_X13Y122_AQ),
.I1(CLBLM_R_X11Y121_SLICE_X14Y121_BO5),
.I2(CLBLM_L_X8Y122_SLICE_X11Y122_DO6),
.I3(CLBLM_L_X10Y123_SLICE_X12Y123_CO6),
.I4(CLBLM_R_X11Y121_SLICE_X14Y121_BO6),
.I5(CLBLM_L_X8Y120_SLICE_X11Y120_BQ),
.O5(CLBLM_L_X10Y122_SLICE_X12Y122_DO5),
.O6(CLBLM_L_X10Y122_SLICE_X12Y122_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f0a0a005050000)
  ) CLBLM_L_X10Y122_SLICE_X12Y122_CLUT (
.I0(CLBLM_L_X10Y124_SLICE_X12Y124_AQ),
.I1(1'b1),
.I2(CLBLM_R_X7Y124_SLICE_X8Y124_AQ),
.I3(1'b1),
.I4(CLBLM_R_X7Y120_SLICE_X9Y120_A5Q),
.I5(1'b1),
.O5(CLBLM_L_X10Y122_SLICE_X12Y122_CO5),
.O6(CLBLM_L_X10Y122_SLICE_X12Y122_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'he2f3e2c0e2f3e2f3)
  ) CLBLM_L_X10Y122_SLICE_X12Y122_BLUT (
.I0(CLBLM_R_X7Y119_SLICE_X9Y119_DO6),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(CLBLM_L_X10Y119_SLICE_X13Y119_AQ),
.I3(CLBLM_L_X10Y123_SLICE_X12Y123_AO6),
.I4(CLBLM_L_X10Y122_SLICE_X12Y122_CO5),
.I5(CLBLM_L_X8Y122_SLICE_X10Y122_CO6),
.O5(CLBLM_L_X10Y122_SLICE_X12Y122_BO5),
.O6(CLBLM_L_X10Y122_SLICE_X12Y122_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff000000cc00cc)
  ) CLBLM_L_X10Y122_SLICE_X12Y122_ALUT (
.I0(1'b1),
.I1(CLBLM_R_X7Y122_SLICE_X8Y122_CQ),
.I2(1'b1),
.I3(CLBLM_L_X10Y124_SLICE_X13Y124_BO6),
.I4(CLBLM_L_X10Y118_SLICE_X13Y118_AQ),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLM_L_X10Y122_SLICE_X12Y122_AO5),
.O6(CLBLM_L_X10Y122_SLICE_X12Y122_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y122_SLICE_X13Y122_A5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y124_SLICE_X13Y124_AO6),
.Q(CLBLM_L_X10Y122_SLICE_X13Y122_A5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y122_SLICE_X13Y122_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y122_SLICE_X13Y122_AO6),
.Q(CLBLM_L_X10Y122_SLICE_X13Y122_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y122_SLICE_X13Y122_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y122_SLICE_X13Y122_BO6),
.Q(CLBLM_L_X10Y122_SLICE_X13Y122_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y122_SLICE_X13Y122_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y122_SLICE_X13Y122_CO6),
.Q(CLBLM_L_X10Y122_SLICE_X13Y122_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h3130313333333333)
  ) CLBLM_L_X10Y122_SLICE_X13Y122_DLUT (
.I0(CLBLM_R_X11Y121_SLICE_X14Y121_BO6),
.I1(CLBLM_L_X10Y123_SLICE_X12Y123_CO6),
.I2(CLBLM_L_X8Y122_SLICE_X11Y122_DO6),
.I3(CLBLM_L_X10Y122_SLICE_X13Y122_AQ),
.I4(CLBLM_R_X11Y121_SLICE_X14Y121_BO5),
.I5(CLBLM_L_X8Y121_SLICE_X11Y121_AQ),
.O5(CLBLM_L_X10Y122_SLICE_X13Y122_DO5),
.O6(CLBLM_L_X10Y122_SLICE_X13Y122_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h90ff000090ff90ff)
  ) CLBLM_L_X10Y122_SLICE_X13Y122_CLUT (
.I0(CLBLM_R_X11Y122_SLICE_X14Y122_BO6),
.I1(CLBLM_L_X10Y122_SLICE_X13Y122_CQ),
.I2(CLBLM_L_X10Y124_SLICE_X13Y124_BO5),
.I3(CLBLM_L_X10Y124_SLICE_X13Y124_AO5),
.I4(CLBLM_L_X10Y119_SLICE_X12Y119_AQ),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLM_L_X10Y122_SLICE_X13Y122_CO5),
.O6(CLBLM_L_X10Y122_SLICE_X13Y122_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h88220802ffff0f0f)
  ) CLBLM_L_X10Y122_SLICE_X13Y122_BLUT (
.I0(CLBLM_L_X10Y124_SLICE_X13Y124_BO5),
.I1(CLBLM_L_X10Y122_SLICE_X13Y122_BQ),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLM_L_X10Y122_SLICE_X13Y122_DO6),
.I4(CLBLM_R_X7Y120_SLICE_X9Y120_DQ),
.I5(CLBLM_L_X10Y124_SLICE_X13Y124_AO5),
.O5(CLBLM_L_X10Y122_SLICE_X13Y122_BO5),
.O6(CLBLM_L_X10Y122_SLICE_X13Y122_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h00a200a2f3f3f3f3)
  ) CLBLM_L_X10Y122_SLICE_X13Y122_ALUT (
.I0(CLBLM_L_X10Y124_SLICE_X13Y124_BO5),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(CLBLM_L_X10Y112_SLICE_X13Y112_AQ),
.I3(CLBLM_L_X10Y122_SLICE_X12Y122_DO6),
.I4(1'b1),
.I5(CLBLM_L_X10Y124_SLICE_X13Y124_AO5),
.O5(CLBLM_L_X10Y122_SLICE_X13Y122_AO5),
.O6(CLBLM_L_X10Y122_SLICE_X13Y122_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h5a5a5a5a5aa55aa5)
  ) CLBLM_L_X10Y123_SLICE_X12Y123_DLUT (
.I0(CLBLM_L_X8Y123_SLICE_X10Y123_AQ),
.I1(1'b1),
.I2(CLBLM_L_X10Y121_SLICE_X13Y121_BQ),
.I3(CLBLM_L_X10Y123_SLICE_X12Y123_CO6),
.I4(1'b1),
.I5(CLBLM_L_X10Y123_SLICE_X12Y123_BO6),
.O5(CLBLM_L_X10Y123_SLICE_X12Y123_DO5),
.O6(CLBLM_L_X10Y123_SLICE_X12Y123_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h3333ffff3333fff7)
  ) CLBLM_L_X10Y123_SLICE_X12Y123_CLUT (
.I0(CLBLM_L_X10Y124_SLICE_X12Y124_AQ),
.I1(CLBLM_R_X7Y123_SLICE_X9Y123_BO5),
.I2(CLBLM_R_X5Y120_SLICE_X6Y120_A5Q),
.I3(CLBLM_R_X7Y120_SLICE_X9Y120_A5Q),
.I4(CLBLM_L_X10Y118_SLICE_X12Y118_B5Q),
.I5(CLBLM_R_X7Y124_SLICE_X8Y124_AQ),
.O5(CLBLM_L_X10Y123_SLICE_X12Y123_CO5),
.O6(CLBLM_L_X10Y123_SLICE_X12Y123_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h4100010040000000)
  ) CLBLM_L_X10Y123_SLICE_X12Y123_BLUT (
.I0(CLBLM_L_X8Y122_SLICE_X11Y122_DO6),
.I1(CLBLM_L_X10Y122_SLICE_X13Y122_BQ),
.I2(CLBLM_L_X10Y122_SLICE_X13Y122_AQ),
.I3(CLBLM_L_X8Y121_SLICE_X11Y121_BQ),
.I4(CLBLM_R_X11Y121_SLICE_X14Y121_BO6),
.I5(CLBLM_R_X11Y121_SLICE_X14Y121_BO5),
.O5(CLBLM_L_X10Y123_SLICE_X12Y123_BO5),
.O6(CLBLM_L_X10Y123_SLICE_X12Y123_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000300000200)
  ) CLBLM_L_X10Y123_SLICE_X12Y123_ALUT (
.I0(CLBLM_R_X7Y123_SLICE_X9Y123_BO5),
.I1(CLBLM_R_X7Y124_SLICE_X8Y124_AQ),
.I2(CLBLM_R_X5Y120_SLICE_X6Y120_A5Q),
.I3(CLBLM_L_X10Y124_SLICE_X12Y124_AQ),
.I4(CLBLM_R_X7Y120_SLICE_X9Y120_A5Q),
.I5(1'b1),
.O5(CLBLM_L_X10Y123_SLICE_X12Y123_AO5),
.O6(CLBLM_L_X10Y123_SLICE_X12Y123_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y123_SLICE_X13Y123_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y123_SLICE_X13Y123_AO6),
.Q(CLBLM_L_X10Y123_SLICE_X13Y123_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0c000a0a00000a0a)
  ) CLBLM_L_X10Y123_SLICE_X13Y123_DLUT (
.I0(CLBLM_R_X11Y123_SLICE_X14Y123_AO6),
.I1(CLBLM_L_X10Y122_SLICE_X13Y122_CQ),
.I2(CLBLM_L_X8Y122_SLICE_X11Y122_DO6),
.I3(CLBLM_R_X11Y123_SLICE_X14Y123_BO5),
.I4(CLBLM_L_X10Y123_SLICE_X13Y123_AQ),
.I5(CLBLM_L_X10Y121_SLICE_X13Y121_BQ),
.O5(CLBLM_L_X10Y123_SLICE_X13Y123_DO5),
.O6(CLBLM_L_X10Y123_SLICE_X13Y123_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hcc33fe01cc33cc33)
  ) CLBLM_L_X10Y123_SLICE_X13Y123_CLUT (
.I0(CLBLM_R_X11Y123_SLICE_X14Y123_BO6),
.I1(CLBLM_L_X10Y123_SLICE_X12Y123_CO6),
.I2(CLBLM_R_X11Y123_SLICE_X14Y123_AO6),
.I3(CLBLM_L_X10Y123_SLICE_X13Y123_AQ),
.I4(CLBLM_L_X8Y122_SLICE_X11Y122_DO6),
.I5(CLBLM_L_X8Y121_SLICE_X10Y121_AQ),
.O5(CLBLM_L_X10Y123_SLICE_X13Y123_CO5),
.O6(CLBLM_L_X10Y123_SLICE_X13Y123_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h00000c0f00000f0a)
  ) CLBLM_L_X10Y123_SLICE_X13Y123_BLUT (
.I0(CLBLM_L_X10Y123_SLICE_X12Y123_AO5),
.I1(CLBLM_R_X7Y123_SLICE_X9Y123_CO6),
.I2(RIOB33_X105Y121_IOB_X1Y121_I),
.I3(CLBLM_L_X10Y118_SLICE_X12Y118_B5Q),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(CLBLM_L_X8Y121_SLICE_X10Y121_AQ),
.O5(CLBLM_L_X10Y123_SLICE_X13Y123_BO5),
.O6(CLBLM_L_X10Y123_SLICE_X13Y123_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h33330303bbbb0b0b)
  ) CLBLM_L_X10Y123_SLICE_X13Y123_ALUT (
.I0(CLBLM_L_X10Y124_SLICE_X13Y124_BO5),
.I1(CLBLM_L_X10Y124_SLICE_X13Y124_AO5),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(1'b1),
.I4(CLBLM_L_X10Y120_SLICE_X13Y120_A5Q),
.I5(CLBLM_L_X10Y123_SLICE_X13Y123_CO6),
.O5(CLBLM_L_X10Y123_SLICE_X13Y123_AO5),
.O6(CLBLM_L_X10Y123_SLICE_X13Y123_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y124_SLICE_X12Y124_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y124_SLICE_X12Y124_AO6),
.Q(CLBLM_L_X10Y124_SLICE_X12Y124_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X10Y124_SLICE_X12Y124_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X10Y124_SLICE_X12Y124_DO5),
.O6(CLBLM_L_X10Y124_SLICE_X12Y124_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X10Y124_SLICE_X12Y124_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X10Y124_SLICE_X12Y124_CO5),
.O6(CLBLM_L_X10Y124_SLICE_X12Y124_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X10Y124_SLICE_X12Y124_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X10Y124_SLICE_X12Y124_BO5),
.O6(CLBLM_L_X10Y124_SLICE_X12Y124_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h8888b88b8888b8b8)
  ) CLBLM_L_X10Y124_SLICE_X12Y124_ALUT (
.I0(CLBLM_L_X8Y121_SLICE_X11Y121_DQ),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(CLBLM_L_X10Y124_SLICE_X12Y124_AQ),
.I3(CLBLM_L_X10Y124_SLICE_X13Y124_CO6),
.I4(RIOB33_X105Y121_IOB_X1Y121_I),
.I5(CLBLM_L_X10Y123_SLICE_X13Y123_DO6),
.O5(CLBLM_L_X10Y124_SLICE_X12Y124_AO5),
.O6(CLBLM_L_X10Y124_SLICE_X12Y124_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y124_SLICE_X13Y124_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(LIOB33_X0Y77_IOB_X0Y77_I),
.D(CLBLM_L_X10Y118_SLICE_X12Y118_B5Q),
.Q(CLBLM_L_X10Y124_SLICE_X13Y124_AQ),
.R(CLBLM_R_X11Y123_SLICE_X14Y123_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X10Y124_SLICE_X13Y124_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X10Y124_SLICE_X13Y124_DO5),
.O6(CLBLM_L_X10Y124_SLICE_X13Y124_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hc4f533330ace33dd)
  ) CLBLM_L_X10Y124_SLICE_X13Y124_CLUT (
.I0(CLBLM_R_X5Y120_SLICE_X6Y120_A5Q),
.I1(CLBLM_R_X7Y124_SLICE_X8Y124_AQ),
.I2(CLBLM_L_X10Y118_SLICE_X12Y118_B5Q),
.I3(CLBLM_R_X7Y120_SLICE_X9Y120_A5Q),
.I4(CLBLM_L_X10Y124_SLICE_X12Y124_AQ),
.I5(1'b1),
.O5(CLBLM_L_X10Y124_SLICE_X13Y124_CO5),
.O6(CLBLM_L_X10Y124_SLICE_X13Y124_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000ff0533333332)
  ) CLBLM_L_X10Y124_SLICE_X13Y124_BLUT (
.I0(CLBLM_R_X7Y124_SLICE_X8Y124_AQ),
.I1(CLBLM_L_X10Y123_SLICE_X13Y123_DO6),
.I2(CLBLM_R_X7Y120_SLICE_X9Y120_A5Q),
.I3(CLBLM_R_X5Y120_SLICE_X6Y120_A5Q),
.I4(CLBLM_L_X10Y124_SLICE_X12Y124_AQ),
.I5(1'b1),
.O5(CLBLM_L_X10Y124_SLICE_X13Y124_BO5),
.O6(CLBLM_L_X10Y124_SLICE_X13Y124_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfa50fa5055551111)
  ) CLBLM_L_X10Y124_SLICE_X13Y124_ALUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_L_X10Y123_SLICE_X13Y123_DO6),
.I2(CLBLM_L_X10Y120_SLICE_X13Y120_A5Q),
.I3(CLBLM_L_X10Y120_SLICE_X13Y120_AQ),
.I4(CLBLM_L_X10Y124_SLICE_X13Y124_CO5),
.I5(1'b1),
.O5(CLBLM_L_X10Y124_SLICE_X13Y124_AO5),
.O6(CLBLM_L_X10Y124_SLICE_X13Y124_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y126_SLICE_X12Y126_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y128_SLICE_X14Y128_AO6),
.Q(CLBLM_L_X10Y126_SLICE_X12Y126_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X10Y126_SLICE_X12Y126_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X10Y126_SLICE_X12Y126_DO5),
.O6(CLBLM_L_X10Y126_SLICE_X12Y126_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X10Y126_SLICE_X12Y126_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X10Y126_SLICE_X12Y126_CO5),
.O6(CLBLM_L_X10Y126_SLICE_X12Y126_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X10Y126_SLICE_X12Y126_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X10Y126_SLICE_X12Y126_BO5),
.O6(CLBLM_L_X10Y126_SLICE_X12Y126_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X10Y126_SLICE_X12Y126_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X10Y126_SLICE_X12Y126_AO5),
.O6(CLBLM_L_X10Y126_SLICE_X12Y126_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X10Y126_SLICE_X13Y126_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X10Y126_SLICE_X13Y126_DO5),
.O6(CLBLM_L_X10Y126_SLICE_X13Y126_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X10Y126_SLICE_X13Y126_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X10Y126_SLICE_X13Y126_CO5),
.O6(CLBLM_L_X10Y126_SLICE_X13Y126_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X10Y126_SLICE_X13Y126_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X10Y126_SLICE_X13Y126_BO5),
.O6(CLBLM_L_X10Y126_SLICE_X13Y126_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X10Y126_SLICE_X13Y126_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X10Y126_SLICE_X13Y126_AO5),
.O6(CLBLM_L_X10Y126_SLICE_X13Y126_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y127_SLICE_X12Y127_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y128_SLICE_X13Y128_AO5),
.Q(CLBLM_L_X10Y127_SLICE_X12Y127_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X10Y127_SLICE_X12Y127_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X10Y127_SLICE_X12Y127_DO5),
.O6(CLBLM_L_X10Y127_SLICE_X12Y127_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X10Y127_SLICE_X12Y127_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X10Y127_SLICE_X12Y127_CO5),
.O6(CLBLM_L_X10Y127_SLICE_X12Y127_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X10Y127_SLICE_X12Y127_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X10Y127_SLICE_X12Y127_BO5),
.O6(CLBLM_L_X10Y127_SLICE_X12Y127_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X10Y127_SLICE_X12Y127_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X10Y127_SLICE_X12Y127_AO5),
.O6(CLBLM_L_X10Y127_SLICE_X12Y127_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X10Y127_SLICE_X13Y127_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X10Y127_SLICE_X13Y127_DO5),
.O6(CLBLM_L_X10Y127_SLICE_X13Y127_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X10Y127_SLICE_X13Y127_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X10Y127_SLICE_X13Y127_CO5),
.O6(CLBLM_L_X10Y127_SLICE_X13Y127_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X10Y127_SLICE_X13Y127_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X10Y127_SLICE_X13Y127_BO5),
.O6(CLBLM_L_X10Y127_SLICE_X13Y127_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X10Y127_SLICE_X13Y127_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X10Y127_SLICE_X13Y127_AO5),
.O6(CLBLM_L_X10Y127_SLICE_X13Y127_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X10Y128_SLICE_X12Y128_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X10Y128_SLICE_X12Y128_DO5),
.O6(CLBLM_L_X10Y128_SLICE_X12Y128_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X10Y128_SLICE_X12Y128_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X10Y128_SLICE_X12Y128_CO5),
.O6(CLBLM_L_X10Y128_SLICE_X12Y128_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X10Y128_SLICE_X12Y128_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X10Y128_SLICE_X12Y128_BO5),
.O6(CLBLM_L_X10Y128_SLICE_X12Y128_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X10Y128_SLICE_X12Y128_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X10Y128_SLICE_X12Y128_AO5),
.O6(CLBLM_L_X10Y128_SLICE_X12Y128_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X10Y128_SLICE_X13Y128_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X10Y128_SLICE_X13Y128_DO5),
.O6(CLBLM_L_X10Y128_SLICE_X13Y128_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X10Y128_SLICE_X13Y128_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X10Y128_SLICE_X13Y128_CO5),
.O6(CLBLM_L_X10Y128_SLICE_X13Y128_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X10Y128_SLICE_X13Y128_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X10Y128_SLICE_X13Y128_BO5),
.O6(CLBLM_L_X10Y128_SLICE_X13Y128_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0fff0fff5f5a0a0)
  ) CLBLM_L_X10Y128_SLICE_X13Y128_ALUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(1'b1),
.I2(CLBLM_L_X10Y124_SLICE_X13Y124_AQ),
.I3(RIOB33_X105Y143_IOB_X1Y143_I),
.I4(CLBLM_L_X8Y122_SLICE_X11Y122_A5Q),
.I5(1'b1),
.O5(CLBLM_L_X10Y128_SLICE_X13Y128_AO5),
.O6(CLBLM_L_X10Y128_SLICE_X13Y128_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y115_SLICE_X16Y115_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X12Y115_SLICE_X16Y115_AO6),
.Q(CLBLM_L_X12Y115_SLICE_X16Y115_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y115_SLICE_X16Y115_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X12Y115_SLICE_X16Y115_BO6),
.Q(CLBLM_L_X12Y115_SLICE_X16Y115_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y115_SLICE_X16Y115_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X12Y115_SLICE_X16Y115_CO6),
.Q(CLBLM_L_X12Y115_SLICE_X16Y115_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y115_SLICE_X16Y115_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X12Y115_SLICE_X16Y115_DO6),
.Q(CLBLM_L_X12Y115_SLICE_X16Y115_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hcc55cc00cc50cc00)
  ) CLBLM_L_X12Y115_SLICE_X16Y115_DLUT (
.I0(RIOB33_X105Y117_IOB_X1Y118_I),
.I1(CLBLM_L_X10Y114_SLICE_X13Y114_AQ),
.I2(CLBLM_L_X12Y115_SLICE_X16Y115_DQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLM_R_X3Y118_SLICE_X2Y118_AQ),
.I5(CLBLM_L_X10Y114_SLICE_X13Y114_CQ),
.O5(CLBLM_L_X12Y115_SLICE_X16Y115_DO5),
.O6(CLBLM_L_X12Y115_SLICE_X16Y115_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hff00ff00f0f0e4e4)
  ) CLBLM_L_X12Y115_SLICE_X16Y115_CLUT (
.I0(RIOB33_X105Y117_IOB_X1Y118_I),
.I1(CLBLM_L_X12Y115_SLICE_X16Y115_CQ),
.I2(CLBLM_L_X12Y115_SLICE_X16Y115_DQ),
.I3(CLBLM_L_X12Y115_SLICE_X16Y115_BQ),
.I4(CLBLM_R_X3Y118_SLICE_X2Y118_AQ),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLM_L_X12Y115_SLICE_X16Y115_CO5),
.O6(CLBLM_L_X12Y115_SLICE_X16Y115_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'he4f5e4e4e4f5e4e4)
  ) CLBLM_L_X12Y115_SLICE_X16Y115_BLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_L_X12Y115_SLICE_X16Y115_BQ),
.I2(CLBLM_R_X7Y114_SLICE_X8Y114_AQ),
.I3(CLBLM_R_X7Y128_SLICE_X8Y128_AQ),
.I4(RIOB33_X105Y141_IOB_X1Y142_I),
.I5(1'b1),
.O5(CLBLM_L_X12Y115_SLICE_X16Y115_BO5),
.O6(CLBLM_L_X12Y115_SLICE_X16Y115_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfafffafa50555050)
  ) CLBLM_L_X12Y115_SLICE_X16Y115_ALUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(1'b1),
.I2(CLBLM_L_X12Y115_SLICE_X16Y115_AQ),
.I3(CLBLM_R_X7Y128_SLICE_X8Y128_AQ),
.I4(RIOB33_X105Y141_IOB_X1Y142_I),
.I5(CLBLM_R_X7Y115_SLICE_X9Y115_B5Q),
.O5(CLBLM_L_X12Y115_SLICE_X16Y115_AO5),
.O6(CLBLM_L_X12Y115_SLICE_X16Y115_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X12Y115_SLICE_X17Y115_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X12Y115_SLICE_X17Y115_DO5),
.O6(CLBLM_L_X12Y115_SLICE_X17Y115_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X12Y115_SLICE_X17Y115_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X12Y115_SLICE_X17Y115_CO5),
.O6(CLBLM_L_X12Y115_SLICE_X17Y115_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X12Y115_SLICE_X17Y115_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X12Y115_SLICE_X17Y115_BO5),
.O6(CLBLM_L_X12Y115_SLICE_X17Y115_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X12Y115_SLICE_X17Y115_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X12Y115_SLICE_X17Y115_AO5),
.O6(CLBLM_L_X12Y115_SLICE_X17Y115_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y118_SLICE_X16Y118_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X12Y118_SLICE_X16Y118_AO6),
.Q(CLBLM_L_X12Y118_SLICE_X16Y118_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y118_SLICE_X16Y118_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X12Y118_SLICE_X16Y118_BO6),
.Q(CLBLM_L_X12Y118_SLICE_X16Y118_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X12Y118_SLICE_X16Y118_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X12Y118_SLICE_X16Y118_DO5),
.O6(CLBLM_L_X12Y118_SLICE_X16Y118_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h339c33cc339c339c)
  ) CLBLM_L_X12Y118_SLICE_X16Y118_CLUT (
.I0(CLBLM_R_X11Y118_SLICE_X14Y118_DO5),
.I1(CLBLM_L_X12Y118_SLICE_X16Y118_AQ),
.I2(CLBLM_R_X11Y118_SLICE_X15Y118_CQ),
.I3(CLBLM_L_X12Y119_SLICE_X17Y119_DO6),
.I4(CLBLM_L_X12Y119_SLICE_X16Y119_DO6),
.I5(CLBLM_L_X12Y118_SLICE_X17Y118_AO6),
.O5(CLBLM_L_X12Y118_SLICE_X16Y118_CO5),
.O6(CLBLM_L_X12Y118_SLICE_X16Y118_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf2f3f3f202030302)
  ) CLBLM_L_X12Y118_SLICE_X16Y118_BLUT (
.I0(CLBLM_R_X11Y120_SLICE_X14Y120_AO5),
.I1(CLBLM_L_X12Y120_SLICE_X17Y120_CO5),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLM_L_X12Y119_SLICE_X16Y119_BO6),
.I4(CLBLM_L_X12Y118_SLICE_X16Y118_BQ),
.I5(CLBLM_R_X7Y118_SLICE_X9Y118_CQ),
.O5(CLBLM_L_X12Y118_SLICE_X16Y118_BO5),
.O6(CLBLM_L_X12Y118_SLICE_X16Y118_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hc0cfc0cfc0cac0ca)
  ) CLBLM_L_X12Y118_SLICE_X16Y118_ALUT (
.I0(CLBLM_R_X11Y120_SLICE_X14Y120_AO5),
.I1(CLBLM_R_X11Y118_SLICE_X14Y118_CQ),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLM_L_X12Y120_SLICE_X17Y120_CO5),
.I4(1'b1),
.I5(CLBLM_L_X12Y118_SLICE_X16Y118_CO6),
.O5(CLBLM_L_X12Y118_SLICE_X16Y118_AO5),
.O6(CLBLM_L_X12Y118_SLICE_X16Y118_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X12Y118_SLICE_X17Y118_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X12Y118_SLICE_X17Y118_DO5),
.O6(CLBLM_L_X12Y118_SLICE_X17Y118_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X12Y118_SLICE_X17Y118_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X12Y118_SLICE_X17Y118_CO5),
.O6(CLBLM_L_X12Y118_SLICE_X17Y118_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X12Y118_SLICE_X17Y118_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X12Y118_SLICE_X17Y118_BO5),
.O6(CLBLM_L_X12Y118_SLICE_X17Y118_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h5fffffffffffffff)
  ) CLBLM_L_X12Y118_SLICE_X17Y118_ALUT (
.I0(CLBLM_R_X11Y119_SLICE_X15Y119_AQ),
.I1(1'b1),
.I2(CLBLM_R_X11Y119_SLICE_X15Y119_BQ),
.I3(CLBLM_L_X12Y118_SLICE_X16Y118_BQ),
.I4(CLBLM_R_X13Y119_SLICE_X18Y119_DO6),
.I5(CLBLM_L_X12Y120_SLICE_X17Y120_BQ),
.O5(CLBLM_L_X12Y118_SLICE_X17Y118_AO5),
.O6(CLBLM_L_X12Y118_SLICE_X17Y118_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000001000100)
  ) CLBLM_L_X12Y119_SLICE_X16Y119_DLUT (
.I0(CLBLM_R_X11Y119_SLICE_X15Y119_BQ),
.I1(CLBLM_L_X12Y120_SLICE_X17Y120_BQ),
.I2(CLBLM_R_X11Y119_SLICE_X15Y119_AQ),
.I3(CLBLM_R_X13Y120_SLICE_X18Y120_CO6),
.I4(1'b1),
.I5(CLBLM_L_X12Y118_SLICE_X16Y118_BQ),
.O5(CLBLM_L_X12Y119_SLICE_X16Y119_DO5),
.O6(CLBLM_L_X12Y119_SLICE_X16Y119_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000004)
  ) CLBLM_L_X12Y119_SLICE_X16Y119_CLUT (
.I0(CLBLM_L_X12Y118_SLICE_X16Y118_AQ),
.I1(CLBLM_R_X13Y120_SLICE_X18Y120_CO6),
.I2(CLBLM_L_X12Y120_SLICE_X17Y120_BQ),
.I3(CLBLM_R_X11Y119_SLICE_X15Y119_AQ),
.I4(CLBLM_R_X11Y119_SLICE_X15Y119_BQ),
.I5(CLBLM_L_X12Y118_SLICE_X16Y118_BQ),
.O5(CLBLM_L_X12Y119_SLICE_X16Y119_CO5),
.O6(CLBLM_L_X12Y119_SLICE_X16Y119_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f3f1f1f0f0f0f0)
  ) CLBLM_L_X12Y119_SLICE_X16Y119_BLUT (
.I0(CLBLM_R_X13Y120_SLICE_X18Y120_AO6),
.I1(CLBLM_R_X11Y118_SLICE_X14Y118_DO5),
.I2(CLBLM_L_X12Y119_SLICE_X17Y119_DO6),
.I3(CLBLM_R_X13Y120_SLICE_X18Y120_BO6),
.I4(CLBLM_R_X11Y119_SLICE_X15Y119_BQ),
.I5(CLBLM_L_X10Y118_SLICE_X13Y118_BQ),
.O5(CLBLM_L_X12Y119_SLICE_X16Y119_BO5),
.O6(CLBLM_L_X12Y119_SLICE_X16Y119_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0f0ff0f00b03f4fc)
  ) CLBLM_L_X12Y119_SLICE_X16Y119_ALUT (
.I0(CLBLM_R_X13Y120_SLICE_X18Y120_AO6),
.I1(CLBLM_L_X10Y117_SLICE_X12Y117_BQ),
.I2(CLBLM_L_X12Y119_SLICE_X17Y119_DO6),
.I3(CLBLM_R_X13Y120_SLICE_X18Y120_BO6),
.I4(CLBLM_R_X11Y119_SLICE_X15Y119_BQ),
.I5(CLBLM_R_X11Y118_SLICE_X14Y118_DO5),
.O5(CLBLM_L_X12Y119_SLICE_X16Y119_AO5),
.O6(CLBLM_L_X12Y119_SLICE_X16Y119_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h55ff55fd55ff55ff)
  ) CLBLM_L_X12Y119_SLICE_X17Y119_DLUT (
.I0(CLBLM_L_X10Y116_SLICE_X12Y116_DO5),
.I1(CLBLM_L_X10Y119_SLICE_X13Y119_AQ),
.I2(CLBLM_R_X11Y118_SLICE_X14Y118_BQ),
.I3(CLBLM_R_X7Y120_SLICE_X9Y120_AQ),
.I4(CLBLM_R_X13Y119_SLICE_X18Y119_CQ),
.I5(CLBLM_R_X11Y119_SLICE_X15Y119_CQ),
.O5(CLBLM_L_X12Y119_SLICE_X17Y119_DO5),
.O6(CLBLM_L_X12Y119_SLICE_X17Y119_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h8000000000000000)
  ) CLBLM_L_X12Y119_SLICE_X17Y119_CLUT (
.I0(CLBLM_L_X12Y118_SLICE_X16Y118_AQ),
.I1(CLBLM_R_X11Y119_SLICE_X15Y119_AQ),
.I2(CLBLM_L_X12Y118_SLICE_X16Y118_BQ),
.I3(CLBLM_R_X13Y119_SLICE_X18Y119_DO6),
.I4(CLBLM_L_X12Y120_SLICE_X17Y120_BQ),
.I5(CLBLM_R_X11Y119_SLICE_X15Y119_BQ),
.O5(CLBLM_L_X12Y119_SLICE_X17Y119_CO5),
.O6(CLBLM_L_X12Y119_SLICE_X17Y119_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h00cf00ff00dd00ff)
  ) CLBLM_L_X12Y119_SLICE_X17Y119_BLUT (
.I0(CLBLM_R_X13Y120_SLICE_X18Y120_CO6),
.I1(CLBLM_R_X11Y118_SLICE_X14Y118_DO5),
.I2(CLBLM_R_X13Y119_SLICE_X18Y119_DO6),
.I3(CLBLM_L_X12Y119_SLICE_X17Y119_DO6),
.I4(CLBLM_R_X11Y117_SLICE_X15Y117_AQ),
.I5(CLBLM_R_X11Y119_SLICE_X15Y119_AQ),
.O5(CLBLM_L_X12Y119_SLICE_X17Y119_BO5),
.O6(CLBLM_L_X12Y119_SLICE_X17Y119_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h5f5f1f5f20202020)
  ) CLBLM_L_X12Y119_SLICE_X17Y119_ALUT (
.I0(CLBLM_R_X7Y120_SLICE_X9Y120_AQ),
.I1(CLBLM_R_X13Y119_SLICE_X18Y119_CQ),
.I2(CLBLM_L_X10Y116_SLICE_X12Y116_DO5),
.I3(CLBLM_R_X11Y119_SLICE_X15Y119_CQ),
.I4(CLBLM_L_X12Y120_SLICE_X16Y120_AO5),
.I5(1'b1),
.O5(CLBLM_L_X12Y119_SLICE_X17Y119_AO5),
.O6(CLBLM_L_X12Y119_SLICE_X17Y119_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h55555555a5a6aaaa)
  ) CLBLM_L_X12Y120_SLICE_X16Y120_DLUT (
.I0(CLBLM_L_X12Y121_SLICE_X16Y121_AQ),
.I1(CLBLM_L_X12Y119_SLICE_X16Y119_CO6),
.I2(CLBLM_R_X11Y118_SLICE_X14Y118_DO5),
.I3(CLBLM_L_X12Y119_SLICE_X17Y119_CO6),
.I4(CLBLM_L_X10Y120_SLICE_X12Y120_DQ),
.I5(CLBLM_L_X12Y119_SLICE_X17Y119_DO6),
.O5(CLBLM_L_X12Y120_SLICE_X16Y120_DO5),
.O6(CLBLM_L_X12Y120_SLICE_X16Y120_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h3333cc963333cccc)
  ) CLBLM_L_X12Y120_SLICE_X16Y120_CLUT (
.I0(CLBLM_R_X11Y118_SLICE_X15Y118_AQ),
.I1(CLBLM_L_X12Y120_SLICE_X17Y120_AQ),
.I2(CLBLM_L_X12Y120_SLICE_X17Y120_DO6),
.I3(CLBLM_R_X11Y118_SLICE_X14Y118_DO5),
.I4(CLBLM_L_X12Y119_SLICE_X17Y119_DO6),
.I5(CLBLM_L_X10Y118_SLICE_X13Y118_AQ),
.O5(CLBLM_L_X12Y120_SLICE_X16Y120_CO5),
.O6(CLBLM_L_X12Y120_SLICE_X16Y120_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h00000000effbffff)
  ) CLBLM_L_X12Y120_SLICE_X16Y120_BLUT (
.I0(CLBLM_R_X11Y118_SLICE_X14Y118_DO5),
.I1(CLBLM_L_X12Y120_SLICE_X17Y120_DO6),
.I2(CLBLM_R_X11Y118_SLICE_X15Y118_AQ),
.I3(CLBLM_L_X12Y120_SLICE_X17Y120_AQ),
.I4(CLBLM_R_X11Y117_SLICE_X14Y117_AQ),
.I5(CLBLM_L_X12Y119_SLICE_X17Y119_DO6),
.O5(CLBLM_L_X12Y120_SLICE_X16Y120_BO5),
.O6(CLBLM_L_X12Y120_SLICE_X16Y120_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h3030222230302222)
  ) CLBLM_L_X12Y120_SLICE_X16Y120_ALUT (
.I0(CLBLM_L_X12Y119_SLICE_X16Y119_CO6),
.I1(CLBLM_R_X11Y118_SLICE_X14Y118_DO5),
.I2(CLBLM_L_X12Y119_SLICE_X17Y119_CO6),
.I3(1'b1),
.I4(CLBLM_L_X12Y121_SLICE_X16Y121_AQ),
.I5(1'b1),
.O5(CLBLM_L_X12Y120_SLICE_X16Y120_AO5),
.O6(CLBLM_L_X12Y120_SLICE_X16Y120_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y120_SLICE_X17Y120_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X12Y120_SLICE_X17Y120_AO6),
.Q(CLBLM_L_X12Y120_SLICE_X17Y120_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y120_SLICE_X17Y120_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X12Y120_SLICE_X17Y120_BO6),
.Q(CLBLM_L_X12Y120_SLICE_X17Y120_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hffaa0000000000aa)
  ) CLBLM_L_X12Y120_SLICE_X17Y120_DLUT (
.I0(CLBLM_R_X11Y118_SLICE_X14Y118_BQ),
.I1(1'b1),
.I2(1'b1),
.I3(CLBLM_R_X11Y119_SLICE_X15Y119_CQ),
.I4(CLBLM_L_X10Y119_SLICE_X13Y119_AQ),
.I5(1'b1),
.O5(CLBLM_L_X12Y120_SLICE_X17Y120_DO5),
.O6(CLBLM_L_X12Y120_SLICE_X17Y120_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0f000f0533333332)
  ) CLBLM_L_X12Y120_SLICE_X17Y120_CLUT (
.I0(CLBLM_R_X11Y118_SLICE_X14Y118_BQ),
.I1(CLBLM_L_X12Y120_SLICE_X16Y120_AO5),
.I2(CLBLM_R_X11Y119_SLICE_X15Y119_CQ),
.I3(CLBLM_R_X13Y119_SLICE_X18Y119_CQ),
.I4(CLBLM_L_X10Y119_SLICE_X13Y119_AQ),
.I5(1'b1),
.O5(CLBLM_L_X12Y120_SLICE_X17Y120_CO5),
.O6(CLBLM_L_X12Y120_SLICE_X17Y120_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f0fff900000f09)
  ) CLBLM_L_X12Y120_SLICE_X17Y120_BLUT (
.I0(CLBLM_L_X12Y119_SLICE_X17Y119_BO6),
.I1(CLBLM_L_X12Y120_SLICE_X17Y120_BQ),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLM_R_X11Y120_SLICE_X14Y120_AO5),
.I4(CLBLM_L_X12Y120_SLICE_X17Y120_CO5),
.I5(CLBLM_R_X5Y120_SLICE_X6Y120_BQ),
.O5(CLBLM_L_X12Y120_SLICE_X17Y120_BO5),
.O6(CLBLM_L_X12Y120_SLICE_X17Y120_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f0fffa00000f0a)
  ) CLBLM_L_X12Y120_SLICE_X17Y120_ALUT (
.I0(CLBLM_L_X12Y120_SLICE_X16Y120_CO6),
.I1(1'b1),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLM_R_X11Y120_SLICE_X14Y120_AO5),
.I4(CLBLM_L_X12Y120_SLICE_X17Y120_CO5),
.I5(CLBLM_R_X13Y119_SLICE_X18Y119_BQ),
.O5(CLBLM_L_X12Y120_SLICE_X17Y120_AO5),
.O6(CLBLM_L_X12Y120_SLICE_X17Y120_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y121_SLICE_X16Y121_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X12Y121_SLICE_X16Y121_AO6),
.Q(CLBLM_L_X12Y121_SLICE_X16Y121_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X12Y121_SLICE_X16Y121_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X12Y121_SLICE_X16Y121_DO5),
.O6(CLBLM_L_X12Y121_SLICE_X16Y121_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X12Y121_SLICE_X16Y121_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X12Y121_SLICE_X16Y121_CO5),
.O6(CLBLM_L_X12Y121_SLICE_X16Y121_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X12Y121_SLICE_X16Y121_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X12Y121_SLICE_X16Y121_BO5),
.O6(CLBLM_L_X12Y121_SLICE_X16Y121_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hf000ff0ff000fa0a)
  ) CLBLM_L_X12Y121_SLICE_X16Y121_ALUT (
.I0(CLBLM_L_X12Y120_SLICE_X16Y120_DO6),
.I1(1'b1),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLM_R_X11Y119_SLICE_X15Y119_CQ),
.I4(CLBLM_L_X12Y120_SLICE_X17Y120_CO5),
.I5(CLBLM_R_X11Y120_SLICE_X14Y120_AO5),
.O5(CLBLM_L_X12Y121_SLICE_X16Y121_AO5),
.O6(CLBLM_L_X12Y121_SLICE_X16Y121_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X12Y121_SLICE_X17Y121_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X12Y121_SLICE_X17Y121_DO5),
.O6(CLBLM_L_X12Y121_SLICE_X17Y121_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X12Y121_SLICE_X17Y121_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X12Y121_SLICE_X17Y121_CO5),
.O6(CLBLM_L_X12Y121_SLICE_X17Y121_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X12Y121_SLICE_X17Y121_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X12Y121_SLICE_X17Y121_BO5),
.O6(CLBLM_L_X12Y121_SLICE_X17Y121_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X12Y121_SLICE_X17Y121_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X12Y121_SLICE_X17Y121_AO5),
.O6(CLBLM_L_X12Y121_SLICE_X17Y121_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y110_SLICE_X2Y110_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y111_SLICE_X2Y111_BO6),
.Q(CLBLM_R_X3Y110_SLICE_X2Y110_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y110_SLICE_X2Y110_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y110_SLICE_X2Y110_DO5),
.O6(CLBLM_R_X3Y110_SLICE_X2Y110_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y110_SLICE_X2Y110_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y110_SLICE_X2Y110_CO5),
.O6(CLBLM_R_X3Y110_SLICE_X2Y110_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y110_SLICE_X2Y110_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y110_SLICE_X2Y110_BO5),
.O6(CLBLM_R_X3Y110_SLICE_X2Y110_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y110_SLICE_X2Y110_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y110_SLICE_X2Y110_AO5),
.O6(CLBLM_R_X3Y110_SLICE_X2Y110_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y110_SLICE_X3Y110_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y110_SLICE_X3Y110_AO6),
.Q(CLBLM_R_X3Y110_SLICE_X3Y110_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y110_SLICE_X3Y110_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y110_SLICE_X3Y110_BO6),
.Q(CLBLM_R_X3Y110_SLICE_X3Y110_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y110_SLICE_X3Y110_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y110_SLICE_X3Y110_DO5),
.O6(CLBLM_R_X3Y110_SLICE_X3Y110_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y110_SLICE_X3Y110_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y110_SLICE_X3Y110_CO5),
.O6(CLBLM_R_X3Y110_SLICE_X3Y110_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hffccff4400cc0044)
  ) CLBLM_R_X3Y110_SLICE_X3Y110_BLUT (
.I0(RIOB33_X105Y117_IOB_X1Y118_I),
.I1(CLBLM_R_X3Y110_SLICE_X3Y110_BQ),
.I2(1'b1),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLM_R_X3Y118_SLICE_X2Y118_AQ),
.I5(CLBLM_R_X3Y112_SLICE_X3Y112_CQ),
.O5(CLBLM_R_X3Y110_SLICE_X3Y110_BO5),
.O6(CLBLM_R_X3Y110_SLICE_X3Y110_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hff720072ff500050)
  ) CLBLM_R_X3Y110_SLICE_X3Y110_ALUT (
.I0(CLBLL_L_X4Y111_SLICE_X4Y111_AO5),
.I1(RIOB33_X105Y105_IOB_X1Y105_I),
.I2(CLBLM_R_X3Y110_SLICE_X3Y110_AQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLM_L_X10Y110_SLICE_X13Y110_BQ),
.I5(CLBLL_L_X2Y120_SLICE_X0Y120_CO6),
.O5(CLBLM_R_X3Y110_SLICE_X3Y110_AO5),
.O6(CLBLM_R_X3Y110_SLICE_X3Y110_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y111_SLICE_X2Y111_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y111_SLICE_X2Y111_AO6),
.Q(CLBLM_R_X3Y111_SLICE_X2Y111_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y111_SLICE_X2Y111_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y111_SLICE_X2Y111_DO5),
.O6(CLBLM_R_X3Y111_SLICE_X2Y111_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hf8f8fff88888ff88)
  ) CLBLM_R_X3Y111_SLICE_X2Y111_CLUT (
.I0(CLBLM_R_X3Y120_SLICE_X3Y120_BO6),
.I1(CLBLM_R_X3Y111_SLICE_X3Y111_AO5),
.I2(CLBLM_R_X3Y117_SLICE_X2Y117_BO5),
.I3(CLBLL_L_X4Y120_SLICE_X4Y120_BO6),
.I4(CLBLM_R_X3Y111_SLICE_X2Y111_BO5),
.I5(CLBLL_L_X4Y120_SLICE_X5Y120_DO6),
.O5(CLBLM_R_X3Y111_SLICE_X2Y111_CO5),
.O6(CLBLM_R_X3Y111_SLICE_X2Y111_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hffcc00ccf7f7f7f7)
  ) CLBLM_R_X3Y111_SLICE_X2Y111_BLUT (
.I0(RIOB33_X105Y105_IOB_X1Y105_I),
.I1(CLBLL_L_X4Y121_SLICE_X4Y121_BQ),
.I2(CLBLM_R_X3Y110_SLICE_X2Y110_AQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLM_R_X3Y110_SLICE_X3Y110_AQ),
.I5(1'b1),
.O5(CLBLM_R_X3Y111_SLICE_X2Y111_BO5),
.O6(CLBLM_R_X3Y111_SLICE_X2Y111_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffaaaaaaffa0a0a0)
  ) CLBLM_R_X3Y111_SLICE_X2Y111_ALUT (
.I0(CLBLM_R_X5Y115_SLICE_X6Y115_CO6),
.I1(1'b1),
.I2(CLBLM_R_X3Y111_SLICE_X2Y111_AQ),
.I3(CLBLM_R_X7Y124_SLICE_X8Y124_CQ),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(CLBLL_L_X4Y111_SLICE_X5Y111_A5Q),
.O5(CLBLM_R_X3Y111_SLICE_X2Y111_AO5),
.O6(CLBLM_R_X3Y111_SLICE_X2Y111_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y111_SLICE_X3Y111_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y111_SLICE_X3Y111_AO6),
.Q(CLBLM_R_X3Y111_SLICE_X3Y111_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y111_SLICE_X3Y111_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y111_SLICE_X3Y111_BO6),
.Q(CLBLM_R_X3Y111_SLICE_X3Y111_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h33b300a033330000)
  ) CLBLM_R_X3Y111_SLICE_X3Y111_DLUT (
.I0(CLBLM_R_X3Y115_SLICE_X3Y115_CQ),
.I1(CLBLM_L_X8Y112_SLICE_X11Y112_AQ),
.I2(CLBLL_L_X4Y120_SLICE_X5Y120_DO6),
.I3(CLBLM_R_X7Y115_SLICE_X9Y115_C5Q),
.I4(CLBLL_L_X2Y120_SLICE_X1Y120_DO6),
.I5(RIOB33_X105Y105_IOB_X1Y105_I),
.O5(CLBLM_R_X3Y111_SLICE_X3Y111_DO5),
.O6(CLBLM_R_X3Y111_SLICE_X3Y111_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h1155b1f55555f5f5)
  ) CLBLM_R_X3Y111_SLICE_X3Y111_CLUT (
.I0(RIOB33_X105Y105_IOB_X1Y105_I),
.I1(CLBLM_L_X8Y112_SLICE_X10Y112_CQ),
.I2(CLBLM_R_X3Y116_SLICE_X3Y116_DO6),
.I3(CLBLM_R_X3Y119_SLICE_X2Y119_AO6),
.I4(CLBLM_R_X3Y111_SLICE_X3Y111_DO6),
.I5(CLBLL_L_X2Y112_SLICE_X1Y112_BQ),
.O5(CLBLM_R_X3Y111_SLICE_X3Y111_CO5),
.O6(CLBLM_R_X3Y111_SLICE_X3Y111_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f00000f3fc030c)
  ) CLBLM_R_X3Y111_SLICE_X3Y111_BLUT (
.I0(1'b1),
.I1(CLBLM_R_X3Y111_SLICE_X3Y111_BQ),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLM_R_X3Y113_SLICE_X3Y113_BO6),
.I4(CLBLM_L_X10Y117_SLICE_X13Y117_BQ),
.I5(CLBLM_R_X5Y110_SLICE_X7Y110_BQ),
.O5(CLBLM_R_X3Y111_SLICE_X3Y111_BO5),
.O6(CLBLM_R_X3Y111_SLICE_X3Y111_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfccc3000aa00aa00)
  ) CLBLM_R_X3Y111_SLICE_X3Y111_ALUT (
.I0(CLBLL_L_X2Y113_SLICE_X1Y113_C5Q),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(CLBLM_R_X3Y111_SLICE_X3Y111_AQ),
.I3(RIOB33_X105Y105_IOB_X1Y105_I),
.I4(CLBLL_L_X4Y110_SLICE_X4Y110_DQ),
.I5(1'b1),
.O5(CLBLM_R_X3Y111_SLICE_X3Y111_AO5),
.O6(CLBLM_R_X3Y111_SLICE_X3Y111_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y112_SLICE_X2Y112_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y112_SLICE_X2Y112_AO6),
.Q(CLBLM_R_X3Y112_SLICE_X2Y112_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y112_SLICE_X2Y112_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y112_SLICE_X2Y112_BO6),
.Q(CLBLM_R_X3Y112_SLICE_X2Y112_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'ha2a2aaa2a2a2aaa2)
  ) CLBLM_R_X3Y112_SLICE_X2Y112_DLUT (
.I0(RIOB33_X105Y105_IOB_X1Y105_I),
.I1(CLBLM_R_X7Y120_SLICE_X9Y120_DQ),
.I2(CLBLM_R_X7Y113_SLICE_X9Y113_A5Q),
.I3(CLBLM_R_X3Y115_SLICE_X3Y115_CQ),
.I4(CLBLM_R_X7Y115_SLICE_X9Y115_C5Q),
.I5(1'b1),
.O5(CLBLM_R_X3Y112_SLICE_X2Y112_DO5),
.O6(CLBLM_R_X3Y112_SLICE_X2Y112_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff7555ffff7755)
  ) CLBLM_R_X3Y112_SLICE_X2Y112_CLUT (
.I0(RIOB33_X105Y105_IOB_X1Y105_I),
.I1(CLBLM_R_X7Y113_SLICE_X9Y113_A5Q),
.I2(CLBLM_R_X7Y115_SLICE_X9Y115_C5Q),
.I3(CLBLM_R_X7Y120_SLICE_X9Y120_DQ),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(CLBLM_R_X3Y115_SLICE_X3Y115_CQ),
.O5(CLBLM_R_X3Y112_SLICE_X2Y112_CO5),
.O6(CLBLM_R_X3Y112_SLICE_X2Y112_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hff880088ff280028)
  ) CLBLM_R_X3Y112_SLICE_X2Y112_BLUT (
.I0(CLBLM_R_X3Y112_SLICE_X2Y112_DO6),
.I1(CLBLM_R_X3Y112_SLICE_X2Y112_BQ),
.I2(CLBLM_R_X3Y112_SLICE_X2Y112_AQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLM_R_X11Y116_SLICE_X14Y116_AQ),
.I5(CLBLL_L_X2Y112_SLICE_X1Y112_CO5),
.O5(CLBLM_R_X3Y112_SLICE_X2Y112_BO5),
.O6(CLBLM_R_X3Y112_SLICE_X2Y112_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hcca0cca0cc0acc0a)
  ) CLBLM_R_X3Y112_SLICE_X2Y112_ALUT (
.I0(CLBLM_R_X3Y112_SLICE_X2Y112_DO6),
.I1(CLBLM_R_X7Y110_SLICE_X9Y110_CQ),
.I2(CLBLM_R_X3Y112_SLICE_X2Y112_AQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(1'b1),
.I5(CLBLL_L_X2Y112_SLICE_X1Y112_CO5),
.O5(CLBLM_R_X3Y112_SLICE_X2Y112_AO5),
.O6(CLBLM_R_X3Y112_SLICE_X2Y112_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y112_SLICE_X3Y112_B5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y112_SLICE_X3Y112_BO5),
.Q(CLBLM_R_X3Y112_SLICE_X3Y112_B5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "C5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y112_SLICE_X3Y112_C5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y112_SLICE_X3Y112_CO5),
.Q(CLBLM_R_X3Y112_SLICE_X3Y112_C5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y112_SLICE_X3Y112_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y112_SLICE_X3Y112_AO6),
.Q(CLBLM_R_X3Y112_SLICE_X3Y112_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y112_SLICE_X3Y112_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y112_SLICE_X3Y112_BO6),
.Q(CLBLM_R_X3Y112_SLICE_X3Y112_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y112_SLICE_X3Y112_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y112_SLICE_X3Y112_CO6),
.Q(CLBLM_R_X3Y112_SLICE_X3Y112_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h2222222212222222)
  ) CLBLM_R_X3Y112_SLICE_X3Y112_DLUT (
.I0(CLBLM_R_X3Y112_SLICE_X3Y112_C5Q),
.I1(CLBLM_R_X3Y112_SLICE_X2Y112_CO6),
.I2(CLBLM_R_X3Y112_SLICE_X2Y112_BQ),
.I3(CLBLM_R_X3Y112_SLICE_X2Y112_AQ),
.I4(CLBLL_L_X2Y112_SLICE_X1Y112_A5Q),
.I5(CLBLM_L_X10Y113_SLICE_X13Y113_BO6),
.O5(CLBLM_R_X3Y112_SLICE_X3Y112_DO5),
.O6(CLBLM_R_X3Y112_SLICE_X3Y112_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hee44ee44ffffa0a0)
  ) CLBLM_R_X3Y112_SLICE_X3Y112_CLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_R_X3Y119_SLICE_X2Y119_AO6),
.I2(CLBLL_L_X4Y115_SLICE_X4Y115_AQ),
.I3(CLBLL_L_X2Y112_SLICE_X1Y112_AQ),
.I4(CLBLM_R_X3Y112_SLICE_X3Y112_DO6),
.I5(1'b1),
.O5(CLBLM_R_X3Y112_SLICE_X3Y112_CO5),
.O6(CLBLM_R_X3Y112_SLICE_X3Y112_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hff0a000aaaccaacc)
  ) CLBLM_R_X3Y112_SLICE_X3Y112_BLUT (
.I0(CLBLL_L_X4Y111_SLICE_X5Y111_A5Q),
.I1(CLBLL_L_X2Y112_SLICE_X1Y112_AQ),
.I2(RIOB33_X105Y105_IOB_X1Y105_I),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLM_R_X7Y113_SLICE_X9Y113_AQ),
.I5(1'b1),
.O5(CLBLM_R_X3Y112_SLICE_X3Y112_BO5),
.O6(CLBLM_R_X3Y112_SLICE_X3Y112_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaabefa00001450)
  ) CLBLM_R_X3Y112_SLICE_X3Y112_ALUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_R_X3Y113_SLICE_X3Y113_BO6),
.I2(CLBLM_R_X3Y112_SLICE_X3Y112_AQ),
.I3(CLBLM_R_X3Y111_SLICE_X3Y111_BQ),
.I4(CLBLM_R_X5Y110_SLICE_X7Y110_BQ),
.I5(CLBLM_R_X7Y115_SLICE_X8Y115_CQ),
.O5(CLBLM_R_X3Y112_SLICE_X3Y112_AO5),
.O6(CLBLM_R_X3Y112_SLICE_X3Y112_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y113_SLICE_X2Y113_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y113_SLICE_X2Y113_AO6),
.Q(CLBLM_R_X3Y113_SLICE_X2Y113_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y113_SLICE_X2Y113_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y113_SLICE_X2Y113_BO6),
.Q(CLBLM_R_X3Y113_SLICE_X2Y113_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'ha0a000005555ffff)
  ) CLBLM_R_X3Y113_SLICE_X2Y113_DLUT (
.I0(CLBLM_R_X5Y113_SLICE_X6Y113_BQ),
.I1(1'b1),
.I2(CLBLL_L_X4Y113_SLICE_X4Y113_CO6),
.I3(1'b1),
.I4(CLBLL_L_X4Y113_SLICE_X4Y113_AQ),
.I5(1'b1),
.O5(CLBLM_R_X3Y113_SLICE_X2Y113_DO5),
.O6(CLBLM_R_X3Y113_SLICE_X2Y113_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h8000000088000000)
  ) CLBLM_R_X3Y113_SLICE_X2Y113_CLUT (
.I0(CLBLM_R_X5Y113_SLICE_X6Y113_BQ),
.I1(CLBLL_L_X4Y113_SLICE_X4Y113_CO6),
.I2(CLBLM_R_X3Y114_SLICE_X2Y114_DQ),
.I3(CLBLM_R_X3Y113_SLICE_X2Y113_BQ),
.I4(CLBLL_L_X4Y113_SLICE_X4Y113_AQ),
.I5(1'b1),
.O5(CLBLM_R_X3Y113_SLICE_X2Y113_CO5),
.O6(CLBLM_R_X3Y113_SLICE_X2Y113_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f0f0fe0000000e)
  ) CLBLM_R_X3Y113_SLICE_X2Y113_BLUT (
.I0(CLBLM_R_X3Y113_SLICE_X2Y113_DO6),
.I1(CLBLM_R_X3Y113_SLICE_X2Y113_BQ),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLM_R_X5Y110_SLICE_X7Y110_BQ),
.I4(CLBLM_R_X3Y113_SLICE_X2Y113_CO5),
.I5(CLBLM_L_X8Y112_SLICE_X10Y112_CQ),
.O5(CLBLM_R_X3Y113_SLICE_X2Y113_BO5),
.O6(CLBLM_R_X3Y113_SLICE_X2Y113_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffc00fcffa800a8)
  ) CLBLM_R_X3Y113_SLICE_X2Y113_ALUT (
.I0(RIOB33_X105Y117_IOB_X1Y118_I),
.I1(CLBLM_R_X5Y112_SLICE_X6Y112_DO6),
.I2(CLBLM_R_X3Y113_SLICE_X2Y113_AQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLM_R_X3Y112_SLICE_X2Y112_BQ),
.I5(CLBLM_R_X3Y118_SLICE_X2Y118_AQ),
.O5(CLBLM_R_X3Y113_SLICE_X2Y113_AO5),
.O6(CLBLM_R_X3Y113_SLICE_X2Y113_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y113_SLICE_X3Y113_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y113_SLICE_X3Y113_AO6),
.Q(CLBLM_R_X3Y113_SLICE_X3Y113_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h7f770f00ff77ff00)
  ) CLBLM_R_X3Y113_SLICE_X3Y113_DLUT (
.I0(CLBLM_R_X3Y111_SLICE_X3Y111_BQ),
.I1(CLBLM_R_X3Y112_SLICE_X3Y112_AQ),
.I2(CLBLM_R_X3Y114_SLICE_X2Y114_DQ),
.I3(CLBLM_R_X3Y113_SLICE_X2Y113_DO5),
.I4(CLBLM_R_X3Y113_SLICE_X3Y113_BO5),
.I5(CLBLM_R_X3Y113_SLICE_X2Y113_BQ),
.O5(CLBLM_R_X3Y113_SLICE_X3Y113_DO5),
.O6(CLBLM_R_X3Y113_SLICE_X3Y113_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffbfffffffff)
  ) CLBLM_R_X3Y113_SLICE_X3Y113_CLUT (
.I0(CLBLM_R_X3Y112_SLICE_X3Y112_AQ),
.I1(CLBLM_R_X3Y117_SLICE_X3Y117_C5Q),
.I2(CLBLM_R_X3Y114_SLICE_X2Y114_DQ),
.I3(CLBLM_R_X3Y113_SLICE_X2Y113_DO5),
.I4(CLBLM_R_X3Y113_SLICE_X3Y113_BO5),
.I5(CLBLM_R_X3Y113_SLICE_X2Y113_BQ),
.O5(CLBLM_R_X3Y113_SLICE_X3Y113_CO5),
.O6(CLBLM_R_X3Y113_SLICE_X3Y113_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h202000000f0fffff)
  ) CLBLM_R_X3Y113_SLICE_X3Y113_BLUT (
.I0(RIOB33_X105Y117_IOB_X1Y118_I),
.I1(CLBLM_R_X3Y118_SLICE_X2Y118_AQ),
.I2(CLBLL_L_X4Y118_SLICE_X5Y118_AQ),
.I3(1'b1),
.I4(CLBLM_R_X5Y116_SLICE_X6Y116_BQ),
.I5(1'b1),
.O5(CLBLM_R_X3Y113_SLICE_X3Y113_BO5),
.O6(CLBLM_R_X3Y113_SLICE_X3Y113_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hccfe0032fefe3232)
  ) CLBLM_R_X3Y113_SLICE_X3Y113_ALUT (
.I0(CLBLM_R_X3Y114_SLICE_X2Y114_DQ),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(CLBLM_R_X3Y113_SLICE_X3Y113_AQ),
.I3(CLBLL_L_X2Y112_SLICE_X1Y112_BQ),
.I4(CLBLM_R_X3Y117_SLICE_X3Y117_C5Q),
.I5(CLBLM_L_X8Y112_SLICE_X10Y112_CQ),
.O5(CLBLM_R_X3Y113_SLICE_X3Y113_AO5),
.O6(CLBLM_R_X3Y113_SLICE_X3Y113_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y114_SLICE_X2Y114_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y114_SLICE_X2Y114_AO6),
.Q(CLBLM_R_X3Y114_SLICE_X2Y114_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y114_SLICE_X2Y114_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y114_SLICE_X2Y114_BO6),
.Q(CLBLM_R_X3Y114_SLICE_X2Y114_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y114_SLICE_X2Y114_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y114_SLICE_X2Y114_CO6),
.Q(CLBLM_R_X3Y114_SLICE_X2Y114_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y114_SLICE_X2Y114_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y114_SLICE_X2Y114_DO6),
.Q(CLBLM_R_X3Y114_SLICE_X2Y114_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff003200000032)
  ) CLBLM_R_X3Y114_SLICE_X2Y114_DLUT (
.I0(CLBLM_R_X3Y113_SLICE_X2Y113_CO5),
.I1(CLBLM_R_X3Y113_SLICE_X2Y113_CO6),
.I2(CLBLM_R_X3Y114_SLICE_X2Y114_DQ),
.I3(CLBLM_R_X5Y110_SLICE_X7Y110_BQ),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(CLBLL_L_X4Y118_SLICE_X5Y118_AQ),
.O5(CLBLM_R_X3Y114_SLICE_X2Y114_DO5),
.O6(CLBLM_R_X3Y114_SLICE_X2Y114_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'haaef00cfaaeb00c3)
  ) CLBLM_R_X3Y114_SLICE_X2Y114_CLUT (
.I0(CLBLM_R_X7Y123_SLICE_X8Y123_AQ),
.I1(CLBLM_R_X3Y114_SLICE_X2Y114_CQ),
.I2(CLBLM_R_X5Y111_SLICE_X7Y111_DO6),
.I3(CLBLM_R_X3Y114_SLICE_X2Y114_AO5),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(CLBLL_L_X2Y114_SLICE_X1Y114_BO5),
.O5(CLBLM_R_X3Y114_SLICE_X2Y114_CO5),
.O6(CLBLM_R_X3Y114_SLICE_X2Y114_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffcccf000f000)
  ) CLBLM_R_X3Y114_SLICE_X2Y114_BLUT (
.I0(1'b1),
.I1(CLBLM_R_X3Y114_SLICE_X2Y114_BQ),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLM_R_X3Y114_SLICE_X2Y114_CQ),
.I4(CLBLM_R_X3Y112_SLICE_X3Y112_BQ),
.I5(CLBLM_R_X5Y115_SLICE_X6Y115_CO6),
.O5(CLBLM_R_X3Y114_SLICE_X2Y114_BO5),
.O6(CLBLM_R_X3Y114_SLICE_X2Y114_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hc0c0d1c0eeffeeff)
  ) CLBLM_R_X3Y114_SLICE_X2Y114_ALUT (
.I0(CLBLM_R_X5Y115_SLICE_X7Y115_AQ),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(CLBLM_R_X11Y115_SLICE_X15Y115_AQ),
.I3(RIOB33_X105Y105_IOB_X1Y105_I),
.I4(CLBLL_L_X2Y114_SLICE_X1Y114_BO6),
.I5(1'b1),
.O5(CLBLM_R_X3Y114_SLICE_X2Y114_AO5),
.O6(CLBLM_R_X3Y114_SLICE_X2Y114_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y114_SLICE_X3Y114_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y114_SLICE_X3Y114_AO6),
.Q(CLBLM_R_X3Y114_SLICE_X3Y114_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y114_SLICE_X3Y114_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y114_SLICE_X3Y114_BO6),
.Q(CLBLM_R_X3Y114_SLICE_X3Y114_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y114_SLICE_X3Y114_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y114_SLICE_X3Y114_CO6),
.Q(CLBLM_R_X3Y114_SLICE_X3Y114_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hff0f0f0fff0f0f0f)
  ) CLBLM_R_X3Y114_SLICE_X3Y114_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(RIOB33_X105Y121_IOB_X1Y121_I),
.I3(CLBLM_R_X3Y114_SLICE_X3Y114_AQ),
.I4(CLBLM_R_X7Y115_SLICE_X8Y115_CQ),
.I5(1'b1),
.O5(CLBLM_R_X3Y114_SLICE_X3Y114_DO5),
.O6(CLBLM_R_X3Y114_SLICE_X3Y114_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hff55ef45ba10aa00)
  ) CLBLM_R_X3Y114_SLICE_X3Y114_CLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_L_X10Y113_SLICE_X13Y113_BO6),
.I2(CLBLM_R_X7Y119_SLICE_X8Y119_D5Q),
.I3(CLBLM_R_X11Y113_SLICE_X15Y113_BQ),
.I4(CLBLM_R_X3Y114_SLICE_X3Y114_CQ),
.I5(CLBLM_R_X5Y116_SLICE_X6Y116_BQ),
.O5(CLBLM_R_X3Y114_SLICE_X3Y114_CO5),
.O6(CLBLM_R_X3Y114_SLICE_X3Y114_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'ha0a0aca0a0a0a0a0)
  ) CLBLM_R_X3Y114_SLICE_X3Y114_BLUT (
.I0(CLBLL_L_X4Y119_SLICE_X4Y119_DQ),
.I1(CLBLM_R_X3Y117_SLICE_X3Y117_BQ),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLM_R_X3Y115_SLICE_X2Y115_BQ),
.I4(CLBLM_R_X3Y113_SLICE_X3Y113_CO6),
.I5(CLBLM_R_X3Y111_SLICE_X3Y111_BQ),
.O5(CLBLM_R_X3Y114_SLICE_X3Y114_BO5),
.O6(CLBLM_R_X3Y114_SLICE_X3Y114_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hb8b8b8bbb8b8b888)
  ) CLBLM_R_X3Y114_SLICE_X3Y114_ALUT (
.I0(CLBLM_R_X3Y114_SLICE_X3Y114_CQ),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(CLBLL_L_X4Y114_SLICE_X4Y114_DO6),
.I3(RIOB33_X105Y117_IOB_X1Y118_I),
.I4(CLBLM_R_X3Y118_SLICE_X2Y118_AQ),
.I5(CLBLM_R_X3Y114_SLICE_X3Y114_AQ),
.O5(CLBLM_R_X3Y114_SLICE_X3Y114_AO5),
.O6(CLBLM_R_X3Y114_SLICE_X3Y114_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y115_SLICE_X2Y115_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y115_SLICE_X2Y115_AO6),
.Q(CLBLM_R_X3Y115_SLICE_X2Y115_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y115_SLICE_X2Y115_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y115_SLICE_X2Y115_BO6),
.Q(CLBLM_R_X3Y115_SLICE_X2Y115_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y115_SLICE_X2Y115_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y115_SLICE_X2Y115_CO6),
.Q(CLBLM_R_X3Y115_SLICE_X2Y115_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y115_SLICE_X2Y115_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y115_SLICE_X2Y115_DO6),
.Q(CLBLM_R_X3Y115_SLICE_X2Y115_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hd8d8ddddd888dd88)
  ) CLBLM_R_X3Y115_SLICE_X2Y115_DLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_R_X3Y113_SLICE_X2Y113_BQ),
.I2(CLBLM_L_X10Y113_SLICE_X13Y113_BO6),
.I3(CLBLM_R_X3Y115_SLICE_X2Y115_DQ),
.I4(CLBLM_R_X7Y119_SLICE_X8Y119_D5Q),
.I5(CLBLM_R_X5Y113_SLICE_X6Y113_BQ),
.O5(CLBLM_R_X3Y115_SLICE_X2Y115_DO5),
.O6(CLBLM_R_X3Y115_SLICE_X2Y115_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hafaa0500aeaa0400)
  ) CLBLM_R_X3Y115_SLICE_X2Y115_CLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_R_X3Y115_SLICE_X2Y115_CQ),
.I2(RIOB33_X105Y117_IOB_X1Y118_I),
.I3(CLBLM_R_X3Y118_SLICE_X2Y118_AQ),
.I4(CLBLM_R_X7Y121_SLICE_X8Y121_C5Q),
.I5(CLBLM_R_X11Y115_SLICE_X14Y115_BQ),
.O5(CLBLM_R_X3Y115_SLICE_X2Y115_CO5),
.O6(CLBLM_R_X3Y115_SLICE_X2Y115_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f30003f0fc000c)
  ) CLBLM_R_X3Y115_SLICE_X2Y115_BLUT (
.I0(1'b1),
.I1(CLBLM_R_X3Y115_SLICE_X2Y115_BQ),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLM_R_X5Y110_SLICE_X7Y110_BQ),
.I4(CLBLM_R_X3Y118_SLICE_X3Y118_AQ),
.I5(CLBLM_R_X3Y113_SLICE_X2Y113_CO6),
.O5(CLBLM_R_X3Y115_SLICE_X2Y115_BO5),
.O6(CLBLM_R_X3Y115_SLICE_X2Y115_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfff0ffcc00f000cc)
  ) CLBLM_R_X3Y115_SLICE_X2Y115_ALUT (
.I0(1'b1),
.I1(CLBLL_L_X4Y112_SLICE_X4Y112_BQ),
.I2(CLBLM_R_X3Y115_SLICE_X2Y115_AQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLM_R_X5Y115_SLICE_X6Y115_CO5),
.I5(CLBLM_R_X3Y115_SLICE_X2Y115_DQ),
.O5(CLBLM_R_X3Y115_SLICE_X2Y115_AO5),
.O6(CLBLM_R_X3Y115_SLICE_X2Y115_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y115_SLICE_X3Y115_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y115_SLICE_X3Y115_AO6),
.Q(CLBLM_R_X3Y115_SLICE_X3Y115_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y115_SLICE_X3Y115_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y115_SLICE_X3Y115_BO6),
.Q(CLBLM_R_X3Y115_SLICE_X3Y115_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y115_SLICE_X3Y115_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y115_SLICE_X3Y115_CO6),
.Q(CLBLM_R_X3Y115_SLICE_X3Y115_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y115_SLICE_X3Y115_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y115_SLICE_X3Y115_DO6),
.Q(CLBLM_R_X3Y115_SLICE_X3Y115_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hc0c0c5c5c5c5c0c0)
  ) CLBLM_R_X3Y115_SLICE_X3Y115_DLUT (
.I0(RIOB33_X105Y105_IOB_X1Y105_I),
.I1(CLBLM_R_X3Y117_SLICE_X3Y117_A5Q),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(1'b1),
.I4(CLBLM_R_X3Y114_SLICE_X3Y114_DO6),
.I5(CLBLL_L_X4Y112_SLICE_X4Y112_BQ),
.O5(CLBLM_R_X3Y115_SLICE_X3Y115_DO5),
.O6(CLBLM_R_X3Y115_SLICE_X3Y115_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'he4a0a0a0a0a0a0a0)
  ) CLBLM_R_X3Y115_SLICE_X3Y115_CLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_R_X3Y112_SLICE_X2Y112_BQ),
.I2(CLBLL_L_X4Y115_SLICE_X4Y115_C5Q),
.I3(CLBLM_R_X3Y112_SLICE_X3Y112_C5Q),
.I4(CLBLL_L_X2Y112_SLICE_X1Y112_A5Q),
.I5(CLBLM_R_X3Y112_SLICE_X2Y112_AQ),
.O5(CLBLM_R_X3Y115_SLICE_X3Y115_CO5),
.O6(CLBLM_R_X3Y115_SLICE_X3Y115_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffc00fc00fc00)
  ) CLBLM_R_X3Y115_SLICE_X3Y115_BLUT (
.I0(1'b1),
.I1(CLBLM_R_X3Y115_SLICE_X3Y115_BQ),
.I2(CLBLL_L_X4Y111_SLICE_X5Y111_BQ),
.I3(CLBLM_R_X5Y115_SLICE_X6Y115_CO6),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(CLBLM_R_X3Y116_SLICE_X3Y116_A5Q),
.O5(CLBLM_R_X3Y115_SLICE_X3Y115_BO5),
.O6(CLBLM_R_X3Y115_SLICE_X3Y115_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hbbfb1151aaea0040)
  ) CLBLM_R_X3Y115_SLICE_X3Y115_ALUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLL_L_X4Y111_SLICE_X4Y111_AO5),
.I2(CLBLM_R_X3Y120_SLICE_X3Y120_BO6),
.I3(RIOB33_X105Y105_IOB_X1Y105_I),
.I4(CLBLL_L_X4Y112_SLICE_X4Y112_BQ),
.I5(CLBLM_R_X3Y115_SLICE_X3Y115_AQ),
.O5(CLBLM_R_X3Y115_SLICE_X3Y115_AO5),
.O6(CLBLM_R_X3Y115_SLICE_X3Y115_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y116_SLICE_X2Y116_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y116_SLICE_X2Y116_AO6),
.Q(CLBLM_R_X3Y116_SLICE_X2Y116_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y116_SLICE_X2Y116_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y116_SLICE_X2Y116_BO6),
.Q(CLBLM_R_X3Y116_SLICE_X2Y116_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h000c004c00000000)
  ) CLBLM_R_X3Y116_SLICE_X2Y116_DLUT (
.I0(CLBLL_L_X2Y113_SLICE_X1Y113_C5Q),
.I1(CLBLL_L_X2Y114_SLICE_X1Y114_BO5),
.I2(RIOB33_X105Y105_IOB_X1Y105_I),
.I3(CLBLM_L_X8Y116_SLICE_X10Y116_AO6),
.I4(CLBLM_R_X3Y117_SLICE_X2Y117_BO5),
.I5(CLBLM_R_X5Y111_SLICE_X7Y111_DO6),
.O5(CLBLM_R_X3Y116_SLICE_X2Y116_DO5),
.O6(CLBLM_R_X3Y116_SLICE_X2Y116_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff0f2fffff0f3f)
  ) CLBLM_R_X3Y116_SLICE_X2Y116_CLUT (
.I0(CLBLM_R_X3Y110_SLICE_X2Y110_AQ),
.I1(LIOB33_X0Y53_IOB_X0Y53_I),
.I2(RIOB33_X105Y105_IOB_X1Y105_I),
.I3(CLBLM_R_X3Y117_SLICE_X3Y117_A5Q),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(CLBLL_L_X4Y121_SLICE_X4Y121_BQ),
.O5(CLBLM_R_X3Y116_SLICE_X2Y116_CO5),
.O6(CLBLM_R_X3Y116_SLICE_X2Y116_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfefeaaaafcfc0000)
  ) CLBLM_R_X3Y116_SLICE_X2Y116_BLUT (
.I0(CLBLL_L_X4Y116_SLICE_X4Y116_CQ),
.I1(CLBLM_R_X3Y116_SLICE_X2Y116_BQ),
.I2(CLBLM_R_X5Y111_SLICE_X6Y111_CQ),
.I3(1'b1),
.I4(CLBLM_R_X5Y115_SLICE_X6Y115_CO6),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLM_R_X3Y116_SLICE_X2Y116_BO5),
.O6(CLBLM_R_X3Y116_SLICE_X2Y116_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfbfbf1fb0b0b010b)
  ) CLBLM_R_X3Y116_SLICE_X2Y116_ALUT (
.I0(RIOB33_X105Y105_IOB_X1Y105_I),
.I1(LIOB33_X0Y53_IOB_X0Y53_I),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLL_L_X4Y121_SLICE_X4Y121_BQ),
.I4(CLBLM_R_X3Y110_SLICE_X2Y110_AQ),
.I5(CLBLM_R_X11Y115_SLICE_X14Y115_BQ),
.O5(CLBLM_R_X3Y116_SLICE_X2Y116_AO5),
.O6(CLBLM_R_X3Y116_SLICE_X2Y116_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y116_SLICE_X3Y116_A5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y116_SLICE_X13Y116_AO6),
.Q(CLBLM_R_X3Y116_SLICE_X3Y116_A5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y116_SLICE_X3Y116_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y116_SLICE_X3Y116_AO6),
.Q(CLBLM_R_X3Y116_SLICE_X3Y116_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y116_SLICE_X3Y116_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y116_SLICE_X3Y116_BO6),
.Q(CLBLM_R_X3Y116_SLICE_X3Y116_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y116_SLICE_X3Y116_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y116_SLICE_X3Y116_CO6),
.Q(CLBLM_R_X3Y116_SLICE_X3Y116_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h2a3f2a3f2a3f2a3f)
  ) CLBLM_R_X3Y116_SLICE_X3Y116_DLUT (
.I0(CLBLL_L_X2Y119_SLICE_X0Y119_BO6),
.I1(CLBLM_R_X7Y113_SLICE_X9Y113_A5Q),
.I2(CLBLM_R_X3Y120_SLICE_X3Y120_BO6),
.I3(CLBLM_R_X5Y124_SLICE_X6Y124_CQ),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y116_SLICE_X3Y116_DO5),
.O6(CLBLM_R_X3Y116_SLICE_X3Y116_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaacfc0aaaacfc0)
  ) CLBLM_R_X3Y116_SLICE_X3Y116_CLUT (
.I0(CLBLL_L_X4Y114_SLICE_X5Y114_AQ),
.I1(CLBLM_R_X3Y116_SLICE_X3Y116_CQ),
.I2(CLBLM_R_X3Y116_SLICE_X2Y116_DO6),
.I3(CLBLM_R_X5Y119_SLICE_X6Y119_B5Q),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(1'b1),
.O5(CLBLM_R_X3Y116_SLICE_X3Y116_CO5),
.O6(CLBLM_R_X3Y116_SLICE_X3Y116_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfafa0a0af0f00000)
  ) CLBLM_R_X3Y116_SLICE_X3Y116_BLUT (
.I0(RIOB33_X105Y105_IOB_X1Y105_I),
.I1(1'b1),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(1'b1),
.I4(CLBLL_L_X2Y117_SLICE_X1Y117_AQ),
.I5(CLBLM_R_X5Y115_SLICE_X7Y115_BQ),
.O5(CLBLM_R_X3Y116_SLICE_X3Y116_BO5),
.O6(CLBLM_R_X3Y116_SLICE_X3Y116_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hbb11aa00ba10aa00)
  ) CLBLM_R_X3Y116_SLICE_X3Y116_ALUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(RIOB33_X105Y117_IOB_X1Y118_I),
.I2(CLBLM_R_X3Y116_SLICE_X3Y116_AQ),
.I3(CLBLL_L_X4Y121_SLICE_X4Y121_BQ),
.I4(CLBLM_R_X3Y118_SLICE_X2Y118_AQ),
.I5(CLBLM_R_X11Y113_SLICE_X14Y113_BQ),
.O5(CLBLM_R_X3Y116_SLICE_X3Y116_AO5),
.O6(CLBLM_R_X3Y116_SLICE_X3Y116_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y117_SLICE_X2Y117_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y117_SLICE_X2Y117_AO6),
.Q(CLBLM_R_X3Y117_SLICE_X2Y117_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h050d050d000c000c)
  ) CLBLM_R_X3Y117_SLICE_X2Y117_DLUT (
.I0(CLBLL_L_X2Y120_SLICE_X1Y120_AO6),
.I1(CLBLL_L_X4Y114_SLICE_X4Y114_AQ),
.I2(CLBLM_R_X3Y122_SLICE_X3Y122_AO6),
.I3(CLBLL_L_X2Y121_SLICE_X1Y121_BO6),
.I4(1'b1),
.I5(CLBLM_R_X3Y114_SLICE_X2Y114_BQ),
.O5(CLBLM_R_X3Y117_SLICE_X2Y117_DO5),
.O6(CLBLM_R_X3Y117_SLICE_X2Y117_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h00000000000c000a)
  ) CLBLM_R_X3Y117_SLICE_X2Y117_CLUT (
.I0(CLBLM_R_X5Y116_SLICE_X6Y116_AQ),
.I1(CLBLM_R_X3Y114_SLICE_X3Y114_CQ),
.I2(CLBLM_R_X3Y122_SLICE_X3Y122_AO5),
.I3(CLBLL_L_X2Y120_SLICE_X1Y120_AO6),
.I4(RIOB33_X105Y135_IOB_X1Y136_I),
.I5(RIOB33_X105Y135_IOB_X1Y135_I),
.O5(CLBLM_R_X3Y117_SLICE_X2Y117_CO5),
.O6(CLBLM_R_X3Y117_SLICE_X2Y117_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hae00ff000c0c0c0c)
  ) CLBLM_R_X3Y117_SLICE_X2Y117_BLUT (
.I0(CLBLL_L_X2Y113_SLICE_X1Y113_C5Q),
.I1(CLBLL_L_X2Y117_SLICE_X0Y117_A5Q),
.I2(CLBLM_R_X7Y121_SLICE_X8Y121_C5Q),
.I3(RIOB33_X105Y105_IOB_X1Y105_I),
.I4(CLBLM_R_X5Y115_SLICE_X7Y115_AQ),
.I5(1'b1),
.O5(CLBLM_R_X3Y117_SLICE_X2Y117_BO5),
.O6(CLBLM_R_X3Y117_SLICE_X2Y117_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hccccaaffcccca0f0)
  ) CLBLM_R_X3Y117_SLICE_X2Y117_ALUT (
.I0(CLBLM_L_X10Y113_SLICE_X13Y113_BO6),
.I1(CLBLM_R_X7Y128_SLICE_X8Y128_AQ),
.I2(CLBLM_R_X3Y117_SLICE_X2Y117_AQ),
.I3(CLBLM_R_X7Y119_SLICE_X8Y119_D5Q),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(CLBLM_R_X3Y114_SLICE_X2Y114_DQ),
.O5(CLBLM_R_X3Y117_SLICE_X2Y117_AO5),
.O6(CLBLM_R_X3Y117_SLICE_X2Y117_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y117_SLICE_X3Y117_A5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y117_SLICE_X3Y117_AO5),
.Q(CLBLM_R_X3Y117_SLICE_X3Y117_A5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y117_SLICE_X3Y117_B5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y117_SLICE_X3Y117_BO5),
.Q(CLBLM_R_X3Y117_SLICE_X3Y117_B5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "C5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y117_SLICE_X3Y117_C5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y117_SLICE_X3Y117_CO5),
.Q(CLBLM_R_X3Y117_SLICE_X3Y117_C5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y117_SLICE_X3Y117_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y117_SLICE_X3Y117_AO6),
.Q(CLBLM_R_X3Y117_SLICE_X3Y117_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y117_SLICE_X3Y117_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y117_SLICE_X3Y117_BO6),
.Q(CLBLM_R_X3Y117_SLICE_X3Y117_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y117_SLICE_X3Y117_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y117_SLICE_X3Y117_CO6),
.Q(CLBLM_R_X3Y117_SLICE_X3Y117_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000003202)
  ) CLBLM_R_X3Y117_SLICE_X3Y117_DLUT (
.I0(CLBLM_R_X3Y115_SLICE_X3Y115_BQ),
.I1(CLBLM_R_X3Y122_SLICE_X3Y122_AO5),
.I2(RIOB33_X105Y135_IOB_X1Y136_I),
.I3(CLBLM_R_X3Y117_SLICE_X2Y117_AQ),
.I4(CLBLL_L_X2Y121_SLICE_X1Y121_BO5),
.I5(RIOB33_X105Y135_IOB_X1Y135_I),
.O5(CLBLM_R_X3Y117_SLICE_X3Y117_DO5),
.O6(CLBLM_R_X3Y117_SLICE_X3Y117_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hff003333f0f04444)
  ) CLBLM_R_X3Y117_SLICE_X3Y117_CLUT (
.I0(CLBLM_R_X3Y117_SLICE_X3Y117_C5Q),
.I1(RIOB33_X105Y119_IOB_X1Y119_I),
.I2(CLBLM_L_X8Y114_SLICE_X10Y114_C5Q),
.I3(CLBLM_R_X5Y114_SLICE_X6Y114_CQ),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(1'b1),
.O5(CLBLM_R_X3Y117_SLICE_X3Y117_CO5),
.O6(CLBLM_R_X3Y117_SLICE_X3Y117_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f02222ff00f5f5)
  ) CLBLM_R_X3Y117_SLICE_X3Y117_BLUT (
.I0(RIOB33_X105Y119_IOB_X1Y119_I),
.I1(CLBLM_R_X3Y117_SLICE_X3Y117_BQ),
.I2(CLBLM_R_X3Y117_SLICE_X3Y117_CQ),
.I3(CLBLM_R_X3Y112_SLICE_X2Y112_AQ),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(1'b1),
.O5(CLBLM_R_X3Y117_SLICE_X3Y117_BO5),
.O6(CLBLM_R_X3Y117_SLICE_X3Y117_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfff00f00acacacac)
  ) CLBLM_R_X3Y117_SLICE_X3Y117_ALUT (
.I0(CLBLM_R_X5Y116_SLICE_X7Y116_A5Q),
.I1(CLBLM_R_X3Y116_SLICE_X2Y116_AQ),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLM_R_X7Y121_SLICE_X8Y121_AQ),
.I4(CLBLM_R_X3Y117_SLICE_X2Y117_AQ),
.I5(1'b1),
.O5(CLBLM_R_X3Y117_SLICE_X3Y117_AO5),
.O6(CLBLM_R_X3Y117_SLICE_X3Y117_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y118_SLICE_X2Y118_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y118_SLICE_X2Y118_AO6),
.Q(CLBLM_R_X3Y118_SLICE_X2Y118_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hff77ff33ff55ff00)
  ) CLBLM_R_X3Y118_SLICE_X2Y118_DLUT (
.I0(CLBLL_L_X4Y120_SLICE_X5Y120_BO6),
.I1(CLBLL_L_X2Y119_SLICE_X1Y119_AO5),
.I2(1'b1),
.I3(CLBLM_R_X3Y118_SLICE_X2Y118_CO6),
.I4(CLBLM_R_X5Y115_SLICE_X6Y115_AQ),
.I5(CLBLL_L_X2Y112_SLICE_X1Y112_A5Q),
.O5(CLBLM_R_X3Y118_SLICE_X2Y118_DO5),
.O6(CLBLM_R_X3Y118_SLICE_X2Y118_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0050005000ff0050)
  ) CLBLM_R_X3Y118_SLICE_X2Y118_CLUT (
.I0(CLBLL_L_X2Y121_SLICE_X1Y121_BO5),
.I1(1'b1),
.I2(CLBLL_L_X4Y118_SLICE_X4Y118_AQ),
.I3(CLBLM_R_X3Y122_SLICE_X3Y122_AO6),
.I4(CLBLL_L_X4Y119_SLICE_X4Y119_AQ),
.I5(CLBLL_L_X2Y121_SLICE_X1Y121_BO6),
.O5(CLBLM_R_X3Y118_SLICE_X2Y118_CO5),
.O6(CLBLM_R_X3Y118_SLICE_X2Y118_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000005000404)
  ) CLBLM_R_X3Y118_SLICE_X2Y118_BLUT (
.I0(CLBLM_R_X3Y122_SLICE_X3Y122_AO5),
.I1(CLBLM_R_X5Y118_SLICE_X7Y118_AQ),
.I2(RIOB33_X105Y135_IOB_X1Y135_I),
.I3(CLBLL_L_X4Y118_SLICE_X5Y118_CQ),
.I4(RIOB33_X105Y135_IOB_X1Y136_I),
.I5(CLBLL_L_X2Y120_SLICE_X1Y120_AO6),
.O5(CLBLM_R_X3Y118_SLICE_X2Y118_BO5),
.O6(CLBLM_R_X3Y118_SLICE_X2Y118_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hff000000ff040004)
  ) CLBLM_R_X3Y118_SLICE_X2Y118_ALUT (
.I0(RIOB33_X105Y117_IOB_X1Y118_I),
.I1(RIOB33_X105Y119_IOB_X1Y119_I),
.I2(CLBLM_R_X3Y118_SLICE_X2Y118_AQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLL_L_X4Y118_SLICE_X4Y118_AQ),
.I5(CLBLM_R_X3Y117_SLICE_X3Y117_CQ),
.O5(CLBLM_R_X3Y118_SLICE_X2Y118_AO5),
.O6(CLBLM_R_X3Y118_SLICE_X2Y118_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y118_SLICE_X3Y118_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y118_SLICE_X3Y118_AO6),
.Q(CLBLM_R_X3Y118_SLICE_X3Y118_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h00cc00ccaaeeaaee)
  ) CLBLM_R_X3Y118_SLICE_X3Y118_DLUT (
.I0(CLBLL_L_X2Y115_SLICE_X1Y115_AQ),
.I1(CLBLM_L_X10Y114_SLICE_X13Y114_D5Q),
.I2(1'b1),
.I3(CLBLL_L_X4Y121_SLICE_X4Y121_CO6),
.I4(1'b1),
.I5(CLBLM_R_X3Y121_SLICE_X2Y121_AO5),
.O5(CLBLM_R_X3Y118_SLICE_X3Y118_DO5),
.O6(CLBLM_R_X3Y118_SLICE_X3Y118_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0faf0faf00aa00aa)
  ) CLBLM_R_X3Y118_SLICE_X3Y118_CLUT (
.I0(CLBLM_R_X3Y115_SLICE_X3Y115_AQ),
.I1(1'b1),
.I2(CLBLL_L_X2Y120_SLICE_X0Y120_AO5),
.I3(CLBLM_R_X3Y121_SLICE_X2Y121_AO6),
.I4(1'b1),
.I5(CLBLM_R_X3Y118_SLICE_X3Y118_AQ),
.O5(CLBLM_R_X3Y118_SLICE_X3Y118_CO5),
.O6(CLBLM_R_X3Y118_SLICE_X3Y118_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h4400404000000000)
  ) CLBLM_R_X3Y118_SLICE_X3Y118_BLUT (
.I0(CLBLM_R_X3Y121_SLICE_X3Y121_CO6),
.I1(RIOB33_X105Y133_IOB_X1Y133_I),
.I2(CLBLL_L_X4Y117_SLICE_X5Y117_AQ),
.I3(CLBLM_R_X3Y110_SLICE_X3Y110_AQ),
.I4(RIOB33_X105Y131_IOB_X1Y131_I),
.I5(RIOB33_X105Y133_IOB_X1Y134_I),
.O5(CLBLM_R_X3Y118_SLICE_X3Y118_BO5),
.O6(CLBLM_R_X3Y118_SLICE_X3Y118_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfbf8fbf80b080b08)
  ) CLBLM_R_X3Y118_SLICE_X3Y118_ALUT (
.I0(CLBLL_L_X4Y117_SLICE_X5Y117_DQ),
.I1(CLBLM_R_X11Y121_SLICE_X14Y121_CO6),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLM_R_X3Y118_SLICE_X3Y118_AQ),
.I4(1'b1),
.I5(CLBLL_L_X2Y112_SLICE_X1Y112_A5Q),
.O5(CLBLM_R_X3Y118_SLICE_X3Y118_AO5),
.O6(CLBLM_R_X3Y118_SLICE_X3Y118_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h00000000000e0002)
  ) CLBLM_R_X3Y119_SLICE_X2Y119_DLUT (
.I0(CLBLM_R_X3Y115_SLICE_X2Y115_AQ),
.I1(RIOB33_X105Y135_IOB_X1Y136_I),
.I2(RIOB33_X105Y135_IOB_X1Y135_I),
.I3(CLBLM_R_X3Y122_SLICE_X3Y122_AO5),
.I4(RIOB33_X105Y111_IOB_X1Y111_I),
.I5(CLBLL_L_X2Y121_SLICE_X1Y121_BO6),
.O5(CLBLM_R_X3Y119_SLICE_X2Y119_DO5),
.O6(CLBLM_R_X3Y119_SLICE_X2Y119_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hfcfcf0fcfefefafe)
  ) CLBLM_R_X3Y119_SLICE_X2Y119_CLUT (
.I0(LIOB33_X0Y67_IOB_X0Y67_I),
.I1(CLBLM_R_X3Y112_SLICE_X3Y112_CQ),
.I2(CLBLL_L_X4Y122_SLICE_X4Y122_DO6),
.I3(RIOB33_X105Y137_IOB_X1Y137_I),
.I4(RIOB33_X105Y129_IOB_X1Y129_I),
.I5(CLBLL_L_X2Y121_SLICE_X0Y121_AO6),
.O5(CLBLM_R_X3Y119_SLICE_X2Y119_CO5),
.O6(CLBLM_R_X3Y119_SLICE_X2Y119_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h7f5f77553f0f3300)
  ) CLBLM_R_X3Y119_SLICE_X2Y119_BLUT (
.I0(CLBLL_L_X2Y121_SLICE_X1Y121_AO6),
.I1(CLBLL_L_X2Y122_SLICE_X0Y122_AO6),
.I2(CLBLL_L_X2Y120_SLICE_X0Y120_AO6),
.I3(RIOB33_X105Y111_IOB_X1Y112_I),
.I4(CLBLM_R_X3Y119_SLICE_X3Y119_AQ),
.I5(CLBLL_L_X4Y115_SLICE_X5Y115_DQ),
.O5(CLBLM_R_X3Y119_SLICE_X2Y119_BO5),
.O6(CLBLM_R_X3Y119_SLICE_X2Y119_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffffffffffff4)
  ) CLBLM_R_X3Y119_SLICE_X2Y119_ALUT (
.I0(CLBLL_L_X2Y119_SLICE_X1Y119_AO6),
.I1(CLBLL_L_X2Y120_SLICE_X1Y120_CO6),
.I2(CLBLM_R_X5Y118_SLICE_X6Y118_DO6),
.I3(CLBLM_R_X3Y119_SLICE_X2Y119_BO6),
.I4(CLBLM_R_X3Y118_SLICE_X2Y118_BO6),
.I5(CLBLM_R_X3Y119_SLICE_X2Y119_CO6),
.O5(CLBLM_R_X3Y119_SLICE_X2Y119_AO5),
.O6(CLBLM_R_X3Y119_SLICE_X2Y119_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y119_SLICE_X3Y119_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y119_SLICE_X3Y119_AO6),
.Q(CLBLM_R_X3Y119_SLICE_X3Y119_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h000000cc0000f0fc)
  ) CLBLM_R_X3Y119_SLICE_X3Y119_DLUT (
.I0(1'b1),
.I1(CLBLM_R_X3Y112_SLICE_X3Y112_C5Q),
.I2(RIOB33_X105Y109_IOB_X1Y109_I),
.I3(CLBLL_L_X2Y120_SLICE_X1Y120_AO6),
.I4(CLBLM_R_X3Y124_SLICE_X2Y124_AO6),
.I5(CLBLL_L_X2Y121_SLICE_X1Y121_BO6),
.O5(CLBLM_R_X3Y119_SLICE_X3Y119_DO5),
.O6(CLBLM_R_X3Y119_SLICE_X3Y119_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h5dff5d5d0cff0c0c)
  ) CLBLM_R_X3Y119_SLICE_X3Y119_CLUT (
.I0(CLBLL_L_X4Y120_SLICE_X5Y120_BO5),
.I1(CLBLM_L_X8Y119_SLICE_X11Y119_AQ),
.I2(CLBLL_L_X2Y120_SLICE_X0Y120_AO5),
.I3(CLBLM_R_X3Y121_SLICE_X2Y121_AO5),
.I4(CLBLM_R_X3Y113_SLICE_X3Y113_AQ),
.I5(CLBLM_R_X5Y122_SLICE_X7Y122_BQ),
.O5(CLBLM_R_X3Y119_SLICE_X3Y119_CO5),
.O6(CLBLM_R_X3Y119_SLICE_X3Y119_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0005000400010000)
  ) CLBLM_R_X3Y119_SLICE_X3Y119_BLUT (
.I0(CLBLL_L_X2Y122_SLICE_X1Y122_DO6),
.I1(RIOB33_X105Y131_IOB_X1Y131_I),
.I2(CLBLM_R_X3Y122_SLICE_X3Y122_AO6),
.I3(RIOB33_X105Y131_IOB_X1Y132_I),
.I4(CLBLM_R_X5Y122_SLICE_X7Y122_BQ),
.I5(CLBLM_L_X8Y119_SLICE_X11Y119_AQ),
.O5(CLBLM_R_X3Y119_SLICE_X3Y119_BO5),
.O6(CLBLM_R_X3Y119_SLICE_X3Y119_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000fffa000000fa)
  ) CLBLM_R_X3Y119_SLICE_X3Y119_ALUT (
.I0(CLBLL_L_X4Y113_SLICE_X5Y113_CQ),
.I1(1'b1),
.I2(CLBLM_R_X3Y119_SLICE_X3Y119_AQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLM_R_X5Y115_SLICE_X6Y115_CO6),
.I5(CLBLL_L_X4Y123_SLICE_X4Y123_BQ),
.O5(CLBLM_R_X3Y119_SLICE_X3Y119_AO5),
.O6(CLBLM_R_X3Y119_SLICE_X3Y119_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0fffafff0f0fafa)
  ) CLBLM_R_X3Y120_SLICE_X2Y120_DLUT (
.I0(CLBLM_R_X3Y111_SLICE_X2Y111_AQ),
.I1(1'b1),
.I2(CLBLM_R_X3Y119_SLICE_X2Y119_DO6),
.I3(CLBLL_L_X4Y120_SLICE_X5Y120_BO6),
.I4(CLBLM_R_X3Y122_SLICE_X2Y122_BO5),
.I5(CLBLM_R_X3Y116_SLICE_X2Y116_BQ),
.O5(CLBLM_R_X3Y120_SLICE_X2Y120_DO5),
.O6(CLBLM_R_X3Y120_SLICE_X2Y120_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h002f002f00220022)
  ) CLBLM_R_X3Y120_SLICE_X2Y120_CLUT (
.I0(CLBLM_R_X3Y111_SLICE_X2Y111_AQ),
.I1(CLBLL_L_X2Y120_SLICE_X1Y120_AO6),
.I2(CLBLL_L_X2Y121_SLICE_X0Y121_BO6),
.I3(CLBLM_R_X3Y122_SLICE_X3Y122_AO6),
.I4(1'b1),
.I5(CLBLM_R_X3Y116_SLICE_X2Y116_BQ),
.O5(CLBLM_R_X3Y120_SLICE_X2Y120_CO5),
.O6(CLBLM_R_X3Y120_SLICE_X2Y120_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hcfdf0055cfcf0000)
  ) CLBLM_R_X3Y120_SLICE_X2Y120_BLUT (
.I0(CLBLM_R_X3Y124_SLICE_X2Y124_AO5),
.I1(RIOB33_X105Y129_IOB_X1Y129_I),
.I2(RIOB33_X105Y137_IOB_X1Y137_I),
.I3(CLBLL_L_X2Y121_SLICE_X1Y121_BO6),
.I4(CLBLM_R_X3Y112_SLICE_X3Y112_CQ),
.I5(LIOB33_X0Y67_IOB_X0Y67_I),
.O5(CLBLM_R_X3Y120_SLICE_X2Y120_BO5),
.O6(CLBLM_R_X3Y120_SLICE_X2Y120_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffffffffafffe)
  ) CLBLM_R_X3Y120_SLICE_X2Y120_ALUT (
.I0(CLBLL_L_X4Y122_SLICE_X4Y122_DO6),
.I1(CLBLL_L_X4Y115_SLICE_X5Y115_DQ),
.I2(CLBLM_R_X3Y120_SLICE_X3Y120_AO6),
.I3(CLBLM_R_X3Y120_SLICE_X2Y120_BO6),
.I4(CLBLL_L_X2Y121_SLICE_X1Y121_AO6),
.I5(CLBLM_R_X3Y118_SLICE_X2Y118_BO6),
.O5(CLBLM_R_X3Y120_SLICE_X2Y120_AO5),
.O6(CLBLM_R_X3Y120_SLICE_X2Y120_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hdcdcdcdcffffdcdc)
  ) CLBLM_R_X3Y120_SLICE_X3Y120_DLUT (
.I0(CLBLL_L_X2Y121_SLICE_X1Y121_AO6),
.I1(CLBLM_R_X3Y119_SLICE_X3Y119_DO6),
.I2(CLBLM_R_X3Y115_SLICE_X2Y115_DQ),
.I3(1'b1),
.I4(CLBLM_R_X5Y120_SLICE_X7Y120_BQ),
.I5(CLBLL_L_X2Y120_SLICE_X0Y120_AO6),
.O5(CLBLM_R_X3Y120_SLICE_X3Y120_DO5),
.O6(CLBLM_R_X3Y120_SLICE_X3Y120_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0202020203030000)
  ) CLBLM_R_X3Y120_SLICE_X3Y120_CLUT (
.I0(CLBLM_R_X3Y112_SLICE_X2Y112_BQ),
.I1(CLBLL_L_X4Y122_SLICE_X4Y122_AO6),
.I2(CLBLM_R_X3Y124_SLICE_X2Y124_AO6),
.I3(1'b1),
.I4(CLBLL_L_X4Y114_SLICE_X4Y114_CQ),
.I5(RIOB33_X105Y131_IOB_X1Y131_I),
.O5(CLBLM_R_X3Y120_SLICE_X3Y120_CO5),
.O6(CLBLM_R_X3Y120_SLICE_X3Y120_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffffffffffffe)
  ) CLBLM_R_X3Y120_SLICE_X3Y120_BLUT (
.I0(CLBLM_R_X3Y118_SLICE_X3Y118_DO6),
.I1(CLBLL_L_X4Y120_SLICE_X5Y120_CO6),
.I2(CLBLL_L_X2Y121_SLICE_X1Y121_CO6),
.I3(CLBLM_R_X3Y120_SLICE_X3Y120_DO6),
.I4(CLBLM_R_X3Y122_SLICE_X2Y122_DO6),
.I5(CLBLM_R_X3Y118_SLICE_X3Y118_CO6),
.O5(CLBLM_R_X3Y120_SLICE_X3Y120_BO5),
.O6(CLBLM_R_X3Y120_SLICE_X3Y120_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000011011000)
  ) CLBLM_R_X3Y120_SLICE_X3Y120_ALUT (
.I0(CLBLM_R_X3Y122_SLICE_X3Y122_AO5),
.I1(CLBLL_L_X2Y121_SLICE_X1Y121_BO6),
.I2(RIOB33_X105Y135_IOB_X1Y136_I),
.I3(RIOB33_X105Y111_IOB_X1Y112_I),
.I4(CLBLM_R_X3Y119_SLICE_X3Y119_AQ),
.I5(RIOB33_X105Y135_IOB_X1Y135_I),
.O5(CLBLM_R_X3Y120_SLICE_X3Y120_AO5),
.O6(CLBLM_R_X3Y120_SLICE_X3Y120_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0008000000000000)
  ) CLBLM_R_X3Y121_SLICE_X2Y121_DLUT (
.I0(CLBLM_R_X3Y122_SLICE_X2Y122_AO6),
.I1(CLBLL_L_X4Y121_SLICE_X4Y121_CO5),
.I2(CLBLM_R_X3Y122_SLICE_X2Y122_BO6),
.I3(CLBLL_L_X4Y121_SLICE_X5Y121_BO6),
.I4(CLBLL_L_X2Y120_SLICE_X0Y120_AO6),
.I5(CLBLM_R_X3Y123_SLICE_X3Y123_BO6),
.O5(CLBLM_R_X3Y121_SLICE_X2Y121_DO5),
.O6(CLBLM_R_X3Y121_SLICE_X2Y121_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hfefefffeffffffff)
  ) CLBLM_R_X3Y121_SLICE_X2Y121_CLUT (
.I0(CLBLM_R_X5Y118_SLICE_X6Y118_DO6),
.I1(CLBLM_R_X3Y121_SLICE_X3Y121_AO6),
.I2(CLBLM_R_X3Y120_SLICE_X2Y120_AO6),
.I3(CLBLL_L_X2Y121_SLICE_X1Y121_DO6),
.I4(CLBLL_L_X4Y122_SLICE_X5Y122_DO6),
.I5(CLBLM_R_X3Y121_SLICE_X2Y121_BO6),
.O5(CLBLM_R_X3Y121_SLICE_X2Y121_CO5),
.O6(CLBLM_R_X3Y121_SLICE_X2Y121_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffefffffffffff)
  ) CLBLM_R_X3Y121_SLICE_X2Y121_BLUT (
.I0(CLBLM_R_X3Y122_SLICE_X2Y122_CO6),
.I1(CLBLL_L_X4Y121_SLICE_X4Y121_DO6),
.I2(CLBLM_R_X3Y122_SLICE_X2Y122_AO6),
.I3(CLBLL_L_X2Y121_SLICE_X1Y121_AO6),
.I4(CLBLL_L_X2Y119_SLICE_X1Y119_AO6),
.I5(CLBLM_R_X3Y121_SLICE_X2Y121_AO5),
.O5(CLBLM_R_X3Y121_SLICE_X2Y121_BO5),
.O6(CLBLM_R_X3Y121_SLICE_X2Y121_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hbfffffffffffbfff)
  ) CLBLM_R_X3Y121_SLICE_X2Y121_ALUT (
.I0(CLBLM_R_X3Y124_SLICE_X2Y124_AO6),
.I1(RIOB33_X105Y131_IOB_X1Y132_I),
.I2(RIOB33_X105Y133_IOB_X1Y134_I),
.I3(RIOB33_X105Y133_IOB_X1Y133_I),
.I4(RIOB33_X105Y131_IOB_X1Y131_I),
.I5(1'b1),
.O5(CLBLM_R_X3Y121_SLICE_X2Y121_AO5),
.O6(CLBLM_R_X3Y121_SLICE_X2Y121_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hffaeffaeffffffae)
  ) CLBLM_R_X3Y121_SLICE_X3Y121_DLUT (
.I0(CLBLM_L_X8Y122_SLICE_X10Y122_BO6),
.I1(CLBLM_R_X5Y120_SLICE_X7Y120_CQ),
.I2(CLBLM_R_X3Y123_SLICE_X3Y123_BO5),
.I3(CLBLM_R_X3Y117_SLICE_X3Y117_DO6),
.I4(LIOB33_X0Y65_IOB_X0Y66_I),
.I5(CLBLL_L_X2Y121_SLICE_X0Y121_AO6),
.O5(CLBLM_R_X3Y121_SLICE_X3Y121_DO5),
.O6(CLBLM_R_X3Y121_SLICE_X3Y121_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffffffffdfff)
  ) CLBLM_R_X3Y121_SLICE_X3Y121_CLUT (
.I0(RIOB33_X105Y131_IOB_X1Y132_I),
.I1(RIOB33_X105Y129_IOB_X1Y129_I),
.I2(RIOB33_X105Y135_IOB_X1Y136_I),
.I3(RIOB33_X105Y137_IOB_X1Y137_I),
.I4(RIOB33_X105Y129_IOB_X1Y130_I),
.I5(RIOB33_X105Y135_IOB_X1Y135_I),
.O5(CLBLM_R_X3Y121_SLICE_X3Y121_CO5),
.O6(CLBLM_R_X3Y121_SLICE_X3Y121_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff0404ffff5504)
  ) CLBLM_R_X3Y121_SLICE_X3Y121_BLUT (
.I0(CLBLM_R_X3Y124_SLICE_X2Y124_AO5),
.I1(CLBLM_R_X5Y120_SLICE_X7Y120_CQ),
.I2(CLBLL_L_X2Y121_SLICE_X1Y121_BO5),
.I3(LIOB33_X0Y65_IOB_X0Y66_I),
.I4(CLBLM_L_X8Y122_SLICE_X10Y122_BO6),
.I5(CLBLL_L_X2Y121_SLICE_X1Y121_BO6),
.O5(CLBLM_R_X3Y121_SLICE_X3Y121_BO5),
.O6(CLBLM_R_X3Y121_SLICE_X3Y121_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffffffffffffe)
  ) CLBLM_R_X3Y121_SLICE_X3Y121_ALUT (
.I0(CLBLM_R_X3Y117_SLICE_X3Y117_DO6),
.I1(CLBLM_R_X3Y122_SLICE_X3Y122_BO6),
.I2(CLBLM_R_X3Y119_SLICE_X3Y119_BO6),
.I3(CLBLM_R_X3Y121_SLICE_X3Y121_BO6),
.I4(CLBLM_R_X3Y120_SLICE_X2Y120_CO6),
.I5(CLBLM_R_X3Y119_SLICE_X2Y119_DO6),
.O5(CLBLM_R_X3Y121_SLICE_X3Y121_AO5),
.O6(CLBLM_R_X3Y121_SLICE_X3Y121_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffefffffffefe)
  ) CLBLM_R_X3Y122_SLICE_X2Y122_DLUT (
.I0(CLBLL_L_X2Y121_SLICE_X0Y121_DO6),
.I1(CLBLL_L_X2Y122_SLICE_X1Y122_CO6),
.I2(CLBLM_R_X3Y122_SLICE_X3Y122_DO6),
.I3(CLBLM_R_X3Y122_SLICE_X2Y122_AO5),
.I4(CLBLM_R_X5Y122_SLICE_X6Y122_DO6),
.I5(LIOB33_X0Y57_IOB_X0Y58_I),
.O5(CLBLM_R_X3Y122_SLICE_X2Y122_DO5),
.O6(CLBLM_R_X3Y122_SLICE_X2Y122_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hf1f1f3fff1f1f3f3)
  ) CLBLM_R_X3Y122_SLICE_X2Y122_CLUT (
.I0(CLBLL_L_X2Y121_SLICE_X0Y121_BO6),
.I1(CLBLM_R_X3Y122_SLICE_X3Y122_AO6),
.I2(CLBLL_L_X4Y121_SLICE_X5Y121_BO6),
.I3(CLBLM_R_X3Y124_SLICE_X2Y124_AO5),
.I4(CLBLL_L_X4Y122_SLICE_X4Y122_AO6),
.I5(RIOB33_X105Y131_IOB_X1Y131_I),
.O5(CLBLM_R_X3Y122_SLICE_X2Y122_CO5),
.O6(CLBLM_R_X3Y122_SLICE_X2Y122_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h00030400fffdffff)
  ) CLBLM_R_X3Y122_SLICE_X2Y122_BLUT (
.I0(RIOB33_X105Y131_IOB_X1Y131_I),
.I1(RIOB33_X105Y133_IOB_X1Y133_I),
.I2(CLBLM_R_X3Y122_SLICE_X3Y122_AO6),
.I3(RIOB33_X105Y131_IOB_X1Y132_I),
.I4(RIOB33_X105Y133_IOB_X1Y134_I),
.I5(1'b1),
.O5(CLBLM_R_X3Y122_SLICE_X2Y122_BO5),
.O6(CLBLM_R_X3Y122_SLICE_X2Y122_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hebefbffbfbffffff)
  ) CLBLM_R_X3Y122_SLICE_X2Y122_ALUT (
.I0(CLBLM_R_X3Y124_SLICE_X2Y124_AO5),
.I1(RIOB33_X105Y133_IOB_X1Y134_I),
.I2(RIOB33_X105Y133_IOB_X1Y133_I),
.I3(RIOB33_X105Y131_IOB_X1Y131_I),
.I4(RIOB33_X105Y131_IOB_X1Y132_I),
.I5(1'b1),
.O5(CLBLM_R_X3Y122_SLICE_X2Y122_AO5),
.O6(CLBLM_R_X3Y122_SLICE_X2Y122_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaa2222afaa2f22)
  ) CLBLM_R_X3Y122_SLICE_X3Y122_DLUT (
.I0(CLBLM_R_X5Y122_SLICE_X7Y122_AQ),
.I1(RIOB33_X105Y137_IOB_X1Y137_I),
.I2(CLBLL_L_X2Y121_SLICE_X0Y121_BO6),
.I3(RIOB33_X105Y117_IOB_X1Y117_I),
.I4(RIOB33_X105Y129_IOB_X1Y129_I),
.I5(CLBLM_R_X3Y124_SLICE_X2Y124_AO6),
.O5(CLBLM_R_X3Y122_SLICE_X3Y122_DO5),
.O6(CLBLM_R_X3Y122_SLICE_X3Y122_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff575503000300)
  ) CLBLM_R_X3Y122_SLICE_X3Y122_CLUT (
.I0(RIOB33_X105Y137_IOB_X1Y137_I),
.I1(CLBLL_L_X2Y121_SLICE_X1Y121_BO6),
.I2(CLBLM_R_X3Y124_SLICE_X2Y124_AO5),
.I3(LIOB33_X0Y61_IOB_X0Y62_I),
.I4(RIOB33_X105Y129_IOB_X1Y129_I),
.I5(CLBLM_R_X5Y120_SLICE_X6Y120_AQ),
.O5(CLBLM_R_X3Y122_SLICE_X3Y122_CO5),
.O6(CLBLM_R_X3Y122_SLICE_X3Y122_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0020000000000000)
  ) CLBLM_R_X3Y122_SLICE_X3Y122_BLUT (
.I0(CLBLM_R_X3Y113_SLICE_X3Y113_AQ),
.I1(RIOB33_X105Y131_IOB_X1Y131_I),
.I2(RIOB33_X105Y133_IOB_X1Y134_I),
.I3(CLBLM_R_X3Y124_SLICE_X2Y124_AO6),
.I4(RIOB33_X105Y133_IOB_X1Y133_I),
.I5(RIOB33_X105Y131_IOB_X1Y132_I),
.O5(CLBLM_R_X3Y122_SLICE_X3Y122_BO5),
.O6(CLBLM_R_X3Y122_SLICE_X3Y122_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffefffafffaff)
  ) CLBLM_R_X3Y122_SLICE_X3Y122_ALUT (
.I0(RIOB33_X105Y129_IOB_X1Y129_I),
.I1(RIOB33_X105Y135_IOB_X1Y135_I),
.I2(RIOB33_X105Y129_IOB_X1Y130_I),
.I3(RIOB33_X105Y137_IOB_X1Y137_I),
.I4(RIOB33_X105Y135_IOB_X1Y136_I),
.I5(1'b1),
.O5(CLBLM_R_X3Y122_SLICE_X3Y122_AO5),
.O6(CLBLM_R_X3Y122_SLICE_X3Y122_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000300000000202)
  ) CLBLM_R_X3Y123_SLICE_X2Y123_DLUT (
.I0(CLBLM_R_X3Y123_SLICE_X3Y123_AQ),
.I1(CLBLM_R_X3Y124_SLICE_X2Y124_AO5),
.I2(RIOB33_X105Y131_IOB_X1Y131_I),
.I3(LIOB33_X0Y57_IOB_X0Y57_I),
.I4(CLBLM_R_X3Y124_SLICE_X2Y124_BO5),
.I5(RIOB33_X105Y131_IOB_X1Y132_I),
.O5(CLBLM_R_X3Y123_SLICE_X2Y123_DO5),
.O6(CLBLM_R_X3Y123_SLICE_X2Y123_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0009000100080000)
  ) CLBLM_R_X3Y123_SLICE_X2Y123_CLUT (
.I0(RIOB33_X105Y131_IOB_X1Y132_I),
.I1(RIOB33_X105Y131_IOB_X1Y131_I),
.I2(CLBLM_R_X3Y124_SLICE_X2Y124_BO5),
.I3(CLBLM_R_X3Y124_SLICE_X2Y124_AO5),
.I4(LIOB33_X0Y55_IOB_X0Y55_I),
.I5(CLBLL_L_X4Y119_SLICE_X4Y119_DQ),
.O5(CLBLM_R_X3Y123_SLICE_X2Y123_CO5),
.O6(CLBLM_R_X3Y123_SLICE_X2Y123_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffffffffffff2)
  ) CLBLM_R_X3Y123_SLICE_X2Y123_BLUT (
.I0(CLBLL_L_X2Y117_SLICE_X0Y117_AQ),
.I1(CLBLM_R_X3Y123_SLICE_X3Y123_BO6),
.I2(CLBLL_L_X2Y122_SLICE_X1Y122_AO6),
.I3(CLBLM_R_X3Y123_SLICE_X3Y123_CO6),
.I4(CLBLM_R_X3Y123_SLICE_X2Y123_AO6),
.I5(CLBLM_R_X3Y123_SLICE_X2Y123_CO6),
.O5(CLBLM_R_X3Y123_SLICE_X2Y123_BO5),
.O6(CLBLM_R_X3Y123_SLICE_X2Y123_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hf000f0f0f222f2f2)
  ) CLBLM_R_X3Y123_SLICE_X2Y123_ALUT (
.I0(RIOB33_X105Y115_IOB_X1Y115_I),
.I1(CLBLL_L_X2Y121_SLICE_X0Y121_BO6),
.I2(CLBLM_R_X7Y119_SLICE_X8Y119_C5Q),
.I3(RIOB33_X105Y129_IOB_X1Y129_I),
.I4(RIOB33_X105Y137_IOB_X1Y137_I),
.I5(CLBLM_R_X3Y124_SLICE_X2Y124_AO6),
.O5(CLBLM_R_X3Y123_SLICE_X2Y123_AO5),
.O6(CLBLM_R_X3Y123_SLICE_X2Y123_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y123_SLICE_X3Y123_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y123_SLICE_X3Y123_AO6),
.Q(CLBLM_R_X3Y123_SLICE_X3Y123_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffefffefffffffe)
  ) CLBLM_R_X3Y123_SLICE_X3Y123_DLUT (
.I0(CLBLM_R_X3Y124_SLICE_X3Y124_AO6),
.I1(CLBLL_L_X4Y123_SLICE_X4Y123_DO6),
.I2(CLBLM_R_X3Y123_SLICE_X2Y123_DO6),
.I3(CLBLM_R_X3Y122_SLICE_X3Y122_CO6),
.I4(CLBLL_L_X2Y117_SLICE_X1Y117_BQ),
.I5(CLBLM_R_X3Y123_SLICE_X3Y123_BO6),
.O5(CLBLM_R_X3Y123_SLICE_X3Y123_DO5),
.O6(CLBLM_R_X3Y123_SLICE_X3Y123_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000020000000)
  ) CLBLM_R_X3Y123_SLICE_X3Y123_CLUT (
.I0(RIOB33_X105Y133_IOB_X1Y134_I),
.I1(CLBLM_R_X3Y124_SLICE_X2Y124_AO5),
.I2(CLBLM_R_X7Y120_SLICE_X8Y120_CQ),
.I3(RIOB33_X105Y133_IOB_X1Y133_I),
.I4(RIOB33_X105Y131_IOB_X1Y131_I),
.I5(RIOB33_X105Y131_IOB_X1Y132_I),
.O5(CLBLM_R_X3Y123_SLICE_X3Y123_CO5),
.O6(CLBLM_R_X3Y123_SLICE_X3Y123_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffdfffffffeff)
  ) CLBLM_R_X3Y123_SLICE_X3Y123_BLUT (
.I0(RIOB33_X105Y131_IOB_X1Y131_I),
.I1(RIOB33_X105Y133_IOB_X1Y133_I),
.I2(CLBLM_R_X3Y124_SLICE_X2Y124_AO5),
.I3(RIOB33_X105Y133_IOB_X1Y134_I),
.I4(RIOB33_X105Y131_IOB_X1Y132_I),
.I5(1'b1),
.O5(CLBLM_R_X3Y123_SLICE_X3Y123_BO5),
.O6(CLBLM_R_X3Y123_SLICE_X3Y123_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfff000f0ffcc00cc)
  ) CLBLM_R_X3Y123_SLICE_X3Y123_ALUT (
.I0(1'b1),
.I1(CLBLM_R_X3Y117_SLICE_X3Y117_AQ),
.I2(CLBLM_R_X3Y123_SLICE_X3Y123_AQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLM_R_X7Y124_SLICE_X8Y124_BQ),
.I5(CLBLM_R_X3Y116_SLICE_X2Y116_DO6),
.O5(CLBLM_R_X3Y123_SLICE_X3Y123_AO5),
.O6(CLBLM_R_X3Y123_SLICE_X3Y123_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y124_SLICE_X2Y124_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y124_SLICE_X2Y124_DO5),
.O6(CLBLM_R_X3Y124_SLICE_X2Y124_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y124_SLICE_X2Y124_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y124_SLICE_X2Y124_CO5),
.O6(CLBLM_R_X3Y124_SLICE_X2Y124_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hffccffffccffccff)
  ) CLBLM_R_X3Y124_SLICE_X2Y124_BLUT (
.I0(1'b1),
.I1(RIOB33_X105Y133_IOB_X1Y133_I),
.I2(1'b1),
.I3(RIOB33_X105Y133_IOB_X1Y134_I),
.I4(RIOB33_X105Y131_IOB_X1Y132_I),
.I5(1'b1),
.O5(CLBLM_R_X3Y124_SLICE_X2Y124_BO5),
.O6(CLBLM_R_X3Y124_SLICE_X2Y124_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffbffffffbff)
  ) CLBLM_R_X3Y124_SLICE_X2Y124_ALUT (
.I0(RIOB33_X105Y129_IOB_X1Y129_I),
.I1(RIOB33_X105Y137_IOB_X1Y137_I),
.I2(RIOB33_X105Y135_IOB_X1Y136_I),
.I3(RIOB33_X105Y135_IOB_X1Y135_I),
.I4(RIOB33_X105Y129_IOB_X1Y130_I),
.I5(1'b1),
.O5(CLBLM_R_X3Y124_SLICE_X2Y124_AO5),
.O6(CLBLM_R_X3Y124_SLICE_X2Y124_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y124_SLICE_X3Y124_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y124_SLICE_X3Y124_DO5),
.O6(CLBLM_R_X3Y124_SLICE_X3Y124_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y124_SLICE_X3Y124_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y124_SLICE_X3Y124_CO5),
.O6(CLBLM_R_X3Y124_SLICE_X3Y124_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y124_SLICE_X3Y124_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y124_SLICE_X3Y124_BO5),
.O6(CLBLM_R_X3Y124_SLICE_X3Y124_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000080000)
  ) CLBLM_R_X3Y124_SLICE_X3Y124_ALUT (
.I0(RIOB33_X105Y115_IOB_X1Y116_I),
.I1(RIOB33_X105Y133_IOB_X1Y133_I),
.I2(CLBLM_R_X3Y124_SLICE_X2Y124_AO6),
.I3(RIOB33_X105Y133_IOB_X1Y134_I),
.I4(RIOB33_X105Y131_IOB_X1Y132_I),
.I5(RIOB33_X105Y131_IOB_X1Y131_I),
.O5(CLBLM_R_X3Y124_SLICE_X3Y124_AO5),
.O6(CLBLM_R_X3Y124_SLICE_X3Y124_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y109_SLICE_X6Y109_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y109_SLICE_X6Y109_AO6),
.Q(CLBLM_R_X5Y109_SLICE_X6Y109_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y109_SLICE_X6Y109_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y109_SLICE_X6Y109_BO6),
.Q(CLBLM_R_X5Y109_SLICE_X6Y109_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y109_SLICE_X6Y109_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y109_SLICE_X6Y109_CO6),
.Q(CLBLM_R_X5Y109_SLICE_X6Y109_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X5Y109_SLICE_X6Y109_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y109_SLICE_X6Y109_DO5),
.O6(CLBLM_R_X5Y109_SLICE_X6Y109_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hffefbaaa55451000)
  ) CLBLM_R_X5Y109_SLICE_X6Y109_CLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_R_X3Y118_SLICE_X2Y118_AQ),
.I2(RIOB33_X105Y117_IOB_X1Y118_I),
.I3(CLBLM_R_X5Y110_SLICE_X6Y110_CO6),
.I4(CLBLM_R_X5Y109_SLICE_X6Y109_CQ),
.I5(CLBLM_L_X10Y110_SLICE_X12Y110_BQ),
.O5(CLBLM_R_X5Y109_SLICE_X6Y109_CO5),
.O6(CLBLM_R_X5Y109_SLICE_X6Y109_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'haca0aca0acacacac)
  ) CLBLM_R_X5Y109_SLICE_X6Y109_BLUT (
.I0(CLBLM_R_X3Y117_SLICE_X3Y117_B5Q),
.I1(CLBLM_R_X5Y109_SLICE_X6Y109_BQ),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLM_R_X3Y118_SLICE_X2Y118_AQ),
.I4(1'b1),
.I5(RIOB33_X105Y117_IOB_X1Y118_I),
.O5(CLBLM_R_X5Y109_SLICE_X6Y109_BO5),
.O6(CLBLM_R_X5Y109_SLICE_X6Y109_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hb888b888b8b8b8b8)
  ) CLBLM_R_X5Y109_SLICE_X6Y109_ALUT (
.I0(CLBLM_R_X5Y109_SLICE_X6Y109_CQ),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(CLBLM_R_X5Y109_SLICE_X6Y109_AQ),
.I3(CLBLM_R_X3Y118_SLICE_X2Y118_AQ),
.I4(1'b1),
.I5(RIOB33_X105Y117_IOB_X1Y118_I),
.O5(CLBLM_R_X5Y109_SLICE_X6Y109_AO5),
.O6(CLBLM_R_X5Y109_SLICE_X6Y109_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y109_SLICE_X7Y109_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y109_SLICE_X7Y109_AO6),
.Q(CLBLM_R_X5Y109_SLICE_X7Y109_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X5Y109_SLICE_X7Y109_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y109_SLICE_X7Y109_DO5),
.O6(CLBLM_R_X5Y109_SLICE_X7Y109_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X5Y109_SLICE_X7Y109_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y109_SLICE_X7Y109_CO5),
.O6(CLBLM_R_X5Y109_SLICE_X7Y109_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X5Y109_SLICE_X7Y109_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y109_SLICE_X7Y109_BO5),
.O6(CLBLM_R_X5Y109_SLICE_X7Y109_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff000054005400)
  ) CLBLM_R_X5Y109_SLICE_X7Y109_ALUT (
.I0(RIOB33_X105Y117_IOB_X1Y118_I),
.I1(CLBLM_R_X5Y112_SLICE_X7Y112_AO6),
.I2(CLBLM_R_X5Y109_SLICE_X7Y109_AQ),
.I3(CLBLM_R_X3Y118_SLICE_X2Y118_AQ),
.I4(CLBLM_R_X5Y109_SLICE_X6Y109_AQ),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLM_R_X5Y109_SLICE_X7Y109_AO5),
.O6(CLBLM_R_X5Y109_SLICE_X7Y109_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y110_SLICE_X6Y110_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y110_SLICE_X6Y110_AO6),
.Q(CLBLM_R_X5Y110_SLICE_X6Y110_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h1310131010131013)
  ) CLBLM_R_X5Y110_SLICE_X6Y110_DLUT (
.I0(CLBLM_R_X5Y111_SLICE_X6Y111_C5Q),
.I1(CLBLM_R_X5Y110_SLICE_X6Y110_AQ),
.I2(CLBLM_R_X5Y111_SLICE_X7Y111_DO6),
.I3(CLBLM_R_X7Y111_SLICE_X9Y111_BO5),
.I4(1'b1),
.I5(CLBLM_R_X5Y114_SLICE_X6Y114_DQ),
.O5(CLBLM_R_X5Y110_SLICE_X6Y110_DO5),
.O6(CLBLM_R_X5Y110_SLICE_X6Y110_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffffffffff3ff)
  ) CLBLM_R_X5Y110_SLICE_X6Y110_CLUT (
.I0(1'b1),
.I1(CLBLM_R_X5Y111_SLICE_X7Y111_CO5),
.I2(CLBLL_L_X2Y120_SLICE_X0Y120_CO6),
.I3(CLBLM_R_X3Y120_SLICE_X3Y120_BO6),
.I4(CLBLM_R_X5Y117_SLICE_X7Y117_DO6),
.I5(CLBLL_L_X4Y120_SLICE_X5Y120_AO6),
.O5(CLBLM_R_X5Y110_SLICE_X6Y110_CO5),
.O6(CLBLM_R_X5Y110_SLICE_X6Y110_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hff0f0000ffee0000)
  ) CLBLM_R_X5Y110_SLICE_X6Y110_BLUT (
.I0(CLBLL_L_X2Y120_SLICE_X1Y120_DO6),
.I1(CLBLM_R_X5Y117_SLICE_X7Y117_DO6),
.I2(CLBLM_R_X5Y109_SLICE_X6Y109_CQ),
.I3(CLBLM_R_X7Y112_SLICE_X8Y112_BQ),
.I4(RIOB33_X105Y121_IOB_X1Y121_I),
.I5(CLBLL_L_X4Y110_SLICE_X5Y110_DO6),
.O5(CLBLM_R_X5Y110_SLICE_X6Y110_BO5),
.O6(CLBLM_R_X5Y110_SLICE_X6Y110_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff550500005505)
  ) CLBLM_R_X5Y110_SLICE_X6Y110_ALUT (
.I0(CLBLM_R_X5Y110_SLICE_X6Y110_DO6),
.I1(1'b1),
.I2(RIOB33_X105Y141_IOB_X1Y142_I),
.I3(CLBLM_R_X7Y128_SLICE_X8Y128_AQ),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(CLBLM_R_X5Y111_SLICE_X6Y111_CQ),
.O5(CLBLM_R_X5Y110_SLICE_X6Y110_AO5),
.O6(CLBLM_R_X5Y110_SLICE_X6Y110_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y110_SLICE_X7Y110_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y110_SLICE_X7Y110_AO6),
.Q(CLBLM_R_X5Y110_SLICE_X7Y110_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y110_SLICE_X7Y110_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y110_SLICE_X7Y110_BO6),
.Q(CLBLM_R_X5Y110_SLICE_X7Y110_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y110_SLICE_X7Y110_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y110_SLICE_X7Y110_CO6),
.Q(CLBLM_R_X5Y110_SLICE_X7Y110_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000ff4f55505550)
  ) CLBLM_R_X5Y110_SLICE_X7Y110_DLUT (
.I0(CLBLM_R_X3Y120_SLICE_X3Y120_BO6),
.I1(RIOB33_X105Y105_IOB_X1Y105_I),
.I2(CLBLM_R_X7Y109_SLICE_X8Y109_AQ),
.I3(CLBLM_R_X5Y116_SLICE_X7Y116_CQ),
.I4(CLBLM_R_X5Y110_SLICE_X7Y110_AQ),
.I5(1'b1),
.O5(CLBLM_R_X5Y110_SLICE_X7Y110_DO5),
.O6(CLBLM_R_X5Y110_SLICE_X7Y110_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'haaeeaaee00440044)
  ) CLBLM_R_X5Y110_SLICE_X7Y110_CLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_R_X7Y112_SLICE_X8Y112_BQ),
.I2(1'b1),
.I3(RIOB33_X105Y105_IOB_X1Y105_I),
.I4(1'b1),
.I5(CLBLL_L_X2Y114_SLICE_X1Y114_AQ),
.O5(CLBLM_R_X5Y110_SLICE_X7Y110_CO5),
.O6(CLBLM_R_X5Y110_SLICE_X7Y110_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hafafacacafa0aca0)
  ) CLBLM_R_X5Y110_SLICE_X7Y110_BLUT (
.I0(CLBLM_R_X7Y110_SLICE_X8Y110_BQ),
.I1(CLBLM_R_X5Y110_SLICE_X7Y110_BQ),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLM_R_X3Y118_SLICE_X2Y118_AQ),
.I4(CLBLM_R_X3Y117_SLICE_X3Y117_B5Q),
.I5(RIOB33_X105Y117_IOB_X1Y118_I),
.O5(CLBLM_R_X5Y110_SLICE_X7Y110_BO5),
.O6(CLBLM_R_X5Y110_SLICE_X7Y110_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hff0004040000fcfc)
  ) CLBLM_R_X5Y110_SLICE_X7Y110_ALUT (
.I0(CLBLM_R_X5Y110_SLICE_X7Y110_DO6),
.I1(CLBLM_R_X3Y118_SLICE_X2Y118_AQ),
.I2(RIOB33_X105Y117_IOB_X1Y118_I),
.I3(CLBLM_L_X8Y112_SLICE_X11Y112_AQ),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(1'b1),
.O5(CLBLM_R_X5Y110_SLICE_X7Y110_AO5),
.O6(CLBLM_R_X5Y110_SLICE_X7Y110_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y111_SLICE_X6Y111_C5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y111_SLICE_X6Y111_CO5),
.Q(CLBLM_R_X5Y111_SLICE_X6Y111_C5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y111_SLICE_X6Y111_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y111_SLICE_X6Y111_AO6),
.Q(CLBLM_R_X5Y111_SLICE_X6Y111_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y111_SLICE_X6Y111_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y111_SLICE_X6Y111_BO6),
.Q(CLBLM_R_X5Y111_SLICE_X6Y111_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y111_SLICE_X6Y111_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y111_SLICE_X6Y111_CO6),
.Q(CLBLM_R_X5Y111_SLICE_X6Y111_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h2211112244888844)
  ) CLBLM_R_X5Y111_SLICE_X6Y111_DLUT (
.I0(CLBLL_L_X4Y115_SLICE_X4Y115_BQ),
.I1(CLBLM_R_X5Y111_SLICE_X6Y111_CQ),
.I2(1'b1),
.I3(CLBLM_R_X5Y115_SLICE_X6Y115_BQ),
.I4(CLBLM_R_X7Y113_SLICE_X8Y113_AQ),
.I5(RIOB33_X105Y105_IOB_X1Y105_I),
.O5(CLBLM_R_X5Y111_SLICE_X6Y111_DO5),
.O6(CLBLM_R_X5Y111_SLICE_X6Y111_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hf3f3c0c0bb88bb88)
  ) CLBLM_R_X5Y111_SLICE_X6Y111_CLUT (
.I0(CLBLM_R_X5Y110_SLICE_X6Y110_AQ),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(CLBLM_R_X5Y111_SLICE_X6Y111_BQ),
.I3(CLBLL_L_X4Y110_SLICE_X4Y110_A5Q),
.I4(CLBLM_R_X5Y111_SLICE_X6Y111_DO6),
.I5(1'b1),
.O5(CLBLM_R_X5Y111_SLICE_X6Y111_CO5),
.O6(CLBLM_R_X5Y111_SLICE_X6Y111_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hff00ff0009090909)
  ) CLBLM_R_X5Y111_SLICE_X6Y111_BLUT (
.I0(CLBLM_R_X5Y112_SLICE_X6Y112_CO6),
.I1(CLBLM_R_X7Y117_SLICE_X8Y117_CQ),
.I2(RIOB33_X105Y105_IOB_X1Y105_I),
.I3(CLBLM_R_X7Y110_SLICE_X9Y110_AQ),
.I4(1'b1),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLM_R_X5Y111_SLICE_X6Y111_BO5),
.O6(CLBLM_R_X5Y111_SLICE_X6Y111_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff000075307530)
  ) CLBLM_R_X5Y111_SLICE_X6Y111_ALUT (
.I0(CLBLM_R_X5Y115_SLICE_X6Y115_DO6),
.I1(RIOB33_X105Y105_IOB_X1Y105_I),
.I2(CLBLM_R_X5Y111_SLICE_X6Y111_AQ),
.I3(CLBLL_L_X4Y111_SLICE_X5Y111_CO6),
.I4(CLBLM_L_X10Y110_SLICE_X13Y110_AQ),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLM_R_X5Y111_SLICE_X6Y111_AO5),
.O6(CLBLM_R_X5Y111_SLICE_X6Y111_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y111_SLICE_X7Y111_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y111_SLICE_X7Y111_AO6),
.Q(CLBLM_R_X5Y111_SLICE_X7Y111_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y111_SLICE_X7Y111_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y111_SLICE_X7Y111_BO6),
.Q(CLBLM_R_X5Y111_SLICE_X7Y111_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hccccccccccccddcc)
  ) CLBLM_R_X5Y111_SLICE_X7Y111_DLUT (
.I0(CLBLL_L_X4Y120_SLICE_X5Y120_AO6),
.I1(CLBLM_R_X5Y119_SLICE_X7Y119_CO6),
.I2(1'b1),
.I3(CLBLM_R_X5Y111_SLICE_X7Y111_CO6),
.I4(CLBLL_L_X2Y120_SLICE_X1Y120_DO6),
.I5(CLBLM_R_X3Y119_SLICE_X2Y119_AO6),
.O5(CLBLM_R_X5Y111_SLICE_X7Y111_DO5),
.O6(CLBLM_R_X5Y111_SLICE_X7Y111_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h000003000a0a0a0a)
  ) CLBLM_R_X5Y111_SLICE_X7Y111_CLUT (
.I0(RIOB33_X105Y105_IOB_X1Y105_I),
.I1(CLBLL_L_X2Y120_SLICE_X0Y120_CO6),
.I2(CLBLL_L_X4Y120_SLICE_X5Y120_DO6),
.I3(CLBLL_L_X2Y119_SLICE_X0Y119_BO6),
.I4(CLBLM_R_X3Y120_SLICE_X3Y120_BO6),
.I5(1'b1),
.O5(CLBLM_R_X5Y111_SLICE_X7Y111_CO5),
.O6(CLBLM_R_X5Y111_SLICE_X7Y111_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hffdededeff000000)
  ) CLBLM_R_X5Y111_SLICE_X7Y111_BLUT (
.I0(CLBLM_R_X5Y113_SLICE_X7Y113_CO6),
.I1(CLBLM_R_X5Y111_SLICE_X7Y111_BQ),
.I2(CLBLM_R_X5Y110_SLICE_X6Y110_BO6),
.I3(CLBLL_L_X4Y110_SLICE_X4Y110_CQ),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(CLBLM_R_X5Y110_SLICE_X7Y110_AO5),
.O5(CLBLM_R_X5Y111_SLICE_X7Y111_BO5),
.O6(CLBLM_R_X5Y111_SLICE_X7Y111_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hff00eeeeff00e0e0)
  ) CLBLM_R_X5Y111_SLICE_X7Y111_ALUT (
.I0(RIOB33_X105Y117_IOB_X1Y118_I),
.I1(CLBLM_R_X3Y118_SLICE_X2Y118_AQ),
.I2(CLBLM_R_X5Y111_SLICE_X7Y111_AQ),
.I3(CLBLM_R_X7Y110_SLICE_X8Y110_AQ),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(CLBLM_R_X5Y112_SLICE_X7Y112_CO6),
.O5(CLBLM_R_X5Y111_SLICE_X7Y111_AO5),
.O6(CLBLM_R_X5Y111_SLICE_X7Y111_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y112_SLICE_X6Y112_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y112_SLICE_X6Y112_AO6),
.Q(CLBLM_R_X5Y112_SLICE_X6Y112_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffa9a90000a9a9)
  ) CLBLM_R_X5Y112_SLICE_X6Y112_DLUT (
.I0(CLBLM_R_X7Y110_SLICE_X9Y110_CQ),
.I1(CLBLM_R_X5Y113_SLICE_X6Y113_DO5),
.I2(CLBLL_L_X4Y121_SLICE_X4Y121_AQ),
.I3(1'b1),
.I4(RIOB33_X105Y121_IOB_X1Y121_I),
.I5(CLBLM_R_X5Y119_SLICE_X6Y119_BQ),
.O5(CLBLM_R_X5Y112_SLICE_X6Y112_DO5),
.O6(CLBLM_R_X5Y112_SLICE_X6Y112_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0f0f0f0b5f5f5fdb)
  ) CLBLM_R_X5Y112_SLICE_X6Y112_CLUT (
.I0(CLBLL_L_X4Y111_SLICE_X5Y111_AQ),
.I1(CLBLM_R_X5Y114_SLICE_X7Y114_AQ),
.I2(RIOB33_X105Y121_IOB_X1Y121_I),
.I3(CLBLM_R_X7Y120_SLICE_X9Y120_CQ),
.I4(CLBLM_R_X5Y114_SLICE_X7Y114_BO5),
.I5(CLBLM_L_X8Y115_SLICE_X10Y115_CQ),
.O5(CLBLM_R_X5Y112_SLICE_X6Y112_CO5),
.O6(CLBLM_R_X5Y112_SLICE_X6Y112_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hff55aa0057575757)
  ) CLBLM_R_X5Y112_SLICE_X6Y112_BLUT (
.I0(RIOB33_X105Y121_IOB_X1Y121_I),
.I1(CLBLM_R_X5Y119_SLICE_X6Y119_BQ),
.I2(CLBLM_R_X5Y112_SLICE_X6Y112_AQ),
.I3(CLBLM_L_X8Y115_SLICE_X10Y115_CQ),
.I4(CLBLM_R_X5Y111_SLICE_X7Y111_AQ),
.I5(1'b1),
.O5(CLBLM_R_X5Y112_SLICE_X6Y112_BO5),
.O6(CLBLM_R_X5Y112_SLICE_X6Y112_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfcecffee30203322)
  ) CLBLM_R_X5Y112_SLICE_X6Y112_ALUT (
.I0(CLBLM_R_X3Y118_SLICE_X2Y118_AQ),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(CLBLM_R_X5Y112_SLICE_X6Y112_AQ),
.I3(RIOB33_X105Y117_IOB_X1Y118_I),
.I4(CLBLM_R_X5Y112_SLICE_X6Y112_CO6),
.I5(CLBLM_R_X5Y125_SLICE_X6Y125_A5Q),
.O5(CLBLM_R_X5Y112_SLICE_X6Y112_AO5),
.O6(CLBLM_R_X5Y112_SLICE_X6Y112_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000001101)
  ) CLBLM_R_X5Y112_SLICE_X7Y112_DLUT (
.I0(RIOB33_X105Y117_IOB_X1Y118_I),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(CLBLM_R_X7Y109_SLICE_X8Y109_AQ),
.I3(RIOB33_X105Y105_IOB_X1Y105_I),
.I4(CLBLM_R_X3Y118_SLICE_X2Y118_AQ),
.I5(CLBLM_R_X5Y116_SLICE_X7Y116_CQ),
.O5(CLBLM_R_X5Y112_SLICE_X7Y112_DO5),
.O6(CLBLM_R_X5Y112_SLICE_X7Y112_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hfdce0000ffcc0000)
  ) CLBLM_R_X5Y112_SLICE_X7Y112_CLUT (
.I0(CLBLM_R_X5Y114_SLICE_X7Y114_AQ),
.I1(CLBLM_R_X7Y118_SLICE_X9Y118_CQ),
.I2(CLBLM_R_X7Y120_SLICE_X9Y120_CQ),
.I3(CLBLM_R_X5Y115_SLICE_X7Y115_A5Q),
.I4(RIOB33_X105Y121_IOB_X1Y121_I),
.I5(CLBLM_R_X5Y114_SLICE_X7Y114_BO6),
.O5(CLBLM_R_X5Y112_SLICE_X7Y112_CO5),
.O6(CLBLM_R_X5Y112_SLICE_X7Y112_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000aaaa000088a0)
  ) CLBLM_R_X5Y112_SLICE_X7Y112_BLUT (
.I0(CLBLM_R_X5Y112_SLICE_X7Y112_DO6),
.I1(CLBLM_L_X8Y115_SLICE_X10Y115_CQ),
.I2(CLBLM_R_X5Y111_SLICE_X7Y111_AQ),
.I3(RIOB33_X105Y121_IOB_X1Y121_I),
.I4(CLBLM_R_X5Y110_SLICE_X7Y110_DO5),
.I5(CLBLM_R_X5Y112_SLICE_X7Y112_AO5),
.O5(CLBLM_R_X5Y112_SLICE_X7Y112_BO5),
.O6(CLBLM_R_X5Y112_SLICE_X7Y112_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfff00d00000f000f)
  ) CLBLM_R_X5Y112_SLICE_X7Y112_ALUT (
.I0(RIOB33_X105Y105_IOB_X1Y105_I),
.I1(CLBLM_R_X3Y119_SLICE_X2Y119_AO6),
.I2(CLBLM_R_X5Y116_SLICE_X7Y116_CQ),
.I3(CLBLM_R_X7Y109_SLICE_X8Y109_AQ),
.I4(CLBLM_R_X7Y113_SLICE_X8Y113_BO6),
.I5(1'b1),
.O5(CLBLM_R_X5Y112_SLICE_X7Y112_AO5),
.O6(CLBLM_R_X5Y112_SLICE_X7Y112_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y113_SLICE_X6Y113_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y113_SLICE_X6Y113_AO6),
.Q(CLBLM_R_X5Y113_SLICE_X6Y113_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y113_SLICE_X6Y113_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y113_SLICE_X6Y113_BO6),
.Q(CLBLM_R_X5Y113_SLICE_X6Y113_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y113_SLICE_X6Y113_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y113_SLICE_X6Y113_CO6),
.Q(CLBLM_R_X5Y113_SLICE_X6Y113_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0002fffdffcfffcf)
  ) CLBLM_R_X5Y113_SLICE_X6Y113_DLUT (
.I0(CLBLL_L_X4Y121_SLICE_X4Y121_AQ),
.I1(CLBLM_R_X7Y120_SLICE_X9Y120_CQ),
.I2(CLBLL_L_X4Y114_SLICE_X4Y114_BQ),
.I3(CLBLM_R_X5Y114_SLICE_X7Y114_AQ),
.I4(CLBLM_R_X7Y119_SLICE_X8Y119_DQ),
.I5(1'b1),
.O5(CLBLM_R_X5Y113_SLICE_X6Y113_DO5),
.O6(CLBLM_R_X5Y113_SLICE_X6Y113_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f000aaf0f00088)
  ) CLBLM_R_X5Y113_SLICE_X6Y113_CLUT (
.I0(CLBLM_R_X3Y118_SLICE_X2Y118_AQ),
.I1(CLBLM_R_X5Y113_SLICE_X6Y113_CQ),
.I2(CLBLM_R_X5Y113_SLICE_X6Y113_AQ),
.I3(RIOB33_X105Y117_IOB_X1Y118_I),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(CLBLM_L_X8Y113_SLICE_X11Y113_CQ),
.O5(CLBLM_R_X5Y113_SLICE_X6Y113_CO5),
.O6(CLBLM_R_X5Y113_SLICE_X6Y113_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff060c0000060c)
  ) CLBLM_R_X5Y113_SLICE_X6Y113_BLUT (
.I0(CLBLL_L_X4Y113_SLICE_X4Y113_CO6),
.I1(CLBLM_R_X5Y113_SLICE_X6Y113_BQ),
.I2(CLBLM_R_X5Y110_SLICE_X7Y110_BQ),
.I3(CLBLL_L_X4Y113_SLICE_X4Y113_AQ),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(CLBLM_R_X7Y113_SLICE_X9Y113_BQ),
.O5(CLBLM_R_X5Y113_SLICE_X6Y113_BO5),
.O6(CLBLM_R_X5Y113_SLICE_X6Y113_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hccccccccfafafa00)
  ) CLBLM_R_X5Y113_SLICE_X6Y113_ALUT (
.I0(CLBLM_R_X5Y114_SLICE_X7Y114_DO6),
.I1(CLBLM_L_X8Y121_SLICE_X11Y121_BQ),
.I2(CLBLM_R_X5Y113_SLICE_X6Y113_AQ),
.I3(RIOB33_X105Y117_IOB_X1Y118_I),
.I4(CLBLM_R_X3Y118_SLICE_X2Y118_AQ),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLM_R_X5Y113_SLICE_X6Y113_AO5),
.O6(CLBLM_R_X5Y113_SLICE_X6Y113_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y113_SLICE_X7Y113_A5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y113_SLICE_X7Y113_AO5),
.Q(CLBLM_R_X5Y113_SLICE_X7Y113_A5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y113_SLICE_X7Y113_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y113_SLICE_X7Y113_AO6),
.Q(CLBLM_R_X5Y113_SLICE_X7Y113_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h3333333333333332)
  ) CLBLM_R_X5Y113_SLICE_X7Y113_DLUT (
.I0(CLBLM_R_X3Y111_SLICE_X3Y111_AQ),
.I1(CLBLM_R_X5Y117_SLICE_X7Y117_BQ),
.I2(CLBLM_R_X7Y119_SLICE_X8Y119_DQ),
.I3(CLBLM_R_X7Y111_SLICE_X8Y111_DO6),
.I4(CLBLM_R_X5Y113_SLICE_X7Y113_BO6),
.I5(CLBLL_L_X4Y116_SLICE_X4Y116_BQ),
.O5(CLBLM_R_X5Y113_SLICE_X7Y113_DO5),
.O6(CLBLM_R_X5Y113_SLICE_X7Y113_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h695a69a5c3f0c30f)
  ) CLBLM_R_X5Y113_SLICE_X7Y113_CLUT (
.I0(CLBLL_L_X4Y112_SLICE_X4Y112_DO6),
.I1(CLBLM_R_X5Y117_SLICE_X7Y117_BQ),
.I2(CLBLM_L_X8Y112_SLICE_X10Y112_CQ),
.I3(CLBLM_R_X7Y119_SLICE_X8Y119_CQ),
.I4(CLBLM_R_X5Y113_SLICE_X7Y113_DO6),
.I5(CLBLM_R_X5Y114_SLICE_X7Y114_BO6),
.O5(CLBLM_R_X5Y113_SLICE_X7Y113_CO5),
.O6(CLBLM_R_X5Y113_SLICE_X7Y113_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffffffffffffe)
  ) CLBLM_R_X5Y113_SLICE_X7Y113_BLUT (
.I0(CLBLM_R_X7Y122_SLICE_X8Y122_DQ),
.I1(CLBLM_R_X7Y109_SLICE_X8Y109_CQ),
.I2(CLBLM_R_X5Y113_SLICE_X7Y113_AQ),
.I3(CLBLM_R_X5Y121_SLICE_X7Y121_AQ),
.I4(CLBLL_L_X4Y111_SLICE_X5Y111_AQ),
.I5(CLBLL_L_X4Y111_SLICE_X4Y111_DQ),
.O5(CLBLM_R_X5Y113_SLICE_X7Y113_BO5),
.O6(CLBLM_R_X5Y113_SLICE_X7Y113_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hea40ea40f5f5a0a0)
  ) CLBLM_R_X5Y113_SLICE_X7Y113_ALUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(RIOB33_X105Y105_IOB_X1Y105_I),
.I2(CLBLM_R_X5Y113_SLICE_X7Y113_AQ),
.I3(CLBLM_L_X8Y112_SLICE_X10Y112_AQ),
.I4(CLBLM_R_X3Y114_SLICE_X3Y114_BQ),
.I5(1'b1),
.O5(CLBLM_R_X5Y113_SLICE_X7Y113_AO5),
.O6(CLBLM_R_X5Y113_SLICE_X7Y113_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y114_SLICE_X6Y114_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y114_SLICE_X6Y114_AO6),
.Q(CLBLM_R_X5Y114_SLICE_X6Y114_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y114_SLICE_X6Y114_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y114_SLICE_X6Y114_BO6),
.Q(CLBLM_R_X5Y114_SLICE_X6Y114_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y114_SLICE_X6Y114_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y114_SLICE_X6Y114_CO6),
.Q(CLBLM_R_X5Y114_SLICE_X6Y114_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y114_SLICE_X6Y114_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y114_SLICE_X6Y114_DO6),
.Q(CLBLM_R_X5Y114_SLICE_X6Y114_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaa0000fefe5454)
  ) CLBLM_R_X5Y114_SLICE_X6Y114_DLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_L_X10Y115_SLICE_X12Y115_BQ),
.I2(CLBLM_R_X5Y114_SLICE_X6Y114_DQ),
.I3(1'b1),
.I4(CLBLL_L_X4Y114_SLICE_X4Y114_CQ),
.I5(CLBLM_R_X5Y111_SLICE_X7Y111_DO6),
.O5(CLBLM_R_X5Y114_SLICE_X6Y114_DO5),
.O6(CLBLM_R_X5Y114_SLICE_X6Y114_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff000044114411)
  ) CLBLM_R_X5Y114_SLICE_X6Y114_CLUT (
.I0(RIOB33_X105Y105_IOB_X1Y105_I),
.I1(CLBLM_R_X7Y115_SLICE_X8Y115_BQ),
.I2(1'b1),
.I3(CLBLM_R_X5Y112_SLICE_X6Y112_BO5),
.I4(CLBLM_R_X5Y117_SLICE_X6Y117_CQ),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLM_R_X5Y114_SLICE_X6Y114_CO5),
.O6(CLBLM_R_X5Y114_SLICE_X6Y114_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hcc00cf03cc00fc30)
  ) CLBLM_R_X5Y114_SLICE_X6Y114_BLUT (
.I0(1'b1),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(CLBLL_L_X4Y111_SLICE_X4Y111_CQ),
.I3(CLBLM_R_X5Y118_SLICE_X6Y118_BQ),
.I4(RIOB33_X105Y105_IOB_X1Y105_I),
.I5(CLBLL_L_X4Y114_SLICE_X4Y114_DO6),
.O5(CLBLM_R_X5Y114_SLICE_X6Y114_BO5),
.O6(CLBLM_R_X5Y114_SLICE_X6Y114_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaafcfcaaaafc00)
  ) CLBLM_R_X5Y114_SLICE_X6Y114_ALUT (
.I0(CLBLL_L_X4Y119_SLICE_X4Y119_B5Q),
.I1(CLBLM_R_X5Y113_SLICE_X6Y113_CQ),
.I2(CLBLM_R_X5Y114_SLICE_X6Y114_AQ),
.I3(RIOB33_X105Y117_IOB_X1Y118_I),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(CLBLM_R_X3Y118_SLICE_X2Y118_AQ),
.O5(CLBLM_R_X5Y114_SLICE_X6Y114_AO5),
.O6(CLBLM_R_X5Y114_SLICE_X6Y114_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y114_SLICE_X7Y114_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y114_SLICE_X7Y114_AO6),
.Q(CLBLM_R_X5Y114_SLICE_X7Y114_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hf606fa0afa0afa0a)
  ) CLBLM_R_X5Y114_SLICE_X7Y114_DLUT (
.I0(CLBLM_R_X5Y121_SLICE_X7Y121_AQ),
.I1(CLBLM_R_X7Y120_SLICE_X9Y120_CQ),
.I2(RIOB33_X105Y121_IOB_X1Y121_I),
.I3(CLBLM_R_X7Y115_SLICE_X8Y115_CQ),
.I4(CLBLM_R_X5Y114_SLICE_X7Y114_AQ),
.I5(CLBLM_R_X5Y114_SLICE_X7Y114_BO6),
.O5(CLBLM_R_X5Y114_SLICE_X7Y114_DO5),
.O6(CLBLM_R_X5Y114_SLICE_X7Y114_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'he0c0c0c0e0e0e0e0)
  ) CLBLM_R_X5Y114_SLICE_X7Y114_CLUT (
.I0(CLBLL_L_X4Y120_SLICE_X4Y120_BO6),
.I1(CLBLM_R_X5Y112_SLICE_X7Y112_AO5),
.I2(CLBLM_R_X5Y112_SLICE_X7Y112_DO6),
.I3(CLBLM_R_X7Y115_SLICE_X8Y115_CQ),
.I4(CLBLM_R_X3Y114_SLICE_X3Y114_AQ),
.I5(RIOB33_X105Y121_IOB_X1Y121_I),
.O5(CLBLM_R_X5Y114_SLICE_X7Y114_CO5),
.O6(CLBLM_R_X5Y114_SLICE_X7Y114_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h00003333ccccffff)
  ) CLBLM_R_X5Y114_SLICE_X7Y114_BLUT (
.I0(1'b1),
.I1(CLBLL_L_X4Y114_SLICE_X4Y114_BQ),
.I2(1'b1),
.I3(1'b1),
.I4(CLBLL_L_X4Y121_SLICE_X4Y121_AQ),
.I5(1'b1),
.O5(CLBLM_R_X5Y114_SLICE_X7Y114_BO5),
.O6(CLBLM_R_X5Y114_SLICE_X7Y114_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hcc00cc00cca0cca0)
  ) CLBLM_R_X5Y114_SLICE_X7Y114_ALUT (
.I0(CLBLM_R_X5Y114_SLICE_X7Y114_AQ),
.I1(CLBLL_L_X4Y111_SLICE_X4Y111_DQ),
.I2(RIOB33_X105Y105_IOB_X1Y105_I),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(1'b1),
.I5(CLBLL_L_X4Y115_SLICE_X4Y115_CQ),
.O5(CLBLM_R_X5Y114_SLICE_X7Y114_AO5),
.O6(CLBLM_R_X5Y114_SLICE_X7Y114_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y115_SLICE_X6Y115_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y115_SLICE_X6Y115_AO6),
.Q(CLBLM_R_X5Y115_SLICE_X6Y115_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y115_SLICE_X6Y115_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y115_SLICE_X6Y115_BO6),
.Q(CLBLM_R_X5Y115_SLICE_X6Y115_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff7fffffffffff)
  ) CLBLM_R_X5Y115_SLICE_X6Y115_DLUT (
.I0(CLBLL_L_X4Y115_SLICE_X4Y115_DQ),
.I1(CLBLM_R_X5Y114_SLICE_X6Y114_CQ),
.I2(CLBLM_R_X7Y116_SLICE_X8Y116_BQ),
.I3(CLBLL_L_X4Y115_SLICE_X5Y115_BQ),
.I4(RIOB33_X105Y105_IOB_X1Y105_I),
.I5(CLBLM_R_X7Y115_SLICE_X8Y115_BQ),
.O5(CLBLM_R_X5Y115_SLICE_X6Y115_DO5),
.O6(CLBLM_R_X5Y115_SLICE_X6Y115_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h50504050f0f0c0f0)
  ) CLBLM_R_X5Y115_SLICE_X6Y115_CLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_R_X5Y121_SLICE_X6Y121_AQ),
.I2(RIOB33_X105Y105_IOB_X1Y105_I),
.I3(CLBLM_R_X7Y114_SLICE_X8Y114_BQ),
.I4(RIOB33_X105Y121_IOB_X1Y121_I),
.I5(1'b1),
.O5(CLBLM_R_X5Y115_SLICE_X6Y115_CO5),
.O6(CLBLM_R_X5Y115_SLICE_X6Y115_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h88888d8d8d8d8888)
  ) CLBLM_R_X5Y115_SLICE_X6Y115_BLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_L_X8Y115_SLICE_X11Y115_C5Q),
.I2(RIOB33_X105Y105_IOB_X1Y105_I),
.I3(1'b1),
.I4(CLBLM_R_X7Y113_SLICE_X8Y113_AQ),
.I5(CLBLM_R_X7Y115_SLICE_X8Y115_DO6),
.O5(CLBLM_R_X5Y115_SLICE_X6Y115_BO5),
.O6(CLBLM_R_X5Y115_SLICE_X6Y115_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hbb88b8b8bb88b8b8)
  ) CLBLM_R_X5Y115_SLICE_X6Y115_ALUT (
.I0(CLBLM_R_X7Y115_SLICE_X9Y115_DQ),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(CLBLM_R_X5Y115_SLICE_X6Y115_AQ),
.I3(CLBLM_R_X7Y115_SLICE_X8Y115_BQ),
.I4(CLBLM_R_X5Y115_SLICE_X6Y115_CO5),
.I5(1'b1),
.O5(CLBLM_R_X5Y115_SLICE_X6Y115_AO5),
.O6(CLBLM_R_X5Y115_SLICE_X6Y115_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y115_SLICE_X7Y115_A5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y115_SLICE_X7Y115_AO5),
.Q(CLBLM_R_X5Y115_SLICE_X7Y115_A5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y115_SLICE_X7Y115_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y115_SLICE_X7Y115_AO6),
.Q(CLBLM_R_X5Y115_SLICE_X7Y115_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y115_SLICE_X7Y115_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y115_SLICE_X7Y115_BO6),
.Q(CLBLM_R_X5Y115_SLICE_X7Y115_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000ffff0000fd55)
  ) CLBLM_R_X5Y115_SLICE_X7Y115_DLUT (
.I0(CLBLM_R_X5Y115_SLICE_X7Y115_CO5),
.I1(CLBLM_L_X8Y114_SLICE_X10Y114_C5Q),
.I2(CLBLL_L_X4Y115_SLICE_X5Y115_AQ),
.I3(RIOB33_X105Y121_IOB_X1Y121_I),
.I4(CLBLM_R_X5Y112_SLICE_X7Y112_AO5),
.I5(CLBLL_L_X2Y120_SLICE_X0Y120_CO6),
.O5(CLBLM_R_X5Y115_SLICE_X7Y115_DO5),
.O6(CLBLM_R_X5Y115_SLICE_X7Y115_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hfcccfdcd22222222)
  ) CLBLM_R_X5Y115_SLICE_X7Y115_CLUT (
.I0(RIOB33_X105Y105_IOB_X1Y105_I),
.I1(CLBLM_R_X5Y116_SLICE_X7Y116_CQ),
.I2(CLBLM_R_X7Y109_SLICE_X8Y109_AQ),
.I3(CLBLL_L_X4Y113_SLICE_X5Y113_DO6),
.I4(CLBLL_L_X2Y119_SLICE_X0Y119_BO6),
.I5(1'b1),
.O5(CLBLM_R_X5Y115_SLICE_X7Y115_CO5),
.O6(CLBLM_R_X5Y115_SLICE_X7Y115_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaa00f0aaaa00f0)
  ) CLBLM_R_X5Y115_SLICE_X7Y115_BLUT (
.I0(CLBLM_R_X5Y110_SLICE_X7Y110_AQ),
.I1(1'b1),
.I2(CLBLM_R_X5Y119_SLICE_X6Y119_BQ),
.I3(RIOB33_X105Y105_IOB_X1Y105_I),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(1'b1),
.O5(CLBLM_R_X5Y115_SLICE_X7Y115_BO5),
.O6(CLBLM_R_X5Y115_SLICE_X7Y115_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hacacacacc0cfc0c0)
  ) CLBLM_R_X5Y115_SLICE_X7Y115_ALUT (
.I0(CLBLM_R_X7Y115_SLICE_X9Y115_CQ),
.I1(CLBLM_L_X8Y117_SLICE_X11Y117_AQ),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(RIOB33_X105Y105_IOB_X1Y105_I),
.I4(CLBLM_R_X5Y115_SLICE_X7Y115_A5Q),
.I5(1'b1),
.O5(CLBLM_R_X5Y115_SLICE_X7Y115_AO5),
.O6(CLBLM_R_X5Y115_SLICE_X7Y115_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y116_SLICE_X6Y116_A5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y116_SLICE_X6Y116_CO6),
.Q(CLBLM_R_X5Y116_SLICE_X6Y116_A5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y116_SLICE_X6Y116_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y116_SLICE_X6Y116_AO6),
.Q(CLBLM_R_X5Y116_SLICE_X6Y116_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y116_SLICE_X6Y116_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y116_SLICE_X6Y116_BO6),
.Q(CLBLM_R_X5Y116_SLICE_X6Y116_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y116_SLICE_X6Y116_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y116_SLICE_X6Y116_DO6),
.Q(CLBLM_R_X5Y116_SLICE_X6Y116_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hcc00cc55cc00ccaa)
  ) CLBLM_R_X5Y116_SLICE_X6Y116_DLUT (
.I0(CLBLM_R_X5Y116_SLICE_X6Y116_CO5),
.I1(CLBLM_R_X5Y116_SLICE_X6Y116_AQ),
.I2(1'b1),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(RIOB33_X105Y105_IOB_X1Y105_I),
.I5(CLBLM_R_X7Y116_SLICE_X8Y116_BQ),
.O5(CLBLM_R_X5Y116_SLICE_X6Y116_DO5),
.O6(CLBLM_R_X5Y116_SLICE_X6Y116_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaaff00e0e0e0e0)
  ) CLBLM_R_X5Y116_SLICE_X6Y116_CLUT (
.I0(CLBLL_L_X4Y115_SLICE_X5Y115_AQ),
.I1(CLBLM_L_X8Y114_SLICE_X10Y114_C5Q),
.I2(RIOB33_X105Y121_IOB_X1Y121_I),
.I3(CLBLM_R_X5Y123_SLICE_X7Y123_AQ),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(1'b1),
.O5(CLBLM_R_X5Y116_SLICE_X6Y116_CO5),
.O6(CLBLM_R_X5Y116_SLICE_X6Y116_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf1f40104f4f40404)
  ) CLBLM_R_X5Y116_SLICE_X6Y116_BLUT (
.I0(CLBLM_R_X5Y110_SLICE_X7Y110_BQ),
.I1(CLBLM_R_X5Y116_SLICE_X6Y116_BQ),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLL_L_X4Y118_SLICE_X5Y118_AQ),
.I4(CLBLM_L_X10Y114_SLICE_X13Y114_D5Q),
.I5(CLBLM_R_X5Y116_SLICE_X7Y116_BO5),
.O5(CLBLM_R_X5Y116_SLICE_X6Y116_BO5),
.O6(CLBLM_R_X5Y116_SLICE_X6Y116_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hccccff00ccccf0f0)
  ) CLBLM_R_X5Y116_SLICE_X6Y116_ALUT (
.I0(1'b1),
.I1(CLBLM_L_X8Y119_SLICE_X10Y119_AQ),
.I2(CLBLM_R_X5Y116_SLICE_X6Y116_AQ),
.I3(CLBLL_L_X4Y111_SLICE_X4Y111_CQ),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(CLBLM_R_X5Y115_SLICE_X6Y115_CO5),
.O5(CLBLM_R_X5Y116_SLICE_X6Y116_AO5),
.O6(CLBLM_R_X5Y116_SLICE_X6Y116_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y116_SLICE_X7Y116_A5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y116_SLICE_X7Y116_BO6),
.Q(CLBLM_R_X5Y116_SLICE_X7Y116_A5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y116_SLICE_X7Y116_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y116_SLICE_X7Y116_AO6),
.Q(CLBLM_R_X5Y116_SLICE_X7Y116_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y116_SLICE_X7Y116_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y116_SLICE_X7Y116_CO6),
.Q(CLBLM_R_X5Y116_SLICE_X7Y116_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h000f002d000f000f)
  ) CLBLM_R_X5Y116_SLICE_X7Y116_DLUT (
.I0(CLBLL_L_X4Y121_SLICE_X4Y121_AQ),
.I1(CLBLM_R_X7Y120_SLICE_X9Y120_CQ),
.I2(CLBLM_R_X7Y111_SLICE_X8Y111_AQ),
.I3(CLBLM_R_X5Y116_SLICE_X7Y116_A5Q),
.I4(CLBLM_R_X5Y114_SLICE_X7Y114_AQ),
.I5(CLBLL_L_X4Y114_SLICE_X4Y114_BQ),
.O5(CLBLM_R_X5Y116_SLICE_X7Y116_DO5),
.O6(CLBLM_R_X5Y116_SLICE_X7Y116_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffe0f0ef0f40004)
  ) CLBLM_R_X5Y116_SLICE_X7Y116_CLUT (
.I0(CLBLM_R_X3Y118_SLICE_X2Y118_AQ),
.I1(CLBLM_R_X5Y116_SLICE_X7Y116_CQ),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(RIOB33_X105Y117_IOB_X1Y118_I),
.I4(CLBLM_R_X7Y124_SLICE_X8Y124_A5Q),
.I5(CLBLM_R_X5Y110_SLICE_X7Y110_BQ),
.O5(CLBLM_R_X5Y116_SLICE_X7Y116_CO5),
.O6(CLBLM_R_X5Y116_SLICE_X7Y116_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hd1d1d1c00000ff00)
  ) CLBLM_R_X5Y116_SLICE_X7Y116_BLUT (
.I0(CLBLM_R_X5Y116_SLICE_X7Y116_DO6),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(CLBLM_R_X5Y123_SLICE_X6Y123_AQ),
.I3(RIOB33_X105Y117_IOB_X1Y118_I),
.I4(CLBLM_R_X3Y118_SLICE_X2Y118_AQ),
.I5(1'b1),
.O5(CLBLM_R_X5Y116_SLICE_X7Y116_BO5),
.O6(CLBLM_R_X5Y116_SLICE_X7Y116_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hdd88dd88d8d8d8d8)
  ) CLBLM_R_X5Y116_SLICE_X7Y116_ALUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_R_X7Y113_SLICE_X8Y113_AQ),
.I2(CLBLM_R_X5Y116_SLICE_X7Y116_AQ),
.I3(CLBLM_L_X10Y116_SLICE_X13Y116_AQ),
.I4(1'b1),
.I5(CLBLM_R_X5Y115_SLICE_X6Y115_CO5),
.O5(CLBLM_R_X5Y116_SLICE_X7Y116_AO5),
.O6(CLBLM_R_X5Y116_SLICE_X7Y116_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y117_SLICE_X6Y117_D5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y117_SLICE_X6Y117_DO5),
.Q(CLBLM_R_X5Y117_SLICE_X6Y117_D5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y117_SLICE_X6Y117_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y117_SLICE_X6Y117_AO6),
.Q(CLBLM_R_X5Y117_SLICE_X6Y117_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y117_SLICE_X6Y117_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y117_SLICE_X6Y117_BO6),
.Q(CLBLM_R_X5Y117_SLICE_X6Y117_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y117_SLICE_X6Y117_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y117_SLICE_X6Y117_CO6),
.Q(CLBLM_R_X5Y117_SLICE_X6Y117_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y117_SLICE_X6Y117_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y117_SLICE_X6Y117_DO6),
.Q(CLBLM_R_X5Y117_SLICE_X6Y117_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hf5f5a0a0ff55aa00)
  ) CLBLM_R_X5Y117_SLICE_X6Y117_DLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(1'b1),
.I2(CLBLM_R_X5Y113_SLICE_X6Y113_CQ),
.I3(CLBLM_R_X5Y121_SLICE_X6Y121_BQ),
.I4(RIOB33_X105Y101_IOB_X1Y101_I),
.I5(1'b1),
.O5(CLBLM_R_X5Y117_SLICE_X6Y117_DO5),
.O6(CLBLM_R_X5Y117_SLICE_X6Y117_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'haa00fe54fe54fe54)
  ) CLBLM_R_X5Y117_SLICE_X6Y117_CLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_R_X5Y117_SLICE_X6Y117_CQ),
.I2(CLBLL_L_X4Y118_SLICE_X5Y118_AQ),
.I3(CLBLM_L_X10Y123_SLICE_X13Y123_AQ),
.I4(CLBLM_L_X8Y112_SLICE_X10Y112_CQ),
.I5(CLBLL_L_X2Y112_SLICE_X1Y112_BQ),
.O5(CLBLM_R_X5Y117_SLICE_X6Y117_CO5),
.O6(CLBLM_R_X5Y117_SLICE_X6Y117_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff0f0ffffd0f0d)
  ) CLBLM_R_X5Y117_SLICE_X6Y117_BLUT (
.I0(RIOB33_X105Y135_IOB_X1Y136_I),
.I1(CLBLM_L_X8Y121_SLICE_X10Y121_DO6),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(RIOB33_X105Y135_IOB_X1Y135_I),
.I4(CLBLM_R_X3Y111_SLICE_X3Y111_AQ),
.I5(RIOB33_X105Y131_IOB_X1Y131_I),
.O5(CLBLM_R_X5Y117_SLICE_X6Y117_BO5),
.O6(CLBLM_R_X5Y117_SLICE_X6Y117_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hba10fe54ba10ba10)
  ) CLBLM_R_X5Y117_SLICE_X6Y117_ALUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLL_L_X4Y111_SLICE_X4Y111_AO5),
.I2(CLBLM_R_X5Y117_SLICE_X6Y117_AQ),
.I3(CLBLL_L_X4Y110_SLICE_X5Y110_BQ),
.I4(RIOB33_X105Y105_IOB_X1Y105_I),
.I5(CLBLL_L_X4Y120_SLICE_X4Y120_AO6),
.O5(CLBLM_R_X5Y117_SLICE_X6Y117_AO5),
.O6(CLBLM_R_X5Y117_SLICE_X6Y117_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y117_SLICE_X7Y117_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y117_SLICE_X7Y117_AO6),
.Q(CLBLM_R_X5Y117_SLICE_X7Y117_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y117_SLICE_X7Y117_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y117_SLICE_X7Y117_BO6),
.Q(CLBLM_R_X5Y117_SLICE_X7Y117_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000030000000300)
  ) CLBLM_R_X5Y117_SLICE_X7Y117_DLUT (
.I0(1'b1),
.I1(RIOB33_X105Y135_IOB_X1Y135_I),
.I2(RIOB33_X105Y135_IOB_X1Y136_I),
.I3(RIOB33_X105Y131_IOB_X1Y131_I),
.I4(CLBLM_L_X8Y121_SLICE_X10Y121_DO6),
.I5(1'b1),
.O5(CLBLM_R_X5Y117_SLICE_X7Y117_DO5),
.O6(CLBLM_R_X5Y117_SLICE_X7Y117_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffffffff0004)
  ) CLBLM_R_X5Y117_SLICE_X7Y117_CLUT (
.I0(CLBLL_L_X4Y120_SLICE_X5Y120_AO6),
.I1(CLBLM_R_X5Y111_SLICE_X7Y111_CO6),
.I2(CLBLL_L_X2Y120_SLICE_X1Y120_DO6),
.I3(CLBLM_R_X3Y119_SLICE_X2Y119_AO6),
.I4(CLBLM_R_X7Y120_SLICE_X9Y120_D5Q),
.I5(CLBLM_R_X5Y118_SLICE_X7Y118_DO6),
.O5(CLBLM_R_X5Y117_SLICE_X7Y117_CO5),
.O6(CLBLM_R_X5Y117_SLICE_X7Y117_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hff0c000cff0c000c)
  ) CLBLM_R_X5Y117_SLICE_X7Y117_BLUT (
.I0(1'b1),
.I1(CLBLM_R_X5Y117_SLICE_X7Y117_BQ),
.I2(RIOB33_X105Y105_IOB_X1Y105_I),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLM_L_X12Y118_SLICE_X16Y118_BQ),
.I5(1'b1),
.O5(CLBLM_R_X5Y117_SLICE_X7Y117_BO5),
.O6(CLBLM_R_X5Y117_SLICE_X7Y117_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfbf80b08fff00f00)
  ) CLBLM_R_X5Y117_SLICE_X7Y117_ALUT (
.I0(CLBLM_R_X5Y117_SLICE_X7Y117_AQ),
.I1(CLBLL_L_X2Y112_SLICE_X1Y112_BQ),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLM_R_X3Y112_SLICE_X3Y112_AQ),
.I4(CLBLM_R_X5Y123_SLICE_X7Y123_AQ),
.I5(CLBLM_L_X8Y112_SLICE_X10Y112_CQ),
.O5(CLBLM_R_X5Y117_SLICE_X7Y117_AO5),
.O6(CLBLM_R_X5Y117_SLICE_X7Y117_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y118_SLICE_X6Y118_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y118_SLICE_X6Y118_AO6),
.Q(CLBLM_R_X5Y118_SLICE_X6Y118_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y118_SLICE_X6Y118_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y118_SLICE_X6Y118_BO6),
.Q(CLBLM_R_X5Y118_SLICE_X6Y118_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y118_SLICE_X6Y118_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y118_SLICE_X6Y118_CO6),
.Q(CLBLM_R_X5Y118_SLICE_X6Y118_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0aceffff0ace0ace)
  ) CLBLM_R_X5Y118_SLICE_X6Y118_DLUT (
.I0(CLBLM_R_X7Y117_SLICE_X9Y117_CQ),
.I1(CLBLM_R_X5Y117_SLICE_X6Y117_CQ),
.I2(CLBLM_R_X3Y121_SLICE_X2Y121_AO5),
.I3(CLBLM_R_X3Y121_SLICE_X2Y121_AO6),
.I4(CLBLL_L_X2Y120_SLICE_X0Y120_AO5),
.I5(CLBLL_L_X4Y117_SLICE_X5Y117_CQ),
.O5(CLBLM_R_X5Y118_SLICE_X6Y118_DO5),
.O6(CLBLM_R_X5Y118_SLICE_X6Y118_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hcc00cc00ee22ec20)
  ) CLBLM_R_X5Y118_SLICE_X6Y118_CLUT (
.I0(CLBLM_R_X3Y118_SLICE_X2Y118_AQ),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(CLBLM_R_X5Y110_SLICE_X6Y110_AQ),
.I3(CLBLM_R_X5Y122_SLICE_X7Y122_A5Q),
.I4(CLBLM_R_X5Y118_SLICE_X6Y118_CQ),
.I5(RIOB33_X105Y117_IOB_X1Y118_I),
.O5(CLBLM_R_X5Y118_SLICE_X6Y118_CO5),
.O6(CLBLM_R_X5Y118_SLICE_X6Y118_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfafafafc0a0a0a0c)
  ) CLBLM_R_X5Y118_SLICE_X6Y118_BLUT (
.I0(CLBLM_R_X5Y118_SLICE_X6Y118_CQ),
.I1(CLBLM_R_X5Y118_SLICE_X6Y118_BQ),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(RIOB33_X105Y117_IOB_X1Y118_I),
.I4(CLBLM_R_X3Y118_SLICE_X2Y118_AQ),
.I5(CLBLM_R_X3Y116_SLICE_X3Y116_CQ),
.O5(CLBLM_R_X5Y118_SLICE_X6Y118_BO5),
.O6(CLBLM_R_X5Y118_SLICE_X6Y118_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff50d8000050d8)
  ) CLBLM_R_X5Y118_SLICE_X6Y118_ALUT (
.I0(CLBLL_L_X4Y111_SLICE_X4Y111_AO5),
.I1(CLBLL_L_X4Y120_SLICE_X4Y120_BO6),
.I2(CLBLM_R_X5Y118_SLICE_X6Y118_AQ),
.I3(RIOB33_X105Y105_IOB_X1Y105_I),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(CLBLM_R_X7Y120_SLICE_X9Y120_A5Q),
.O5(CLBLM_R_X5Y118_SLICE_X6Y118_AO5),
.O6(CLBLM_R_X5Y118_SLICE_X6Y118_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y118_SLICE_X7Y118_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y118_SLICE_X7Y118_AO6),
.Q(CLBLM_R_X5Y118_SLICE_X7Y118_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffffffffffffd)
  ) CLBLM_R_X5Y118_SLICE_X7Y118_DLUT (
.I0(RIOB33_X105Y105_IOB_X1Y105_I),
.I1(CLBLM_R_X5Y122_SLICE_X7Y122_A5Q),
.I2(CLBLM_L_X8Y119_SLICE_X11Y119_C5Q),
.I3(CLBLM_R_X5Y121_SLICE_X7Y121_A5Q),
.I4(CLBLM_R_X5Y118_SLICE_X7Y118_BO5),
.I5(CLBLM_R_X3Y117_SLICE_X3Y117_AQ),
.O5(CLBLM_R_X5Y118_SLICE_X7Y118_DO5),
.O6(CLBLM_R_X5Y118_SLICE_X7Y118_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hc0c4c4c4c0cccccc)
  ) CLBLM_R_X5Y118_SLICE_X7Y118_CLUT (
.I0(CLBLL_L_X4Y120_SLICE_X4Y120_AO6),
.I1(CLBLM_R_X3Y113_SLICE_X3Y113_DO6),
.I2(CLBLM_R_X5Y120_SLICE_X7Y120_DO6),
.I3(CLBLL_L_X4Y120_SLICE_X4Y120_BO6),
.I4(CLBLM_R_X3Y120_SLICE_X3Y120_BO6),
.I5(CLBLL_L_X2Y120_SLICE_X0Y120_CO6),
.O5(CLBLM_R_X5Y118_SLICE_X7Y118_CO5),
.O6(CLBLM_R_X5Y118_SLICE_X7Y118_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffffefffefffe)
  ) CLBLM_R_X5Y118_SLICE_X7Y118_BLUT (
.I0(CLBLL_L_X4Y119_SLICE_X4Y119_B5Q),
.I1(CLBLM_R_X5Y116_SLICE_X6Y116_A5Q),
.I2(CLBLM_R_X5Y119_SLICE_X6Y119_B5Q),
.I3(CLBLM_R_X5Y125_SLICE_X6Y125_A5Q),
.I4(CLBLM_R_X3Y117_SLICE_X3Y117_AQ),
.I5(1'b1),
.O5(CLBLM_R_X5Y118_SLICE_X7Y118_BO5),
.O6(CLBLM_R_X5Y118_SLICE_X7Y118_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffcfcfcff000000)
  ) CLBLM_R_X5Y118_SLICE_X7Y118_ALUT (
.I0(1'b1),
.I1(CLBLM_R_X5Y114_SLICE_X6Y114_BQ),
.I2(CLBLM_R_X5Y118_SLICE_X7Y118_AQ),
.I3(CLBLM_R_X7Y118_SLICE_X8Y118_DQ),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(CLBLM_R_X5Y115_SLICE_X6Y115_CO6),
.O5(CLBLM_R_X5Y118_SLICE_X7Y118_AO5),
.O6(CLBLM_R_X5Y118_SLICE_X7Y118_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y119_SLICE_X6Y119_B5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y119_SLICE_X6Y119_BO5),
.Q(CLBLM_R_X5Y119_SLICE_X6Y119_B5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y119_SLICE_X6Y119_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y119_SLICE_X6Y119_AO6),
.Q(CLBLM_R_X5Y119_SLICE_X6Y119_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y119_SLICE_X6Y119_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y119_SLICE_X6Y119_BO6),
.Q(CLBLM_R_X5Y119_SLICE_X6Y119_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y119_SLICE_X6Y119_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y119_SLICE_X6Y119_CO6),
.Q(CLBLM_R_X5Y119_SLICE_X6Y119_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000800)
  ) CLBLM_R_X5Y119_SLICE_X6Y119_DLUT (
.I0(RIOB33_X105Y131_IOB_X1Y132_I),
.I1(RIOB33_X105Y131_IOB_X1Y131_I),
.I2(RIOB33_X105Y133_IOB_X1Y134_I),
.I3(CLBLM_L_X8Y118_SLICE_X10Y118_D5Q),
.I4(RIOB33_X105Y133_IOB_X1Y133_I),
.I5(CLBLM_R_X3Y122_SLICE_X3Y122_AO6),
.O5(CLBLM_R_X5Y119_SLICE_X6Y119_DO5),
.O6(CLBLM_R_X5Y119_SLICE_X6Y119_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f0f0f0ffcc0000)
  ) CLBLM_R_X5Y119_SLICE_X6Y119_CLUT (
.I0(1'b1),
.I1(CLBLM_R_X5Y119_SLICE_X6Y119_CQ),
.I2(CLBLM_R_X5Y115_SLICE_X6Y115_AQ),
.I3(CLBLM_L_X8Y119_SLICE_X11Y119_C5Q),
.I4(CLBLM_R_X3Y116_SLICE_X2Y116_DO6),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLM_R_X5Y119_SLICE_X6Y119_CO5),
.O6(CLBLM_R_X5Y119_SLICE_X6Y119_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf000fa0acfc0cfc0)
  ) CLBLM_R_X5Y119_SLICE_X6Y119_BLUT (
.I0(CLBLM_R_X7Y120_SLICE_X8Y120_DQ),
.I1(CLBLL_L_X4Y118_SLICE_X5Y118_BQ),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLM_R_X7Y121_SLICE_X9Y121_BQ),
.I4(RIOB33_X105Y105_IOB_X1Y105_I),
.I5(1'b1),
.O5(CLBLM_R_X5Y119_SLICE_X6Y119_BO5),
.O6(CLBLM_R_X5Y119_SLICE_X6Y119_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'heefaeefaeefaeeaa)
  ) CLBLM_R_X5Y119_SLICE_X6Y119_ALUT (
.I0(CLBLM_R_X5Y114_SLICE_X7Y114_CO6),
.I1(CLBLM_R_X5Y121_SLICE_X6Y121_A5Q),
.I2(CLBLM_R_X5Y119_SLICE_X6Y119_AQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLM_R_X3Y118_SLICE_X2Y118_AQ),
.I5(RIOB33_X105Y117_IOB_X1Y118_I),
.O5(CLBLM_R_X5Y119_SLICE_X6Y119_AO5),
.O6(CLBLM_R_X5Y119_SLICE_X6Y119_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffff0f0fffff0f0)
  ) CLBLM_R_X5Y119_SLICE_X7Y119_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(CLBLM_R_X5Y122_SLICE_X7Y122_A5Q),
.I3(1'b1),
.I4(CLBLM_R_X5Y121_SLICE_X7Y121_A5Q),
.I5(1'b1),
.O5(CLBLM_R_X5Y119_SLICE_X7Y119_DO5),
.O6(CLBLM_R_X5Y119_SLICE_X7Y119_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffffffffffaff)
  ) CLBLM_R_X5Y119_SLICE_X7Y119_CLUT (
.I0(CLBLM_R_X7Y120_SLICE_X9Y120_D5Q),
.I1(1'b1),
.I2(CLBLM_R_X5Y119_SLICE_X6Y119_B5Q),
.I3(RIOB33_X105Y105_IOB_X1Y105_I),
.I4(CLBLM_R_X5Y121_SLICE_X7Y121_A5Q),
.I5(CLBLM_R_X5Y119_SLICE_X7Y119_BO6),
.O5(CLBLM_R_X5Y119_SLICE_X7Y119_CO5),
.O6(CLBLM_R_X5Y119_SLICE_X7Y119_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffffffffffffe)
  ) CLBLM_R_X5Y119_SLICE_X7Y119_BLUT (
.I0(CLBLL_L_X4Y119_SLICE_X4Y119_B5Q),
.I1(CLBLM_R_X5Y122_SLICE_X7Y122_A5Q),
.I2(CLBLM_R_X3Y117_SLICE_X3Y117_AQ),
.I3(CLBLM_R_X5Y125_SLICE_X6Y125_A5Q),
.I4(CLBLM_R_X5Y116_SLICE_X6Y116_A5Q),
.I5(CLBLM_L_X8Y119_SLICE_X11Y119_C5Q),
.O5(CLBLM_R_X5Y119_SLICE_X7Y119_BO5),
.O6(CLBLM_R_X5Y119_SLICE_X7Y119_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffffffffffef)
  ) CLBLM_R_X5Y119_SLICE_X7Y119_ALUT (
.I0(CLBLM_R_X5Y119_SLICE_X7Y119_DO6),
.I1(CLBLM_R_X5Y118_SLICE_X7Y118_BO6),
.I2(RIOB33_X105Y105_IOB_X1Y105_I),
.I3(CLBLM_R_X7Y120_SLICE_X9Y120_D5Q),
.I4(CLBLL_L_X2Y119_SLICE_X1Y119_BO6),
.I5(CLBLM_L_X8Y119_SLICE_X11Y119_C5Q),
.O5(CLBLM_R_X5Y119_SLICE_X7Y119_AO5),
.O6(CLBLM_R_X5Y119_SLICE_X7Y119_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y120_SLICE_X6Y120_A5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y120_SLICE_X6Y120_AO5),
.Q(CLBLM_R_X5Y120_SLICE_X6Y120_A5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y120_SLICE_X6Y120_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y120_SLICE_X6Y120_AO6),
.Q(CLBLM_R_X5Y120_SLICE_X6Y120_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y120_SLICE_X6Y120_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y120_SLICE_X6Y120_BO6),
.Q(CLBLM_R_X5Y120_SLICE_X6Y120_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0a0a0a0aff0aff0a)
  ) CLBLM_R_X5Y120_SLICE_X6Y120_DLUT (
.I0(CLBLM_R_X5Y120_SLICE_X7Y120_AQ),
.I1(1'b1),
.I2(CLBLL_L_X2Y120_SLICE_X0Y120_AO5),
.I3(CLBLM_R_X7Y112_SLICE_X8Y112_CQ),
.I4(1'b1),
.I5(CLBLM_R_X3Y121_SLICE_X2Y121_AO6),
.O5(CLBLM_R_X5Y120_SLICE_X6Y120_DO5),
.O6(CLBLM_R_X5Y120_SLICE_X6Y120_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h5f0f55005f0f5500)
  ) CLBLM_R_X5Y120_SLICE_X6Y120_CLUT (
.I0(CLBLM_R_X3Y121_SLICE_X2Y121_AO5),
.I1(1'b1),
.I2(CLBLL_L_X2Y120_SLICE_X0Y120_AO5),
.I3(CLBLM_R_X5Y117_SLICE_X7Y117_AQ),
.I4(CLBLM_L_X8Y118_SLICE_X10Y118_AQ),
.I5(1'b1),
.O5(CLBLM_R_X5Y120_SLICE_X6Y120_CO5),
.O6(CLBLM_R_X5Y120_SLICE_X6Y120_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfff00f00fcfc0c0c)
  ) CLBLM_R_X5Y120_SLICE_X6Y120_BLUT (
.I0(1'b1),
.I1(CLBLM_R_X5Y120_SLICE_X6Y120_BQ),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLM_R_X7Y116_SLICE_X8Y116_BQ),
.I4(CLBLL_L_X4Y117_SLICE_X5Y117_AQ),
.I5(CLBLM_R_X5Y115_SLICE_X6Y115_CO5),
.O5(CLBLM_R_X5Y120_SLICE_X6Y120_BO5),
.O6(CLBLM_R_X5Y120_SLICE_X6Y120_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfff000f0eeaaeeaa)
  ) CLBLM_R_X5Y120_SLICE_X6Y120_ALUT (
.I0(CLBLM_R_X7Y122_SLICE_X9Y122_CO6),
.I1(CLBLM_R_X5Y119_SLICE_X6Y119_CQ),
.I2(CLBLL_L_X4Y120_SLICE_X4Y120_BO6),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLM_R_X7Y109_SLICE_X8Y109_AQ),
.I5(1'b1),
.O5(CLBLM_R_X5Y120_SLICE_X6Y120_AO5),
.O6(CLBLM_R_X5Y120_SLICE_X6Y120_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y120_SLICE_X7Y120_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y120_SLICE_X7Y120_AO6),
.Q(CLBLM_R_X5Y120_SLICE_X7Y120_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y120_SLICE_X7Y120_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y120_SLICE_X7Y120_BO6),
.Q(CLBLM_R_X5Y120_SLICE_X7Y120_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y120_SLICE_X7Y120_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y120_SLICE_X7Y120_CO6),
.Q(CLBLM_R_X5Y120_SLICE_X7Y120_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h31f531f566999966)
  ) CLBLM_R_X5Y120_SLICE_X7Y120_DLUT (
.I0(CLBLM_R_X3Y119_SLICE_X2Y119_AO6),
.I1(CLBLL_L_X4Y120_SLICE_X5Y120_DO6),
.I2(CLBLL_L_X2Y119_SLICE_X0Y119_BO6),
.I3(CLBLL_L_X2Y120_SLICE_X1Y120_DO6),
.I4(CLBLM_R_X3Y120_SLICE_X3Y120_BO6),
.I5(1'b1),
.O5(CLBLM_R_X5Y120_SLICE_X7Y120_DO5),
.O6(CLBLM_R_X5Y120_SLICE_X7Y120_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaafefe00005454)
  ) CLBLM_R_X5Y120_SLICE_X7Y120_CLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_R_X5Y120_SLICE_X7Y120_CQ),
.I2(CLBLM_R_X5Y121_SLICE_X7Y121_A5Q),
.I3(1'b1),
.I4(CLBLM_R_X3Y116_SLICE_X2Y116_DO6),
.I5(CLBLM_L_X10Y120_SLICE_X12Y120_CQ),
.O5(CLBLM_R_X5Y120_SLICE_X7Y120_CO5),
.O6(CLBLM_R_X5Y120_SLICE_X7Y120_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfff0fcfc0f000c0c)
  ) CLBLM_R_X5Y120_SLICE_X7Y120_BLUT (
.I0(1'b1),
.I1(CLBLM_R_X5Y120_SLICE_X7Y120_BQ),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLM_R_X7Y113_SLICE_X8Y113_AQ),
.I4(CLBLM_R_X5Y115_SLICE_X6Y115_CO5),
.I5(CLBLL_L_X4Y119_SLICE_X4Y119_CQ),
.O5(CLBLM_R_X5Y120_SLICE_X7Y120_BO5),
.O6(CLBLM_R_X5Y120_SLICE_X7Y120_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaaf3f3aaaac0c0)
  ) CLBLM_R_X5Y120_SLICE_X7Y120_ALUT (
.I0(CLBLM_R_X7Y121_SLICE_X8Y121_BQ),
.I1(CLBLM_R_X11Y121_SLICE_X14Y121_CO6),
.I2(CLBLM_R_X5Y120_SLICE_X7Y120_AQ),
.I3(1'b1),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(CLBLM_L_X8Y115_SLICE_X10Y115_AQ),
.O5(CLBLM_R_X5Y120_SLICE_X7Y120_AO5),
.O6(CLBLM_R_X5Y120_SLICE_X7Y120_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y121_SLICE_X6Y121_A5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y123_SLICE_X6Y123_DO6),
.Q(CLBLM_R_X5Y121_SLICE_X6Y121_A5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y121_SLICE_X6Y121_B5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y121_SLICE_X6Y121_CO6),
.Q(CLBLM_R_X5Y121_SLICE_X6Y121_B5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y121_SLICE_X6Y121_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y121_SLICE_X6Y121_AO6),
.Q(CLBLM_R_X5Y121_SLICE_X6Y121_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y121_SLICE_X6Y121_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y121_SLICE_X6Y121_BO6),
.Q(CLBLM_R_X5Y121_SLICE_X6Y121_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffcceefffffcfe)
  ) CLBLM_R_X5Y121_SLICE_X6Y121_DLUT (
.I0(CLBLM_R_X5Y117_SLICE_X6Y117_AQ),
.I1(CLBLM_R_X5Y121_SLICE_X7Y121_CO6),
.I2(CLBLM_R_X5Y111_SLICE_X6Y111_AQ),
.I3(CLBLM_R_X3Y121_SLICE_X2Y121_AO6),
.I4(CLBLM_R_X5Y121_SLICE_X7Y121_BO6),
.I5(CLBLL_L_X4Y121_SLICE_X4Y121_CO6),
.O5(CLBLM_R_X5Y121_SLICE_X6Y121_DO5),
.O6(CLBLM_R_X5Y121_SLICE_X6Y121_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'haf0faa0088888888)
  ) CLBLM_R_X5Y121_SLICE_X6Y121_CLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_R_X11Y121_SLICE_X14Y121_AQ),
.I2(CLBLM_R_X3Y116_SLICE_X2Y116_CO6),
.I3(CLBLM_R_X5Y120_SLICE_X6Y120_AQ),
.I4(CLBLM_R_X5Y121_SLICE_X6Y121_B5Q),
.I5(1'b1),
.O5(CLBLM_R_X5Y121_SLICE_X6Y121_CO5),
.O6(CLBLM_R_X5Y121_SLICE_X6Y121_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaafcfcaaaa0c0c)
  ) CLBLM_R_X5Y121_SLICE_X6Y121_BLUT (
.I0(CLBLM_R_X7Y122_SLICE_X9Y122_A5Q),
.I1(CLBLM_R_X5Y121_SLICE_X6Y121_BQ),
.I2(CLBLM_R_X5Y115_SLICE_X6Y115_CO5),
.I3(1'b1),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(CLBLL_L_X4Y115_SLICE_X5Y115_BQ),
.O5(CLBLM_R_X5Y121_SLICE_X6Y121_BO5),
.O6(CLBLM_R_X5Y121_SLICE_X6Y121_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'haaf0aa00aafcaa00)
  ) CLBLM_R_X5Y121_SLICE_X6Y121_ALUT (
.I0(CLBLM_R_X5Y117_SLICE_X6Y117_AQ),
.I1(CLBLM_R_X7Y114_SLICE_X8Y114_BQ),
.I2(CLBLM_R_X5Y121_SLICE_X6Y121_AQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(RIOB33_X105Y105_IOB_X1Y105_I),
.I5(RIOB33_X105Y121_IOB_X1Y121_I),
.O5(CLBLM_R_X5Y121_SLICE_X6Y121_AO5),
.O6(CLBLM_R_X5Y121_SLICE_X6Y121_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y121_SLICE_X7Y121_A5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y121_SLICE_X7Y121_AO5),
.Q(CLBLM_R_X5Y121_SLICE_X7Y121_A5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y121_SLICE_X7Y121_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y121_SLICE_X7Y121_AO6),
.Q(CLBLM_R_X5Y121_SLICE_X7Y121_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h15ff15ff3fff3fff)
  ) CLBLM_R_X5Y121_SLICE_X7Y121_DLUT (
.I0(CLBLM_R_X5Y123_SLICE_X7Y123_AQ),
.I1(CLBLM_R_X7Y121_SLICE_X9Y121_BQ),
.I2(CLBLM_R_X7Y121_SLICE_X8Y121_AQ),
.I3(CLBLM_R_X5Y123_SLICE_X6Y123_CQ),
.I4(1'b1),
.I5(CLBLM_R_X5Y123_SLICE_X6Y123_BQ),
.O5(CLBLM_R_X5Y121_SLICE_X7Y121_DO5),
.O6(CLBLM_R_X5Y121_SLICE_X7Y121_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000200000000)
  ) CLBLM_R_X5Y121_SLICE_X7Y121_CLUT (
.I0(CLBLM_R_X5Y121_SLICE_X6Y121_AQ),
.I1(RIOB33_X105Y133_IOB_X1Y133_I),
.I2(RIOB33_X105Y133_IOB_X1Y134_I),
.I3(CLBLM_R_X3Y122_SLICE_X3Y122_AO6),
.I4(RIOB33_X105Y131_IOB_X1Y131_I),
.I5(RIOB33_X105Y131_IOB_X1Y132_I),
.O5(CLBLM_R_X5Y121_SLICE_X7Y121_CO5),
.O6(CLBLM_R_X5Y121_SLICE_X7Y121_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000040000)
  ) CLBLM_R_X5Y121_SLICE_X7Y121_BLUT (
.I0(RIOB33_X105Y131_IOB_X1Y131_I),
.I1(RIOB33_X105Y133_IOB_X1Y133_I),
.I2(RIOB33_X105Y133_IOB_X1Y134_I),
.I3(RIOB33_X105Y131_IOB_X1Y132_I),
.I4(CLBLM_L_X8Y118_SLICE_X10Y118_BQ),
.I5(CLBLM_R_X3Y122_SLICE_X3Y122_AO6),
.O5(CLBLM_R_X5Y121_SLICE_X7Y121_BO5),
.O6(CLBLM_R_X5Y121_SLICE_X7Y121_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'haa00aaf0f0ccf0cc)
  ) CLBLM_R_X5Y121_SLICE_X7Y121_ALUT (
.I0(CLBLM_R_X5Y122_SLICE_X7Y122_DQ),
.I1(CLBLM_R_X5Y123_SLICE_X6Y123_BQ),
.I2(CLBLM_R_X5Y121_SLICE_X7Y121_AQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(RIOB33_X105Y105_IOB_X1Y105_I),
.I5(1'b1),
.O5(CLBLM_R_X5Y121_SLICE_X7Y121_AO5),
.O6(CLBLM_R_X5Y121_SLICE_X7Y121_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y122_SLICE_X6Y122_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y122_SLICE_X6Y122_AO6),
.Q(CLBLM_R_X5Y122_SLICE_X6Y122_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y122_SLICE_X6Y122_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y122_SLICE_X6Y122_BO6),
.Q(CLBLM_R_X5Y122_SLICE_X6Y122_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000040400005504)
  ) CLBLM_R_X5Y122_SLICE_X6Y122_DLUT (
.I0(CLBLM_R_X3Y122_SLICE_X3Y122_AO6),
.I1(CLBLM_R_X7Y118_SLICE_X8Y118_AQ),
.I2(CLBLL_L_X4Y123_SLICE_X5Y123_AO6),
.I3(CLBLM_R_X11Y121_SLICE_X14Y121_AQ),
.I4(RIOB33_X105Y131_IOB_X1Y131_I),
.I5(CLBLM_R_X3Y124_SLICE_X2Y124_BO6),
.O5(CLBLM_R_X5Y122_SLICE_X6Y122_DO5),
.O6(CLBLM_R_X5Y122_SLICE_X6Y122_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h1010000015100500)
  ) CLBLM_R_X5Y122_SLICE_X6Y122_CLUT (
.I0(CLBLM_R_X3Y122_SLICE_X3Y122_AO6),
.I1(CLBLL_L_X4Y123_SLICE_X5Y123_AO6),
.I2(RIOB33_X105Y131_IOB_X1Y131_I),
.I3(CLBLM_R_X13Y119_SLICE_X18Y119_BQ),
.I4(CLBLM_R_X7Y123_SLICE_X8Y123_CQ),
.I5(CLBLM_R_X3Y124_SLICE_X2Y124_BO6),
.O5(CLBLM_R_X5Y122_SLICE_X6Y122_CO5),
.O6(CLBLM_R_X5Y122_SLICE_X6Y122_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf505f505f404f404)
  ) CLBLM_R_X5Y122_SLICE_X6Y122_BLUT (
.I0(CLBLM_R_X3Y116_SLICE_X2Y116_DO6),
.I1(CLBLM_R_X5Y122_SLICE_X6Y122_BQ),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLM_L_X8Y120_SLICE_X10Y120_D5Q),
.I4(1'b1),
.I5(CLBLM_R_X5Y125_SLICE_X6Y125_A5Q),
.O5(CLBLM_R_X5Y122_SLICE_X6Y122_BO5),
.O6(CLBLM_R_X5Y122_SLICE_X6Y122_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hccfc00f00000aaaa)
  ) CLBLM_R_X5Y122_SLICE_X6Y122_ALUT (
.I0(RIOB33_X105Y121_IOB_X1Y121_I),
.I1(CLBLM_L_X8Y121_SLICE_X11Y121_AQ),
.I2(CLBLM_R_X5Y122_SLICE_X6Y122_AQ),
.I3(CLBLM_R_X3Y116_SLICE_X2Y116_CO6),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(1'b1),
.O5(CLBLM_R_X5Y122_SLICE_X6Y122_AO5),
.O6(CLBLM_R_X5Y122_SLICE_X6Y122_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y122_SLICE_X7Y122_A5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y122_SLICE_X7Y122_AO5),
.Q(CLBLM_R_X5Y122_SLICE_X7Y122_A5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y122_SLICE_X7Y122_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y122_SLICE_X7Y122_AO6),
.Q(CLBLM_R_X5Y122_SLICE_X7Y122_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y122_SLICE_X7Y122_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y122_SLICE_X7Y122_BO6),
.Q(CLBLM_R_X5Y122_SLICE_X7Y122_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y122_SLICE_X7Y122_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y122_SLICE_X7Y122_CO6),
.Q(CLBLM_R_X5Y122_SLICE_X7Y122_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y122_SLICE_X7Y122_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y122_SLICE_X7Y122_DO6),
.Q(CLBLM_R_X5Y122_SLICE_X7Y122_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hd8ddd8ddd888d888)
  ) CLBLM_R_X5Y122_SLICE_X7Y122_DLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_L_X10Y126_SLICE_X12Y126_AQ),
.I2(CLBLM_R_X5Y122_SLICE_X7Y122_DQ),
.I3(CLBLM_R_X3Y116_SLICE_X2Y116_DO6),
.I4(1'b1),
.I5(CLBLM_R_X7Y120_SLICE_X9Y120_D5Q),
.O5(CLBLM_R_X5Y122_SLICE_X7Y122_DO5),
.O6(CLBLM_R_X5Y122_SLICE_X7Y122_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hafae0504afae0504)
  ) CLBLM_R_X5Y122_SLICE_X7Y122_CLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_R_X5Y122_SLICE_X7Y122_CQ),
.I2(CLBLM_R_X3Y116_SLICE_X2Y116_DO6),
.I3(CLBLM_R_X5Y122_SLICE_X7Y122_A5Q),
.I4(CLBLM_L_X10Y122_SLICE_X12Y122_BQ),
.I5(1'b1),
.O5(CLBLM_R_X5Y122_SLICE_X7Y122_CO5),
.O6(CLBLM_R_X5Y122_SLICE_X7Y122_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f00000f0f0eeee)
  ) CLBLM_R_X5Y122_SLICE_X7Y122_BLUT (
.I0(CLBLM_L_X8Y121_SLICE_X11Y121_DQ),
.I1(CLBLM_R_X5Y122_SLICE_X7Y122_BQ),
.I2(CLBLM_R_X5Y122_SLICE_X7Y122_AQ),
.I3(1'b1),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(CLBLM_R_X11Y121_SLICE_X14Y121_CO6),
.O5(CLBLM_R_X5Y122_SLICE_X7Y122_BO5),
.O6(CLBLM_R_X5Y122_SLICE_X7Y122_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfc0cfc0cfff00f00)
  ) CLBLM_R_X5Y122_SLICE_X7Y122_ALUT (
.I0(1'b1),
.I1(CLBLM_R_X3Y120_SLICE_X3Y120_BO6),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLM_L_X8Y120_SLICE_X10Y120_CQ),
.I4(CLBLL_L_X4Y119_SLICE_X4Y119_C5Q),
.I5(1'b1),
.O5(CLBLM_R_X5Y122_SLICE_X7Y122_AO5),
.O6(CLBLM_R_X5Y122_SLICE_X7Y122_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y123_SLICE_X6Y123_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y123_SLICE_X6Y123_AO6),
.Q(CLBLM_R_X5Y123_SLICE_X6Y123_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y123_SLICE_X6Y123_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y123_SLICE_X6Y123_BO6),
.Q(CLBLM_R_X5Y123_SLICE_X6Y123_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y123_SLICE_X6Y123_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y123_SLICE_X6Y123_CO6),
.Q(CLBLM_R_X5Y123_SLICE_X6Y123_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0fff00080808080)
  ) CLBLM_R_X5Y123_SLICE_X6Y123_DLUT (
.I0(CLBLM_R_X5Y123_SLICE_X7Y123_AQ),
.I1(CLBLM_R_X7Y121_SLICE_X8Y121_DO6),
.I2(CLBLM_R_X5Y123_SLICE_X6Y123_BQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(RIOB33_X105Y127_IOB_X1Y127_I),
.I5(1'b1),
.O5(CLBLM_R_X5Y123_SLICE_X6Y123_DO5),
.O6(CLBLM_R_X5Y123_SLICE_X6Y123_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hb3b3a0a0ececa0a0)
  ) CLBLM_R_X5Y123_SLICE_X6Y123_CLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_R_X5Y123_SLICE_X6Y123_CQ),
.I2(CLBLM_R_X3Y115_SLICE_X2Y115_BQ),
.I3(1'b1),
.I4(CLBLM_R_X7Y122_SLICE_X9Y122_BO6),
.I5(CLBLM_R_X5Y123_SLICE_X6Y123_DO5),
.O5(CLBLM_R_X5Y123_SLICE_X6Y123_CO5),
.O6(CLBLM_R_X5Y123_SLICE_X6Y123_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hdc50fcf0eca0cc00)
  ) CLBLM_R_X5Y123_SLICE_X6Y123_BLUT (
.I0(CLBLM_R_X7Y121_SLICE_X8Y121_DO6),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(CLBLM_R_X7Y122_SLICE_X9Y122_BO6),
.I3(CLBLL_L_X4Y115_SLICE_X5Y115_BQ),
.I4(CLBLM_R_X5Y123_SLICE_X7Y123_AQ),
.I5(CLBLM_R_X5Y123_SLICE_X6Y123_BQ),
.O5(CLBLM_R_X5Y123_SLICE_X6Y123_BO5),
.O6(CLBLM_R_X5Y123_SLICE_X6Y123_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hff48ffc04848c0c0)
  ) CLBLM_R_X5Y123_SLICE_X6Y123_ALUT (
.I0(CLBLM_R_X5Y125_SLICE_X6Y125_BO5),
.I1(CLBLM_R_X7Y124_SLICE_X8Y124_DO5),
.I2(CLBLM_R_X5Y123_SLICE_X6Y123_AQ),
.I3(CLBLM_R_X3Y117_SLICE_X3Y117_AQ),
.I4(CLBLL_L_X4Y123_SLICE_X4Y123_BQ),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLM_R_X5Y123_SLICE_X6Y123_AO5),
.O6(CLBLM_R_X5Y123_SLICE_X6Y123_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y123_SLICE_X7Y123_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y123_SLICE_X7Y123_AO6),
.Q(CLBLM_R_X5Y123_SLICE_X7Y123_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X5Y123_SLICE_X7Y123_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y123_SLICE_X7Y123_DO5),
.O6(CLBLM_R_X5Y123_SLICE_X7Y123_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X5Y123_SLICE_X7Y123_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y123_SLICE_X7Y123_CO5),
.O6(CLBLM_R_X5Y123_SLICE_X7Y123_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X5Y123_SLICE_X7Y123_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y123_SLICE_X7Y123_BO5),
.O6(CLBLM_R_X5Y123_SLICE_X7Y123_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hafaa0f00faaaf000)
  ) CLBLM_R_X5Y123_SLICE_X7Y123_ALUT (
.I0(CLBLM_R_X7Y123_SLICE_X8Y123_CQ),
.I1(1'b1),
.I2(CLBLM_R_X5Y123_SLICE_X7Y123_AQ),
.I3(CLBLM_R_X7Y122_SLICE_X9Y122_BO6),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(CLBLM_R_X7Y121_SLICE_X8Y121_DO6),
.O5(CLBLM_R_X5Y123_SLICE_X7Y123_AO5),
.O6(CLBLM_R_X5Y123_SLICE_X7Y123_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y124_SLICE_X6Y124_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y124_SLICE_X6Y124_AO6),
.Q(CLBLM_R_X5Y124_SLICE_X6Y124_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y124_SLICE_X6Y124_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y124_SLICE_X6Y124_BO6),
.Q(CLBLM_R_X5Y124_SLICE_X6Y124_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y124_SLICE_X6Y124_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y124_SLICE_X6Y124_CO6),
.Q(CLBLM_R_X5Y124_SLICE_X6Y124_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X5Y124_SLICE_X6Y124_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y124_SLICE_X6Y124_DO5),
.O6(CLBLM_R_X5Y124_SLICE_X6Y124_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hbefa1450fafa5050)
  ) CLBLM_R_X5Y124_SLICE_X6Y124_CLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLL_L_X4Y123_SLICE_X4Y123_BQ),
.I2(CLBLL_L_X4Y119_SLICE_X4Y119_C5Q),
.I3(CLBLM_R_X5Y125_SLICE_X6Y125_BO5),
.I4(CLBLM_R_X5Y116_SLICE_X6Y116_BQ),
.I5(CLBLM_R_X5Y123_SLICE_X6Y123_AQ),
.O5(CLBLM_R_X5Y124_SLICE_X6Y124_CO5),
.O6(CLBLM_R_X5Y124_SLICE_X6Y124_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaa030caaaa0000)
  ) CLBLM_R_X5Y124_SLICE_X6Y124_BLUT (
.I0(CLBLM_R_X5Y111_SLICE_X6Y111_AQ),
.I1(CLBLM_R_X5Y124_SLICE_X6Y124_BQ),
.I2(CLBLL_L_X4Y119_SLICE_X4Y119_C5Q),
.I3(CLBLM_R_X5Y125_SLICE_X6Y125_CO5),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(RIOB33_X105Y105_IOB_X1Y105_I),
.O5(CLBLM_R_X5Y124_SLICE_X6Y124_BO5),
.O6(CLBLM_R_X5Y124_SLICE_X6Y124_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hcccccccc05005000)
  ) CLBLM_R_X5Y124_SLICE_X6Y124_ALUT (
.I0(CLBLL_L_X4Y119_SLICE_X4Y119_C5Q),
.I1(CLBLM_L_X10Y122_SLICE_X13Y122_BQ),
.I2(CLBLM_R_X5Y124_SLICE_X6Y124_AQ),
.I3(RIOB33_X105Y105_IOB_X1Y105_I),
.I4(CLBLM_R_X5Y125_SLICE_X6Y125_DO6),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLM_R_X5Y124_SLICE_X6Y124_AO5),
.O6(CLBLM_R_X5Y124_SLICE_X6Y124_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X5Y124_SLICE_X7Y124_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y124_SLICE_X7Y124_DO5),
.O6(CLBLM_R_X5Y124_SLICE_X7Y124_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X5Y124_SLICE_X7Y124_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y124_SLICE_X7Y124_CO5),
.O6(CLBLM_R_X5Y124_SLICE_X7Y124_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X5Y124_SLICE_X7Y124_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y124_SLICE_X7Y124_BO5),
.O6(CLBLM_R_X5Y124_SLICE_X7Y124_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X5Y124_SLICE_X7Y124_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y124_SLICE_X7Y124_AO5),
.O6(CLBLM_R_X5Y124_SLICE_X7Y124_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y125_SLICE_X6Y125_A5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y125_SLICE_X6Y125_BO6),
.Q(CLBLM_R_X5Y125_SLICE_X6Y125_A5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y125_SLICE_X6Y125_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y125_SLICE_X6Y125_AO6),
.Q(CLBLM_R_X5Y125_SLICE_X6Y125_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h8000000000000000)
  ) CLBLM_R_X5Y125_SLICE_X6Y125_DLUT (
.I0(CLBLL_L_X4Y123_SLICE_X4Y123_AQ),
.I1(CLBLM_R_X5Y125_SLICE_X6Y125_AQ),
.I2(CLBLM_R_X7Y124_SLICE_X8Y124_A5Q),
.I3(CLBLM_R_X7Y124_SLICE_X8Y124_CQ),
.I4(CLBLM_R_X7Y124_SLICE_X8Y124_BQ),
.I5(CLBLM_R_X5Y124_SLICE_X6Y124_BQ),
.O5(CLBLM_R_X5Y125_SLICE_X6Y125_DO5),
.O6(CLBLM_R_X5Y125_SLICE_X6Y125_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h8000000088000000)
  ) CLBLM_R_X5Y125_SLICE_X6Y125_CLUT (
.I0(CLBLL_L_X4Y123_SLICE_X4Y123_AQ),
.I1(CLBLM_R_X7Y124_SLICE_X8Y124_A5Q),
.I2(CLBLM_R_X5Y124_SLICE_X6Y124_BQ),
.I3(CLBLM_R_X7Y124_SLICE_X8Y124_CQ),
.I4(CLBLM_R_X7Y124_SLICE_X8Y124_BQ),
.I5(1'b1),
.O5(CLBLM_R_X5Y125_SLICE_X6Y125_CO5),
.O6(CLBLM_R_X5Y125_SLICE_X6Y125_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf5a0f5a0c0c00000)
  ) CLBLM_R_X5Y125_SLICE_X6Y125_BLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_R_X5Y124_SLICE_X6Y124_AQ),
.I2(CLBLM_R_X5Y125_SLICE_X6Y125_AQ),
.I3(CLBLM_R_X5Y123_SLICE_X6Y123_CQ),
.I4(CLBLM_R_X5Y125_SLICE_X6Y125_CO6),
.I5(1'b1),
.O5(CLBLM_R_X5Y125_SLICE_X6Y125_BO5),
.O6(CLBLM_R_X5Y125_SLICE_X6Y125_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h888d888888d88888)
  ) CLBLM_R_X5Y125_SLICE_X6Y125_ALUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_L_X8Y119_SLICE_X10Y119_A5Q),
.I2(CLBLM_R_X5Y125_SLICE_X6Y125_AQ),
.I3(CLBLL_L_X4Y119_SLICE_X4Y119_C5Q),
.I4(RIOB33_X105Y105_IOB_X1Y105_I),
.I5(CLBLM_R_X5Y125_SLICE_X6Y125_CO6),
.O5(CLBLM_R_X5Y125_SLICE_X6Y125_AO5),
.O6(CLBLM_R_X5Y125_SLICE_X6Y125_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X5Y125_SLICE_X7Y125_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y125_SLICE_X7Y125_DO5),
.O6(CLBLM_R_X5Y125_SLICE_X7Y125_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X5Y125_SLICE_X7Y125_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y125_SLICE_X7Y125_CO5),
.O6(CLBLM_R_X5Y125_SLICE_X7Y125_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X5Y125_SLICE_X7Y125_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y125_SLICE_X7Y125_BO5),
.O6(CLBLM_R_X5Y125_SLICE_X7Y125_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X5Y125_SLICE_X7Y125_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y125_SLICE_X7Y125_AO5),
.O6(CLBLM_R_X5Y125_SLICE_X7Y125_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y109_SLICE_X8Y109_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y109_SLICE_X8Y109_AO6),
.Q(CLBLM_R_X7Y109_SLICE_X8Y109_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y109_SLICE_X8Y109_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y109_SLICE_X8Y109_BO6),
.Q(CLBLM_R_X7Y109_SLICE_X8Y109_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y109_SLICE_X8Y109_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y109_SLICE_X8Y109_CO6),
.Q(CLBLM_R_X7Y109_SLICE_X8Y109_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X7Y109_SLICE_X8Y109_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y109_SLICE_X8Y109_DO5),
.O6(CLBLM_R_X7Y109_SLICE_X8Y109_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaaaaaa0000cccc)
  ) CLBLM_R_X7Y109_SLICE_X8Y109_CLUT (
.I0(CLBLM_R_X5Y111_SLICE_X6Y111_C5Q),
.I1(CLBLM_R_X7Y109_SLICE_X8Y109_CQ),
.I2(1'b1),
.I3(1'b1),
.I4(RIOB33_X105Y105_IOB_X1Y105_I),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLM_R_X7Y109_SLICE_X8Y109_CO5),
.O6(CLBLM_R_X7Y109_SLICE_X8Y109_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'he2c0e2c0e2c0e2c0)
  ) CLBLM_R_X7Y109_SLICE_X8Y109_BLUT (
.I0(RIOB33_X105Y105_IOB_X1Y105_I),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(CLBLM_R_X5Y109_SLICE_X7Y109_AQ),
.I3(CLBLM_R_X5Y110_SLICE_X7Y110_CQ),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y109_SLICE_X8Y109_BO5),
.O6(CLBLM_R_X7Y109_SLICE_X8Y109_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'haa00aa00aa30aa30)
  ) CLBLM_R_X7Y109_SLICE_X8Y109_ALUT (
.I0(CLBLM_R_X7Y109_SLICE_X8Y109_CQ),
.I1(RIOB33_X105Y117_IOB_X1Y118_I),
.I2(CLBLM_R_X7Y109_SLICE_X8Y109_AQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(1'b1),
.I5(CLBLM_R_X3Y118_SLICE_X2Y118_AQ),
.O5(CLBLM_R_X7Y109_SLICE_X8Y109_AO5),
.O6(CLBLM_R_X7Y109_SLICE_X8Y109_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X7Y109_SLICE_X9Y109_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y109_SLICE_X9Y109_DO5),
.O6(CLBLM_R_X7Y109_SLICE_X9Y109_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X7Y109_SLICE_X9Y109_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y109_SLICE_X9Y109_CO5),
.O6(CLBLM_R_X7Y109_SLICE_X9Y109_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X7Y109_SLICE_X9Y109_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y109_SLICE_X9Y109_BO5),
.O6(CLBLM_R_X7Y109_SLICE_X9Y109_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X7Y109_SLICE_X9Y109_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y109_SLICE_X9Y109_AO5),
.O6(CLBLM_R_X7Y109_SLICE_X9Y109_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y110_SLICE_X8Y110_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y110_SLICE_X8Y110_AO6),
.Q(CLBLM_R_X7Y110_SLICE_X8Y110_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y110_SLICE_X8Y110_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y110_SLICE_X8Y110_BO6),
.Q(CLBLM_R_X7Y110_SLICE_X8Y110_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y110_SLICE_X8Y110_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y110_SLICE_X8Y110_CO6),
.Q(CLBLM_R_X7Y110_SLICE_X8Y110_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff800000000888)
  ) CLBLM_R_X7Y110_SLICE_X8Y110_DLUT (
.I0(CLBLM_L_X10Y112_SLICE_X13Y112_CQ),
.I1(CLBLM_R_X7Y110_SLICE_X8Y110_CQ),
.I2(CLBLL_L_X4Y110_SLICE_X5Y110_AQ),
.I3(CLBLM_L_X8Y110_SLICE_X10Y110_BQ),
.I4(CLBLM_R_X5Y111_SLICE_X7Y111_DO6),
.I5(1'b1),
.O5(CLBLM_R_X7Y110_SLICE_X8Y110_DO5),
.O6(CLBLM_R_X7Y110_SLICE_X8Y110_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'haa00aa00ea40ba10)
  ) CLBLM_R_X7Y110_SLICE_X8Y110_CLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_R_X7Y110_SLICE_X8Y110_CQ),
.I2(RIOB33_X105Y105_IOB_X1Y105_I),
.I3(CLBLM_L_X8Y113_SLICE_X11Y113_CQ),
.I4(CLBLM_R_X7Y110_SLICE_X8Y110_DO6),
.I5(CLBLM_L_X8Y118_SLICE_X10Y118_DQ),
.O5(CLBLM_R_X7Y110_SLICE_X8Y110_CO5),
.O6(CLBLM_R_X7Y110_SLICE_X8Y110_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf000f000fe0ef000)
  ) CLBLM_R_X7Y110_SLICE_X8Y110_BLUT (
.I0(CLBLM_R_X7Y111_SLICE_X8Y111_CQ),
.I1(CLBLM_R_X7Y110_SLICE_X8Y110_BQ),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLM_R_X7Y115_SLICE_X8Y115_BQ),
.I4(CLBLM_R_X3Y118_SLICE_X2Y118_AQ),
.I5(RIOB33_X105Y117_IOB_X1Y118_I),
.O5(CLBLM_R_X7Y110_SLICE_X8Y110_BO5),
.O6(CLBLM_R_X7Y110_SLICE_X8Y110_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffccd80000ccd8)
  ) CLBLM_R_X7Y110_SLICE_X8Y110_ALUT (
.I0(RIOB33_X105Y117_IOB_X1Y118_I),
.I1(CLBLM_R_X7Y110_SLICE_X8Y110_BQ),
.I2(CLBLM_R_X7Y110_SLICE_X8Y110_AQ),
.I3(CLBLM_R_X3Y118_SLICE_X2Y118_AQ),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(CLBLM_R_X7Y118_SLICE_X8Y118_CQ),
.O5(CLBLM_R_X7Y110_SLICE_X8Y110_AO5),
.O6(CLBLM_R_X7Y110_SLICE_X8Y110_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y110_SLICE_X9Y110_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y110_SLICE_X9Y110_AO6),
.Q(CLBLM_R_X7Y110_SLICE_X9Y110_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y110_SLICE_X9Y110_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y110_SLICE_X9Y110_BO6),
.Q(CLBLM_R_X7Y110_SLICE_X9Y110_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y110_SLICE_X9Y110_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y110_SLICE_X9Y110_CO6),
.Q(CLBLM_R_X7Y110_SLICE_X9Y110_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X7Y110_SLICE_X9Y110_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y110_SLICE_X9Y110_DO5),
.O6(CLBLM_R_X7Y110_SLICE_X9Y110_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hff00ffcc000000cc)
  ) CLBLM_R_X7Y110_SLICE_X9Y110_CLUT (
.I0(1'b1),
.I1(CLBLM_R_X7Y110_SLICE_X9Y110_CQ),
.I2(1'b1),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(RIOB33_X105Y105_IOB_X1Y105_I),
.I5(CLBLM_R_X7Y115_SLICE_X9Y115_BQ),
.O5(CLBLM_R_X7Y110_SLICE_X9Y110_CO5),
.O6(CLBLM_R_X7Y110_SLICE_X9Y110_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf5f5f4f405050404)
  ) CLBLM_R_X7Y110_SLICE_X9Y110_BLUT (
.I0(CLBLM_R_X5Y111_SLICE_X7Y111_DO6),
.I1(CLBLM_R_X7Y110_SLICE_X9Y110_BQ),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(1'b1),
.I4(CLBLM_L_X8Y117_SLICE_X10Y117_AQ),
.I5(CLBLM_R_X5Y116_SLICE_X7Y116_CQ),
.O5(CLBLM_R_X7Y110_SLICE_X9Y110_BO5),
.O6(CLBLM_R_X7Y110_SLICE_X9Y110_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfefefecc32323200)
  ) CLBLM_R_X7Y110_SLICE_X9Y110_ALUT (
.I0(CLBLM_L_X10Y112_SLICE_X12Y112_DQ),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(CLBLM_R_X7Y110_SLICE_X9Y110_AQ),
.I3(CLBLM_R_X3Y118_SLICE_X2Y118_AQ),
.I4(RIOB33_X105Y117_IOB_X1Y118_I),
.I5(CLBLM_R_X5Y113_SLICE_X7Y113_A5Q),
.O5(CLBLM_R_X7Y110_SLICE_X9Y110_AO5),
.O6(CLBLM_R_X7Y110_SLICE_X9Y110_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y111_SLICE_X8Y111_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y111_SLICE_X8Y111_AO6),
.Q(CLBLM_R_X7Y111_SLICE_X8Y111_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y111_SLICE_X8Y111_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y111_SLICE_X8Y111_BO6),
.Q(CLBLM_R_X7Y111_SLICE_X8Y111_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y111_SLICE_X8Y111_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y111_SLICE_X8Y111_CO6),
.Q(CLBLM_R_X7Y111_SLICE_X8Y111_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffffffffcfffc)
  ) CLBLM_R_X7Y111_SLICE_X8Y111_DLUT (
.I0(1'b1),
.I1(CLBLM_R_X7Y110_SLICE_X9Y110_CQ),
.I2(CLBLM_R_X7Y111_SLICE_X8Y111_BQ),
.I3(CLBLM_R_X5Y115_SLICE_X7Y115_A5Q),
.I4(1'b1),
.I5(CLBLM_R_X7Y111_SLICE_X8Y111_AQ),
.O5(CLBLM_R_X7Y111_SLICE_X8Y111_DO5),
.O6(CLBLM_R_X7Y111_SLICE_X8Y111_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hb1a0b1a0b1b1b1b1)
  ) CLBLM_R_X7Y111_SLICE_X8Y111_CLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_R_X7Y111_SLICE_X9Y111_CO6),
.I2(CLBLM_R_X7Y111_SLICE_X8Y111_BQ),
.I3(CLBLM_R_X7Y128_SLICE_X8Y128_AQ),
.I4(1'b1),
.I5(RIOB33_X105Y141_IOB_X1Y142_I),
.O5(CLBLM_R_X7Y111_SLICE_X8Y111_CO5),
.O6(CLBLM_R_X7Y111_SLICE_X8Y111_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'haaccaaccaa00aa00)
  ) CLBLM_R_X7Y111_SLICE_X8Y111_BLUT (
.I0(CLBLM_R_X3Y115_SLICE_X3Y115_DQ),
.I1(RIOB33_X105Y105_IOB_X1Y105_I),
.I2(1'b1),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(1'b1),
.I5(CLBLM_R_X7Y111_SLICE_X8Y111_BQ),
.O5(CLBLM_R_X7Y111_SLICE_X8Y111_BO5),
.O6(CLBLM_R_X7Y111_SLICE_X8Y111_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfccc3000fccc3000)
  ) CLBLM_R_X7Y111_SLICE_X8Y111_ALUT (
.I0(1'b1),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(CLBLM_R_X7Y111_SLICE_X8Y111_AQ),
.I3(RIOB33_X105Y105_IOB_X1Y105_I),
.I4(CLBLM_R_X5Y111_SLICE_X7Y111_AQ),
.I5(1'b1),
.O5(CLBLM_R_X7Y111_SLICE_X8Y111_AO5),
.O6(CLBLM_R_X7Y111_SLICE_X8Y111_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h5a785a785a785a78)
  ) CLBLM_R_X7Y111_SLICE_X9Y111_DLUT (
.I0(CLBLM_R_X7Y110_SLICE_X9Y110_AQ),
.I1(CLBLM_R_X5Y117_SLICE_X7Y117_DO6),
.I2(CLBLM_R_X5Y114_SLICE_X6Y114_AQ),
.I3(CLBLM_R_X3Y119_SLICE_X2Y119_AO6),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y111_SLICE_X9Y111_DO5),
.O6(CLBLM_R_X7Y111_SLICE_X9Y111_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h00330000003300ff)
  ) CLBLM_R_X7Y111_SLICE_X9Y111_CLUT (
.I0(1'b1),
.I1(CLBLL_L_X4Y119_SLICE_X4Y119_CQ),
.I2(1'b1),
.I3(CLBLM_R_X7Y111_SLICE_X8Y111_CQ),
.I4(CLBLM_R_X5Y111_SLICE_X7Y111_DO6),
.I5(CLBLM_R_X7Y111_SLICE_X9Y111_BO6),
.O5(CLBLM_R_X7Y111_SLICE_X9Y111_CO5),
.O6(CLBLM_R_X7Y111_SLICE_X9Y111_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hcccccc9c00a00000)
  ) CLBLM_R_X7Y111_SLICE_X9Y111_BLUT (
.I0(CLBLL_L_X4Y110_SLICE_X5Y110_AQ),
.I1(CLBLM_L_X8Y117_SLICE_X11Y117_BQ),
.I2(CLBLM_L_X10Y112_SLICE_X13Y112_CQ),
.I3(CLBLM_L_X8Y110_SLICE_X10Y110_BQ),
.I4(CLBLM_R_X7Y110_SLICE_X8Y110_CQ),
.I5(1'b1),
.O5(CLBLM_R_X7Y111_SLICE_X9Y111_BO5),
.O6(CLBLM_R_X7Y111_SLICE_X9Y111_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h00550055fffffefe)
  ) CLBLM_R_X7Y111_SLICE_X9Y111_ALUT (
.I0(CLBLM_R_X3Y119_SLICE_X2Y119_AO6),
.I1(CLBLL_L_X4Y120_SLICE_X4Y120_BO6),
.I2(CLBLL_L_X2Y120_SLICE_X1Y120_DO6),
.I3(CLBLM_R_X5Y117_SLICE_X7Y117_DO6),
.I4(CLBLL_L_X4Y120_SLICE_X4Y120_AO6),
.I5(1'b1),
.O5(CLBLM_R_X7Y111_SLICE_X9Y111_AO5),
.O6(CLBLM_R_X7Y111_SLICE_X9Y111_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y112_SLICE_X8Y112_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y112_SLICE_X8Y112_AO6),
.Q(CLBLM_R_X7Y112_SLICE_X8Y112_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y112_SLICE_X8Y112_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y112_SLICE_X8Y112_BO6),
.Q(CLBLM_R_X7Y112_SLICE_X8Y112_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y112_SLICE_X8Y112_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y112_SLICE_X8Y112_CO6),
.Q(CLBLM_R_X7Y112_SLICE_X8Y112_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'he200e000e000e000)
  ) CLBLM_R_X7Y112_SLICE_X8Y112_DLUT (
.I0(CLBLM_R_X7Y109_SLICE_X8Y109_AQ),
.I1(CLBLM_R_X5Y116_SLICE_X7Y116_CQ),
.I2(CLBLM_R_X7Y115_SLICE_X8Y115_DO6),
.I3(CLBLM_R_X5Y110_SLICE_X7Y110_AO5),
.I4(RIOB33_X105Y105_IOB_X1Y105_I),
.I5(CLBLL_L_X2Y120_SLICE_X0Y120_CO6),
.O5(CLBLM_R_X7Y112_SLICE_X8Y112_DO5),
.O6(CLBLM_R_X7Y112_SLICE_X8Y112_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff5ccc00005ccc)
  ) CLBLM_R_X7Y112_SLICE_X8Y112_CLUT (
.I0(CLBLM_R_X5Y111_SLICE_X7Y111_CO5),
.I1(CLBLM_R_X7Y112_SLICE_X8Y112_CQ),
.I2(CLBLM_R_X3Y118_SLICE_X2Y118_AQ),
.I3(RIOB33_X105Y117_IOB_X1Y118_I),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(CLBLL_L_X2Y112_SLICE_X1Y112_BQ),
.O5(CLBLM_R_X7Y112_SLICE_X8Y112_CO5),
.O6(CLBLM_R_X7Y112_SLICE_X8Y112_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hff00ff0001016868)
  ) CLBLM_R_X7Y112_SLICE_X8Y112_BLUT (
.I0(CLBLM_R_X7Y113_SLICE_X9Y113_DO6),
.I1(CLBLM_R_X7Y112_SLICE_X8Y112_BQ),
.I2(CLBLM_R_X7Y109_SLICE_X8Y109_BQ),
.I3(CLBLM_R_X5Y115_SLICE_X7Y115_A5Q),
.I4(RIOB33_X105Y105_IOB_X1Y105_I),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLM_R_X7Y112_SLICE_X8Y112_BO5),
.O6(CLBLM_R_X7Y112_SLICE_X8Y112_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff000022202220)
  ) CLBLM_R_X7Y112_SLICE_X8Y112_ALUT (
.I0(CLBLM_R_X3Y118_SLICE_X2Y118_AQ),
.I1(RIOB33_X105Y117_IOB_X1Y118_I),
.I2(CLBLM_R_X7Y112_SLICE_X8Y112_AQ),
.I3(CLBLM_R_X7Y112_SLICE_X9Y112_BQ),
.I4(CLBLM_R_X3Y112_SLICE_X3Y112_BQ),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLM_R_X7Y112_SLICE_X8Y112_AO5),
.O6(CLBLM_R_X7Y112_SLICE_X8Y112_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y112_SLICE_X9Y112_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y112_SLICE_X9Y112_AO6),
.Q(CLBLM_R_X7Y112_SLICE_X9Y112_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y112_SLICE_X9Y112_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y112_SLICE_X9Y112_BO6),
.Q(CLBLM_R_X7Y112_SLICE_X9Y112_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y112_SLICE_X9Y112_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y112_SLICE_X9Y112_CO6),
.Q(CLBLM_R_X7Y112_SLICE_X9Y112_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hccddccddccddffff)
  ) CLBLM_R_X7Y112_SLICE_X9Y112_DLUT (
.I0(CLBLM_R_X7Y109_SLICE_X8Y109_AQ),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(1'b1),
.I3(CLBLM_R_X5Y116_SLICE_X7Y116_CQ),
.I4(CLBLM_R_X3Y118_SLICE_X2Y118_AQ),
.I5(RIOB33_X105Y117_IOB_X1Y118_I),
.O5(CLBLM_R_X7Y112_SLICE_X9Y112_DO5),
.O6(CLBLM_R_X7Y112_SLICE_X9Y112_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hff0fff0c000f000c)
  ) CLBLM_R_X7Y112_SLICE_X9Y112_CLUT (
.I0(1'b1),
.I1(CLBLM_R_X7Y112_SLICE_X9Y112_CQ),
.I2(CLBLM_R_X5Y111_SLICE_X7Y111_DO6),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLM_L_X10Y115_SLICE_X12Y115_AQ),
.I5(CLBLM_R_X3Y115_SLICE_X3Y115_CQ),
.O5(CLBLM_R_X7Y112_SLICE_X9Y112_CO5),
.O6(CLBLM_R_X7Y112_SLICE_X9Y112_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hff00ff0022223333)
  ) CLBLM_R_X7Y112_SLICE_X9Y112_BLUT (
.I0(CLBLM_R_X7Y128_SLICE_X8Y128_AQ),
.I1(CLBLM_L_X8Y112_SLICE_X11Y112_CO6),
.I2(1'b1),
.I3(CLBLM_R_X5Y122_SLICE_X7Y122_BQ),
.I4(RIOB33_X105Y141_IOB_X1Y142_I),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLM_R_X7Y112_SLICE_X9Y112_BO5),
.O6(CLBLM_R_X7Y112_SLICE_X9Y112_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hccccccccfffa0050)
  ) CLBLM_R_X7Y112_SLICE_X9Y112_ALUT (
.I0(CLBLM_R_X3Y118_SLICE_X2Y118_AQ),
.I1(CLBLM_R_X7Y110_SLICE_X9Y110_BQ),
.I2(CLBLM_R_X7Y112_SLICE_X9Y112_AQ),
.I3(RIOB33_X105Y117_IOB_X1Y118_I),
.I4(CLBLM_R_X7Y112_SLICE_X8Y112_AQ),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLM_R_X7Y112_SLICE_X9Y112_AO5),
.O6(CLBLM_R_X7Y112_SLICE_X9Y112_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y113_SLICE_X8Y113_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y113_SLICE_X8Y113_AO6),
.Q(CLBLM_R_X7Y113_SLICE_X8Y113_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hfdff111100000000)
  ) CLBLM_R_X7Y113_SLICE_X8Y113_DLUT (
.I0(CLBLM_R_X7Y109_SLICE_X8Y109_AQ),
.I1(CLBLM_R_X5Y116_SLICE_X7Y116_CQ),
.I2(CLBLL_L_X4Y120_SLICE_X4Y120_AO6),
.I3(RIOB33_X105Y105_IOB_X1Y105_I),
.I4(CLBLM_R_X7Y113_SLICE_X8Y113_BO5),
.I5(CLBLM_R_X5Y110_SLICE_X7Y110_AO5),
.O5(CLBLM_R_X7Y113_SLICE_X8Y113_DO5),
.O6(CLBLM_R_X7Y113_SLICE_X8Y113_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h2022eeee00000000)
  ) CLBLM_R_X7Y113_SLICE_X8Y113_CLUT (
.I0(CLBLM_R_X7Y109_SLICE_X8Y109_AQ),
.I1(CLBLM_R_X5Y116_SLICE_X7Y116_CQ),
.I2(CLBLL_L_X2Y120_SLICE_X1Y120_DO6),
.I3(RIOB33_X105Y105_IOB_X1Y105_I),
.I4(CLBLM_R_X5Y112_SLICE_X6Y112_BO5),
.I5(CLBLM_R_X5Y110_SLICE_X7Y110_AO5),
.O5(CLBLM_R_X7Y113_SLICE_X8Y113_CO5),
.O6(CLBLM_R_X7Y113_SLICE_X8Y113_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaaa0a0dd88dd88)
  ) CLBLM_R_X7Y113_SLICE_X8Y113_BLUT (
.I0(RIOB33_X105Y121_IOB_X1Y121_I),
.I1(CLBLM_R_X7Y118_SLICE_X9Y118_CQ),
.I2(CLBLM_L_X8Y120_SLICE_X11Y120_CQ),
.I3(CLBLM_R_X7Y113_SLICE_X9Y113_BQ),
.I4(CLBLM_R_X7Y114_SLICE_X8Y114_AQ),
.I5(1'b1),
.O5(CLBLM_R_X7Y113_SLICE_X8Y113_BO5),
.O6(CLBLM_R_X7Y113_SLICE_X8Y113_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff000000660066)
  ) CLBLM_R_X7Y113_SLICE_X8Y113_ALUT (
.I0(CLBLM_R_X7Y113_SLICE_X8Y113_BO5),
.I1(CLBLM_R_X3Y115_SLICE_X3Y115_DQ),
.I2(1'b1),
.I3(RIOB33_X105Y105_IOB_X1Y105_I),
.I4(CLBLM_L_X8Y116_SLICE_X11Y116_A5Q),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLM_R_X7Y113_SLICE_X8Y113_AO5),
.O6(CLBLM_R_X7Y113_SLICE_X8Y113_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y113_SLICE_X9Y113_A5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y113_SLICE_X9Y113_AO5),
.Q(CLBLM_R_X7Y113_SLICE_X9Y113_A5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y113_SLICE_X9Y113_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y113_SLICE_X9Y113_AO6),
.Q(CLBLM_R_X7Y113_SLICE_X9Y113_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y113_SLICE_X9Y113_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y113_SLICE_X9Y113_BO6),
.Q(CLBLM_R_X7Y113_SLICE_X9Y113_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hff0000ffff0f00f0)
  ) CLBLM_R_X7Y113_SLICE_X9Y113_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(CLBLM_R_X7Y114_SLICE_X8Y114_CO6),
.I3(CLBLM_R_X11Y116_SLICE_X14Y116_DQ),
.I4(CLBLM_L_X8Y112_SLICE_X10Y112_DQ),
.I5(CLBLM_R_X7Y112_SLICE_X8Y112_BQ),
.O5(CLBLM_R_X7Y113_SLICE_X9Y113_DO5),
.O6(CLBLM_R_X7Y113_SLICE_X9Y113_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000f0a00000f3b3)
  ) CLBLM_R_X7Y113_SLICE_X9Y113_CLUT (
.I0(CLBLM_R_X5Y113_SLICE_X6Y113_AQ),
.I1(CLBLM_R_X5Y116_SLICE_X7Y116_CQ),
.I2(RIOB33_X105Y121_IOB_X1Y121_I),
.I3(CLBLM_R_X3Y116_SLICE_X3Y116_BQ),
.I4(CLBLM_R_X7Y112_SLICE_X9Y112_DO6),
.I5(CLBLM_R_X5Y111_SLICE_X7Y111_CO5),
.O5(CLBLM_R_X7Y113_SLICE_X9Y113_CO5),
.O6(CLBLM_R_X7Y113_SLICE_X9Y113_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf5f5f5fc0505050c)
  ) CLBLM_R_X7Y113_SLICE_X9Y113_BLUT (
.I0(CLBLM_R_X5Y113_SLICE_X6Y113_DO6),
.I1(CLBLM_R_X7Y113_SLICE_X9Y113_BQ),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLM_R_X3Y118_SLICE_X2Y118_AQ),
.I4(RIOB33_X105Y117_IOB_X1Y118_I),
.I5(CLBLM_R_X11Y117_SLICE_X14Y117_CQ),
.O5(CLBLM_R_X7Y113_SLICE_X9Y113_BO5),
.O6(CLBLM_R_X7Y113_SLICE_X9Y113_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hee44ee44a0a0f5f5)
  ) CLBLM_R_X7Y113_SLICE_X9Y113_ALUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLL_L_X2Y120_SLICE_X0Y120_CO6),
.I2(CLBLM_R_X11Y114_SLICE_X14Y114_BQ),
.I3(CLBLM_L_X8Y114_SLICE_X10Y114_AQ),
.I4(CLBLM_L_X10Y113_SLICE_X13Y113_BO6),
.I5(1'b1),
.O5(CLBLM_R_X7Y113_SLICE_X9Y113_AO5),
.O6(CLBLM_R_X7Y113_SLICE_X9Y113_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y114_SLICE_X8Y114_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y114_SLICE_X8Y114_AO6),
.Q(CLBLM_R_X7Y114_SLICE_X8Y114_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y114_SLICE_X8Y114_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y114_SLICE_X8Y114_BO6),
.Q(CLBLM_R_X7Y114_SLICE_X8Y114_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hfabafafa000c0000)
  ) CLBLM_R_X7Y114_SLICE_X8Y114_DLUT (
.I0(CLBLM_R_X3Y116_SLICE_X3Y116_BQ),
.I1(CLBLM_R_X7Y120_SLICE_X9Y120_CQ),
.I2(CLBLM_R_X7Y122_SLICE_X8Y122_DQ),
.I3(CLBLM_R_X5Y114_SLICE_X7Y114_BO5),
.I4(CLBLM_R_X5Y114_SLICE_X7Y114_AQ),
.I5(RIOB33_X105Y121_IOB_X1Y121_I),
.O5(CLBLM_R_X7Y114_SLICE_X8Y114_DO5),
.O6(CLBLM_R_X7Y114_SLICE_X8Y114_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffffffffffffe)
  ) CLBLM_R_X7Y114_SLICE_X8Y114_CLUT (
.I0(CLBLM_R_X3Y116_SLICE_X3Y116_BQ),
.I1(CLBLM_R_X7Y114_SLICE_X9Y114_AO6),
.I2(CLBLM_R_X7Y118_SLICE_X9Y118_CQ),
.I3(CLBLM_L_X8Y114_SLICE_X11Y114_DO6),
.I4(CLBLM_L_X8Y115_SLICE_X10Y115_CQ),
.I5(CLBLL_L_X4Y115_SLICE_X4Y115_C5Q),
.O5(CLBLM_R_X7Y114_SLICE_X8Y114_CO5),
.O6(CLBLM_R_X7Y114_SLICE_X8Y114_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f00000f0f80008)
  ) CLBLM_R_X7Y114_SLICE_X8Y114_BLUT (
.I0(CLBLM_L_X10Y115_SLICE_X12Y115_CQ),
.I1(CLBLM_R_X7Y112_SLICE_X8Y112_BQ),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(RIOB33_X105Y105_IOB_X1Y105_I),
.I4(CLBLM_R_X5Y109_SLICE_X6Y109_BQ),
.I5(CLBLM_R_X7Y114_SLICE_X8Y114_CO6),
.O5(CLBLM_R_X7Y114_SLICE_X8Y114_BO5),
.O6(CLBLM_R_X7Y114_SLICE_X8Y114_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff0000fac8fac8)
  ) CLBLM_R_X7Y114_SLICE_X8Y114_ALUT (
.I0(CLBLM_R_X7Y114_SLICE_X8Y114_DO6),
.I1(CLBLM_R_X3Y118_SLICE_X2Y118_AQ),
.I2(CLBLM_R_X7Y114_SLICE_X8Y114_AQ),
.I3(RIOB33_X105Y117_IOB_X1Y118_I),
.I4(CLBLM_L_X8Y120_SLICE_X10Y120_BQ),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLM_R_X7Y114_SLICE_X8Y114_AO5),
.O6(CLBLM_R_X7Y114_SLICE_X8Y114_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffffffefefefe)
  ) CLBLM_R_X7Y114_SLICE_X9Y114_DLUT (
.I0(CLBLM_R_X7Y120_SLICE_X8Y120_DQ),
.I1(CLBLM_R_X11Y116_SLICE_X14Y116_DQ),
.I2(CLBLM_L_X8Y114_SLICE_X10Y114_B5Q),
.I3(1'b1),
.I4(1'b1),
.I5(CLBLM_R_X5Y110_SLICE_X7Y110_CQ),
.O5(CLBLM_R_X7Y114_SLICE_X9Y114_DO5),
.O6(CLBLM_R_X7Y114_SLICE_X9Y114_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffffffefefefe)
  ) CLBLM_R_X7Y114_SLICE_X9Y114_CLUT (
.I0(CLBLM_L_X8Y114_SLICE_X10Y114_C5Q),
.I1(CLBLM_L_X8Y112_SLICE_X10Y112_DQ),
.I2(CLBLM_L_X8Y114_SLICE_X10Y114_BQ),
.I3(1'b1),
.I4(1'b1),
.I5(CLBLM_R_X7Y119_SLICE_X9Y119_CQ),
.O5(CLBLM_R_X7Y114_SLICE_X9Y114_CO5),
.O6(CLBLM_R_X7Y114_SLICE_X9Y114_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffffffefefefe)
  ) CLBLM_R_X7Y114_SLICE_X9Y114_BLUT (
.I0(CLBLM_R_X7Y115_SLICE_X8Y115_CQ),
.I1(CLBLL_L_X4Y114_SLICE_X5Y114_AQ),
.I2(CLBLM_R_X7Y109_SLICE_X8Y109_BQ),
.I3(1'b1),
.I4(1'b1),
.I5(CLBLM_L_X8Y114_SLICE_X11Y114_BQ),
.O5(CLBLM_R_X7Y114_SLICE_X9Y114_BO5),
.O6(CLBLM_R_X7Y114_SLICE_X9Y114_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffffffffffffe)
  ) CLBLM_R_X7Y114_SLICE_X9Y114_ALUT (
.I0(CLBLM_R_X7Y114_SLICE_X9Y114_DO6),
.I1(CLBLL_L_X4Y115_SLICE_X5Y115_CQ),
.I2(CLBLM_R_X5Y115_SLICE_X7Y115_BQ),
.I3(CLBLM_R_X7Y114_SLICE_X9Y114_BO6),
.I4(CLBLM_R_X5Y119_SLICE_X6Y119_BQ),
.I5(CLBLM_R_X7Y114_SLICE_X9Y114_CO6),
.O5(CLBLM_R_X7Y114_SLICE_X9Y114_AO5),
.O6(CLBLM_R_X7Y114_SLICE_X9Y114_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y115_SLICE_X8Y115_A5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y117_SLICE_X10Y117_DO6),
.Q(CLBLM_R_X7Y115_SLICE_X8Y115_A5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y115_SLICE_X8Y115_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y115_SLICE_X8Y115_AO6),
.Q(CLBLM_R_X7Y115_SLICE_X8Y115_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y115_SLICE_X8Y115_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y115_SLICE_X8Y115_BO6),
.Q(CLBLM_R_X7Y115_SLICE_X8Y115_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y115_SLICE_X8Y115_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y115_SLICE_X8Y115_CO6),
.Q(CLBLM_R_X7Y115_SLICE_X8Y115_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hccc0ccc0cccc8888)
  ) CLBLM_R_X7Y115_SLICE_X8Y115_DLUT (
.I0(CLBLM_L_X8Y114_SLICE_X10Y114_BQ),
.I1(RIOB33_X105Y121_IOB_X1Y121_I),
.I2(CLBLM_R_X5Y111_SLICE_X7Y111_BQ),
.I3(CLBLL_L_X4Y114_SLICE_X5Y114_AQ),
.I4(CLBLM_R_X5Y116_SLICE_X7Y116_A5Q),
.I5(1'b1),
.O5(CLBLM_R_X7Y115_SLICE_X8Y115_DO5),
.O6(CLBLM_R_X7Y115_SLICE_X8Y115_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hf5f5a0a0a0a0a0a0)
  ) CLBLM_R_X7Y115_SLICE_X8Y115_CLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(1'b1),
.I2(CLBLM_R_X7Y122_SLICE_X8Y122_BQ),
.I3(1'b1),
.I4(RIOB33_X105Y105_IOB_X1Y105_I),
.I5(CLBLL_L_X4Y115_SLICE_X4Y115_C5Q),
.O5(CLBLM_R_X7Y115_SLICE_X8Y115_CO5),
.O6(CLBLM_R_X7Y115_SLICE_X8Y115_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf1f10101f4f40404)
  ) CLBLM_R_X7Y115_SLICE_X8Y115_BLUT (
.I0(RIOB33_X105Y105_IOB_X1Y105_I),
.I1(CLBLM_R_X7Y113_SLICE_X8Y113_BO6),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(1'b1),
.I4(CLBLM_R_X7Y115_SLICE_X9Y115_AQ),
.I5(CLBLL_L_X4Y115_SLICE_X5Y115_BQ),
.O5(CLBLM_R_X7Y115_SLICE_X8Y115_BO5),
.O6(CLBLM_R_X7Y115_SLICE_X8Y115_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffcff30ffecff20)
  ) CLBLM_R_X7Y115_SLICE_X8Y115_ALUT (
.I0(CLBLM_R_X3Y118_SLICE_X2Y118_AQ),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(CLBLM_R_X7Y115_SLICE_X8Y115_AQ),
.I3(CLBLM_R_X5Y114_SLICE_X7Y114_CO6),
.I4(CLBLM_R_X5Y119_SLICE_X6Y119_BQ),
.I5(RIOB33_X105Y117_IOB_X1Y118_I),
.O5(CLBLM_R_X7Y115_SLICE_X8Y115_AO5),
.O6(CLBLM_R_X7Y115_SLICE_X8Y115_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y115_SLICE_X9Y115_B5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y115_SLICE_X9Y115_BO5),
.Q(CLBLM_R_X7Y115_SLICE_X9Y115_B5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "C5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y115_SLICE_X9Y115_C5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y115_SLICE_X9Y115_CO5),
.Q(CLBLM_R_X7Y115_SLICE_X9Y115_C5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y115_SLICE_X9Y115_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y115_SLICE_X9Y115_AO6),
.Q(CLBLM_R_X7Y115_SLICE_X9Y115_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y115_SLICE_X9Y115_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y115_SLICE_X9Y115_BO6),
.Q(CLBLM_R_X7Y115_SLICE_X9Y115_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y115_SLICE_X9Y115_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y115_SLICE_X9Y115_CO6),
.Q(CLBLM_R_X7Y115_SLICE_X9Y115_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y115_SLICE_X9Y115_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y115_SLICE_X9Y115_DO6),
.Q(CLBLM_R_X7Y115_SLICE_X9Y115_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h888d888d88888888)
  ) CLBLM_R_X7Y115_SLICE_X9Y115_DLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_L_X8Y123_SLICE_X11Y123_A5Q),
.I2(RIOB33_X105Y105_IOB_X1Y105_I),
.I3(CLBLM_R_X7Y114_SLICE_X8Y114_CO6),
.I4(1'b1),
.I5(CLBLM_R_X7Y112_SLICE_X8Y112_BQ),
.O5(CLBLM_R_X7Y115_SLICE_X9Y115_DO5),
.O6(CLBLM_R_X7Y115_SLICE_X9Y115_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hafafa0a0cfc0cfc0)
  ) CLBLM_R_X7Y115_SLICE_X9Y115_CLUT (
.I0(CLBLM_R_X7Y115_SLICE_X8Y115_AQ),
.I1(CLBLM_R_X7Y115_SLICE_X8Y115_A5Q),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLM_R_X3Y115_SLICE_X3Y115_CQ),
.I4(RIOB33_X105Y103_IOB_X1Y103_I),
.I5(1'b1),
.O5(CLBLM_R_X7Y115_SLICE_X9Y115_CO5),
.O6(CLBLM_R_X7Y115_SLICE_X9Y115_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfff00f00cacacaca)
  ) CLBLM_R_X7Y115_SLICE_X9Y115_BLUT (
.I0(CLBLM_R_X7Y117_SLICE_X8Y117_A5Q),
.I1(CLBLM_R_X3Y115_SLICE_X3Y115_BQ),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLM_R_X7Y115_SLICE_X8Y115_A5Q),
.I4(CLBLM_R_X5Y118_SLICE_X7Y118_AQ),
.I5(1'b1),
.O5(CLBLM_R_X7Y115_SLICE_X9Y115_BO5),
.O6(CLBLM_R_X7Y115_SLICE_X9Y115_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaa00fcaaaa00fc)
  ) CLBLM_R_X7Y115_SLICE_X9Y115_ALUT (
.I0(CLBLM_R_X7Y112_SLICE_X8Y112_AQ),
.I1(CLBLM_R_X7Y117_SLICE_X9Y117_BQ),
.I2(CLBLM_R_X7Y115_SLICE_X9Y115_AQ),
.I3(CLBLM_R_X5Y117_SLICE_X7Y117_CO6),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(1'b1),
.O5(CLBLM_R_X7Y115_SLICE_X9Y115_AO5),
.O6(CLBLM_R_X7Y115_SLICE_X9Y115_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y116_SLICE_X8Y116_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y116_SLICE_X8Y116_AO6),
.Q(CLBLM_R_X7Y116_SLICE_X8Y116_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y116_SLICE_X8Y116_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y116_SLICE_X8Y116_BO6),
.Q(CLBLM_R_X7Y116_SLICE_X8Y116_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y116_SLICE_X8Y116_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y116_SLICE_X8Y116_CO6),
.Q(CLBLM_R_X7Y116_SLICE_X8Y116_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hffaeffaeff04ff04)
  ) CLBLM_R_X7Y116_SLICE_X8Y116_DLUT (
.I0(CLBLM_R_X7Y109_SLICE_X8Y109_AQ),
.I1(CLBLL_L_X4Y120_SLICE_X4Y120_AO6),
.I2(RIOB33_X105Y105_IOB_X1Y105_I),
.I3(CLBLM_R_X5Y116_SLICE_X7Y116_CQ),
.I4(1'b1),
.I5(CLBLM_R_X7Y115_SLICE_X8Y115_DO5),
.O5(CLBLM_R_X7Y116_SLICE_X8Y116_DO5),
.O6(CLBLM_R_X7Y116_SLICE_X8Y116_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hff000000ff00eeee)
  ) CLBLM_R_X7Y116_SLICE_X8Y116_CLUT (
.I0(CLBLM_R_X11Y115_SLICE_X15Y115_CQ),
.I1(CLBLM_R_X7Y116_SLICE_X8Y116_CQ),
.I2(1'b1),
.I3(CLBLM_R_X5Y116_SLICE_X6Y116_A5Q),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(CLBLM_R_X5Y111_SLICE_X7Y111_DO6),
.O5(CLBLM_R_X7Y116_SLICE_X8Y116_CO5),
.O6(CLBLM_R_X7Y116_SLICE_X8Y116_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'ha0a0a3aca0a0a3ac)
  ) CLBLM_R_X7Y116_SLICE_X8Y116_BLUT (
.I0(CLBLM_L_X8Y120_SLICE_X10Y120_A5Q),
.I1(CLBLL_L_X4Y116_SLICE_X5Y116_DQ),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLM_R_X7Y115_SLICE_X8Y115_DO5),
.I4(RIOB33_X105Y105_IOB_X1Y105_I),
.I5(1'b1),
.O5(CLBLM_R_X7Y116_SLICE_X8Y116_BO5),
.O6(CLBLM_R_X7Y116_SLICE_X8Y116_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hcccc00facccc00fa)
  ) CLBLM_R_X7Y116_SLICE_X8Y116_ALUT (
.I0(CLBLM_R_X7Y117_SLICE_X8Y117_BQ),
.I1(CLBLM_L_X8Y116_SLICE_X11Y116_AQ),
.I2(CLBLM_R_X7Y116_SLICE_X8Y116_AQ),
.I3(CLBLM_R_X5Y117_SLICE_X7Y117_CO6),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(1'b1),
.O5(CLBLM_R_X7Y116_SLICE_X8Y116_AO5),
.O6(CLBLM_R_X7Y116_SLICE_X8Y116_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y116_SLICE_X9Y116_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y116_SLICE_X9Y116_AO6),
.Q(CLBLM_R_X7Y116_SLICE_X9Y116_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffeeffffffee)
  ) CLBLM_R_X7Y116_SLICE_X9Y116_DLUT (
.I0(CLBLM_R_X7Y115_SLICE_X9Y115_AQ),
.I1(CLBLM_R_X7Y117_SLICE_X9Y117_AQ),
.I2(1'b1),
.I3(CLBLM_R_X7Y116_SLICE_X8Y116_CQ),
.I4(CLBLM_R_X7Y116_SLICE_X9Y116_AQ),
.I5(1'b1),
.O5(CLBLM_R_X7Y116_SLICE_X9Y116_DO5),
.O6(CLBLM_R_X7Y116_SLICE_X9Y116_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'ha3f3a3f3a303a303)
  ) CLBLM_R_X7Y116_SLICE_X9Y116_CLUT (
.I0(CLBLM_R_X7Y116_SLICE_X8Y116_AQ),
.I1(CLBLM_L_X10Y114_SLICE_X13Y114_DQ),
.I2(CLBLL_L_X2Y114_SLICE_X1Y114_BO5),
.I3(CLBLM_L_X8Y116_SLICE_X11Y116_DQ),
.I4(1'b1),
.I5(CLBLM_R_X7Y116_SLICE_X9Y116_BO6),
.O5(CLBLM_R_X7Y116_SLICE_X9Y116_CO5),
.O6(CLBLM_R_X7Y116_SLICE_X9Y116_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000ffff0000ffef)
  ) CLBLM_R_X7Y116_SLICE_X9Y116_BLUT (
.I0(CLBLM_R_X7Y116_SLICE_X9Y116_DO6),
.I1(CLBLM_R_X7Y117_SLICE_X9Y117_BQ),
.I2(CLBLM_L_X8Y116_SLICE_X10Y116_BO6),
.I3(CLBLM_L_X8Y116_SLICE_X11Y116_BQ),
.I4(CLBLM_R_X7Y116_SLICE_X8Y116_AQ),
.I5(CLBLM_R_X7Y117_SLICE_X8Y117_BQ),
.O5(CLBLM_R_X7Y116_SLICE_X9Y116_BO5),
.O6(CLBLM_R_X7Y116_SLICE_X9Y116_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hf202f202f303f303)
  ) CLBLM_R_X7Y116_SLICE_X9Y116_ALUT (
.I0(CLBLM_R_X7Y116_SLICE_X9Y116_AQ),
.I1(CLBLM_R_X5Y119_SLICE_X7Y119_AO6),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLM_R_X7Y119_SLICE_X8Y119_AQ),
.I4(1'b1),
.I5(CLBLM_R_X7Y116_SLICE_X9Y116_CO6),
.O5(CLBLM_R_X7Y116_SLICE_X9Y116_AO5),
.O6(CLBLM_R_X7Y116_SLICE_X9Y116_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y117_SLICE_X8Y117_A5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y117_SLICE_X8Y117_DO6),
.Q(CLBLM_R_X7Y117_SLICE_X8Y117_A5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y117_SLICE_X8Y117_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y117_SLICE_X8Y117_AO6),
.Q(CLBLM_R_X7Y117_SLICE_X8Y117_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y117_SLICE_X8Y117_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y117_SLICE_X8Y117_BO6),
.Q(CLBLM_R_X7Y117_SLICE_X8Y117_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y117_SLICE_X8Y117_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y117_SLICE_X8Y117_CO6),
.Q(CLBLM_R_X7Y117_SLICE_X8Y117_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hfe54aa00fcfc0000)
  ) CLBLM_R_X7Y117_SLICE_X8Y117_DLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_L_X8Y115_SLICE_X10Y115_CQ),
.I2(CLBLM_R_X7Y117_SLICE_X8Y117_AQ),
.I3(CLBLM_L_X8Y118_SLICE_X10Y118_D5Q),
.I4(RIOB33_X105Y121_IOB_X1Y121_I),
.I5(1'b1),
.O5(CLBLM_R_X7Y117_SLICE_X8Y117_DO5),
.O6(CLBLM_R_X7Y117_SLICE_X8Y117_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaaaffa00000550)
  ) CLBLM_R_X7Y117_SLICE_X8Y117_CLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(1'b1),
.I2(CLBLL_L_X2Y113_SLICE_X1Y113_BQ),
.I3(CLBLM_R_X7Y114_SLICE_X8Y114_DO6),
.I4(RIOB33_X105Y105_IOB_X1Y105_I),
.I5(CLBLM_L_X8Y119_SLICE_X11Y119_AQ),
.O5(CLBLM_R_X7Y117_SLICE_X8Y117_CO5),
.O6(CLBLM_R_X7Y117_SLICE_X8Y117_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'haa0faa0caa0faa0c)
  ) CLBLM_R_X7Y117_SLICE_X8Y117_BLUT (
.I0(CLBLM_R_X5Y117_SLICE_X6Y117_DQ),
.I1(CLBLM_R_X7Y117_SLICE_X8Y117_BQ),
.I2(CLBLM_R_X5Y117_SLICE_X7Y117_CO6),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLM_R_X7Y115_SLICE_X9Y115_AQ),
.I5(1'b1),
.O5(CLBLM_R_X7Y117_SLICE_X8Y117_BO5),
.O6(CLBLM_R_X7Y117_SLICE_X8Y117_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffcecccccfcec)
  ) CLBLM_R_X7Y117_SLICE_X8Y117_ALUT (
.I0(CLBLM_R_X3Y118_SLICE_X2Y118_AQ),
.I1(CLBLM_R_X5Y112_SLICE_X7Y112_BO6),
.I2(CLBLM_R_X7Y117_SLICE_X8Y117_AQ),
.I3(RIOB33_X105Y117_IOB_X1Y118_I),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(CLBLL_L_X4Y117_SLICE_X5Y117_BQ),
.O5(CLBLM_R_X7Y117_SLICE_X8Y117_AO5),
.O6(CLBLM_R_X7Y117_SLICE_X8Y117_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y117_SLICE_X9Y117_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y117_SLICE_X9Y117_AO6),
.Q(CLBLM_R_X7Y117_SLICE_X9Y117_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y117_SLICE_X9Y117_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y117_SLICE_X9Y117_BO6),
.Q(CLBLM_R_X7Y117_SLICE_X9Y117_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y117_SLICE_X9Y117_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y117_SLICE_X9Y117_CO6),
.Q(CLBLM_R_X7Y117_SLICE_X9Y117_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y117_SLICE_X9Y117_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y117_SLICE_X9Y117_DO6),
.Q(CLBLM_R_X7Y117_SLICE_X9Y117_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hfefedcdc32321010)
  ) CLBLM_R_X7Y117_SLICE_X9Y117_DLUT (
.I0(CLBLM_R_X5Y115_SLICE_X6Y115_CO5),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(CLBLM_R_X7Y117_SLICE_X9Y117_DQ),
.I3(1'b1),
.I4(CLBLL_L_X2Y113_SLICE_X1Y113_BQ),
.I5(CLBLM_L_X8Y115_SLICE_X11Y115_AQ),
.O5(CLBLM_R_X7Y117_SLICE_X9Y117_DO5),
.O6(CLBLM_R_X7Y117_SLICE_X9Y117_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hff000e0eff00eeee)
  ) CLBLM_R_X7Y117_SLICE_X9Y117_CLUT (
.I0(CLBLM_R_X3Y115_SLICE_X2Y115_BQ),
.I1(CLBLM_R_X7Y117_SLICE_X9Y117_CQ),
.I2(CLBLM_L_X8Y112_SLICE_X10Y112_CQ),
.I3(CLBLM_R_X11Y117_SLICE_X15Y117_AQ),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(CLBLL_L_X2Y112_SLICE_X1Y112_BQ),
.O5(CLBLM_R_X7Y117_SLICE_X9Y117_CO5),
.O6(CLBLM_R_X7Y117_SLICE_X9Y117_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaa0000aaaafcfc)
  ) CLBLM_R_X7Y117_SLICE_X9Y117_BLUT (
.I0(CLBLM_R_X5Y121_SLICE_X7Y121_A5Q),
.I1(CLBLM_R_X7Y117_SLICE_X9Y117_BQ),
.I2(CLBLM_R_X7Y117_SLICE_X9Y117_AQ),
.I3(1'b1),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(CLBLM_R_X5Y117_SLICE_X7Y117_CO6),
.O5(CLBLM_R_X7Y117_SLICE_X9Y117_BO5),
.O6(CLBLM_R_X7Y117_SLICE_X9Y117_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff555000005550)
  ) CLBLM_R_X7Y117_SLICE_X9Y117_ALUT (
.I0(CLBLM_R_X5Y117_SLICE_X7Y117_CO6),
.I1(1'b1),
.I2(CLBLM_R_X7Y117_SLICE_X9Y117_AQ),
.I3(CLBLM_R_X7Y116_SLICE_X8Y116_CQ),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(CLBLM_L_X10Y122_SLICE_X13Y122_A5Q),
.O5(CLBLM_R_X7Y117_SLICE_X9Y117_AO5),
.O6(CLBLM_R_X7Y117_SLICE_X9Y117_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y118_SLICE_X8Y118_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y118_SLICE_X8Y118_AO6),
.Q(CLBLM_R_X7Y118_SLICE_X8Y118_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y118_SLICE_X8Y118_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y118_SLICE_X8Y118_BO6),
.Q(CLBLM_R_X7Y118_SLICE_X8Y118_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y118_SLICE_X8Y118_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y118_SLICE_X8Y118_CO6),
.Q(CLBLM_R_X7Y118_SLICE_X8Y118_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y118_SLICE_X8Y118_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y118_SLICE_X8Y118_DO6),
.Q(CLBLM_R_X7Y118_SLICE_X8Y118_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hffaafafaffaaeaea)
  ) CLBLM_R_X7Y118_SLICE_X8Y118_DLUT (
.I0(CLBLM_R_X7Y113_SLICE_X8Y113_CO6),
.I1(RIOB33_X105Y117_IOB_X1Y118_I),
.I2(CLBLM_R_X7Y118_SLICE_X8Y118_DQ),
.I3(CLBLM_R_X5Y117_SLICE_X6Y117_D5Q),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(CLBLM_R_X3Y118_SLICE_X2Y118_AQ),
.O5(CLBLM_R_X7Y118_SLICE_X8Y118_DO5),
.O6(CLBLM_R_X7Y118_SLICE_X8Y118_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hff540054ff540054)
  ) CLBLM_R_X7Y118_SLICE_X8Y118_CLUT (
.I0(CLBLM_R_X5Y115_SLICE_X6Y115_CO5),
.I1(CLBLM_R_X7Y118_SLICE_X8Y118_CQ),
.I2(CLBLM_R_X5Y116_SLICE_X6Y116_DQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLM_L_X8Y116_SLICE_X10Y116_AQ),
.I5(1'b1),
.O5(CLBLM_R_X7Y118_SLICE_X8Y118_CO5),
.O6(CLBLM_R_X7Y118_SLICE_X8Y118_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hacacafafacaca0a0)
  ) CLBLM_R_X7Y118_SLICE_X8Y118_BLUT (
.I0(CLBLM_R_X5Y116_SLICE_X6Y116_DQ),
.I1(CLBLM_R_X7Y118_SLICE_X8Y118_BQ),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(1'b1),
.I4(CLBLM_R_X5Y115_SLICE_X6Y115_CO5),
.I5(CLBLM_R_X7Y119_SLICE_X9Y119_AQ),
.O5(CLBLM_R_X7Y118_SLICE_X8Y118_BO5),
.O6(CLBLM_R_X7Y118_SLICE_X8Y118_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hcccc0000ccccfff0)
  ) CLBLM_R_X7Y118_SLICE_X8Y118_ALUT (
.I0(1'b1),
.I1(CLBLL_L_X4Y114_SLICE_X4Y114_BQ),
.I2(CLBLM_R_X7Y118_SLICE_X8Y118_AQ),
.I3(CLBLM_L_X8Y119_SLICE_X11Y119_BQ),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(CLBLM_R_X11Y121_SLICE_X14Y121_CO6),
.O5(CLBLM_R_X7Y118_SLICE_X8Y118_AO5),
.O6(CLBLM_R_X7Y118_SLICE_X8Y118_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y118_SLICE_X9Y118_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y118_SLICE_X9Y118_AO6),
.Q(CLBLM_R_X7Y118_SLICE_X9Y118_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y118_SLICE_X9Y118_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y118_SLICE_X9Y118_BO6),
.Q(CLBLM_R_X7Y118_SLICE_X9Y118_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y118_SLICE_X9Y118_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y118_SLICE_X9Y118_CO6),
.Q(CLBLM_R_X7Y118_SLICE_X9Y118_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000100000000)
  ) CLBLM_R_X7Y118_SLICE_X9Y118_DLUT (
.I0(CLBLM_R_X7Y116_SLICE_X9Y116_BO6),
.I1(CLBLL_L_X4Y120_SLICE_X4Y120_BO6),
.I2(CLBLL_L_X4Y121_SLICE_X4Y121_CO6),
.I3(CLBLM_L_X10Y118_SLICE_X13Y118_DO6),
.I4(CLBLM_L_X8Y116_SLICE_X11Y116_DQ),
.I5(CLBLM_R_X5Y110_SLICE_X7Y110_DO5),
.O5(CLBLM_R_X7Y118_SLICE_X9Y118_DO5),
.O6(CLBLM_R_X7Y118_SLICE_X9Y118_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hff00ff00c0c0c0c0)
  ) CLBLM_R_X7Y118_SLICE_X9Y118_CLUT (
.I0(1'b1),
.I1(CLBLM_L_X8Y114_SLICE_X11Y114_BQ),
.I2(RIOB33_X105Y105_IOB_X1Y105_I),
.I3(CLBLM_R_X7Y118_SLICE_X9Y118_BQ),
.I4(1'b1),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLM_R_X7Y118_SLICE_X9Y118_CO5),
.O6(CLBLM_R_X7Y118_SLICE_X9Y118_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hffeecceeffcccccc)
  ) CLBLM_R_X7Y118_SLICE_X9Y118_BLUT (
.I0(RIOB33_X105Y105_IOB_X1Y105_I),
.I1(CLBLM_L_X10Y118_SLICE_X12Y118_CO6),
.I2(1'b1),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLM_R_X7Y117_SLICE_X9Y117_AQ),
.I5(CLBLM_R_X7Y118_SLICE_X9Y118_BQ),
.O5(CLBLM_R_X7Y118_SLICE_X9Y118_BO5),
.O6(CLBLM_R_X7Y118_SLICE_X9Y118_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfb0bf101fb0bfb0b)
  ) CLBLM_R_X7Y118_SLICE_X9Y118_ALUT (
.I0(RIOB33_X105Y105_IOB_X1Y105_I),
.I1(CLBLM_R_X7Y113_SLICE_X9Y113_A5Q),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLM_L_X10Y127_SLICE_X12Y127_AQ),
.I4(CLBLM_R_X7Y115_SLICE_X9Y115_C5Q),
.I5(CLBLM_R_X3Y115_SLICE_X3Y115_CQ),
.O5(CLBLM_R_X7Y118_SLICE_X9Y118_AO5),
.O6(CLBLM_R_X7Y118_SLICE_X9Y118_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y119_SLICE_X8Y119_C5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y119_SLICE_X8Y119_CO5),
.Q(CLBLM_R_X7Y119_SLICE_X8Y119_C5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y119_SLICE_X8Y119_D5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y119_SLICE_X8Y119_DO5),
.Q(CLBLM_R_X7Y119_SLICE_X8Y119_D5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y119_SLICE_X8Y119_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y119_SLICE_X8Y119_AO6),
.Q(CLBLM_R_X7Y119_SLICE_X8Y119_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y119_SLICE_X8Y119_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y119_SLICE_X8Y119_BO6),
.Q(CLBLM_R_X7Y119_SLICE_X8Y119_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y119_SLICE_X8Y119_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y119_SLICE_X8Y119_CO6),
.Q(CLBLM_R_X7Y119_SLICE_X8Y119_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y119_SLICE_X8Y119_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y119_SLICE_X8Y119_DO6),
.Q(CLBLM_R_X7Y119_SLICE_X8Y119_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hdc10dc10f3f3c0c0)
  ) CLBLM_R_X7Y119_SLICE_X8Y119_DLUT (
.I0(RIOB33_X105Y105_IOB_X1Y105_I),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(CLBLM_R_X7Y119_SLICE_X8Y119_DQ),
.I3(CLBLM_R_X11Y122_SLICE_X14Y122_AQ),
.I4(CLBLM_R_X7Y118_SLICE_X9Y118_AQ),
.I5(1'b1),
.O5(CLBLM_R_X7Y119_SLICE_X8Y119_DO5),
.O6(CLBLM_R_X7Y119_SLICE_X8Y119_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'haa00ee44d8d8d8d8)
  ) CLBLM_R_X7Y119_SLICE_X8Y119_CLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_R_X7Y119_SLICE_X8Y119_CQ),
.I2(CLBLL_L_X4Y120_SLICE_X4Y120_AO6),
.I3(CLBLM_L_X8Y119_SLICE_X11Y119_BQ),
.I4(RIOB33_X105Y105_IOB_X1Y105_I),
.I5(1'b1),
.O5(CLBLM_R_X7Y119_SLICE_X8Y119_CO5),
.O6(CLBLM_R_X7Y119_SLICE_X8Y119_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf1f4f1f401040104)
  ) CLBLM_R_X7Y119_SLICE_X8Y119_BLUT (
.I0(RIOB33_X105Y105_IOB_X1Y105_I),
.I1(CLBLM_R_X7Y117_SLICE_X8Y117_DO5),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLM_R_X7Y119_SLICE_X9Y119_BQ),
.I4(1'b1),
.I5(CLBLM_L_X10Y122_SLICE_X12Y122_AQ),
.O5(CLBLM_R_X7Y119_SLICE_X8Y119_BO5),
.O6(CLBLM_R_X7Y119_SLICE_X8Y119_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffc00fcff300030)
  ) CLBLM_R_X7Y119_SLICE_X8Y119_ALUT (
.I0(1'b1),
.I1(CLBLM_R_X11Y121_SLICE_X14Y121_CO6),
.I2(CLBLM_R_X7Y119_SLICE_X8Y119_AQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLM_R_X7Y120_SLICE_X8Y120_AQ),
.I5(CLBLM_L_X10Y118_SLICE_X13Y118_CQ),
.O5(CLBLM_R_X7Y119_SLICE_X8Y119_AO5),
.O6(CLBLM_R_X7Y119_SLICE_X8Y119_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y119_SLICE_X9Y119_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y119_SLICE_X9Y119_AO6),
.Q(CLBLM_R_X7Y119_SLICE_X9Y119_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y119_SLICE_X9Y119_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y119_SLICE_X9Y119_BO6),
.Q(CLBLM_R_X7Y119_SLICE_X9Y119_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y119_SLICE_X9Y119_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y119_SLICE_X9Y119_CO6),
.Q(CLBLM_R_X7Y119_SLICE_X9Y119_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h000055ff0000fcfc)
  ) CLBLM_R_X7Y119_SLICE_X9Y119_DLUT (
.I0(CLBLM_R_X3Y115_SLICE_X2Y115_BQ),
.I1(CLBLM_R_X7Y118_SLICE_X8Y118_DQ),
.I2(CLBLM_R_X5Y110_SLICE_X7Y110_AQ),
.I3(CLBLL_L_X2Y120_SLICE_X0Y120_CO6),
.I4(CLBLM_R_X3Y117_SLICE_X3Y117_BQ),
.I5(1'b1),
.O5(CLBLM_R_X7Y119_SLICE_X9Y119_DO5),
.O6(CLBLM_R_X7Y119_SLICE_X9Y119_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hcececece02020202)
  ) CLBLM_R_X7Y119_SLICE_X9Y119_CLUT (
.I0(CLBLM_L_X8Y114_SLICE_X10Y114_C5Q),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(RIOB33_X105Y105_IOB_X1Y105_I),
.I3(1'b1),
.I4(1'b1),
.I5(CLBLM_R_X5Y120_SLICE_X7Y120_CQ),
.O5(CLBLM_R_X7Y119_SLICE_X9Y119_CO5),
.O6(CLBLM_R_X7Y119_SLICE_X9Y119_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf1f40104f1f40104)
  ) CLBLM_R_X7Y119_SLICE_X9Y119_BLUT (
.I0(RIOB33_X105Y105_IOB_X1Y105_I),
.I1(CLBLM_L_X10Y118_SLICE_X13Y118_CQ),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLM_L_X8Y117_SLICE_X10Y117_DO5),
.I4(CLBLM_R_X5Y119_SLICE_X6Y119_AQ),
.I5(1'b1),
.O5(CLBLM_R_X7Y119_SLICE_X9Y119_BO5),
.O6(CLBLM_R_X7Y119_SLICE_X9Y119_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hcc55cc55cc00cc00)
  ) CLBLM_R_X7Y119_SLICE_X9Y119_ALUT (
.I0(RIOB33_X105Y105_IOB_X1Y105_I),
.I1(CLBLM_L_X10Y118_SLICE_X13Y118_CQ),
.I2(1'b1),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(1'b1),
.I5(CLBLM_L_X8Y120_SLICE_X10Y120_BQ),
.O5(CLBLM_R_X7Y119_SLICE_X9Y119_AO5),
.O6(CLBLM_R_X7Y119_SLICE_X9Y119_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y120_SLICE_X8Y120_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y120_SLICE_X8Y120_AO6),
.Q(CLBLM_R_X7Y120_SLICE_X8Y120_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y120_SLICE_X8Y120_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y120_SLICE_X8Y120_BO6),
.Q(CLBLM_R_X7Y120_SLICE_X8Y120_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y120_SLICE_X8Y120_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y120_SLICE_X8Y120_CO6),
.Q(CLBLM_R_X7Y120_SLICE_X8Y120_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y120_SLICE_X8Y120_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y120_SLICE_X8Y120_DO6),
.Q(CLBLM_R_X7Y120_SLICE_X8Y120_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaafafa00005050)
  ) CLBLM_R_X7Y120_SLICE_X8Y120_DLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(1'b1),
.I2(CLBLM_L_X8Y120_SLICE_X11Y120_CQ),
.I3(1'b1),
.I4(RIOB33_X105Y105_IOB_X1Y105_I),
.I5(CLBLM_R_X7Y123_SLICE_X9Y123_AQ),
.O5(CLBLM_R_X7Y120_SLICE_X8Y120_DO5),
.O6(CLBLM_R_X7Y120_SLICE_X8Y120_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'haaeeaaee00cc00cc)
  ) CLBLM_R_X7Y120_SLICE_X8Y120_CLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_R_X7Y120_SLICE_X8Y120_CQ),
.I2(1'b1),
.I3(CLBLM_R_X3Y116_SLICE_X2Y116_CO6),
.I4(1'b1),
.I5(CLBLM_R_X7Y120_SLICE_X9Y120_BQ),
.O5(CLBLM_R_X7Y120_SLICE_X8Y120_CO5),
.O6(CLBLM_R_X7Y120_SLICE_X8Y120_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffc0c0000fc0c)
  ) CLBLM_R_X7Y120_SLICE_X8Y120_BLUT (
.I0(1'b1),
.I1(CLBLM_R_X7Y120_SLICE_X8Y120_BQ),
.I2(CLBLM_R_X5Y115_SLICE_X6Y115_CO5),
.I3(CLBLM_L_X8Y120_SLICE_X10Y120_BQ),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(CLBLM_L_X8Y117_SLICE_X10Y117_CQ),
.O5(CLBLM_R_X7Y120_SLICE_X8Y120_BO5),
.O6(CLBLM_R_X7Y120_SLICE_X8Y120_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f00000fafb0a0b)
  ) CLBLM_R_X7Y120_SLICE_X8Y120_ALUT (
.I0(CLBLM_R_X5Y120_SLICE_X6Y120_A5Q),
.I1(CLBLM_R_X7Y124_SLICE_X8Y124_AQ),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLM_R_X7Y120_SLICE_X9Y120_A5Q),
.I4(CLBLM_R_X3Y110_SLICE_X2Y110_AQ),
.I5(CLBLM_L_X10Y124_SLICE_X12Y124_AQ),
.O5(CLBLM_R_X7Y120_SLICE_X8Y120_AO5),
.O6(CLBLM_R_X7Y120_SLICE_X8Y120_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y120_SLICE_X9Y120_A5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y120_SLICE_X9Y120_AO5),
.Q(CLBLM_R_X7Y120_SLICE_X9Y120_A5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y120_SLICE_X9Y120_D5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y120_SLICE_X9Y120_DO5),
.Q(CLBLM_R_X7Y120_SLICE_X9Y120_D5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y120_SLICE_X9Y120_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y120_SLICE_X9Y120_AO6),
.Q(CLBLM_R_X7Y120_SLICE_X9Y120_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y120_SLICE_X9Y120_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y120_SLICE_X9Y120_BO6),
.Q(CLBLM_R_X7Y120_SLICE_X9Y120_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y120_SLICE_X9Y120_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y120_SLICE_X9Y120_CO6),
.Q(CLBLM_R_X7Y120_SLICE_X9Y120_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y120_SLICE_X9Y120_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y120_SLICE_X9Y120_DO6),
.Q(CLBLM_R_X7Y120_SLICE_X9Y120_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hcfcfc0c0afa0afa0)
  ) CLBLM_R_X7Y120_SLICE_X9Y120_DLUT (
.I0(CLBLM_L_X10Y118_SLICE_X12Y118_AQ),
.I1(CLBLM_L_X10Y124_SLICE_X12Y124_AQ),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLM_R_X7Y121_SLICE_X8Y121_BQ),
.I4(CLBLM_L_X8Y119_SLICE_X10Y119_AQ),
.I5(1'b1),
.O5(CLBLM_R_X7Y120_SLICE_X9Y120_DO5),
.O6(CLBLM_R_X7Y120_SLICE_X9Y120_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f0f0f000cc0000)
  ) CLBLM_R_X7Y120_SLICE_X9Y120_CLUT (
.I0(1'b1),
.I1(CLBLM_R_X7Y120_SLICE_X9Y120_CQ),
.I2(CLBLM_L_X8Y120_SLICE_X10Y120_AQ),
.I3(CLBLL_L_X4Y115_SLICE_X4Y115_CQ),
.I4(RIOB33_X105Y105_IOB_X1Y105_I),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLM_R_X7Y120_SLICE_X9Y120_CO5),
.O6(CLBLM_R_X7Y120_SLICE_X9Y120_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f05544f0f00000)
  ) CLBLM_R_X7Y120_SLICE_X9Y120_BLUT (
.I0(RIOB33_X105Y117_IOB_X1Y118_I),
.I1(CLBLM_R_X7Y120_SLICE_X9Y120_BQ),
.I2(CLBLL_L_X4Y113_SLICE_X5Y113_BQ),
.I3(CLBLM_L_X10Y118_SLICE_X12Y118_AQ),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(CLBLM_R_X3Y118_SLICE_X2Y118_AQ),
.O5(CLBLM_R_X7Y120_SLICE_X9Y120_BO5),
.O6(CLBLM_R_X7Y120_SLICE_X9Y120_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'heaeaeaeafffff000)
  ) CLBLM_R_X7Y120_SLICE_X9Y120_ALUT (
.I0(CLBLM_R_X11Y120_SLICE_X14Y120_CO6),
.I1(CLBLM_R_X7Y117_SLICE_X8Y117_AQ),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLM_R_X7Y117_SLICE_X9Y117_BQ),
.I4(CLBLM_R_X7Y122_SLICE_X9Y122_DO6),
.I5(1'b1),
.O5(CLBLM_R_X7Y120_SLICE_X9Y120_AO5),
.O6(CLBLM_R_X7Y120_SLICE_X9Y120_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y121_SLICE_X8Y121_C5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y121_SLICE_X8Y121_CO5),
.Q(CLBLM_R_X7Y121_SLICE_X8Y121_C5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y121_SLICE_X8Y121_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y121_SLICE_X8Y121_AO6),
.Q(CLBLM_R_X7Y121_SLICE_X8Y121_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y121_SLICE_X8Y121_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y121_SLICE_X8Y121_BO6),
.Q(CLBLM_R_X7Y121_SLICE_X8Y121_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y121_SLICE_X8Y121_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y121_SLICE_X8Y121_CO6),
.Q(CLBLM_R_X7Y121_SLICE_X8Y121_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h8000000000000000)
  ) CLBLM_R_X7Y121_SLICE_X8Y121_DLUT (
.I0(CLBLM_R_X7Y121_SLICE_X9Y121_AQ),
.I1(CLBLM_R_X7Y121_SLICE_X9Y121_A5Q),
.I2(CLBLM_R_X7Y121_SLICE_X8Y121_BQ),
.I3(CLBLM_L_X8Y120_SLICE_X10Y120_CQ),
.I4(CLBLM_R_X7Y121_SLICE_X8Y121_AQ),
.I5(CLBLM_R_X7Y121_SLICE_X9Y121_BQ),
.O5(CLBLM_R_X7Y121_SLICE_X8Y121_DO5),
.O6(CLBLM_R_X7Y121_SLICE_X8Y121_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hccffcc00aaf0aaf0)
  ) CLBLM_R_X7Y121_SLICE_X8Y121_CLUT (
.I0(CLBLM_R_X7Y127_SLICE_X8Y127_AQ),
.I1(CLBLM_L_X8Y121_SLICE_X10Y121_AQ),
.I2(CLBLL_L_X2Y117_SLICE_X0Y117_A5Q),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLM_R_X7Y122_SLICE_X9Y122_A5Q),
.I5(1'b1),
.O5(CLBLM_R_X7Y121_SLICE_X8Y121_CO5),
.O6(CLBLM_R_X7Y121_SLICE_X8Y121_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf6f06600fcf0cc00)
  ) CLBLM_R_X7Y121_SLICE_X8Y121_BLUT (
.I0(CLBLM_R_X7Y121_SLICE_X9Y121_A5Q),
.I1(CLBLM_R_X7Y121_SLICE_X8Y121_BQ),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLM_R_X7Y122_SLICE_X9Y122_BO6),
.I4(CLBLM_R_X5Y117_SLICE_X7Y117_AQ),
.I5(CLBLM_L_X8Y120_SLICE_X10Y120_CQ),
.O5(CLBLM_R_X7Y121_SLICE_X8Y121_BO5),
.O6(CLBLM_R_X7Y121_SLICE_X8Y121_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff3c003c003c00)
  ) CLBLM_R_X7Y121_SLICE_X8Y121_ALUT (
.I0(1'b1),
.I1(CLBLM_R_X7Y121_SLICE_X9Y121_DO5),
.I2(CLBLM_R_X7Y121_SLICE_X8Y121_AQ),
.I3(CLBLM_R_X7Y122_SLICE_X9Y122_BO6),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(CLBLL_L_X4Y121_SLICE_X5Y121_AQ),
.O5(CLBLM_R_X7Y121_SLICE_X8Y121_AO5),
.O6(CLBLM_R_X7Y121_SLICE_X8Y121_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y121_SLICE_X9Y121_A5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y121_SLICE_X9Y121_CO6),
.Q(CLBLM_R_X7Y121_SLICE_X9Y121_A5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y121_SLICE_X9Y121_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y121_SLICE_X9Y121_AO6),
.Q(CLBLM_R_X7Y121_SLICE_X9Y121_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y121_SLICE_X9Y121_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y121_SLICE_X9Y121_BO6),
.Q(CLBLM_R_X7Y121_SLICE_X9Y121_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hf1f3f5ff88000000)
  ) CLBLM_R_X7Y121_SLICE_X9Y121_DLUT (
.I0(CLBLM_L_X8Y120_SLICE_X10Y120_CQ),
.I1(CLBLM_R_X7Y121_SLICE_X8Y121_BQ),
.I2(CLBLM_R_X5Y121_SLICE_X7Y121_DO6),
.I3(CLBLM_R_X7Y121_SLICE_X9Y121_A5Q),
.I4(CLBLM_R_X7Y121_SLICE_X9Y121_AQ),
.I5(1'b1),
.O5(CLBLM_R_X7Y121_SLICE_X9Y121_DO5),
.O6(CLBLM_R_X7Y121_SLICE_X9Y121_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hef45fe54f0f00000)
  ) CLBLM_R_X7Y121_SLICE_X9Y121_CLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_L_X8Y133_SLICE_X11Y133_AO6),
.I2(CLBLM_R_X7Y121_SLICE_X9Y121_A5Q),
.I3(CLBLM_L_X8Y118_SLICE_X10Y118_CQ),
.I4(CLBLM_L_X8Y120_SLICE_X10Y120_CQ),
.I5(1'b1),
.O5(CLBLM_R_X7Y121_SLICE_X9Y121_CO5),
.O6(CLBLM_R_X7Y121_SLICE_X9Y121_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'ha0a0a0a0a3acacac)
  ) CLBLM_R_X7Y121_SLICE_X9Y121_BLUT (
.I0(CLBLM_L_X8Y115_SLICE_X11Y115_CQ),
.I1(CLBLM_R_X7Y121_SLICE_X9Y121_BQ),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLM_R_X7Y121_SLICE_X9Y121_DO5),
.I4(CLBLM_R_X7Y121_SLICE_X8Y121_AQ),
.I5(CLBLM_L_X8Y133_SLICE_X11Y133_AO6),
.O5(CLBLM_R_X7Y121_SLICE_X9Y121_BO5),
.O6(CLBLM_R_X7Y121_SLICE_X9Y121_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'habbababa01101010)
  ) CLBLM_R_X7Y121_SLICE_X9Y121_ALUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_L_X8Y133_SLICE_X11Y133_AO6),
.I2(CLBLM_R_X7Y121_SLICE_X9Y121_AQ),
.I3(CLBLM_R_X7Y121_SLICE_X8Y121_BQ),
.I4(CLBLM_R_X7Y121_SLICE_X9Y121_CO5),
.I5(CLBLL_L_X4Y115_SLICE_X4Y115_CQ),
.O5(CLBLM_R_X7Y121_SLICE_X9Y121_AO5),
.O6(CLBLM_R_X7Y121_SLICE_X9Y121_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y122_SLICE_X8Y122_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y122_SLICE_X8Y122_AO6),
.Q(CLBLM_R_X7Y122_SLICE_X8Y122_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y122_SLICE_X8Y122_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y122_SLICE_X8Y122_BO6),
.Q(CLBLM_R_X7Y122_SLICE_X8Y122_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y122_SLICE_X8Y122_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y122_SLICE_X8Y122_CO6),
.Q(CLBLM_R_X7Y122_SLICE_X8Y122_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y122_SLICE_X8Y122_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y122_SLICE_X8Y122_DO6),
.Q(CLBLM_R_X7Y122_SLICE_X8Y122_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h88888888d8d8d8d8)
  ) CLBLM_R_X7Y122_SLICE_X8Y122_DLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_R_X7Y122_SLICE_X8Y122_AQ),
.I2(CLBLM_R_X7Y122_SLICE_X8Y122_DQ),
.I3(1'b1),
.I4(1'b1),
.I5(RIOB33_X105Y105_IOB_X1Y105_I),
.O5(CLBLM_R_X7Y122_SLICE_X8Y122_DO5),
.O6(CLBLM_R_X7Y122_SLICE_X8Y122_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f0f0f055005500)
  ) CLBLM_R_X7Y122_SLICE_X8Y122_CLUT (
.I0(CLBLM_L_X10Y124_SLICE_X13Y124_BO6),
.I1(1'b1),
.I2(CLBLM_L_X8Y118_SLICE_X10Y118_BQ),
.I3(CLBLM_R_X7Y122_SLICE_X8Y122_BQ),
.I4(1'b1),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLM_R_X7Y122_SLICE_X8Y122_CO5),
.O6(CLBLM_R_X7Y122_SLICE_X8Y122_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff00000c0c0c0c)
  ) CLBLM_R_X7Y122_SLICE_X8Y122_BLUT (
.I0(1'b1),
.I1(CLBLM_R_X7Y123_SLICE_X8Y123_BQ),
.I2(CLBLM_L_X10Y124_SLICE_X13Y124_BO6),
.I3(1'b1),
.I4(CLBLM_R_X7Y112_SLICE_X9Y112_CQ),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLM_R_X7Y122_SLICE_X8Y122_BO5),
.O6(CLBLM_R_X7Y122_SLICE_X8Y122_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hff000c0cff000c0c)
  ) CLBLM_R_X7Y122_SLICE_X8Y122_ALUT (
.I0(1'b1),
.I1(CLBLM_L_X10Y122_SLICE_X12Y122_AQ),
.I2(CLBLM_L_X10Y124_SLICE_X13Y124_BO6),
.I3(CLBLM_R_X5Y122_SLICE_X6Y122_BQ),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(1'b1),
.O5(CLBLM_R_X7Y122_SLICE_X8Y122_AO5),
.O6(CLBLM_R_X7Y122_SLICE_X8Y122_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y122_SLICE_X9Y122_A5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y122_SLICE_X9Y122_AO5),
.Q(CLBLM_R_X7Y122_SLICE_X9Y122_A5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y122_SLICE_X9Y122_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y122_SLICE_X9Y122_AO6),
.Q(CLBLM_R_X7Y122_SLICE_X9Y122_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y122_SLICE_X9Y122_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y122_SLICE_X9Y122_BO5),
.Q(CLBLM_R_X7Y122_SLICE_X9Y122_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h6f006f0030003100)
  ) CLBLM_R_X7Y122_SLICE_X9Y122_DLUT (
.I0(CLBLM_R_X7Y124_SLICE_X8Y124_AQ),
.I1(CLBLM_L_X10Y124_SLICE_X12Y124_AQ),
.I2(CLBLM_L_X10Y123_SLICE_X13Y123_DO6),
.I3(CLBLM_R_X5Y122_SLICE_X6Y122_AO5),
.I4(CLBLM_R_X5Y120_SLICE_X6Y120_A5Q),
.I5(CLBLM_R_X7Y120_SLICE_X9Y120_A5Q),
.O5(CLBLM_R_X7Y122_SLICE_X9Y122_DO5),
.O6(CLBLM_R_X7Y122_SLICE_X9Y122_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h4044cccc88880000)
  ) CLBLM_R_X7Y122_SLICE_X9Y122_CLUT (
.I0(CLBLM_L_X10Y118_SLICE_X12Y118_B5Q),
.I1(CLBLM_R_X5Y122_SLICE_X6Y122_AO5),
.I2(CLBLM_L_X10Y123_SLICE_X13Y123_DO6),
.I3(CLBLM_L_X10Y124_SLICE_X12Y124_AQ),
.I4(CLBLM_R_X7Y123_SLICE_X9Y123_BO5),
.I5(CLBLM_R_X5Y120_SLICE_X6Y120_A5Q),
.O5(CLBLM_R_X7Y122_SLICE_X9Y122_CO5),
.O6(CLBLM_R_X7Y122_SLICE_X9Y122_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h08080000f3f00300)
  ) CLBLM_R_X7Y122_SLICE_X9Y122_BLUT (
.I0(CLBLM_L_X8Y120_SLICE_X10Y120_A5Q),
.I1(RIOB33_X105Y105_IOB_X1Y105_I),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLM_R_X3Y112_SLICE_X3Y112_BQ),
.I4(CLBLM_L_X8Y120_SLICE_X11Y120_C5Q),
.I5(1'b1),
.O5(CLBLM_R_X7Y122_SLICE_X9Y122_BO5),
.O6(CLBLM_R_X7Y122_SLICE_X9Y122_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hafafa0a0ff0ff000)
  ) CLBLM_R_X7Y122_SLICE_X9Y122_ALUT (
.I0(CLBLL_L_X2Y117_SLICE_X0Y117_CQ),
.I1(1'b1),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLM_L_X10Y122_SLICE_X13Y122_AQ),
.I4(RIOB33_X105Y143_IOB_X1Y144_I),
.I5(1'b1),
.O5(CLBLM_R_X7Y122_SLICE_X9Y122_AO5),
.O6(CLBLM_R_X7Y122_SLICE_X9Y122_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y123_SLICE_X8Y123_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y123_SLICE_X8Y123_AO6),
.Q(CLBLM_R_X7Y123_SLICE_X8Y123_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y123_SLICE_X8Y123_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y123_SLICE_X8Y123_BO6),
.Q(CLBLM_R_X7Y123_SLICE_X8Y123_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y123_SLICE_X8Y123_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y123_SLICE_X8Y123_CO6),
.Q(CLBLM_R_X7Y123_SLICE_X8Y123_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X7Y123_SLICE_X8Y123_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y123_SLICE_X8Y123_DO5),
.O6(CLBLM_R_X7Y123_SLICE_X8Y123_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hf5f5a0a0e4e4e4e4)
  ) CLBLM_R_X7Y123_SLICE_X8Y123_CLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_R_X7Y123_SLICE_X8Y123_CQ),
.I2(CLBLM_R_X7Y123_SLICE_X8Y123_BQ),
.I3(1'b1),
.I4(CLBLM_L_X10Y126_SLICE_X12Y126_AQ),
.I5(CLBLM_R_X11Y121_SLICE_X14Y121_CO6),
.O5(CLBLM_R_X7Y123_SLICE_X8Y123_CO5),
.O6(CLBLM_R_X7Y123_SLICE_X8Y123_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hff0fff0fff0ff000)
  ) CLBLM_R_X7Y123_SLICE_X8Y123_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLM_R_X7Y119_SLICE_X8Y119_C5Q),
.I4(CLBLM_L_X10Y124_SLICE_X13Y124_BO6),
.I5(CLBLM_R_X7Y122_SLICE_X8Y122_AQ),
.O5(CLBLM_R_X7Y123_SLICE_X8Y123_BO5),
.O6(CLBLM_R_X7Y123_SLICE_X8Y123_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'heaeaaeea40400440)
  ) CLBLM_R_X7Y123_SLICE_X8Y123_ALUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_R_X7Y123_SLICE_X9Y123_BO6),
.I2(CLBLM_R_X7Y123_SLICE_X8Y123_AQ),
.I3(CLBLM_R_X7Y122_SLICE_X8Y122_AQ),
.I4(CLBLM_R_X7Y123_SLICE_X9Y123_AQ),
.I5(CLBLM_R_X7Y120_SLICE_X8Y120_BQ),
.O5(CLBLM_R_X7Y123_SLICE_X8Y123_AO5),
.O6(CLBLM_R_X7Y123_SLICE_X8Y123_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y123_SLICE_X9Y123_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y123_SLICE_X9Y123_AO6),
.Q(CLBLM_R_X7Y123_SLICE_X9Y123_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000044444444)
  ) CLBLM_R_X7Y123_SLICE_X9Y123_DLUT (
.I0(CLBLM_R_X7Y123_SLICE_X8Y123_AQ),
.I1(CLBLM_R_X7Y122_SLICE_X8Y122_AQ),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(CLBLM_R_X7Y123_SLICE_X9Y123_AQ),
.O5(CLBLM_R_X7Y123_SLICE_X9Y123_DO5),
.O6(CLBLM_R_X7Y123_SLICE_X9Y123_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000001000)
  ) CLBLM_R_X7Y123_SLICE_X9Y123_CLUT (
.I0(CLBLM_R_X7Y123_SLICE_X8Y123_AQ),
.I1(CLBLM_R_X7Y123_SLICE_X9Y123_AQ),
.I2(CLBLM_R_X7Y122_SLICE_X8Y122_AQ),
.I3(CLBLM_L_X10Y118_SLICE_X12Y118_B5Q),
.I4(CLBLM_R_X7Y124_SLICE_X9Y124_AQ),
.I5(CLBLM_R_X5Y120_SLICE_X6Y120_A5Q),
.O5(CLBLM_R_X7Y123_SLICE_X9Y123_CO5),
.O6(CLBLM_R_X7Y123_SLICE_X9Y123_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h00ff00fd00000202)
  ) CLBLM_R_X7Y123_SLICE_X9Y123_BLUT (
.I0(CLBLM_R_X7Y122_SLICE_X8Y122_AQ),
.I1(CLBLM_R_X7Y124_SLICE_X9Y124_AQ),
.I2(CLBLM_R_X7Y123_SLICE_X9Y123_AQ),
.I3(CLBLM_L_X10Y123_SLICE_X12Y123_AO6),
.I4(CLBLM_R_X7Y123_SLICE_X8Y123_AQ),
.I5(1'b1),
.O5(CLBLM_R_X7Y123_SLICE_X9Y123_BO5),
.O6(CLBLM_R_X7Y123_SLICE_X9Y123_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hbeaa1400beaa1400)
  ) CLBLM_R_X7Y123_SLICE_X9Y123_ALUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_R_X7Y122_SLICE_X8Y122_AQ),
.I2(CLBLM_R_X7Y123_SLICE_X9Y123_AQ),
.I3(CLBLM_R_X7Y123_SLICE_X9Y123_BO6),
.I4(CLBLM_R_X7Y118_SLICE_X8Y118_BQ),
.I5(1'b1),
.O5(CLBLM_R_X7Y123_SLICE_X9Y123_AO5),
.O6(CLBLM_R_X7Y123_SLICE_X9Y123_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y124_SLICE_X8Y124_A5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y124_SLICE_X8Y124_DO6),
.Q(CLBLM_R_X7Y124_SLICE_X8Y124_A5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y124_SLICE_X8Y124_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y124_SLICE_X8Y124_AO6),
.Q(CLBLM_R_X7Y124_SLICE_X8Y124_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y124_SLICE_X8Y124_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y124_SLICE_X8Y124_BO6),
.Q(CLBLM_R_X7Y124_SLICE_X8Y124_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y124_SLICE_X8Y124_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y124_SLICE_X8Y124_CO6),
.Q(CLBLM_R_X7Y124_SLICE_X8Y124_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaa000c00000c0c)
  ) CLBLM_R_X7Y124_SLICE_X8Y124_DLUT (
.I0(CLBLM_R_X7Y124_SLICE_X9Y124_AQ),
.I1(RIOB33_X105Y105_IOB_X1Y105_I),
.I2(CLBLL_L_X4Y119_SLICE_X4Y119_C5Q),
.I3(CLBLM_R_X7Y124_SLICE_X8Y124_A5Q),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(1'b1),
.O5(CLBLM_R_X7Y124_SLICE_X8Y124_DO5),
.O6(CLBLM_R_X7Y124_SLICE_X8Y124_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hab01aa00ae04aa00)
  ) CLBLM_R_X7Y124_SLICE_X8Y124_CLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_R_X7Y124_SLICE_X8Y124_CQ),
.I2(CLBLL_L_X4Y119_SLICE_X4Y119_C5Q),
.I3(CLBLM_R_X7Y122_SLICE_X8Y122_CQ),
.I4(RIOB33_X105Y105_IOB_X1Y105_I),
.I5(CLBLM_R_X7Y125_SLICE_X8Y125_AO6),
.O5(CLBLM_R_X7Y124_SLICE_X8Y124_CO5),
.O6(CLBLM_R_X7Y124_SLICE_X8Y124_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf101f000f404f000)
  ) CLBLM_R_X7Y124_SLICE_X8Y124_BLUT (
.I0(CLBLL_L_X4Y119_SLICE_X4Y119_C5Q),
.I1(CLBLM_R_X7Y124_SLICE_X8Y124_BQ),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLM_R_X7Y116_SLICE_X8Y116_CQ),
.I4(RIOB33_X105Y105_IOB_X1Y105_I),
.I5(CLBLM_R_X7Y124_SLICE_X8Y124_A5Q),
.O5(CLBLM_R_X7Y124_SLICE_X8Y124_BO5),
.O6(CLBLM_R_X7Y124_SLICE_X8Y124_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaa3300aaaa3030)
  ) CLBLM_R_X7Y124_SLICE_X8Y124_ALUT (
.I0(CLBLM_R_X5Y124_SLICE_X6Y124_AQ),
.I1(RIOB33_X105Y121_IOB_X1Y121_I),
.I2(CLBLM_R_X7Y124_SLICE_X8Y124_AQ),
.I3(CLBLM_R_X7Y120_SLICE_X9Y120_A5Q),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(CLBLM_L_X10Y123_SLICE_X13Y123_DO6),
.O5(CLBLM_R_X7Y124_SLICE_X8Y124_AO5),
.O6(CLBLM_R_X7Y124_SLICE_X8Y124_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y124_SLICE_X9Y124_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y124_SLICE_X9Y124_AO6),
.Q(CLBLM_R_X7Y124_SLICE_X9Y124_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X7Y124_SLICE_X9Y124_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y124_SLICE_X9Y124_DO5),
.O6(CLBLM_R_X7Y124_SLICE_X9Y124_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X7Y124_SLICE_X9Y124_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y124_SLICE_X9Y124_CO5),
.O6(CLBLM_R_X7Y124_SLICE_X9Y124_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X7Y124_SLICE_X9Y124_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y124_SLICE_X9Y124_BO5),
.O6(CLBLM_R_X7Y124_SLICE_X9Y124_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hff00ffffff005a5a)
  ) CLBLM_R_X7Y124_SLICE_X9Y124_ALUT (
.I0(CLBLM_R_X7Y123_SLICE_X9Y123_DO6),
.I1(1'b1),
.I2(CLBLM_R_X7Y124_SLICE_X9Y124_AQ),
.I3(CLBLM_R_X5Y114_SLICE_X6Y114_BQ),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(CLBLM_L_X10Y123_SLICE_X12Y123_AO6),
.O5(CLBLM_R_X7Y124_SLICE_X9Y124_AO5),
.O6(CLBLM_R_X7Y124_SLICE_X9Y124_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X7Y125_SLICE_X8Y125_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y125_SLICE_X8Y125_DO5),
.O6(CLBLM_R_X7Y125_SLICE_X8Y125_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X7Y125_SLICE_X8Y125_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y125_SLICE_X8Y125_CO5),
.O6(CLBLM_R_X7Y125_SLICE_X8Y125_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X7Y125_SLICE_X8Y125_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y125_SLICE_X8Y125_BO5),
.O6(CLBLM_R_X7Y125_SLICE_X8Y125_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hcc000000cc000000)
  ) CLBLM_R_X7Y125_SLICE_X8Y125_ALUT (
.I0(1'b1),
.I1(CLBLM_R_X7Y124_SLICE_X8Y124_A5Q),
.I2(1'b1),
.I3(CLBLL_L_X4Y123_SLICE_X4Y123_AQ),
.I4(CLBLM_R_X7Y124_SLICE_X8Y124_BQ),
.I5(1'b1),
.O5(CLBLM_R_X7Y125_SLICE_X8Y125_AO5),
.O6(CLBLM_R_X7Y125_SLICE_X8Y125_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X7Y125_SLICE_X9Y125_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y125_SLICE_X9Y125_DO5),
.O6(CLBLM_R_X7Y125_SLICE_X9Y125_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X7Y125_SLICE_X9Y125_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y125_SLICE_X9Y125_CO5),
.O6(CLBLM_R_X7Y125_SLICE_X9Y125_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X7Y125_SLICE_X9Y125_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y125_SLICE_X9Y125_BO5),
.O6(CLBLM_R_X7Y125_SLICE_X9Y125_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X7Y125_SLICE_X9Y125_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y125_SLICE_X9Y125_AO5),
.O6(CLBLM_R_X7Y125_SLICE_X9Y125_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y127_SLICE_X8Y127_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y128_SLICE_X10Y128_AO6),
.Q(CLBLM_R_X7Y127_SLICE_X8Y127_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X7Y127_SLICE_X8Y127_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y127_SLICE_X8Y127_DO5),
.O6(CLBLM_R_X7Y127_SLICE_X8Y127_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X7Y127_SLICE_X8Y127_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y127_SLICE_X8Y127_CO5),
.O6(CLBLM_R_X7Y127_SLICE_X8Y127_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X7Y127_SLICE_X8Y127_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y127_SLICE_X8Y127_BO5),
.O6(CLBLM_R_X7Y127_SLICE_X8Y127_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X7Y127_SLICE_X8Y127_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y127_SLICE_X8Y127_AO5),
.O6(CLBLM_R_X7Y127_SLICE_X8Y127_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X7Y127_SLICE_X9Y127_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y127_SLICE_X9Y127_DO5),
.O6(CLBLM_R_X7Y127_SLICE_X9Y127_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X7Y127_SLICE_X9Y127_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y127_SLICE_X9Y127_CO5),
.O6(CLBLM_R_X7Y127_SLICE_X9Y127_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X7Y127_SLICE_X9Y127_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y127_SLICE_X9Y127_BO5),
.O6(CLBLM_R_X7Y127_SLICE_X9Y127_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X7Y127_SLICE_X9Y127_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y127_SLICE_X9Y127_AO5),
.O6(CLBLM_R_X7Y127_SLICE_X9Y127_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y128_SLICE_X8Y128_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y128_SLICE_X8Y128_AO6),
.Q(CLBLM_R_X7Y128_SLICE_X8Y128_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X7Y128_SLICE_X8Y128_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y128_SLICE_X8Y128_DO5),
.O6(CLBLM_R_X7Y128_SLICE_X8Y128_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X7Y128_SLICE_X8Y128_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y128_SLICE_X8Y128_CO5),
.O6(CLBLM_R_X7Y128_SLICE_X8Y128_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X7Y128_SLICE_X8Y128_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y128_SLICE_X8Y128_BO5),
.O6(CLBLM_R_X7Y128_SLICE_X8Y128_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hcccca0aa00aa00aa)
  ) CLBLM_R_X7Y128_SLICE_X8Y128_ALUT (
.I0(CLBLM_L_X8Y120_SLICE_X10Y120_A5Q),
.I1(CLBLM_L_X8Y117_SLICE_X11Y117_BQ),
.I2(CLBLM_R_X7Y128_SLICE_X8Y128_AQ),
.I3(RIOB33_X105Y141_IOB_X1Y142_I),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(1'b1),
.O5(CLBLM_R_X7Y128_SLICE_X8Y128_AO5),
.O6(CLBLM_R_X7Y128_SLICE_X8Y128_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X7Y128_SLICE_X9Y128_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y128_SLICE_X9Y128_DO5),
.O6(CLBLM_R_X7Y128_SLICE_X9Y128_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X7Y128_SLICE_X9Y128_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y128_SLICE_X9Y128_CO5),
.O6(CLBLM_R_X7Y128_SLICE_X9Y128_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X7Y128_SLICE_X9Y128_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y128_SLICE_X9Y128_BO5),
.O6(CLBLM_R_X7Y128_SLICE_X9Y128_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X7Y128_SLICE_X9Y128_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y128_SLICE_X9Y128_AO5),
.O6(CLBLM_R_X7Y128_SLICE_X9Y128_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X7Y151_SLICE_X8Y151_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y151_SLICE_X8Y151_DO5),
.O6(CLBLM_R_X7Y151_SLICE_X8Y151_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X7Y151_SLICE_X8Y151_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y151_SLICE_X8Y151_CO5),
.O6(CLBLM_R_X7Y151_SLICE_X8Y151_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X7Y151_SLICE_X8Y151_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y151_SLICE_X8Y151_BO5),
.O6(CLBLM_R_X7Y151_SLICE_X8Y151_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h00000000ffffffff)
  ) CLBLM_R_X7Y151_SLICE_X8Y151_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(CLBLM_R_X5Y113_SLICE_X7Y113_A5Q),
.O5(CLBLM_R_X7Y151_SLICE_X8Y151_AO5),
.O6(CLBLM_R_X7Y151_SLICE_X8Y151_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X7Y151_SLICE_X9Y151_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y151_SLICE_X9Y151_DO5),
.O6(CLBLM_R_X7Y151_SLICE_X9Y151_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X7Y151_SLICE_X9Y151_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y151_SLICE_X9Y151_CO5),
.O6(CLBLM_R_X7Y151_SLICE_X9Y151_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X7Y151_SLICE_X9Y151_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y151_SLICE_X9Y151_BO5),
.O6(CLBLM_R_X7Y151_SLICE_X9Y151_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X7Y151_SLICE_X9Y151_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y151_SLICE_X9Y151_AO5),
.O6(CLBLM_R_X7Y151_SLICE_X9Y151_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y113_SLICE_X14Y113_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y113_SLICE_X14Y113_AO6),
.Q(CLBLM_R_X11Y113_SLICE_X14Y113_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y113_SLICE_X14Y113_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y113_SLICE_X14Y113_BO6),
.Q(CLBLM_R_X11Y113_SLICE_X14Y113_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffffafffffffa)
  ) CLBLM_R_X11Y113_SLICE_X14Y113_DLUT (
.I0(CLBLM_L_X8Y113_SLICE_X11Y113_BQ),
.I1(1'b1),
.I2(CLBLM_L_X10Y112_SLICE_X13Y112_BQ),
.I3(CLBLM_L_X8Y111_SLICE_X10Y111_AQ),
.I4(CLBLM_R_X11Y114_SLICE_X14Y114_CQ),
.I5(1'b1),
.O5(CLBLM_R_X11Y113_SLICE_X14Y113_DO5),
.O6(CLBLM_R_X11Y113_SLICE_X14Y113_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0404150415150415)
  ) CLBLM_R_X11Y113_SLICE_X14Y113_CLUT (
.I0(CLBLM_R_X11Y113_SLICE_X14Y113_BQ),
.I1(CLBLM_R_X5Y111_SLICE_X7Y111_DO6),
.I2(CLBLM_L_X10Y122_SLICE_X13Y122_A5Q),
.I3(CLBLM_L_X10Y112_SLICE_X13Y112_CQ),
.I4(CLBLM_L_X10Y113_SLICE_X12Y113_AO5),
.I5(CLBLM_R_X11Y117_SLICE_X14Y117_BQ),
.O5(CLBLM_R_X11Y113_SLICE_X14Y113_CO5),
.O6(CLBLM_R_X11Y113_SLICE_X14Y113_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h88888888bbbb88bb)
  ) CLBLM_R_X11Y113_SLICE_X14Y113_BLUT (
.I0(CLBLM_R_X11Y114_SLICE_X14Y114_CQ),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(1'b1),
.I3(RIOB33_X105Y141_IOB_X1Y142_I),
.I4(CLBLM_R_X7Y128_SLICE_X8Y128_AQ),
.I5(CLBLM_R_X11Y113_SLICE_X14Y113_CO6),
.O5(CLBLM_R_X11Y113_SLICE_X14Y113_BO5),
.O6(CLBLM_R_X11Y113_SLICE_X14Y113_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffa0cc0000a0cc)
  ) CLBLM_R_X11Y113_SLICE_X14Y113_ALUT (
.I0(RIOB33_X105Y105_IOB_X1Y105_I),
.I1(CLBLM_L_X8Y112_SLICE_X10Y112_AQ),
.I2(CLBLM_R_X11Y113_SLICE_X14Y113_AQ),
.I3(CLBLM_L_X10Y113_SLICE_X12Y113_DO6),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(CLBLM_L_X10Y121_SLICE_X13Y121_AQ),
.O5(CLBLM_R_X11Y113_SLICE_X14Y113_AO5),
.O6(CLBLM_R_X11Y113_SLICE_X14Y113_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y113_SLICE_X15Y113_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y113_SLICE_X15Y113_AO6),
.Q(CLBLM_R_X11Y113_SLICE_X15Y113_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y113_SLICE_X15Y113_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y113_SLICE_X15Y113_BO6),
.Q(CLBLM_R_X11Y113_SLICE_X15Y113_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h00000000ffaaffaa)
  ) CLBLM_R_X11Y113_SLICE_X15Y113_DLUT (
.I0(CLBLM_L_X10Y112_SLICE_X12Y112_BQ),
.I1(1'b1),
.I2(1'b1),
.I3(CLBLM_R_X5Y109_SLICE_X7Y109_AQ),
.I4(1'b1),
.I5(CLBLM_R_X3Y117_SLICE_X3Y117_BQ),
.O5(CLBLM_R_X11Y113_SLICE_X15Y113_DO5),
.O6(CLBLM_R_X11Y113_SLICE_X15Y113_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffccffffffcc)
  ) CLBLM_R_X11Y113_SLICE_X15Y113_CLUT (
.I0(1'b1),
.I1(CLBLM_L_X8Y113_SLICE_X11Y113_AQ),
.I2(1'b1),
.I3(CLBLM_L_X8Y112_SLICE_X10Y112_BQ),
.I4(CLBLM_R_X11Y113_SLICE_X15Y113_AQ),
.I5(1'b1),
.O5(CLBLM_R_X11Y113_SLICE_X15Y113_CO5),
.O6(CLBLM_R_X11Y113_SLICE_X15Y113_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f0f0f088ff8800)
  ) CLBLM_R_X11Y113_SLICE_X15Y113_BLUT (
.I0(RIOB33_X105Y105_IOB_X1Y105_I),
.I1(CLBLM_R_X11Y113_SLICE_X15Y113_BQ),
.I2(CLBLM_L_X12Y115_SLICE_X16Y115_AQ),
.I3(CLBLM_L_X10Y113_SLICE_X12Y113_DO6),
.I4(CLBLM_L_X10Y113_SLICE_X13Y113_AO6),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLM_R_X11Y113_SLICE_X15Y113_BO5),
.O6(CLBLM_R_X11Y113_SLICE_X15Y113_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff0000b380b380)
  ) CLBLM_R_X11Y113_SLICE_X15Y113_ALUT (
.I0(RIOB33_X105Y105_IOB_X1Y105_I),
.I1(CLBLM_L_X10Y113_SLICE_X12Y113_DO6),
.I2(CLBLM_R_X11Y113_SLICE_X15Y113_AQ),
.I3(CLBLM_L_X10Y112_SLICE_X13Y112_BQ),
.I4(CLBLM_R_X11Y119_SLICE_X15Y119_BQ),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLM_R_X11Y113_SLICE_X15Y113_AO5),
.O6(CLBLM_R_X11Y113_SLICE_X15Y113_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y114_SLICE_X14Y114_D5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y114_SLICE_X14Y114_DO5),
.Q(CLBLM_R_X11Y114_SLICE_X14Y114_D5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y114_SLICE_X14Y114_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y114_SLICE_X14Y114_AO6),
.Q(CLBLM_R_X11Y114_SLICE_X14Y114_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y114_SLICE_X14Y114_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y114_SLICE_X14Y114_BO6),
.Q(CLBLM_R_X11Y114_SLICE_X14Y114_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y114_SLICE_X14Y114_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y114_SLICE_X14Y114_CO6),
.Q(CLBLM_R_X11Y114_SLICE_X14Y114_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y114_SLICE_X14Y114_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y114_SLICE_X14Y114_DO6),
.Q(CLBLM_R_X11Y114_SLICE_X14Y114_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f0ff00aaaacccc)
  ) CLBLM_R_X11Y114_SLICE_X14Y114_DLUT (
.I0(CLBLM_L_X10Y114_SLICE_X13Y114_CQ),
.I1(CLBLM_L_X8Y115_SLICE_X10Y115_C5Q),
.I2(CLBLM_R_X11Y114_SLICE_X14Y114_AQ),
.I3(RIOB33_X105Y103_IOB_X1Y104_I),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(1'b1),
.O5(CLBLM_R_X11Y114_SLICE_X14Y114_DO5),
.O6(CLBLM_R_X11Y114_SLICE_X14Y114_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f0f0f0ccaa00aa)
  ) CLBLM_R_X11Y114_SLICE_X14Y114_CLUT (
.I0(CLBLM_L_X8Y113_SLICE_X11Y113_AQ),
.I1(CLBLM_R_X11Y114_SLICE_X14Y114_CQ),
.I2(CLBLM_L_X12Y115_SLICE_X16Y115_CQ),
.I3(CLBLM_L_X10Y113_SLICE_X12Y113_DO6),
.I4(RIOB33_X105Y105_IOB_X1Y105_I),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLM_R_X11Y114_SLICE_X14Y114_CO5),
.O6(CLBLM_R_X11Y114_SLICE_X14Y114_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hff880088fff000f0)
  ) CLBLM_R_X11Y114_SLICE_X14Y114_BLUT (
.I0(RIOB33_X105Y105_IOB_X1Y105_I),
.I1(CLBLM_R_X11Y114_SLICE_X14Y114_BQ),
.I2(CLBLM_L_X8Y113_SLICE_X11Y113_BQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLM_L_X10Y120_SLICE_X13Y120_BQ),
.I5(CLBLM_L_X10Y113_SLICE_X12Y113_DO6),
.O5(CLBLM_R_X11Y114_SLICE_X14Y114_BO5),
.O6(CLBLM_R_X11Y114_SLICE_X14Y114_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hec20ec20ff33cc00)
  ) CLBLM_R_X11Y114_SLICE_X14Y114_ALUT (
.I0(RIOB33_X105Y105_IOB_X1Y105_I),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(CLBLM_R_X11Y114_SLICE_X14Y114_AQ),
.I3(CLBLM_R_X11Y117_SLICE_X14Y117_AQ),
.I4(CLBLM_R_X11Y114_SLICE_X14Y114_CQ),
.I5(CLBLM_L_X10Y113_SLICE_X12Y113_DO6),
.O5(CLBLM_R_X11Y114_SLICE_X14Y114_AO5),
.O6(CLBLM_R_X11Y114_SLICE_X14Y114_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X11Y114_SLICE_X15Y114_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X11Y114_SLICE_X15Y114_DO5),
.O6(CLBLM_R_X11Y114_SLICE_X15Y114_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X11Y114_SLICE_X15Y114_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X11Y114_SLICE_X15Y114_CO5),
.O6(CLBLM_R_X11Y114_SLICE_X15Y114_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X11Y114_SLICE_X15Y114_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X11Y114_SLICE_X15Y114_BO5),
.O6(CLBLM_R_X11Y114_SLICE_X15Y114_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X11Y114_SLICE_X15Y114_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X11Y114_SLICE_X15Y114_AO5),
.O6(CLBLM_R_X11Y114_SLICE_X15Y114_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y115_SLICE_X14Y115_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y115_SLICE_X14Y115_AO6),
.Q(CLBLM_R_X11Y115_SLICE_X14Y115_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y115_SLICE_X14Y115_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y115_SLICE_X14Y115_BO6),
.Q(CLBLM_R_X11Y115_SLICE_X14Y115_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y115_SLICE_X14Y115_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y115_SLICE_X14Y115_CO6),
.Q(CLBLM_R_X11Y115_SLICE_X14Y115_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y115_SLICE_X14Y115_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y115_SLICE_X14Y115_DO6),
.Q(CLBLM_R_X11Y115_SLICE_X14Y115_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hffeefeeeddccdccc)
  ) CLBLM_R_X11Y115_SLICE_X14Y115_DLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_R_X7Y113_SLICE_X8Y113_DO6),
.I2(CLBLM_R_X3Y118_SLICE_X2Y118_AQ),
.I3(CLBLM_R_X11Y115_SLICE_X14Y115_DQ),
.I4(RIOB33_X105Y117_IOB_X1Y118_I),
.I5(CLBLM_L_X8Y115_SLICE_X10Y115_C5Q),
.O5(CLBLM_R_X11Y115_SLICE_X14Y115_DO5),
.O6(CLBLM_R_X11Y115_SLICE_X14Y115_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hf000f0aaf000f0ff)
  ) CLBLM_R_X11Y115_SLICE_X14Y115_CLUT (
.I0(CLBLM_R_X7Y128_SLICE_X8Y128_AQ),
.I1(1'b1),
.I2(CLBLM_R_X7Y117_SLICE_X9Y117_CQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLM_L_X10Y115_SLICE_X13Y115_AO6),
.I5(RIOB33_X105Y141_IOB_X1Y142_I),
.O5(CLBLM_R_X11Y115_SLICE_X14Y115_CO5),
.O6(CLBLM_R_X11Y115_SLICE_X14Y115_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hccccfcff00003033)
  ) CLBLM_R_X11Y115_SLICE_X14Y115_BLUT (
.I0(1'b1),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(CLBLM_R_X7Y128_SLICE_X8Y128_AQ),
.I3(RIOB33_X105Y141_IOB_X1Y142_I),
.I4(CLBLM_L_X10Y115_SLICE_X13Y115_BO6),
.I5(CLBLM_R_X11Y115_SLICE_X14Y115_DQ),
.O5(CLBLM_R_X11Y115_SLICE_X14Y115_BO5),
.O6(CLBLM_R_X11Y115_SLICE_X14Y115_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffa0ff8aa0a08a8a)
  ) CLBLM_R_X11Y115_SLICE_X14Y115_ALUT (
.I0(CLBLM_R_X11Y116_SLICE_X14Y116_BO5),
.I1(CLBLM_L_X10Y110_SLICE_X13Y110_CO5),
.I2(CLBLM_R_X11Y115_SLICE_X14Y115_AQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLM_L_X10Y113_SLICE_X12Y113_DO6),
.I5(CLBLM_R_X11Y120_SLICE_X15Y120_CQ),
.O5(CLBLM_R_X11Y115_SLICE_X14Y115_AO5),
.O6(CLBLM_R_X11Y115_SLICE_X14Y115_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y115_SLICE_X15Y115_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y115_SLICE_X15Y115_AO6),
.Q(CLBLM_R_X11Y115_SLICE_X15Y115_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y115_SLICE_X15Y115_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y115_SLICE_X15Y115_BO6),
.Q(CLBLM_R_X11Y115_SLICE_X15Y115_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y115_SLICE_X15Y115_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y115_SLICE_X15Y115_CO6),
.Q(CLBLM_R_X11Y115_SLICE_X15Y115_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y115_SLICE_X15Y115_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y115_SLICE_X15Y115_DO6),
.Q(CLBLM_R_X11Y115_SLICE_X15Y115_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hcccc5555cccc5050)
  ) CLBLM_R_X11Y115_SLICE_X15Y115_DLUT (
.I0(CLBLM_R_X5Y111_SLICE_X7Y111_DO6),
.I1(CLBLM_R_X11Y115_SLICE_X15Y115_CQ),
.I2(CLBLM_R_X11Y115_SLICE_X15Y115_DQ),
.I3(1'b1),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(CLBLM_R_X11Y117_SLICE_X14Y117_BQ),
.O5(CLBLM_R_X11Y115_SLICE_X15Y115_DO5),
.O6(CLBLM_R_X11Y115_SLICE_X15Y115_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f0f0f055445544)
  ) CLBLM_R_X11Y115_SLICE_X15Y115_CLUT (
.I0(CLBLM_R_X5Y111_SLICE_X7Y111_DO6),
.I1(CLBLM_R_X11Y115_SLICE_X15Y115_CQ),
.I2(CLBLM_R_X11Y115_SLICE_X15Y115_BQ),
.I3(CLBLM_L_X10Y115_SLICE_X12Y115_DQ),
.I4(1'b1),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLM_R_X11Y115_SLICE_X15Y115_CO5),
.O6(CLBLM_R_X11Y115_SLICE_X15Y115_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf000f0fff000f0cc)
  ) CLBLM_R_X11Y115_SLICE_X15Y115_BLUT (
.I0(1'b1),
.I1(CLBLM_R_X11Y115_SLICE_X15Y115_DQ),
.I2(CLBLM_L_X8Y113_SLICE_X11Y113_BQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLM_R_X5Y111_SLICE_X7Y111_DO6),
.I5(CLBLM_R_X11Y115_SLICE_X15Y115_BQ),
.O5(CLBLM_R_X11Y115_SLICE_X15Y115_BO5),
.O6(CLBLM_R_X11Y115_SLICE_X15Y115_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffffccf0cca0)
  ) CLBLM_R_X11Y115_SLICE_X15Y115_ALUT (
.I0(CLBLM_R_X3Y118_SLICE_X2Y118_AQ),
.I1(CLBLM_R_X11Y115_SLICE_X15Y115_DQ),
.I2(CLBLM_R_X11Y115_SLICE_X15Y115_AQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(RIOB33_X105Y117_IOB_X1Y118_I),
.I5(CLBLM_R_X5Y112_SLICE_X7Y112_BO6),
.O5(CLBLM_R_X11Y115_SLICE_X15Y115_AO5),
.O6(CLBLM_R_X11Y115_SLICE_X15Y115_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y116_SLICE_X14Y116_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y116_SLICE_X14Y116_AO6),
.Q(CLBLM_R_X11Y116_SLICE_X14Y116_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y116_SLICE_X14Y116_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y116_SLICE_X14Y116_CO6),
.Q(CLBLM_R_X11Y116_SLICE_X14Y116_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y116_SLICE_X14Y116_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y116_SLICE_X14Y116_DO6),
.Q(CLBLM_R_X11Y116_SLICE_X14Y116_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaaaaaa0f000f00)
  ) CLBLM_R_X11Y116_SLICE_X14Y116_DLUT (
.I0(CLBLM_R_X11Y118_SLICE_X15Y118_AQ),
.I1(1'b1),
.I2(RIOB33_X105Y105_IOB_X1Y105_I),
.I3(CLBLL_L_X4Y114_SLICE_X5Y114_AQ),
.I4(1'b1),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLM_R_X11Y116_SLICE_X14Y116_DO5),
.O6(CLBLM_R_X11Y116_SLICE_X14Y116_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f0f0f0002200cc)
  ) CLBLM_R_X11Y116_SLICE_X14Y116_CLUT (
.I0(CLBLM_L_X10Y116_SLICE_X12Y116_BQ),
.I1(CLBLM_R_X11Y116_SLICE_X14Y116_CQ),
.I2(CLBLM_L_X12Y115_SLICE_X16Y115_DQ),
.I3(CLBLM_R_X11Y119_SLICE_X14Y119_AO6),
.I4(CLBLM_L_X10Y116_SLICE_X13Y116_CO5),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLM_R_X11Y116_SLICE_X14Y116_CO5),
.O6(CLBLM_R_X11Y116_SLICE_X14Y116_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hff000a0a00003030)
  ) CLBLM_R_X11Y116_SLICE_X14Y116_BLUT (
.I0(CLBLM_R_X7Y119_SLICE_X9Y119_AQ),
.I1(CLBLM_R_X7Y120_SLICE_X9Y120_DQ),
.I2(RIOB33_X105Y105_IOB_X1Y105_I),
.I3(CLBLM_L_X8Y119_SLICE_X10Y119_CQ),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(1'b1),
.O5(CLBLM_R_X11Y116_SLICE_X14Y116_BO5),
.O6(CLBLM_R_X11Y116_SLICE_X14Y116_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hff000000fffa00fa)
  ) CLBLM_R_X11Y116_SLICE_X14Y116_ALUT (
.I0(CLBLM_L_X10Y119_SLICE_X12Y119_CQ),
.I1(1'b1),
.I2(CLBLM_R_X11Y116_SLICE_X14Y116_AQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLM_L_X10Y116_SLICE_X12Y116_BQ),
.I5(CLBLM_R_X11Y121_SLICE_X14Y121_CO6),
.O5(CLBLM_R_X11Y116_SLICE_X14Y116_AO5),
.O6(CLBLM_R_X11Y116_SLICE_X14Y116_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y116_SLICE_X15Y116_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y116_SLICE_X15Y116_AO6),
.Q(CLBLM_R_X11Y116_SLICE_X15Y116_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X11Y116_SLICE_X15Y116_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X11Y116_SLICE_X15Y116_DO5),
.O6(CLBLM_R_X11Y116_SLICE_X15Y116_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X11Y116_SLICE_X15Y116_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X11Y116_SLICE_X15Y116_CO5),
.O6(CLBLM_R_X11Y116_SLICE_X15Y116_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X11Y116_SLICE_X15Y116_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X11Y116_SLICE_X15Y116_BO5),
.O6(CLBLM_R_X11Y116_SLICE_X15Y116_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffaffeaaafaaaea)
  ) CLBLM_R_X11Y116_SLICE_X15Y116_ALUT (
.I0(CLBLM_R_X7Y113_SLICE_X8Y113_DO6),
.I1(CLBLM_R_X3Y118_SLICE_X2Y118_AQ),
.I2(CLBLM_R_X11Y116_SLICE_X15Y116_AQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(RIOB33_X105Y117_IOB_X1Y118_I),
.I5(CLBLM_R_X11Y119_SLICE_X14Y119_AQ),
.O5(CLBLM_R_X11Y116_SLICE_X15Y116_AO5),
.O6(CLBLM_R_X11Y116_SLICE_X15Y116_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y117_SLICE_X14Y117_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y117_SLICE_X14Y117_AO6),
.Q(CLBLM_R_X11Y117_SLICE_X14Y117_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y117_SLICE_X14Y117_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y117_SLICE_X14Y117_BO6),
.Q(CLBLM_R_X11Y117_SLICE_X14Y117_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y117_SLICE_X14Y117_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y117_SLICE_X14Y117_CO6),
.Q(CLBLM_R_X11Y117_SLICE_X14Y117_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0f0a0f0a0f0f0c0c)
  ) CLBLM_R_X11Y117_SLICE_X14Y117_DLUT (
.I0(CLBLM_R_X11Y115_SLICE_X15Y115_AQ),
.I1(CLBLM_R_X11Y117_SLICE_X14Y117_CQ),
.I2(CLBLM_R_X3Y117_SLICE_X3Y117_BQ),
.I3(CLBLM_L_X8Y117_SLICE_X11Y117_DQ),
.I4(CLBLL_L_X4Y111_SLICE_X4Y111_AQ),
.I5(1'b1),
.O5(CLBLM_R_X11Y117_SLICE_X14Y117_DO5),
.O6(CLBLM_R_X11Y117_SLICE_X14Y117_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hfafafcfcfafafcf0)
  ) CLBLM_R_X11Y117_SLICE_X14Y117_CLUT (
.I0(CLBLM_R_X11Y118_SLICE_X14Y118_AQ),
.I1(CLBLM_R_X11Y117_SLICE_X14Y117_CQ),
.I2(CLBLM_R_X7Y113_SLICE_X9Y113_CO6),
.I3(RIOB33_X105Y117_IOB_X1Y118_I),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(CLBLM_R_X3Y118_SLICE_X2Y118_AQ),
.O5(CLBLM_R_X11Y117_SLICE_X14Y117_CO5),
.O6(CLBLM_R_X11Y117_SLICE_X14Y117_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hff00ff000000eeee)
  ) CLBLM_R_X11Y117_SLICE_X14Y117_BLUT (
.I0(CLBLM_L_X8Y110_SLICE_X10Y110_AQ),
.I1(CLBLM_R_X11Y117_SLICE_X14Y117_BQ),
.I2(1'b1),
.I3(CLBLM_R_X7Y117_SLICE_X8Y117_BQ),
.I4(CLBLM_R_X5Y111_SLICE_X7Y111_DO6),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLM_R_X11Y117_SLICE_X14Y117_BO5),
.O6(CLBLM_R_X11Y117_SLICE_X14Y117_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'haa30aa30aaffaa00)
  ) CLBLM_R_X11Y117_SLICE_X14Y117_ALUT (
.I0(CLBLL_L_X4Y113_SLICE_X4Y113_AQ),
.I1(CLBLM_R_X11Y119_SLICE_X14Y119_AO6),
.I2(CLBLM_R_X11Y117_SLICE_X14Y117_AQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLM_L_X10Y118_SLICE_X13Y118_AQ),
.I5(CLBLM_L_X12Y119_SLICE_X17Y119_AO5),
.O5(CLBLM_R_X11Y117_SLICE_X14Y117_AO5),
.O6(CLBLM_R_X11Y117_SLICE_X14Y117_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y117_SLICE_X15Y117_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y117_SLICE_X15Y117_AO6),
.Q(CLBLM_R_X11Y117_SLICE_X15Y117_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X11Y117_SLICE_X15Y117_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X11Y117_SLICE_X15Y117_DO5),
.O6(CLBLM_R_X11Y117_SLICE_X15Y117_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X11Y117_SLICE_X15Y117_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X11Y117_SLICE_X15Y117_CO5),
.O6(CLBLM_R_X11Y117_SLICE_X15Y117_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X11Y117_SLICE_X15Y117_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X11Y117_SLICE_X15Y117_BO5),
.O6(CLBLM_R_X11Y117_SLICE_X15Y117_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hccfceeee00302222)
  ) CLBLM_R_X11Y117_SLICE_X15Y117_ALUT (
.I0(CLBLM_R_X11Y118_SLICE_X15Y118_BQ),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(CLBLM_R_X11Y117_SLICE_X15Y117_AQ),
.I3(CLBLM_R_X11Y119_SLICE_X14Y119_AO6),
.I4(CLBLM_L_X12Y119_SLICE_X17Y119_AO5),
.I5(CLBLM_L_X8Y117_SLICE_X11Y117_DQ),
.O5(CLBLM_R_X11Y117_SLICE_X15Y117_AO5),
.O6(CLBLM_R_X11Y117_SLICE_X15Y117_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y118_SLICE_X14Y118_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y118_SLICE_X14Y118_AO6),
.Q(CLBLM_R_X11Y118_SLICE_X14Y118_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y118_SLICE_X14Y118_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y118_SLICE_X14Y118_BO6),
.Q(CLBLM_R_X11Y118_SLICE_X14Y118_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y118_SLICE_X14Y118_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y118_SLICE_X14Y118_CO6),
.Q(CLBLM_R_X11Y118_SLICE_X14Y118_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h000f000f5555777f)
  ) CLBLM_R_X11Y118_SLICE_X14Y118_DLUT (
.I0(CLBLM_L_X10Y116_SLICE_X12Y116_DO5),
.I1(CLBLM_R_X11Y118_SLICE_X14Y118_AQ),
.I2(CLBLM_L_X10Y119_SLICE_X13Y119_AQ),
.I3(CLBLM_R_X11Y118_SLICE_X14Y118_BQ),
.I4(CLBLM_R_X11Y120_SLICE_X14Y120_BO5),
.I5(1'b1),
.O5(CLBLM_R_X11Y118_SLICE_X14Y118_DO5),
.O6(CLBLM_R_X11Y118_SLICE_X14Y118_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaa0f0caaaa0000)
  ) CLBLM_R_X11Y118_SLICE_X14Y118_CLUT (
.I0(CLBLM_L_X8Y114_SLICE_X10Y114_BQ),
.I1(CLBLM_R_X11Y118_SLICE_X14Y118_CQ),
.I2(RIOB33_X105Y117_IOB_X1Y118_I),
.I3(CLBLM_R_X5Y115_SLICE_X7Y115_CO6),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(CLBLM_R_X3Y118_SLICE_X2Y118_AQ),
.O5(CLBLM_R_X11Y118_SLICE_X14Y118_CO5),
.O6(CLBLM_R_X11Y118_SLICE_X14Y118_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff000070607060)
  ) CLBLM_R_X11Y118_SLICE_X14Y118_BLUT (
.I0(CLBLM_R_X11Y120_SLICE_X14Y120_DO6),
.I1(CLBLM_R_X11Y118_SLICE_X14Y118_BQ),
.I2(RIOB33_X105Y121_IOB_X1Y121_I),
.I3(CLBLM_R_X11Y119_SLICE_X14Y119_AO6),
.I4(CLBLM_R_X11Y115_SLICE_X14Y115_AQ),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLM_R_X11Y118_SLICE_X14Y118_BO5),
.O6(CLBLM_R_X11Y118_SLICE_X14Y118_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hccffccffcc05ccf0)
  ) CLBLM_R_X11Y118_SLICE_X14Y118_ALUT (
.I0(CLBLM_R_X11Y118_SLICE_X14Y118_DO6),
.I1(CLBLM_R_X3Y116_SLICE_X2Y116_AQ),
.I2(CLBLM_R_X11Y118_SLICE_X14Y118_AQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLM_L_X10Y116_SLICE_X12Y116_DO5),
.I5(CLBLM_R_X11Y119_SLICE_X14Y119_AO6),
.O5(CLBLM_R_X11Y118_SLICE_X14Y118_AO5),
.O6(CLBLM_R_X11Y118_SLICE_X14Y118_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y118_SLICE_X15Y118_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y118_SLICE_X15Y118_AO6),
.Q(CLBLM_R_X11Y118_SLICE_X15Y118_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y118_SLICE_X15Y118_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y118_SLICE_X15Y118_BO6),
.Q(CLBLM_R_X11Y118_SLICE_X15Y118_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y118_SLICE_X15Y118_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y118_SLICE_X15Y118_CO6),
.Q(CLBLM_R_X11Y118_SLICE_X15Y118_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hcfcccfcffcfffcfc)
  ) CLBLM_R_X11Y118_SLICE_X15Y118_DLUT (
.I0(1'b1),
.I1(CLBLM_R_X11Y120_SLICE_X14Y120_AO5),
.I2(CLBLM_L_X12Y119_SLICE_X17Y119_DO6),
.I3(CLBLM_R_X11Y118_SLICE_X14Y118_DO5),
.I4(CLBLM_L_X10Y120_SLICE_X12Y120_CQ),
.I5(CLBLM_R_X11Y118_SLICE_X15Y118_AQ),
.O5(CLBLM_R_X11Y118_SLICE_X15Y118_DO5),
.O6(CLBLM_R_X11Y118_SLICE_X15Y118_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'ha3a3afa0a0a0afa0)
  ) CLBLM_R_X11Y118_SLICE_X15Y118_CLUT (
.I0(CLBLL_L_X4Y114_SLICE_X4Y114_AQ),
.I1(CLBLM_R_X11Y119_SLICE_X14Y119_AO6),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLM_L_X10Y118_SLICE_X13Y118_BQ),
.I4(CLBLM_L_X12Y119_SLICE_X17Y119_AO5),
.I5(CLBLM_R_X11Y118_SLICE_X15Y118_CQ),
.O5(CLBLM_R_X11Y118_SLICE_X15Y118_CO5),
.O6(CLBLM_R_X11Y118_SLICE_X15Y118_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'haa00aaccaaf0aaf0)
  ) CLBLM_R_X11Y118_SLICE_X15Y118_BLUT (
.I0(CLBLM_R_X5Y116_SLICE_X7Y116_AQ),
.I1(CLBLM_R_X11Y118_SLICE_X15Y118_BQ),
.I2(CLBLM_R_X11Y117_SLICE_X14Y117_AQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLM_R_X11Y119_SLICE_X14Y119_AO6),
.I5(CLBLM_L_X12Y119_SLICE_X17Y119_AO5),
.O5(CLBLM_R_X11Y118_SLICE_X15Y118_BO5),
.O6(CLBLM_R_X11Y118_SLICE_X15Y118_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hccee0022ccee0022)
  ) CLBLM_R_X11Y118_SLICE_X15Y118_ALUT (
.I0(CLBLM_R_X11Y118_SLICE_X15Y118_DO6),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(1'b1),
.I3(CLBLM_L_X12Y120_SLICE_X17Y120_CO5),
.I4(CLBLM_L_X8Y117_SLICE_X10Y117_AQ),
.I5(1'b1),
.O5(CLBLM_R_X11Y118_SLICE_X15Y118_AO5),
.O6(CLBLM_R_X11Y118_SLICE_X15Y118_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y119_SLICE_X14Y119_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(LIOB33_X0Y77_IOB_X0Y77_I),
.D(CLBLM_L_X10Y118_SLICE_X13Y118_BQ),
.Q(CLBLM_R_X11Y119_SLICE_X14Y119_AQ),
.R(CLBLM_R_X11Y123_SLICE_X14Y123_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h2020040420a00400)
  ) CLBLM_R_X11Y119_SLICE_X14Y119_DLUT (
.I0(CLBLM_R_X11Y118_SLICE_X15Y118_AQ),
.I1(CLBLM_L_X10Y119_SLICE_X13Y119_AQ),
.I2(CLBLM_R_X11Y120_SLICE_X15Y120_AQ),
.I3(CLBLM_R_X11Y119_SLICE_X15Y119_CQ),
.I4(CLBLM_L_X12Y120_SLICE_X17Y120_AQ),
.I5(CLBLM_R_X11Y118_SLICE_X14Y118_BQ),
.O5(CLBLM_R_X11Y119_SLICE_X14Y119_DO5),
.O6(CLBLM_R_X11Y119_SLICE_X14Y119_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000fff00000eeee)
  ) CLBLM_R_X11Y119_SLICE_X14Y119_CLUT (
.I0(CLBLM_R_X5Y119_SLICE_X6Y119_AQ),
.I1(CLBLM_L_X10Y120_SLICE_X12Y120_AQ),
.I2(CLBLM_R_X11Y115_SLICE_X14Y115_DQ),
.I3(CLBLM_R_X11Y118_SLICE_X14Y118_CQ),
.I4(CLBLM_R_X3Y117_SLICE_X3Y117_BQ),
.I5(1'b1),
.O5(CLBLM_R_X11Y119_SLICE_X14Y119_CO5),
.O6(CLBLM_R_X11Y119_SLICE_X14Y119_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h9199d1dd00002222)
  ) CLBLM_R_X11Y119_SLICE_X14Y119_BLUT (
.I0(CLBLM_L_X10Y119_SLICE_X13Y119_AQ),
.I1(CLBLM_R_X11Y119_SLICE_X15Y119_CQ),
.I2(CLBLM_R_X7Y120_SLICE_X9Y120_AQ),
.I3(CLBLM_R_X13Y119_SLICE_X18Y119_CQ),
.I4(CLBLM_R_X11Y118_SLICE_X14Y118_BQ),
.I5(1'b1),
.O5(CLBLM_R_X11Y119_SLICE_X14Y119_BO5),
.O6(CLBLM_R_X11Y119_SLICE_X14Y119_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000001100000040)
  ) CLBLM_R_X11Y119_SLICE_X14Y119_ALUT (
.I0(CLBLM_L_X10Y119_SLICE_X13Y119_AQ),
.I1(CLBLM_R_X11Y119_SLICE_X15Y119_CQ),
.I2(CLBLM_L_X10Y116_SLICE_X12Y116_DO5),
.I3(CLBLM_R_X13Y119_SLICE_X18Y119_CQ),
.I4(CLBLM_R_X11Y118_SLICE_X14Y118_BQ),
.I5(1'b1),
.O5(CLBLM_R_X11Y119_SLICE_X14Y119_AO5),
.O6(CLBLM_R_X11Y119_SLICE_X14Y119_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y119_SLICE_X15Y119_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y119_SLICE_X15Y119_AO6),
.Q(CLBLM_R_X11Y119_SLICE_X15Y119_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y119_SLICE_X15Y119_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y119_SLICE_X15Y119_BO6),
.Q(CLBLM_R_X11Y119_SLICE_X15Y119_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y119_SLICE_X15Y119_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y119_SLICE_X15Y119_CO6),
.Q(CLBLM_R_X11Y119_SLICE_X15Y119_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hccefffdcccffffcc)
  ) CLBLM_R_X11Y119_SLICE_X15Y119_DLUT (
.I0(CLBLM_R_X11Y118_SLICE_X14Y118_DO5),
.I1(CLBLM_R_X11Y120_SLICE_X14Y120_AO5),
.I2(CLBLM_R_X11Y119_SLICE_X14Y119_DO6),
.I3(CLBLM_L_X12Y119_SLICE_X17Y119_DO6),
.I4(CLBLM_R_X11Y119_SLICE_X15Y119_AQ),
.I5(CLBLM_R_X11Y118_SLICE_X15Y118_BQ),
.O5(CLBLM_R_X11Y119_SLICE_X15Y119_DO5),
.O6(CLBLM_R_X11Y119_SLICE_X15Y119_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff00000c060c06)
  ) CLBLM_R_X11Y119_SLICE_X15Y119_CLUT (
.I0(CLBLM_L_X12Y120_SLICE_X16Y120_AO6),
.I1(CLBLM_R_X11Y119_SLICE_X15Y119_CQ),
.I2(RIOB33_X105Y121_IOB_X1Y121_I),
.I3(CLBLM_R_X11Y119_SLICE_X14Y119_BO6),
.I4(CLBLM_L_X8Y120_SLICE_X11Y120_AQ),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLM_R_X11Y119_SLICE_X15Y119_CO5),
.O6(CLBLM_R_X11Y119_SLICE_X15Y119_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaa3333aaaa3300)
  ) CLBLM_R_X11Y119_SLICE_X15Y119_BLUT (
.I0(CLBLM_R_X5Y118_SLICE_X6Y118_CQ),
.I1(CLBLM_L_X12Y120_SLICE_X17Y120_CO5),
.I2(1'b1),
.I3(CLBLM_L_X12Y119_SLICE_X16Y119_AO6),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(CLBLM_R_X11Y120_SLICE_X14Y120_AO5),
.O5(CLBLM_R_X11Y119_SLICE_X15Y119_BO5),
.O6(CLBLM_R_X11Y119_SLICE_X15Y119_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hff22ff2200220022)
  ) CLBLM_R_X11Y119_SLICE_X15Y119_ALUT (
.I0(CLBLM_R_X11Y119_SLICE_X15Y119_DO6),
.I1(CLBLM_L_X12Y120_SLICE_X17Y120_CO5),
.I2(1'b1),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(1'b1),
.I5(CLBLM_R_X7Y119_SLICE_X9Y119_AQ),
.O5(CLBLM_R_X11Y119_SLICE_X15Y119_AO5),
.O6(CLBLM_R_X11Y119_SLICE_X15Y119_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y120_SLICE_X14Y120_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(LIOB33_X0Y77_IOB_X0Y77_I),
.D(CLBLM_R_X11Y118_SLICE_X14Y118_BQ),
.Q(CLBLM_R_X11Y120_SLICE_X14Y120_AQ),
.R(CLBLM_R_X11Y123_SLICE_X14Y123_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h84408440cccc8440)
  ) CLBLM_R_X11Y120_SLICE_X14Y120_DLUT (
.I0(CLBLM_R_X11Y119_SLICE_X15Y119_CQ),
.I1(CLBLM_L_X12Y120_SLICE_X16Y120_AO6),
.I2(CLBLM_R_X11Y118_SLICE_X14Y118_BQ),
.I3(CLBLM_L_X10Y119_SLICE_X13Y119_AQ),
.I4(CLBLM_R_X11Y120_SLICE_X14Y120_BO5),
.I5(CLBLM_R_X11Y120_SLICE_X15Y120_BQ),
.O5(CLBLM_R_X11Y120_SLICE_X14Y120_DO5),
.O6(CLBLM_R_X11Y120_SLICE_X14Y120_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h00000f0500000e0e)
  ) CLBLM_R_X11Y120_SLICE_X14Y120_CLUT (
.I0(CLBLM_R_X7Y120_SLICE_X9Y120_AQ),
.I1(CLBLM_R_X11Y119_SLICE_X14Y119_AO5),
.I2(RIOB33_X105Y121_IOB_X1Y121_I),
.I3(CLBLM_L_X12Y119_SLICE_X17Y119_AO5),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(CLBLM_L_X10Y120_SLICE_X12Y120_DQ),
.O5(CLBLM_R_X11Y120_SLICE_X14Y120_CO5),
.O6(CLBLM_R_X11Y120_SLICE_X14Y120_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h000800000c0c0000)
  ) CLBLM_R_X11Y120_SLICE_X14Y120_BLUT (
.I0(CLBLM_L_X12Y120_SLICE_X16Y120_AO6),
.I1(CLBLM_R_X13Y119_SLICE_X18Y119_CQ),
.I2(CLBLM_R_X7Y120_SLICE_X9Y120_AQ),
.I3(CLBLM_R_X11Y120_SLICE_X15Y120_BQ),
.I4(CLBLM_R_X11Y119_SLICE_X15Y119_CQ),
.I5(1'b1),
.O5(CLBLM_R_X11Y120_SLICE_X14Y120_BO5),
.O6(CLBLM_R_X11Y120_SLICE_X14Y120_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0c0c0011a2f3aa44)
  ) CLBLM_R_X11Y120_SLICE_X14Y120_ALUT (
.I0(CLBLM_R_X11Y118_SLICE_X14Y118_BQ),
.I1(CLBLM_R_X13Y119_SLICE_X18Y119_CQ),
.I2(CLBLM_R_X7Y120_SLICE_X9Y120_AQ),
.I3(CLBLM_L_X10Y119_SLICE_X13Y119_AQ),
.I4(CLBLM_R_X11Y119_SLICE_X15Y119_CQ),
.I5(1'b1),
.O5(CLBLM_R_X11Y120_SLICE_X14Y120_AO5),
.O6(CLBLM_R_X11Y120_SLICE_X14Y120_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y120_SLICE_X15Y120_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y120_SLICE_X15Y120_AO6),
.Q(CLBLM_R_X11Y120_SLICE_X15Y120_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y120_SLICE_X15Y120_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y120_SLICE_X15Y120_BO6),
.Q(CLBLM_R_X11Y120_SLICE_X15Y120_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y120_SLICE_X15Y120_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y120_SLICE_X15Y120_CO6),
.Q(CLBLM_R_X11Y120_SLICE_X15Y120_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hddccddccd5c0ddcc)
  ) CLBLM_R_X11Y120_SLICE_X15Y120_DLUT (
.I0(CLBLM_R_X11Y120_SLICE_X15Y120_BQ),
.I1(CLBLM_R_X11Y120_SLICE_X15Y120_CQ),
.I2(CLBLM_R_X11Y121_SLICE_X15Y121_AO6),
.I3(CLBLM_L_X12Y120_SLICE_X17Y120_DO5),
.I4(CLBLM_L_X8Y119_SLICE_X10Y119_CQ),
.I5(CLBLM_L_X12Y120_SLICE_X17Y120_CO6),
.O5(CLBLM_R_X11Y120_SLICE_X15Y120_DO5),
.O6(CLBLM_R_X11Y120_SLICE_X15Y120_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaaaaaaf0fff000)
  ) CLBLM_R_X11Y120_SLICE_X15Y120_CLUT (
.I0(CLBLM_L_X12Y121_SLICE_X16Y121_AQ),
.I1(1'b1),
.I2(CLBLM_R_X7Y121_SLICE_X9Y121_DO6),
.I3(CLBLM_R_X11Y119_SLICE_X14Y119_AO6),
.I4(CLBLM_R_X11Y120_SLICE_X15Y120_DO6),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLM_R_X11Y120_SLICE_X15Y120_CO5),
.O6(CLBLM_R_X11Y120_SLICE_X15Y120_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hff55ff55ee44ae04)
  ) CLBLM_R_X11Y120_SLICE_X15Y120_BLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_R_X11Y120_SLICE_X15Y120_BQ),
.I2(CLBLM_R_X11Y120_SLICE_X14Y120_AO6),
.I3(CLBLM_R_X5Y120_SLICE_X7Y120_BQ),
.I4(CLBLM_L_X12Y120_SLICE_X17Y120_CO5),
.I5(CLBLM_R_X11Y120_SLICE_X14Y120_BO6),
.O5(CLBLM_R_X11Y120_SLICE_X15Y120_BO5),
.O6(CLBLM_R_X11Y120_SLICE_X15Y120_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hff00ff0032322323)
  ) CLBLM_R_X11Y120_SLICE_X15Y120_ALUT (
.I0(CLBLM_R_X11Y120_SLICE_X14Y120_AO5),
.I1(CLBLM_L_X12Y120_SLICE_X17Y120_CO5),
.I2(CLBLM_R_X11Y120_SLICE_X15Y120_AQ),
.I3(CLBLM_L_X10Y121_SLICE_X13Y121_CQ),
.I4(CLBLM_L_X12Y120_SLICE_X16Y120_BO6),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLM_R_X11Y120_SLICE_X15Y120_AO5),
.O6(CLBLM_R_X11Y120_SLICE_X15Y120_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y121_SLICE_X14Y121_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y121_SLICE_X14Y121_AO6),
.Q(CLBLM_R_X11Y121_SLICE_X14Y121_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hf30cf00ff30cf00f)
  ) CLBLM_R_X11Y121_SLICE_X14Y121_DLUT (
.I0(1'b1),
.I1(CLBLM_L_X8Y122_SLICE_X11Y122_DO6),
.I2(CLBLM_L_X10Y123_SLICE_X12Y123_CO6),
.I3(CLBLM_L_X10Y121_SLICE_X13Y121_CQ),
.I4(CLBLM_L_X8Y121_SLICE_X11Y121_CQ),
.I5(1'b1),
.O5(CLBLM_R_X11Y121_SLICE_X14Y121_DO5),
.O6(CLBLM_R_X11Y121_SLICE_X14Y121_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h333f3333333f3333)
  ) CLBLM_R_X11Y121_SLICE_X14Y121_CLUT (
.I0(1'b1),
.I1(RIOB33_X105Y105_IOB_X1Y105_I),
.I2(CLBLM_R_X13Y119_SLICE_X18Y119_BQ),
.I3(RIOB33_X105Y121_IOB_X1Y121_I),
.I4(CLBLM_R_X7Y114_SLICE_X8Y114_BQ),
.I5(1'b1),
.O5(CLBLM_R_X11Y121_SLICE_X14Y121_CO5),
.O6(CLBLM_R_X11Y121_SLICE_X14Y121_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h4000000000000002)
  ) CLBLM_R_X11Y121_SLICE_X14Y121_BLUT (
.I0(CLBLM_L_X10Y122_SLICE_X12Y122_CO6),
.I1(CLBLM_L_X10Y121_SLICE_X13Y121_CQ),
.I2(CLBLM_L_X10Y120_SLICE_X13Y120_BQ),
.I3(CLBLM_L_X10Y121_SLICE_X13Y121_AQ),
.I4(CLBLM_L_X10Y120_SLICE_X13Y120_AQ),
.I5(1'b1),
.O5(CLBLM_R_X11Y121_SLICE_X14Y121_BO5),
.O6(CLBLM_R_X11Y121_SLICE_X14Y121_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hcf03cf03cc00cd01)
  ) CLBLM_R_X11Y121_SLICE_X14Y121_ALUT (
.I0(CLBLM_L_X10Y119_SLICE_X13Y119_AQ),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(CLBLM_R_X11Y119_SLICE_X15Y119_CQ),
.I3(CLBLM_R_X7Y120_SLICE_X9Y120_AQ),
.I4(CLBLM_R_X11Y118_SLICE_X14Y118_BQ),
.I5(CLBLM_R_X13Y119_SLICE_X18Y119_CQ),
.O5(CLBLM_R_X11Y121_SLICE_X14Y121_AO5),
.O6(CLBLM_R_X11Y121_SLICE_X14Y121_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X11Y121_SLICE_X15Y121_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X11Y121_SLICE_X15Y121_DO5),
.O6(CLBLM_R_X11Y121_SLICE_X15Y121_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h33ff33ff33ff33ff)
  ) CLBLM_R_X11Y121_SLICE_X15Y121_CLUT (
.I0(1'b1),
.I1(CLBLM_L_X10Y120_SLICE_X13Y120_A5Q),
.I2(1'b1),
.I3(CLBLM_R_X11Y120_SLICE_X15Y120_BQ),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X11Y121_SLICE_X15Y121_CO5),
.O6(CLBLM_R_X11Y121_SLICE_X15Y121_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h000000005f5f5f5f)
  ) CLBLM_R_X11Y121_SLICE_X15Y121_BLUT (
.I0(CLBLM_R_X11Y119_SLICE_X15Y119_CQ),
.I1(1'b1),
.I2(CLBLM_R_X11Y118_SLICE_X14Y118_BQ),
.I3(1'b1),
.I4(1'b1),
.I5(CLBLM_R_X13Y119_SLICE_X18Y119_CQ),
.O5(CLBLM_R_X11Y121_SLICE_X15Y121_BO5),
.O6(CLBLM_R_X11Y121_SLICE_X15Y121_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfff05f50440ff5af)
  ) CLBLM_R_X11Y121_SLICE_X15Y121_ALUT (
.I0(CLBLM_L_X10Y119_SLICE_X13Y119_AQ),
.I1(CLBLM_R_X7Y120_SLICE_X9Y120_AQ),
.I2(CLBLM_R_X11Y118_SLICE_X14Y118_AQ),
.I3(CLBLM_R_X11Y121_SLICE_X15Y121_BO6),
.I4(CLBLM_R_X11Y119_SLICE_X15Y119_CQ),
.I5(CLBLM_R_X11Y121_SLICE_X15Y121_CO6),
.O5(CLBLM_R_X11Y121_SLICE_X15Y121_AO5),
.O6(CLBLM_R_X11Y121_SLICE_X15Y121_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y122_SLICE_X14Y122_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y122_SLICE_X14Y122_AO6),
.Q(CLBLM_R_X11Y122_SLICE_X14Y122_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X11Y122_SLICE_X14Y122_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X11Y122_SLICE_X14Y122_DO5),
.O6(CLBLM_R_X11Y122_SLICE_X14Y122_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X11Y122_SLICE_X14Y122_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X11Y122_SLICE_X14Y122_CO5),
.O6(CLBLM_R_X11Y122_SLICE_X14Y122_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000ffff000047ff)
  ) CLBLM_R_X11Y122_SLICE_X14Y122_BLUT (
.I0(CLBLM_R_X11Y123_SLICE_X14Y123_BO5),
.I1(CLBLM_L_X10Y121_SLICE_X13Y121_BQ),
.I2(CLBLM_R_X11Y123_SLICE_X14Y123_AO5),
.I3(CLBLM_L_X8Y122_SLICE_X11Y122_AQ),
.I4(CLBLM_L_X10Y123_SLICE_X12Y123_CO6),
.I5(CLBLM_L_X8Y122_SLICE_X11Y122_DO6),
.O5(CLBLM_R_X11Y122_SLICE_X14Y122_BO5),
.O6(CLBLM_R_X11Y122_SLICE_X14Y122_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hccf0ccffccf0ccf0)
  ) CLBLM_R_X11Y122_SLICE_X14Y122_ALUT (
.I0(1'b1),
.I1(CLBLM_L_X10Y122_SLICE_X13Y122_CQ),
.I2(CLBLM_R_X11Y122_SLICE_X14Y122_AQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLM_R_X7Y128_SLICE_X8Y128_AQ),
.I5(RIOB33_X105Y141_IOB_X1Y142_I),
.O5(CLBLM_R_X11Y122_SLICE_X14Y122_AO5),
.O6(CLBLM_R_X11Y122_SLICE_X14Y122_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X11Y122_SLICE_X15Y122_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X11Y122_SLICE_X15Y122_DO5),
.O6(CLBLM_R_X11Y122_SLICE_X15Y122_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X11Y122_SLICE_X15Y122_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X11Y122_SLICE_X15Y122_CO5),
.O6(CLBLM_R_X11Y122_SLICE_X15Y122_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X11Y122_SLICE_X15Y122_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X11Y122_SLICE_X15Y122_BO5),
.O6(CLBLM_R_X11Y122_SLICE_X15Y122_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X11Y122_SLICE_X15Y122_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X11Y122_SLICE_X15Y122_AO5),
.O6(CLBLM_R_X11Y122_SLICE_X15Y122_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X11Y123_SLICE_X14Y123_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X11Y123_SLICE_X14Y123_DO5),
.O6(CLBLM_R_X11Y123_SLICE_X14Y123_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h00aa00aa00ff00ff)
  ) CLBLM_R_X11Y123_SLICE_X14Y123_CLUT (
.I0(CLBLM_R_X7Y128_SLICE_X8Y128_AQ),
.I1(1'b1),
.I2(1'b1),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(1'b1),
.I5(RIOB33_X105Y141_IOB_X1Y142_I),
.O5(CLBLM_R_X11Y123_SLICE_X14Y123_CO5),
.O6(CLBLM_R_X11Y123_SLICE_X14Y123_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h8000000080808080)
  ) CLBLM_R_X11Y123_SLICE_X14Y123_BLUT (
.I0(CLBLM_L_X10Y122_SLICE_X13Y122_AQ),
.I1(CLBLM_R_X11Y121_SLICE_X14Y121_BO6),
.I2(CLBLM_L_X10Y122_SLICE_X13Y122_BQ),
.I3(CLBLM_L_X10Y122_SLICE_X13Y122_CQ),
.I4(CLBLM_L_X10Y121_SLICE_X13Y121_BQ),
.I5(1'b1),
.O5(CLBLM_R_X11Y123_SLICE_X14Y123_BO5),
.O6(CLBLM_R_X11Y123_SLICE_X14Y123_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000001010101010)
  ) CLBLM_R_X11Y123_SLICE_X14Y123_ALUT (
.I0(CLBLM_L_X10Y122_SLICE_X13Y122_AQ),
.I1(CLBLM_L_X10Y122_SLICE_X13Y122_BQ),
.I2(CLBLM_R_X11Y121_SLICE_X14Y121_BO5),
.I3(CLBLM_L_X10Y122_SLICE_X13Y122_CQ),
.I4(CLBLM_L_X10Y121_SLICE_X13Y121_BQ),
.I5(1'b1),
.O5(CLBLM_R_X11Y123_SLICE_X14Y123_AO5),
.O6(CLBLM_R_X11Y123_SLICE_X14Y123_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X11Y123_SLICE_X15Y123_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X11Y123_SLICE_X15Y123_DO5),
.O6(CLBLM_R_X11Y123_SLICE_X15Y123_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X11Y123_SLICE_X15Y123_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X11Y123_SLICE_X15Y123_CO5),
.O6(CLBLM_R_X11Y123_SLICE_X15Y123_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X11Y123_SLICE_X15Y123_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X11Y123_SLICE_X15Y123_BO5),
.O6(CLBLM_R_X11Y123_SLICE_X15Y123_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X11Y123_SLICE_X15Y123_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X11Y123_SLICE_X15Y123_AO5),
.O6(CLBLM_R_X11Y123_SLICE_X15Y123_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X11Y128_SLICE_X14Y128_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X11Y128_SLICE_X14Y128_DO5),
.O6(CLBLM_R_X11Y128_SLICE_X14Y128_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X11Y128_SLICE_X14Y128_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X11Y128_SLICE_X14Y128_CO5),
.O6(CLBLM_R_X11Y128_SLICE_X14Y128_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X11Y128_SLICE_X14Y128_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X11Y128_SLICE_X14Y128_BO5),
.O6(CLBLM_R_X11Y128_SLICE_X14Y128_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hbbaa1100ffff0f0f)
  ) CLBLM_R_X11Y128_SLICE_X14Y128_ALUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(RIOB33_X105Y105_IOB_X1Y105_I),
.I2(RIOB33_X105Y143_IOB_X1Y143_I),
.I3(CLBLM_L_X8Y119_SLICE_X11Y119_CQ),
.I4(CLBLM_R_X11Y120_SLICE_X14Y120_AQ),
.I5(1'b1),
.O5(CLBLM_R_X11Y128_SLICE_X14Y128_AO5),
.O6(CLBLM_R_X11Y128_SLICE_X14Y128_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y128_SLICE_X15Y128_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y128_SLICE_X15Y128_AO6),
.Q(CLBLM_R_X11Y128_SLICE_X15Y128_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X11Y128_SLICE_X15Y128_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X11Y128_SLICE_X15Y128_DO5),
.O6(CLBLM_R_X11Y128_SLICE_X15Y128_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X11Y128_SLICE_X15Y128_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X11Y128_SLICE_X15Y128_CO5),
.O6(CLBLM_R_X11Y128_SLICE_X15Y128_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X11Y128_SLICE_X15Y128_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X11Y128_SLICE_X15Y128_BO5),
.O6(CLBLM_R_X11Y128_SLICE_X15Y128_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaaaaaaf0f0fcfc)
  ) CLBLM_R_X11Y128_SLICE_X15Y128_ALUT (
.I0(CLBLM_L_X8Y121_SLICE_X11Y121_CQ),
.I1(RIOB33_X105Y141_IOB_X1Y142_I),
.I2(CLBLM_R_X11Y128_SLICE_X15Y128_AQ),
.I3(1'b1),
.I4(CLBLM_R_X7Y128_SLICE_X8Y128_AQ),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLM_R_X11Y128_SLICE_X15Y128_AO5),
.O6(CLBLM_R_X11Y128_SLICE_X15Y128_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X13Y119_SLICE_X18Y119_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X13Y119_SLICE_X18Y119_AO6),
.Q(CLBLM_R_X13Y119_SLICE_X18Y119_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X13Y119_SLICE_X18Y119_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X13Y119_SLICE_X18Y119_BO6),
.Q(CLBLM_R_X13Y119_SLICE_X18Y119_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X13Y119_SLICE_X18Y119_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X13Y119_SLICE_X18Y119_CO6),
.Q(CLBLM_R_X13Y119_SLICE_X18Y119_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0808000008880000)
  ) CLBLM_R_X13Y119_SLICE_X18Y119_DLUT (
.I0(CLBLM_R_X11Y118_SLICE_X15Y118_AQ),
.I1(CLBLM_L_X12Y120_SLICE_X17Y120_AQ),
.I2(CLBLM_L_X10Y119_SLICE_X13Y119_AQ),
.I3(CLBLM_R_X11Y119_SLICE_X15Y119_CQ),
.I4(CLBLM_R_X11Y120_SLICE_X15Y120_AQ),
.I5(CLBLM_R_X11Y118_SLICE_X14Y118_BQ),
.O5(CLBLM_R_X13Y119_SLICE_X18Y119_DO5),
.O6(CLBLM_R_X13Y119_SLICE_X18Y119_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hf000f606f000f303)
  ) CLBLM_R_X13Y119_SLICE_X18Y119_CLUT (
.I0(CLBLM_R_X11Y120_SLICE_X14Y120_BO6),
.I1(CLBLM_R_X13Y119_SLICE_X18Y119_CQ),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLL_L_X4Y118_SLICE_X5Y118_CQ),
.I4(RIOB33_X105Y121_IOB_X1Y121_I),
.I5(CLBLM_L_X12Y119_SLICE_X17Y119_AO6),
.O5(CLBLM_R_X13Y119_SLICE_X18Y119_CO5),
.O6(CLBLM_R_X13Y119_SLICE_X18Y119_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f088aaf0f08888)
  ) CLBLM_R_X13Y119_SLICE_X18Y119_BLUT (
.I0(RIOB33_X105Y105_IOB_X1Y105_I),
.I1(CLBLM_R_X13Y119_SLICE_X18Y119_BQ),
.I2(CLBLM_R_X11Y117_SLICE_X14Y117_BQ),
.I3(RIOB33_X105Y121_IOB_X1Y121_I),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(CLBLM_R_X7Y114_SLICE_X8Y114_BQ),
.O5(CLBLM_R_X13Y119_SLICE_X18Y119_BO5),
.O6(CLBLM_R_X13Y119_SLICE_X18Y119_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hb8b8bbb8b8b8bbb8)
  ) CLBLM_R_X13Y119_SLICE_X18Y119_ALUT (
.I0(CLBLM_L_X12Y118_SLICE_X16Y118_AQ),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(CLBLM_R_X13Y119_SLICE_X18Y119_AQ),
.I3(RIOB33_X105Y141_IOB_X1Y142_I),
.I4(CLBLM_R_X7Y128_SLICE_X8Y128_AQ),
.I5(1'b1),
.O5(CLBLM_R_X13Y119_SLICE_X18Y119_AO5),
.O6(CLBLM_R_X13Y119_SLICE_X18Y119_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X13Y119_SLICE_X19Y119_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X13Y119_SLICE_X19Y119_DO5),
.O6(CLBLM_R_X13Y119_SLICE_X19Y119_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X13Y119_SLICE_X19Y119_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X13Y119_SLICE_X19Y119_CO5),
.O6(CLBLM_R_X13Y119_SLICE_X19Y119_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X13Y119_SLICE_X19Y119_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X13Y119_SLICE_X19Y119_BO5),
.O6(CLBLM_R_X13Y119_SLICE_X19Y119_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X13Y119_SLICE_X19Y119_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X13Y119_SLICE_X19Y119_AO5),
.O6(CLBLM_R_X13Y119_SLICE_X19Y119_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X13Y120_SLICE_X18Y120_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X13Y120_SLICE_X18Y120_DO5),
.O6(CLBLM_R_X13Y120_SLICE_X18Y120_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000010101000)
  ) CLBLM_R_X13Y120_SLICE_X18Y120_CLUT (
.I0(CLBLM_R_X11Y118_SLICE_X15Y118_AQ),
.I1(CLBLM_R_X11Y120_SLICE_X15Y120_AQ),
.I2(CLBLM_L_X10Y119_SLICE_X13Y119_AQ),
.I3(CLBLM_R_X11Y119_SLICE_X15Y119_CQ),
.I4(CLBLM_R_X11Y118_SLICE_X14Y118_BQ),
.I5(CLBLM_L_X12Y120_SLICE_X17Y120_AQ),
.O5(CLBLM_R_X13Y120_SLICE_X18Y120_CO5),
.O6(CLBLM_R_X13Y120_SLICE_X18Y120_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hff7fffffffffffff)
  ) CLBLM_R_X13Y120_SLICE_X18Y120_BLUT (
.I0(CLBLM_L_X12Y120_SLICE_X17Y120_BQ),
.I1(CLBLM_R_X11Y119_SLICE_X15Y119_AQ),
.I2(CLBLM_R_X11Y118_SLICE_X15Y118_AQ),
.I3(CLBLM_L_X12Y120_SLICE_X17Y120_DO6),
.I4(CLBLM_R_X11Y120_SLICE_X15Y120_AQ),
.I5(CLBLM_L_X12Y120_SLICE_X17Y120_AQ),
.O5(CLBLM_R_X13Y120_SLICE_X18Y120_BO5),
.O6(CLBLM_R_X13Y120_SLICE_X18Y120_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffffeffffffff)
  ) CLBLM_R_X13Y120_SLICE_X18Y120_ALUT (
.I0(CLBLM_L_X12Y120_SLICE_X17Y120_BQ),
.I1(CLBLM_R_X11Y119_SLICE_X15Y119_AQ),
.I2(CLBLM_R_X11Y118_SLICE_X15Y118_AQ),
.I3(CLBLM_L_X12Y120_SLICE_X17Y120_AQ),
.I4(CLBLM_R_X11Y120_SLICE_X15Y120_AQ),
.I5(CLBLM_L_X12Y120_SLICE_X17Y120_DO6),
.O5(CLBLM_R_X13Y120_SLICE_X18Y120_AO5),
.O6(CLBLM_R_X13Y120_SLICE_X18Y120_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X13Y120_SLICE_X19Y120_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X13Y120_SLICE_X19Y120_DO5),
.O6(CLBLM_R_X13Y120_SLICE_X19Y120_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X13Y120_SLICE_X19Y120_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X13Y120_SLICE_X19Y120_CO5),
.O6(CLBLM_R_X13Y120_SLICE_X19Y120_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X13Y120_SLICE_X19Y120_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X13Y120_SLICE_X19Y120_BO5),
.O6(CLBLM_R_X13Y120_SLICE_X19Y120_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X13Y120_SLICE_X19Y120_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X13Y120_SLICE_X19Y120_AO5),
.O6(CLBLM_R_X13Y120_SLICE_X19Y120_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X37Y119_SLICE_X56Y119_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X37Y119_SLICE_X56Y119_DO5),
.O6(CLBLM_R_X37Y119_SLICE_X56Y119_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X37Y119_SLICE_X56Y119_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X37Y119_SLICE_X56Y119_CO5),
.O6(CLBLM_R_X37Y119_SLICE_X56Y119_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X37Y119_SLICE_X56Y119_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X37Y119_SLICE_X56Y119_BO5),
.O6(CLBLM_R_X37Y119_SLICE_X56Y119_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h1100110011001100)
  ) CLBLM_R_X37Y119_SLICE_X56Y119_ALUT (
.I0(RIOB33_X105Y117_IOB_X1Y118_I),
.I1(CLBLM_R_X3Y117_SLICE_X3Y117_CQ),
.I2(1'b1),
.I3(RIOB33_X105Y119_IOB_X1Y119_I),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X37Y119_SLICE_X56Y119_AO5),
.O6(CLBLM_R_X37Y119_SLICE_X56Y119_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X37Y119_SLICE_X57Y119_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X37Y119_SLICE_X57Y119_DO5),
.O6(CLBLM_R_X37Y119_SLICE_X57Y119_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X37Y119_SLICE_X57Y119_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X37Y119_SLICE_X57Y119_CO5),
.O6(CLBLM_R_X37Y119_SLICE_X57Y119_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X37Y119_SLICE_X57Y119_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X37Y119_SLICE_X57Y119_BO5),
.O6(CLBLM_R_X37Y119_SLICE_X57Y119_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X37Y119_SLICE_X57Y119_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X37Y119_SLICE_X57Y119_AO5),
.O6(CLBLM_R_X37Y119_SLICE_X57Y119_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y138_SLICE_X162Y138_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y138_SLICE_X162Y138_DO5),
.O6(CLBLM_R_X103Y138_SLICE_X162Y138_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y138_SLICE_X162Y138_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y138_SLICE_X162Y138_CO5),
.O6(CLBLM_R_X103Y138_SLICE_X162Y138_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y138_SLICE_X162Y138_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y138_SLICE_X162Y138_BO5),
.O6(CLBLM_R_X103Y138_SLICE_X162Y138_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y138_SLICE_X162Y138_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y138_SLICE_X162Y138_AO5),
.O6(CLBLM_R_X103Y138_SLICE_X162Y138_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y138_SLICE_X163Y138_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y138_SLICE_X163Y138_DO5),
.O6(CLBLM_R_X103Y138_SLICE_X163Y138_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y138_SLICE_X163Y138_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y138_SLICE_X163Y138_CO5),
.O6(CLBLM_R_X103Y138_SLICE_X163Y138_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y138_SLICE_X163Y138_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y138_SLICE_X163Y138_BO5),
.O6(CLBLM_R_X103Y138_SLICE_X163Y138_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'haa00aa0000000000)
  ) CLBLM_R_X103Y138_SLICE_X163Y138_ALUT (
.I0(RIOB33_X105Y139_IOB_X1Y139_I),
.I1(1'b1),
.I2(1'b1),
.I3(RIOB33_X105Y137_IOB_X1Y138_I),
.I4(1'b1),
.I5(RIOB33_X105Y105_IOB_X1Y105_I),
.O5(CLBLM_R_X103Y138_SLICE_X163Y138_AO5),
.O6(CLBLM_R_X103Y138_SLICE_X163Y138_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y169_SLICE_X162Y169_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y169_SLICE_X162Y169_DO5),
.O6(CLBLM_R_X103Y169_SLICE_X162Y169_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y169_SLICE_X162Y169_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y169_SLICE_X162Y169_CO5),
.O6(CLBLM_R_X103Y169_SLICE_X162Y169_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y169_SLICE_X162Y169_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y169_SLICE_X162Y169_BO5),
.O6(CLBLM_R_X103Y169_SLICE_X162Y169_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y169_SLICE_X162Y169_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y169_SLICE_X162Y169_AO5),
.O6(CLBLM_R_X103Y169_SLICE_X162Y169_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y169_SLICE_X163Y169_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y169_SLICE_X163Y169_DO5),
.O6(CLBLM_R_X103Y169_SLICE_X163Y169_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y169_SLICE_X163Y169_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y169_SLICE_X163Y169_CO5),
.O6(CLBLM_R_X103Y169_SLICE_X163Y169_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y169_SLICE_X163Y169_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y169_SLICE_X163Y169_BO5),
.O6(CLBLM_R_X103Y169_SLICE_X163Y169_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hafafafafffff0f0f)
  ) CLBLM_R_X103Y169_SLICE_X163Y169_ALUT (
.I0(CLBLM_L_X10Y114_SLICE_X12Y114_AQ),
.I1(1'b1),
.I2(RIOB33_X105Y143_IOB_X1Y143_I),
.I3(1'b1),
.I4(CLBLM_R_X11Y122_SLICE_X14Y122_AQ),
.I5(1'b1),
.O5(CLBLM_R_X103Y169_SLICE_X163Y169_AO5),
.O6(CLBLM_R_X103Y169_SLICE_X163Y169_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y172_SLICE_X162Y172_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y172_SLICE_X162Y172_DO5),
.O6(CLBLM_R_X103Y172_SLICE_X162Y172_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y172_SLICE_X162Y172_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y172_SLICE_X162Y172_CO5),
.O6(CLBLM_R_X103Y172_SLICE_X162Y172_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y172_SLICE_X162Y172_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y172_SLICE_X162Y172_BO5),
.O6(CLBLM_R_X103Y172_SLICE_X162Y172_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y172_SLICE_X162Y172_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y172_SLICE_X162Y172_AO5),
.O6(CLBLM_R_X103Y172_SLICE_X162Y172_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y172_SLICE_X163Y172_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y172_SLICE_X163Y172_DO5),
.O6(CLBLM_R_X103Y172_SLICE_X163Y172_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y172_SLICE_X163Y172_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y172_SLICE_X163Y172_CO5),
.O6(CLBLM_R_X103Y172_SLICE_X163Y172_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y172_SLICE_X163Y172_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y172_SLICE_X163Y172_BO5),
.O6(CLBLM_R_X103Y172_SLICE_X163Y172_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hff55ff55dddddddd)
  ) CLBLM_R_X103Y172_SLICE_X163Y172_ALUT (
.I0(RIOB33_X105Y143_IOB_X1Y143_I),
.I1(CLBLM_L_X8Y116_SLICE_X10Y116_AQ),
.I2(1'b1),
.I3(CLBLM_R_X13Y119_SLICE_X18Y119_AQ),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y172_SLICE_X163Y172_AO5),
.O6(CLBLM_R_X103Y172_SLICE_X163Y172_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y174_SLICE_X162Y174_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y174_SLICE_X162Y174_DO5),
.O6(CLBLM_R_X103Y174_SLICE_X162Y174_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y174_SLICE_X162Y174_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y174_SLICE_X162Y174_CO5),
.O6(CLBLM_R_X103Y174_SLICE_X162Y174_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y174_SLICE_X162Y174_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y174_SLICE_X162Y174_BO5),
.O6(CLBLM_R_X103Y174_SLICE_X162Y174_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y174_SLICE_X162Y174_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y174_SLICE_X162Y174_AO5),
.O6(CLBLM_R_X103Y174_SLICE_X162Y174_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y174_SLICE_X163Y174_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y174_SLICE_X163Y174_DO5),
.O6(CLBLM_R_X103Y174_SLICE_X163Y174_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y174_SLICE_X163Y174_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y174_SLICE_X163Y174_CO5),
.O6(CLBLM_R_X103Y174_SLICE_X163Y174_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y174_SLICE_X163Y174_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y174_SLICE_X163Y174_BO5),
.O6(CLBLM_R_X103Y174_SLICE_X163Y174_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff5555f5f5f5f5)
  ) CLBLM_R_X103Y174_SLICE_X163Y174_ALUT (
.I0(RIOB33_X105Y143_IOB_X1Y143_I),
.I1(1'b1),
.I2(CLBLM_R_X11Y128_SLICE_X15Y128_AQ),
.I3(1'b1),
.I4(CLBLM_L_X12Y115_SLICE_X16Y115_AQ),
.I5(1'b1),
.O5(CLBLM_R_X103Y174_SLICE_X163Y174_AO5),
.O6(CLBLM_R_X103Y174_SLICE_X163Y174_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y177_SLICE_X162Y177_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y177_SLICE_X162Y177_DO5),
.O6(CLBLM_R_X103Y177_SLICE_X162Y177_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y177_SLICE_X162Y177_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y177_SLICE_X162Y177_CO5),
.O6(CLBLM_R_X103Y177_SLICE_X162Y177_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y177_SLICE_X162Y177_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y177_SLICE_X162Y177_BO5),
.O6(CLBLM_R_X103Y177_SLICE_X162Y177_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y177_SLICE_X162Y177_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y177_SLICE_X162Y177_AO5),
.O6(CLBLM_R_X103Y177_SLICE_X162Y177_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y177_SLICE_X163Y177_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y177_SLICE_X163Y177_DO5),
.O6(CLBLM_R_X103Y177_SLICE_X163Y177_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y177_SLICE_X163Y177_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y177_SLICE_X163Y177_CO5),
.O6(CLBLM_R_X103Y177_SLICE_X163Y177_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y177_SLICE_X163Y177_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y177_SLICE_X163Y177_BO5),
.O6(CLBLM_R_X103Y177_SLICE_X163Y177_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff3333f3f3f3f3)
  ) CLBLM_R_X103Y177_SLICE_X163Y177_ALUT (
.I0(1'b1),
.I1(RIOB33_X105Y143_IOB_X1Y143_I),
.I2(CLBLM_R_X11Y119_SLICE_X14Y119_AQ),
.I3(1'b1),
.I4(CLBLM_L_X12Y115_SLICE_X16Y115_BQ),
.I5(1'b1),
.O5(CLBLM_R_X103Y177_SLICE_X163Y177_AO5),
.O6(CLBLM_R_X103Y177_SLICE_X163Y177_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "BUFGCTRL" *)
  BUFGCTRL #(
    .INIT_OUT(0),
    .IS_CE0_INVERTED(0),
    .IS_CE1_INVERTED(1),
    .IS_IGNORE0_INVERTED(1),
    .IS_IGNORE1_INVERTED(0),
    .IS_S0_INVERTED(0),
    .IS_S1_INVERTED(1),
    .PRESELECT_I0("TRUE"),
    .PRESELECT_I1("FALSE")
  ) CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_BUFGCTRL (
.CE0(1'b1),
.CE1(1'b1),
.I0(LIOB33_X0Y77_IOB_X0Y78_I),
.I1(1'b1),
.IGNORE0(1'b1),
.IGNORE1(1'b1),
.O(CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_O),
.S0(1'b1),
.S1(1'b1)
  );


  (* KEEP, DONT_TOUCH, BEL = "BUFHCE" *)
  BUFHCE #(
    .CE_TYPE("SYNC"),
    .INIT_OUT(0),
    .IS_CE_INVERTED(0)
  ) CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_BUFHCE (
.CE(1'b1),
.I(CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_O),
.O(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y51_IOB_X0Y51_IBUF (
.I(LIOB33_X0Y51_IOB_X0Y51_IPAD),
.O(LIOB33_X0Y51_IOB_X0Y51_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y51_IOB_X0Y52_IBUF (
.I(LIOB33_X0Y51_IOB_X0Y52_IPAD),
.O(LIOB33_X0Y51_IOB_X0Y52_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y53_IOB_X0Y53_IBUF (
.I(LIOB33_X0Y53_IOB_X0Y53_IPAD),
.O(LIOB33_X0Y53_IOB_X0Y53_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y53_IOB_X0Y54_IBUF (
.I(LIOB33_X0Y53_IOB_X0Y54_IPAD),
.O(LIOB33_X0Y53_IOB_X0Y54_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y55_IOB_X0Y55_IBUF (
.I(LIOB33_X0Y55_IOB_X0Y55_IPAD),
.O(LIOB33_X0Y55_IOB_X0Y55_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y55_IOB_X0Y56_IBUF (
.I(LIOB33_X0Y55_IOB_X0Y56_IPAD),
.O(LIOB33_X0Y55_IOB_X0Y56_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y57_IOB_X0Y57_IBUF (
.I(LIOB33_X0Y57_IOB_X0Y57_IPAD),
.O(LIOB33_X0Y57_IOB_X0Y57_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y57_IOB_X0Y58_IBUF (
.I(LIOB33_X0Y57_IOB_X0Y58_IPAD),
.O(LIOB33_X0Y57_IOB_X0Y58_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y59_IOB_X0Y59_IBUF (
.I(LIOB33_X0Y59_IOB_X0Y59_IPAD),
.O(LIOB33_X0Y59_IOB_X0Y59_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y59_IOB_X0Y60_IBUF (
.I(LIOB33_X0Y59_IOB_X0Y60_IPAD),
.O(LIOB33_X0Y59_IOB_X0Y60_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y61_IOB_X0Y61_IBUF (
.I(LIOB33_X0Y61_IOB_X0Y61_IPAD),
.O(LIOB33_X0Y61_IOB_X0Y61_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y61_IOB_X0Y62_IBUF (
.I(LIOB33_X0Y61_IOB_X0Y62_IPAD),
.O(LIOB33_X0Y61_IOB_X0Y62_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y63_IOB_X0Y63_IBUF (
.I(LIOB33_X0Y63_IOB_X0Y63_IPAD),
.O(LIOB33_X0Y63_IOB_X0Y63_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y63_IOB_X0Y64_IBUF (
.I(LIOB33_X0Y63_IOB_X0Y64_IPAD),
.O(LIOB33_X0Y63_IOB_X0Y64_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y65_IOB_X0Y65_IBUF (
.I(LIOB33_X0Y65_IOB_X0Y65_IPAD),
.O(LIOB33_X0Y65_IOB_X0Y65_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y65_IOB_X0Y66_IBUF (
.I(LIOB33_X0Y65_IOB_X0Y66_IPAD),
.O(LIOB33_X0Y65_IOB_X0Y66_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y67_IOB_X0Y67_IBUF (
.I(LIOB33_X0Y67_IOB_X0Y67_IPAD),
.O(LIOB33_X0Y67_IOB_X0Y67_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y67_IOB_X0Y68_IBUF (
.I(LIOB33_X0Y67_IOB_X0Y68_IPAD),
.O(LIOB33_X0Y67_IOB_X0Y68_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y69_IOB_X0Y69_IBUF (
.I(LIOB33_X0Y69_IOB_X0Y69_IPAD),
.O(LIOB33_X0Y69_IOB_X0Y69_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y69_IOB_X0Y70_IBUF (
.I(LIOB33_X0Y69_IOB_X0Y70_IPAD),
.O(LIOB33_X0Y69_IOB_X0Y70_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y71_IOB_X0Y71_IBUF (
.I(LIOB33_X0Y71_IOB_X0Y71_IPAD),
.O(LIOB33_X0Y71_IOB_X0Y71_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y71_IOB_X0Y72_IBUF (
.I(LIOB33_X0Y71_IOB_X0Y72_IPAD),
.O(LIOB33_X0Y71_IOB_X0Y72_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y73_IOB_X0Y73_IBUF (
.I(LIOB33_X0Y73_IOB_X0Y73_IPAD),
.O(LIOB33_X0Y73_IOB_X0Y73_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y73_IOB_X0Y74_IBUF (
.I(LIOB33_X0Y73_IOB_X0Y74_IPAD),
.O(LIOB33_X0Y73_IOB_X0Y74_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y75_IOB_X0Y75_IBUF (
.I(LIOB33_X0Y75_IOB_X0Y75_IPAD),
.O(LIOB33_X0Y75_IOB_X0Y75_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y75_IOB_X0Y76_IBUF (
.I(LIOB33_X0Y75_IOB_X0Y76_IPAD),
.O(LIOB33_X0Y75_IOB_X0Y76_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y77_IOB_X0Y77_IBUF (
.I(LIOB33_X0Y77_IOB_X0Y77_IPAD),
.O(LIOB33_X0Y77_IOB_X0Y77_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y77_IOB_X0Y78_IBUF (
.I(LIOB33_X0Y77_IOB_X0Y78_IPAD),
.O(LIOB33_X0Y77_IOB_X0Y78_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y79_IOB_X0Y79_IBUF (
.I(LIOB33_X0Y79_IOB_X0Y79_IPAD),
.O(LIOB33_X0Y79_IOB_X0Y79_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y79_IOB_X0Y80_OBUF (
.I(CLBLL_L_X2Y111_SLICE_X0Y111_AO6),
.O(LIOB33_X0Y79_IOB_X0Y80_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y101_IOB_X0Y101_OBUF (
.I(CLBLL_L_X2Y111_SLICE_X0Y111_CO6),
.O(LIOB33_X0Y101_IOB_X0Y101_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y101_IOB_X0Y102_OBUF (
.I(CLBLL_L_X2Y111_SLICE_X0Y111_AO5),
.O(LIOB33_X0Y101_IOB_X0Y102_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y103_IOB_X0Y103_OBUF (
.I(CLBLL_L_X2Y113_SLICE_X0Y113_AO6),
.O(LIOB33_X0Y103_IOB_X0Y103_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y103_IOB_X0Y104_OBUF (
.I(CLBLL_L_X2Y111_SLICE_X0Y111_CO5),
.O(LIOB33_X0Y103_IOB_X0Y104_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y105_IOB_X0Y105_OBUF (
.I(CLBLL_L_X2Y111_SLICE_X0Y111_DO6),
.O(LIOB33_X0Y105_IOB_X0Y105_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y105_IOB_X0Y106_OBUF (
.I(CLBLL_L_X2Y111_SLICE_X0Y111_DO5),
.O(LIOB33_X0Y105_IOB_X0Y106_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y107_IOB_X0Y107_OBUF (
.I(CLBLL_L_X2Y109_SLICE_X0Y109_AO6),
.O(LIOB33_X0Y107_IOB_X0Y107_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y107_IOB_X0Y108_OBUF (
.I(CLBLL_L_X2Y111_SLICE_X0Y111_BO5),
.O(LIOB33_X0Y107_IOB_X0Y108_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y109_IOB_X0Y109_OBUF (
.I(CLBLL_L_X2Y110_SLICE_X0Y110_AO6),
.O(LIOB33_X0Y109_IOB_X0Y109_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y109_IOB_X0Y110_OBUF (
.I(CLBLL_L_X2Y110_SLICE_X0Y110_AO5),
.O(LIOB33_X0Y109_IOB_X0Y110_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y111_IOB_X0Y111_OBUF (
.I(1'b0),
.O(LIOB33_X0Y111_IOB_X0Y111_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y111_IOB_X0Y112_OBUF (
.I(CLBLM_R_X11Y114_SLICE_X14Y114_D5Q),
.O(LIOB33_X0Y111_IOB_X0Y112_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y113_IOB_X0Y113_OBUF (
.I(RIOB33_X105Y121_IOB_X1Y121_I),
.O(LIOB33_X0Y113_IOB_X0Y113_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y113_IOB_X0Y114_OBUF (
.I(CLBLM_R_X5Y117_SLICE_X6Y117_DQ),
.O(LIOB33_X0Y113_IOB_X0Y114_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y115_IOB_X0Y115_OBUF (
.I(CLBLM_R_X11Y114_SLICE_X14Y114_DQ),
.O(LIOB33_X0Y115_IOB_X0Y115_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y115_IOB_X0Y116_OBUF (
.I(CLBLM_L_X8Y123_SLICE_X11Y123_AQ),
.O(LIOB33_X0Y115_IOB_X0Y116_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y117_IOB_X0Y117_OBUF (
.I(CLBLL_L_X4Y119_SLICE_X4Y119_BQ),
.O(LIOB33_X0Y117_IOB_X0Y117_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y117_IOB_X0Y118_OBUF (
.I(CLBLL_L_X4Y116_SLICE_X4Y116_CQ),
.O(LIOB33_X0Y117_IOB_X0Y118_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y119_IOB_X0Y119_OBUF (
.I(CLBLM_L_X8Y114_SLICE_X10Y114_CQ),
.O(LIOB33_X0Y119_IOB_X0Y119_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y119_IOB_X0Y120_OBUF (
.I(CLBLM_R_X3Y116_SLICE_X3Y116_A5Q),
.O(LIOB33_X0Y119_IOB_X0Y120_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y121_IOB_X0Y121_OBUF (
.I(CLBLM_L_X8Y123_SLICE_X11Y123_A5Q),
.O(LIOB33_X0Y121_IOB_X0Y121_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y121_IOB_X0Y122_OBUF (
.I(CLBLM_R_X5Y121_SLICE_X6Y121_A5Q),
.O(LIOB33_X0Y121_IOB_X0Y122_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y123_IOB_X0Y123_OBUF (
.I(CLBLM_R_X5Y117_SLICE_X6Y117_D5Q),
.O(LIOB33_X0Y123_IOB_X0Y123_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y123_IOB_X0Y124_OBUF (
.I(CLBLL_L_X4Y116_SLICE_X4Y116_C5Q),
.O(LIOB33_X0Y123_IOB_X0Y124_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y125_IOB_X0Y125_OBUF (
.I(CLBLM_R_X7Y115_SLICE_X9Y115_CQ),
.O(LIOB33_X0Y125_IOB_X0Y125_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y125_IOB_X0Y126_OBUF (
.I(CLBLM_R_X5Y124_SLICE_X6Y124_CQ),
.O(LIOB33_X0Y125_IOB_X0Y126_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y127_IOB_X0Y127_OBUF (
.I(CLBLL_L_X4Y121_SLICE_X4Y121_BQ),
.O(LIOB33_X0Y127_IOB_X0Y127_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y127_IOB_X0Y128_OBUF (
.I(CLBLL_L_X2Y117_SLICE_X0Y117_A5Q),
.O(LIOB33_X0Y127_IOB_X0Y128_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y129_IOB_X0Y129_OBUF (
.I(CLBLM_R_X3Y115_SLICE_X3Y115_CQ),
.O(LIOB33_X0Y129_IOB_X0Y129_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y129_IOB_X0Y130_OBUF (
.I(CLBLL_L_X52Y126_SLICE_X78Y126_AO6),
.O(LIOB33_X0Y129_IOB_X0Y130_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y131_IOB_X0Y131_OBUF (
.I(CLBLM_R_X7Y128_SLICE_X8Y128_AO5),
.O(LIOB33_X0Y131_IOB_X0Y131_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y131_IOB_X0Y132_OBUF (
.I(CLBLM_R_X7Y128_SLICE_X8Y128_AQ),
.O(LIOB33_X0Y131_IOB_X0Y132_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y133_IOB_X0Y133_OBUF (
.I(CLBLM_R_X7Y124_SLICE_X8Y124_A5Q),
.O(LIOB33_X0Y133_IOB_X0Y133_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y133_IOB_X0Y134_OBUF (
.I(CLBLM_R_X7Y124_SLICE_X8Y124_BQ),
.O(LIOB33_X0Y133_IOB_X0Y134_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y135_IOB_X0Y135_OBUF (
.I(CLBLL_L_X4Y123_SLICE_X4Y123_AQ),
.O(LIOB33_X0Y135_IOB_X0Y135_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y135_IOB_X0Y136_OBUF (
.I(CLBLM_R_X7Y124_SLICE_X8Y124_CQ),
.O(LIOB33_X0Y135_IOB_X0Y136_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y137_IOB_X0Y137_OBUF (
.I(CLBLM_R_X5Y124_SLICE_X6Y124_BQ),
.O(LIOB33_X0Y137_IOB_X0Y137_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y137_IOB_X0Y138_OBUF (
.I(CLBLM_R_X5Y125_SLICE_X6Y125_AQ),
.O(LIOB33_X0Y137_IOB_X0Y138_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y139_IOB_X0Y139_OBUF (
.I(CLBLM_R_X5Y124_SLICE_X6Y124_AQ),
.O(LIOB33_X0Y139_IOB_X0Y139_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y139_IOB_X0Y140_OBUF (
.I(CLBLL_L_X4Y123_SLICE_X4Y123_BQ),
.O(LIOB33_X0Y139_IOB_X0Y140_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y141_IOB_X0Y141_OBUF (
.I(CLBLM_R_X5Y123_SLICE_X6Y123_AQ),
.O(LIOB33_X0Y141_IOB_X0Y141_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y141_IOB_X0Y142_OBUF (
.I(LIOB33_X0Y53_IOB_X0Y54_I),
.O(LIOB33_X0Y141_IOB_X0Y142_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y143_IOB_X0Y143_OBUF (
.I(LIOB33_X0Y55_IOB_X0Y55_I),
.O(LIOB33_X0Y143_IOB_X0Y143_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y145_IOB_X0Y145_OBUF (
.I(LIOB33_X0Y57_IOB_X0Y58_I),
.O(LIOB33_X0Y145_IOB_X0Y145_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y145_IOB_X0Y146_OBUF (
.I(LIOB33_X0Y59_IOB_X0Y59_I),
.O(LIOB33_X0Y145_IOB_X0Y146_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y147_IOB_X0Y147_OBUF (
.I(LIOB33_X0Y71_IOB_X0Y71_I),
.O(LIOB33_X0Y147_IOB_X0Y147_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y147_IOB_X0Y148_OBUF (
.I(LIOB33_X0Y61_IOB_X0Y61_I),
.O(LIOB33_X0Y147_IOB_X0Y148_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y151_IOB_X0Y151_OBUF (
.I(LIOB33_X0Y65_IOB_X0Y65_I),
.O(LIOB33_X0Y151_IOB_X0Y151_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y151_IOB_X0Y152_OBUF (
.I(LIOB33_X0Y65_IOB_X0Y66_I),
.O(LIOB33_X0Y151_IOB_X0Y152_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y153_IOB_X0Y153_OBUF (
.I(LIOB33_X0Y67_IOB_X0Y67_I),
.O(LIOB33_X0Y153_IOB_X0Y153_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y153_IOB_X0Y154_OBUF (
.I(LIOB33_X0Y67_IOB_X0Y68_I),
.O(LIOB33_X0Y153_IOB_X0Y154_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y155_IOB_X0Y155_OBUF (
.I(LIOB33_X0Y69_IOB_X0Y70_I),
.O(LIOB33_X0Y155_IOB_X0Y155_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y155_IOB_X0Y156_OBUF (
.I(RIOB33_X105Y105_IOB_X1Y106_I),
.O(LIOB33_X0Y155_IOB_X0Y156_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y157_IOB_X0Y157_OBUF (
.I(RIOB33_X105Y115_IOB_X1Y115_I),
.O(LIOB33_X0Y157_IOB_X0Y157_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y157_IOB_X0Y158_OBUF (
.I(RIOB33_X105Y115_IOB_X1Y116_I),
.O(LIOB33_X0Y157_IOB_X0Y158_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y159_IOB_X0Y159_OBUF (
.I(RIOB33_X105Y117_IOB_X1Y117_I),
.O(LIOB33_X0Y159_IOB_X0Y159_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y159_IOB_X0Y160_OBUF (
.I(RIOB33_X105Y107_IOB_X1Y107_I),
.O(LIOB33_X0Y159_IOB_X0Y160_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y161_IOB_X0Y161_OBUF (
.I(RIOB33_X105Y107_IOB_X1Y108_I),
.O(LIOB33_X0Y161_IOB_X0Y161_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y161_IOB_X0Y162_OBUF (
.I(RIOB33_X105Y109_IOB_X1Y109_I),
.O(LIOB33_X0Y161_IOB_X0Y162_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y163_IOB_X0Y163_OBUF (
.I(RIOB33_X105Y109_IOB_X1Y110_I),
.O(LIOB33_X0Y163_IOB_X0Y163_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y163_IOB_X0Y164_OBUF (
.I(RIOB33_X105Y111_IOB_X1Y111_I),
.O(LIOB33_X0Y163_IOB_X0Y164_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y165_IOB_X0Y165_OBUF (
.I(RIOB33_X105Y111_IOB_X1Y112_I),
.O(LIOB33_X0Y165_IOB_X0Y165_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y165_IOB_X0Y166_OBUF (
.I(RIOB33_X105Y113_IOB_X1Y113_I),
.O(LIOB33_X0Y165_IOB_X0Y166_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y167_IOB_X0Y167_OBUF (
.I(RIOB33_X105Y113_IOB_X1Y114_I),
.O(LIOB33_X0Y167_IOB_X0Y167_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y167_IOB_X0Y168_OBUF (
.I(RIOB33_X105Y123_IOB_X1Y123_I),
.O(LIOB33_X0Y167_IOB_X0Y168_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y169_IOB_X0Y169_OBUF (
.I(RIOB33_X105Y121_IOB_X1Y122_I),
.O(LIOB33_X0Y169_IOB_X0Y169_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y169_IOB_X0Y170_OBUF (
.I(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.O(LIOB33_X0Y169_IOB_X0Y170_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y171_IOB_X0Y171_OBUF (
.I(LIOB33_SING_X0Y50_IOB_X0Y50_I),
.O(LIOB33_X0Y171_IOB_X0Y171_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y171_IOB_X0Y172_OBUF (
.I(CLBLM_R_X103Y138_SLICE_X163Y138_AO6),
.O(LIOB33_X0Y171_IOB_X0Y172_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y173_IOB_X0Y173_OBUF (
.I(CLBLM_L_X8Y133_SLICE_X11Y133_AO5),
.O(LIOB33_X0Y173_IOB_X0Y173_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y173_IOB_X0Y174_OBUF (
.I(CLBLM_R_X7Y151_SLICE_X8Y151_AO6),
.O(LIOB33_X0Y173_IOB_X0Y174_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y175_IOB_X0Y175_OBUF (
.I(RIOB33_X105Y127_IOB_X1Y127_I),
.O(LIOB33_X0Y175_IOB_X0Y175_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y175_IOB_X0Y176_OBUF (
.I(RIOB33_X105Y127_IOB_X1Y128_I),
.O(LIOB33_X0Y175_IOB_X0Y176_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y177_IOB_X0Y177_OBUF (
.I(RIOB33_X105Y129_IOB_X1Y129_I),
.O(LIOB33_X0Y177_IOB_X0Y177_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y177_IOB_X0Y178_OBUF (
.I(RIOB33_X105Y129_IOB_X1Y130_I),
.O(LIOB33_X0Y177_IOB_X0Y178_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y179_IOB_X0Y179_OBUF (
.I(RIOB33_X105Y131_IOB_X1Y131_I),
.O(LIOB33_X0Y179_IOB_X0Y179_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y179_IOB_X0Y180_OBUF (
.I(RIOB33_X105Y131_IOB_X1Y132_I),
.O(LIOB33_X0Y179_IOB_X0Y180_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y181_IOB_X0Y181_OBUF (
.I(RIOB33_X105Y133_IOB_X1Y133_I),
.O(LIOB33_X0Y181_IOB_X0Y181_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y181_IOB_X0Y182_OBUF (
.I(RIOB33_X105Y133_IOB_X1Y134_I),
.O(LIOB33_X0Y181_IOB_X0Y182_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y183_IOB_X0Y183_OBUF (
.I(RIOB33_X105Y135_IOB_X1Y135_I),
.O(LIOB33_X0Y183_IOB_X0Y183_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y183_IOB_X0Y184_OBUF (
.I(RIOB33_X105Y135_IOB_X1Y136_I),
.O(LIOB33_X0Y183_IOB_X0Y184_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y185_IOB_X0Y185_OBUF (
.I(RIOB33_X105Y137_IOB_X1Y137_I),
.O(LIOB33_X0Y185_IOB_X0Y185_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y185_IOB_X0Y186_OBUF (
.I(RIOB33_X105Y143_IOB_X1Y143_I),
.O(LIOB33_X0Y185_IOB_X0Y186_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y187_IOB_X0Y187_OBUF (
.I(RIOB33_X105Y143_IOB_X1Y144_I),
.O(LIOB33_X0Y187_IOB_X0Y187_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y187_IOB_X0Y188_OBUF (
.I(RIOB33_X105Y145_IOB_X1Y145_I),
.O(LIOB33_X0Y187_IOB_X0Y188_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y189_IOB_X0Y189_OBUF (
.I(RIOB33_X105Y145_IOB_X1Y146_I),
.O(LIOB33_X0Y189_IOB_X0Y189_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y189_IOB_X0Y190_OBUF (
.I(RIOB33_X105Y147_IOB_X1Y147_I),
.O(LIOB33_X0Y189_IOB_X0Y190_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y191_IOB_X0Y191_OBUF (
.I(RIOB33_X105Y147_IOB_X1Y148_I),
.O(LIOB33_X0Y191_IOB_X0Y191_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y191_IOB_X0Y192_OBUF (
.I(LIOB33_X0Y51_IOB_X0Y52_I),
.O(LIOB33_X0Y191_IOB_X0Y192_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y193_IOB_X0Y193_OBUF (
.I(LIOB33_X0Y55_IOB_X0Y56_I),
.O(LIOB33_X0Y193_IOB_X0Y193_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y193_IOB_X0Y194_OBUF (
.I(LIOB33_X0Y59_IOB_X0Y60_I),
.O(LIOB33_X0Y193_IOB_X0Y194_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y195_IOB_X0Y195_OBUF (
.I(LIOB33_X0Y63_IOB_X0Y64_I),
.O(LIOB33_X0Y195_IOB_X0Y195_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y195_IOB_X0Y196_OBUF (
.I(LIOB33_X0Y69_IOB_X0Y69_I),
.O(LIOB33_X0Y195_IOB_X0Y196_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y197_IOB_X0Y197_OBUF (
.I(LIOB33_X0Y71_IOB_X0Y72_I),
.O(LIOB33_X0Y197_IOB_X0Y197_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y197_IOB_X0Y198_OBUF (
.I(LIOB33_X0Y73_IOB_X0Y73_I),
.O(LIOB33_X0Y197_IOB_X0Y198_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_SING_X0Y50_IOB_X0Y50_IBUF (
.I(LIOB33_SING_X0Y50_IOB_X0Y50_IPAD),
.O(LIOB33_SING_X0Y50_IOB_X0Y50_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_SING_X0Y100_IOB_X0Y100_OBUF (
.I(CLBLL_L_X2Y111_SLICE_X0Y111_BO6),
.O(LIOB33_SING_X0Y100_IOB_X0Y100_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_SING_X0Y149_IOB_X0Y149_OBUF (
.I(LIOB33_X0Y61_IOB_X0Y62_I),
.O(LIOB33_SING_X0Y149_IOB_X0Y149_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_SING_X0Y150_IOB_X0Y150_OBUF (
.I(LIOB33_X0Y63_IOB_X0Y63_I),
.O(LIOB33_SING_X0Y150_IOB_X0Y150_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_SING_X0Y199_IOB_X0Y199_OBUF (
.I(LIOB33_X0Y73_IOB_X0Y74_I),
.O(LIOB33_SING_X0Y199_IOB_X0Y199_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y101_IOB_X1Y101_IBUF (
.I(RIOB33_X105Y101_IOB_X1Y101_IPAD),
.O(RIOB33_X105Y101_IOB_X1Y101_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y101_IOB_X1Y102_IBUF (
.I(RIOB33_X105Y101_IOB_X1Y102_IPAD),
.O(RIOB33_X105Y101_IOB_X1Y102_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y103_IOB_X1Y103_IBUF (
.I(RIOB33_X105Y103_IOB_X1Y103_IPAD),
.O(RIOB33_X105Y103_IOB_X1Y103_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y103_IOB_X1Y104_IBUF (
.I(RIOB33_X105Y103_IOB_X1Y104_IPAD),
.O(RIOB33_X105Y103_IOB_X1Y104_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y105_IOB_X1Y105_IBUF (
.I(RIOB33_X105Y105_IOB_X1Y105_IPAD),
.O(RIOB33_X105Y105_IOB_X1Y105_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y105_IOB_X1Y106_IBUF (
.I(RIOB33_X105Y105_IOB_X1Y106_IPAD),
.O(RIOB33_X105Y105_IOB_X1Y106_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y107_IOB_X1Y107_IBUF (
.I(RIOB33_X105Y107_IOB_X1Y107_IPAD),
.O(RIOB33_X105Y107_IOB_X1Y107_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y107_IOB_X1Y108_IBUF (
.I(RIOB33_X105Y107_IOB_X1Y108_IPAD),
.O(RIOB33_X105Y107_IOB_X1Y108_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y109_IOB_X1Y109_IBUF (
.I(RIOB33_X105Y109_IOB_X1Y109_IPAD),
.O(RIOB33_X105Y109_IOB_X1Y109_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y109_IOB_X1Y110_IBUF (
.I(RIOB33_X105Y109_IOB_X1Y110_IPAD),
.O(RIOB33_X105Y109_IOB_X1Y110_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y111_IOB_X1Y111_IBUF (
.I(RIOB33_X105Y111_IOB_X1Y111_IPAD),
.O(RIOB33_X105Y111_IOB_X1Y111_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y111_IOB_X1Y112_IBUF (
.I(RIOB33_X105Y111_IOB_X1Y112_IPAD),
.O(RIOB33_X105Y111_IOB_X1Y112_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y113_IOB_X1Y113_IBUF (
.I(RIOB33_X105Y113_IOB_X1Y113_IPAD),
.O(RIOB33_X105Y113_IOB_X1Y113_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y113_IOB_X1Y114_IBUF (
.I(RIOB33_X105Y113_IOB_X1Y114_IPAD),
.O(RIOB33_X105Y113_IOB_X1Y114_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y115_IOB_X1Y115_IBUF (
.I(RIOB33_X105Y115_IOB_X1Y115_IPAD),
.O(RIOB33_X105Y115_IOB_X1Y115_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y115_IOB_X1Y116_IBUF (
.I(RIOB33_X105Y115_IOB_X1Y116_IPAD),
.O(RIOB33_X105Y115_IOB_X1Y116_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y117_IOB_X1Y117_IBUF (
.I(RIOB33_X105Y117_IOB_X1Y117_IPAD),
.O(RIOB33_X105Y117_IOB_X1Y117_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y117_IOB_X1Y118_IBUF (
.I(RIOB33_X105Y117_IOB_X1Y118_IPAD),
.O(RIOB33_X105Y117_IOB_X1Y118_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y119_IOB_X1Y119_IBUF (
.I(RIOB33_X105Y119_IOB_X1Y119_IPAD),
.O(RIOB33_X105Y119_IOB_X1Y119_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y119_IOB_X1Y120_IBUF (
.I(RIOB33_X105Y119_IOB_X1Y120_IPAD),
.O(RIOB33_X105Y119_IOB_X1Y120_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y121_IOB_X1Y121_IBUF (
.I(RIOB33_X105Y121_IOB_X1Y121_IPAD),
.O(RIOB33_X105Y121_IOB_X1Y121_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y121_IOB_X1Y122_IBUF (
.I(RIOB33_X105Y121_IOB_X1Y122_IPAD),
.O(RIOB33_X105Y121_IOB_X1Y122_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y123_IOB_X1Y123_IBUF (
.I(RIOB33_X105Y123_IOB_X1Y123_IPAD),
.O(RIOB33_X105Y123_IOB_X1Y123_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y123_IOB_X1Y124_IBUF (
.I(RIOB33_X105Y123_IOB_X1Y124_IPAD),
.O(RIOB33_X105Y123_IOB_X1Y124_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y125_IOB_X1Y125_IBUF (
.I(RIOB33_X105Y125_IOB_X1Y125_IPAD),
.O(RIOB33_X105Y125_IOB_X1Y125_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y125_IOB_X1Y126_IBUF (
.I(RIOB33_X105Y125_IOB_X1Y126_IPAD),
.O(RIOB33_X105Y125_IOB_X1Y126_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y127_IOB_X1Y127_IBUF (
.I(RIOB33_X105Y127_IOB_X1Y127_IPAD),
.O(RIOB33_X105Y127_IOB_X1Y127_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y127_IOB_X1Y128_IBUF (
.I(RIOB33_X105Y127_IOB_X1Y128_IPAD),
.O(RIOB33_X105Y127_IOB_X1Y128_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y129_IOB_X1Y129_IBUF (
.I(RIOB33_X105Y129_IOB_X1Y129_IPAD),
.O(RIOB33_X105Y129_IOB_X1Y129_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y129_IOB_X1Y130_IBUF (
.I(RIOB33_X105Y129_IOB_X1Y130_IPAD),
.O(RIOB33_X105Y129_IOB_X1Y130_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y131_IOB_X1Y131_IBUF (
.I(RIOB33_X105Y131_IOB_X1Y131_IPAD),
.O(RIOB33_X105Y131_IOB_X1Y131_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y131_IOB_X1Y132_IBUF (
.I(RIOB33_X105Y131_IOB_X1Y132_IPAD),
.O(RIOB33_X105Y131_IOB_X1Y132_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y133_IOB_X1Y133_IBUF (
.I(RIOB33_X105Y133_IOB_X1Y133_IPAD),
.O(RIOB33_X105Y133_IOB_X1Y133_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y133_IOB_X1Y134_IBUF (
.I(RIOB33_X105Y133_IOB_X1Y134_IPAD),
.O(RIOB33_X105Y133_IOB_X1Y134_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y135_IOB_X1Y135_IBUF (
.I(RIOB33_X105Y135_IOB_X1Y135_IPAD),
.O(RIOB33_X105Y135_IOB_X1Y135_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y135_IOB_X1Y136_IBUF (
.I(RIOB33_X105Y135_IOB_X1Y136_IPAD),
.O(RIOB33_X105Y135_IOB_X1Y136_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y137_IOB_X1Y137_IBUF (
.I(RIOB33_X105Y137_IOB_X1Y137_IPAD),
.O(RIOB33_X105Y137_IOB_X1Y137_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y137_IOB_X1Y138_IBUF (
.I(RIOB33_X105Y137_IOB_X1Y138_IPAD),
.O(RIOB33_X105Y137_IOB_X1Y138_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y139_IOB_X1Y139_IBUF (
.I(RIOB33_X105Y139_IOB_X1Y139_IPAD),
.O(RIOB33_X105Y139_IOB_X1Y139_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y139_IOB_X1Y140_IBUF (
.I(RIOB33_X105Y139_IOB_X1Y140_IPAD),
.O(RIOB33_X105Y139_IOB_X1Y140_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y141_IOB_X1Y141_IBUF (
.I(RIOB33_X105Y141_IOB_X1Y141_IPAD),
.O(RIOB33_X105Y141_IOB_X1Y141_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y141_IOB_X1Y142_IBUF (
.I(RIOB33_X105Y141_IOB_X1Y142_IPAD),
.O(RIOB33_X105Y141_IOB_X1Y142_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y143_IOB_X1Y143_IBUF (
.I(RIOB33_X105Y143_IOB_X1Y143_IPAD),
.O(RIOB33_X105Y143_IOB_X1Y143_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y143_IOB_X1Y144_IBUF (
.I(RIOB33_X105Y143_IOB_X1Y144_IPAD),
.O(RIOB33_X105Y143_IOB_X1Y144_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y145_IOB_X1Y145_IBUF (
.I(RIOB33_X105Y145_IOB_X1Y145_IPAD),
.O(RIOB33_X105Y145_IOB_X1Y145_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y145_IOB_X1Y146_IBUF (
.I(RIOB33_X105Y145_IOB_X1Y146_IPAD),
.O(RIOB33_X105Y145_IOB_X1Y146_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y147_IOB_X1Y147_IBUF (
.I(RIOB33_X105Y147_IOB_X1Y147_IPAD),
.O(RIOB33_X105Y147_IOB_X1Y147_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y147_IOB_X1Y148_IBUF (
.I(RIOB33_X105Y147_IOB_X1Y148_IPAD),
.O(RIOB33_X105Y147_IOB_X1Y148_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y151_IOB_X1Y151_OBUF (
.I(LIOB33_X0Y75_IOB_X0Y76_I),
.O(RIOB33_X105Y151_IOB_X1Y151_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y151_IOB_X1Y152_OBUF (
.I(RIOB33_SING_X105Y100_IOB_X1Y100_I),
.O(RIOB33_X105Y151_IOB_X1Y152_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y153_IOB_X1Y153_OBUF (
.I(RIOB33_X105Y101_IOB_X1Y101_I),
.O(RIOB33_X105Y153_IOB_X1Y153_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y153_IOB_X1Y154_OBUF (
.I(RIOB33_X105Y101_IOB_X1Y102_I),
.O(RIOB33_X105Y153_IOB_X1Y154_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y155_IOB_X1Y155_OBUF (
.I(RIOB33_X105Y103_IOB_X1Y103_I),
.O(RIOB33_X105Y155_IOB_X1Y155_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y155_IOB_X1Y156_OBUF (
.I(RIOB33_X105Y103_IOB_X1Y104_I),
.O(RIOB33_X105Y155_IOB_X1Y156_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y157_IOB_X1Y157_OBUF (
.I(RIOB33_X105Y125_IOB_X1Y126_I),
.O(RIOB33_X105Y157_IOB_X1Y157_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y157_IOB_X1Y158_OBUF (
.I(CLBLM_R_X37Y119_SLICE_X56Y119_AO6),
.O(RIOB33_X105Y157_IOB_X1Y158_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y159_IOB_X1Y159_OBUF (
.I(CLBLM_R_X11Y113_SLICE_X15Y113_DO6),
.O(RIOB33_X105Y159_IOB_X1Y159_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y159_IOB_X1Y160_OBUF (
.I(CLBLM_R_X11Y119_SLICE_X14Y119_CO6),
.O(RIOB33_X105Y159_IOB_X1Y160_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y161_IOB_X1Y161_OBUF (
.I(CLBLM_R_X11Y119_SLICE_X14Y119_CO5),
.O(RIOB33_X105Y161_IOB_X1Y161_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y161_IOB_X1Y162_OBUF (
.I(CLBLM_R_X11Y117_SLICE_X14Y117_DO6),
.O(RIOB33_X105Y161_IOB_X1Y162_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y163_IOB_X1Y163_OBUF (
.I(CLBLM_R_X11Y117_SLICE_X14Y117_DO5),
.O(RIOB33_X105Y163_IOB_X1Y163_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y163_IOB_X1Y164_OBUF (
.I(CLBLM_R_X7Y119_SLICE_X9Y119_DO5),
.O(RIOB33_X105Y163_IOB_X1Y164_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y165_IOB_X1Y165_OBUF (
.I(RIOB33_X105Y125_IOB_X1Y125_I),
.O(RIOB33_X105Y165_IOB_X1Y165_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y165_IOB_X1Y166_OBUF (
.I(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.O(RIOB33_X105Y165_IOB_X1Y166_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y167_IOB_X1Y167_OBUF (
.I(LIOB33_SING_X0Y50_IOB_X0Y50_I),
.O(RIOB33_X105Y167_IOB_X1Y167_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y167_IOB_X1Y168_OBUF (
.I(CLBLM_R_X7Y151_SLICE_X8Y151_AO6),
.O(RIOB33_X105Y167_IOB_X1Y168_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y169_IOB_X1Y169_OBUF (
.I(CLBLM_R_X103Y169_SLICE_X163Y169_AO6),
.O(RIOB33_X105Y169_IOB_X1Y169_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y169_IOB_X1Y170_OBUF (
.I(CLBLM_R_X103Y169_SLICE_X163Y169_AO5),
.O(RIOB33_X105Y169_IOB_X1Y170_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y171_IOB_X1Y171_OBUF (
.I(CLBLM_L_X8Y128_SLICE_X10Y128_AO5),
.O(RIOB33_X105Y171_IOB_X1Y171_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y171_IOB_X1Y172_OBUF (
.I(CLBLM_R_X103Y172_SLICE_X163Y172_AO6),
.O(RIOB33_X105Y171_IOB_X1Y172_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y173_IOB_X1Y173_OBUF (
.I(CLBLM_R_X103Y172_SLICE_X163Y172_AO5),
.O(RIOB33_X105Y173_IOB_X1Y173_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y173_IOB_X1Y174_OBUF (
.I(CLBLM_R_X103Y174_SLICE_X163Y174_AO6),
.O(RIOB33_X105Y173_IOB_X1Y174_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y175_IOB_X1Y175_OBUF (
.I(CLBLM_L_X10Y128_SLICE_X13Y128_AO6),
.O(RIOB33_X105Y175_IOB_X1Y175_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y175_IOB_X1Y176_OBUF (
.I(CLBLM_R_X103Y174_SLICE_X163Y174_AO5),
.O(RIOB33_X105Y175_IOB_X1Y176_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y177_IOB_X1Y177_OBUF (
.I(CLBLM_R_X103Y177_SLICE_X163Y177_AO6),
.O(RIOB33_X105Y177_IOB_X1Y177_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y177_IOB_X1Y178_OBUF (
.I(CLBLM_R_X103Y177_SLICE_X163Y177_AO5),
.O(RIOB33_X105Y177_IOB_X1Y178_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y179_IOB_X1Y179_OBUF (
.I(CLBLM_R_X11Y128_SLICE_X14Y128_AO5),
.O(RIOB33_X105Y179_IOB_X1Y179_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y179_IOB_X1Y180_OBUF (
.I(CLBLM_R_X11Y113_SLICE_X15Y113_DO6),
.O(RIOB33_X105Y179_IOB_X1Y180_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y181_IOB_X1Y181_OBUF (
.I(CLBLM_R_X11Y119_SLICE_X14Y119_CO6),
.O(RIOB33_X105Y181_IOB_X1Y181_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y181_IOB_X1Y182_OBUF (
.I(CLBLM_R_X11Y119_SLICE_X14Y119_CO5),
.O(RIOB33_X105Y181_IOB_X1Y182_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y183_IOB_X1Y183_OBUF (
.I(CLBLM_R_X11Y117_SLICE_X14Y117_DO6),
.O(RIOB33_X105Y183_IOB_X1Y183_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y183_IOB_X1Y184_OBUF (
.I(CLBLM_R_X11Y117_SLICE_X14Y117_DO5),
.O(RIOB33_X105Y183_IOB_X1Y184_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y185_IOB_X1Y185_OBUF (
.I(CLBLM_R_X7Y119_SLICE_X9Y119_DO5),
.O(RIOB33_X105Y185_IOB_X1Y185_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y185_IOB_X1Y186_OBUF (
.I(CLBLM_L_X12Y115_SLICE_X16Y115_BQ),
.O(RIOB33_X105Y185_IOB_X1Y186_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y187_IOB_X1Y187_OBUF (
.I(CLBLM_L_X10Y114_SLICE_X12Y114_AQ),
.O(RIOB33_X105Y187_IOB_X1Y187_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y187_IOB_X1Y188_OBUF (
.I(CLBLM_R_X11Y122_SLICE_X14Y122_AQ),
.O(RIOB33_X105Y187_IOB_X1Y188_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y189_IOB_X1Y189_OBUF (
.I(CLBLM_L_X8Y122_SLICE_X10Y122_AQ),
.O(RIOB33_X105Y189_IOB_X1Y189_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y189_IOB_X1Y190_OBUF (
.I(CLBLM_R_X13Y119_SLICE_X18Y119_AQ),
.O(RIOB33_X105Y189_IOB_X1Y190_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y191_IOB_X1Y191_OBUF (
.I(CLBLM_L_X8Y116_SLICE_X10Y116_AQ),
.O(RIOB33_X105Y191_IOB_X1Y191_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y191_IOB_X1Y192_OBUF (
.I(CLBLM_L_X12Y115_SLICE_X16Y115_AQ),
.O(RIOB33_X105Y191_IOB_X1Y192_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y193_IOB_X1Y193_OBUF (
.I(CLBLM_L_X10Y124_SLICE_X13Y124_AQ),
.O(RIOB33_X105Y193_IOB_X1Y193_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y193_IOB_X1Y194_OBUF (
.I(CLBLM_R_X11Y128_SLICE_X15Y128_AQ),
.O(RIOB33_X105Y193_IOB_X1Y194_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y195_IOB_X1Y195_OBUF (
.I(CLBLM_R_X11Y119_SLICE_X14Y119_AQ),
.O(RIOB33_X105Y195_IOB_X1Y195_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y195_IOB_X1Y196_OBUF (
.I(CLBLM_R_X11Y120_SLICE_X14Y120_AQ),
.O(RIOB33_X105Y195_IOB_X1Y196_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y197_IOB_X1Y197_OBUF (
.I(CLBLM_L_X8Y122_SLICE_X10Y122_BO5),
.O(RIOB33_X105Y197_IOB_X1Y197_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y197_IOB_X1Y198_OBUF (
.I(CLBLM_L_X8Y122_SLICE_X10Y122_BO5),
.O(RIOB33_X105Y197_IOB_X1Y198_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_SING_X105Y100_IOB_X1Y100_IBUF (
.I(RIOB33_SING_X105Y100_IOB_X1Y100_IPAD),
.O(RIOB33_SING_X105Y100_IOB_X1Y100_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_SING_X105Y149_IOB_X1Y149_IBUF (
.I(RIOB33_SING_X105Y149_IOB_X1Y149_IPAD),
.O(RIOB33_SING_X105Y149_IOB_X1Y149_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_SING_X105Y150_IOB_X1Y150_OBUF (
.I(LIOB33_X0Y75_IOB_X0Y75_I),
.O(RIOB33_SING_X105Y150_IOB_X1Y150_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_SING_X105Y199_IOB_X1Y199_OBUF (
.I(CLBLM_R_X11Y128_SLICE_X15Y128_AQ),
.O(RIOB33_SING_X105Y199_IOB_X1Y199_OPAD)
  );
  assign CLBLL_L_X2Y109_SLICE_X0Y109_A = CLBLL_L_X2Y109_SLICE_X0Y109_AO6;
  assign CLBLL_L_X2Y109_SLICE_X0Y109_B = CLBLL_L_X2Y109_SLICE_X0Y109_BO6;
  assign CLBLL_L_X2Y109_SLICE_X0Y109_C = CLBLL_L_X2Y109_SLICE_X0Y109_CO6;
  assign CLBLL_L_X2Y109_SLICE_X0Y109_D = CLBLL_L_X2Y109_SLICE_X0Y109_DO6;
  assign CLBLL_L_X2Y109_SLICE_X1Y109_A = CLBLL_L_X2Y109_SLICE_X1Y109_AO6;
  assign CLBLL_L_X2Y109_SLICE_X1Y109_B = CLBLL_L_X2Y109_SLICE_X1Y109_BO6;
  assign CLBLL_L_X2Y109_SLICE_X1Y109_C = CLBLL_L_X2Y109_SLICE_X1Y109_CO6;
  assign CLBLL_L_X2Y109_SLICE_X1Y109_D = CLBLL_L_X2Y109_SLICE_X1Y109_DO6;
  assign CLBLL_L_X2Y110_SLICE_X0Y110_A = CLBLL_L_X2Y110_SLICE_X0Y110_AO6;
  assign CLBLL_L_X2Y110_SLICE_X0Y110_B = CLBLL_L_X2Y110_SLICE_X0Y110_BO6;
  assign CLBLL_L_X2Y110_SLICE_X0Y110_C = CLBLL_L_X2Y110_SLICE_X0Y110_CO6;
  assign CLBLL_L_X2Y110_SLICE_X0Y110_D = CLBLL_L_X2Y110_SLICE_X0Y110_DO6;
  assign CLBLL_L_X2Y110_SLICE_X0Y110_AMUX = CLBLL_L_X2Y110_SLICE_X0Y110_AO5;
  assign CLBLL_L_X2Y110_SLICE_X1Y110_A = CLBLL_L_X2Y110_SLICE_X1Y110_AO6;
  assign CLBLL_L_X2Y110_SLICE_X1Y110_B = CLBLL_L_X2Y110_SLICE_X1Y110_BO6;
  assign CLBLL_L_X2Y110_SLICE_X1Y110_C = CLBLL_L_X2Y110_SLICE_X1Y110_CO6;
  assign CLBLL_L_X2Y110_SLICE_X1Y110_D = CLBLL_L_X2Y110_SLICE_X1Y110_DO6;
  assign CLBLL_L_X2Y111_SLICE_X0Y111_A = CLBLL_L_X2Y111_SLICE_X0Y111_AO6;
  assign CLBLL_L_X2Y111_SLICE_X0Y111_B = CLBLL_L_X2Y111_SLICE_X0Y111_BO6;
  assign CLBLL_L_X2Y111_SLICE_X0Y111_C = CLBLL_L_X2Y111_SLICE_X0Y111_CO6;
  assign CLBLL_L_X2Y111_SLICE_X0Y111_D = CLBLL_L_X2Y111_SLICE_X0Y111_DO6;
  assign CLBLL_L_X2Y111_SLICE_X0Y111_AMUX = CLBLL_L_X2Y111_SLICE_X0Y111_AO5;
  assign CLBLL_L_X2Y111_SLICE_X0Y111_BMUX = CLBLL_L_X2Y111_SLICE_X0Y111_BO5;
  assign CLBLL_L_X2Y111_SLICE_X0Y111_CMUX = CLBLL_L_X2Y111_SLICE_X0Y111_CO5;
  assign CLBLL_L_X2Y111_SLICE_X0Y111_DMUX = CLBLL_L_X2Y111_SLICE_X0Y111_DO5;
  assign CLBLL_L_X2Y111_SLICE_X1Y111_A = CLBLL_L_X2Y111_SLICE_X1Y111_AO6;
  assign CLBLL_L_X2Y111_SLICE_X1Y111_B = CLBLL_L_X2Y111_SLICE_X1Y111_BO6;
  assign CLBLL_L_X2Y111_SLICE_X1Y111_C = CLBLL_L_X2Y111_SLICE_X1Y111_CO6;
  assign CLBLL_L_X2Y111_SLICE_X1Y111_D = CLBLL_L_X2Y111_SLICE_X1Y111_DO6;
  assign CLBLL_L_X2Y112_SLICE_X0Y112_A = CLBLL_L_X2Y112_SLICE_X0Y112_AO6;
  assign CLBLL_L_X2Y112_SLICE_X0Y112_B = CLBLL_L_X2Y112_SLICE_X0Y112_BO6;
  assign CLBLL_L_X2Y112_SLICE_X0Y112_C = CLBLL_L_X2Y112_SLICE_X0Y112_CO6;
  assign CLBLL_L_X2Y112_SLICE_X0Y112_D = CLBLL_L_X2Y112_SLICE_X0Y112_DO6;
  assign CLBLL_L_X2Y112_SLICE_X1Y112_A = CLBLL_L_X2Y112_SLICE_X1Y112_AO6;
  assign CLBLL_L_X2Y112_SLICE_X1Y112_B = CLBLL_L_X2Y112_SLICE_X1Y112_BO6;
  assign CLBLL_L_X2Y112_SLICE_X1Y112_C = CLBLL_L_X2Y112_SLICE_X1Y112_CO6;
  assign CLBLL_L_X2Y112_SLICE_X1Y112_D = CLBLL_L_X2Y112_SLICE_X1Y112_DO6;
  assign CLBLL_L_X2Y112_SLICE_X1Y112_AMUX = CLBLL_L_X2Y112_SLICE_X1Y112_A5Q;
  assign CLBLL_L_X2Y112_SLICE_X1Y112_CMUX = CLBLL_L_X2Y112_SLICE_X1Y112_CO5;
  assign CLBLL_L_X2Y113_SLICE_X0Y113_A = CLBLL_L_X2Y113_SLICE_X0Y113_AO6;
  assign CLBLL_L_X2Y113_SLICE_X0Y113_B = CLBLL_L_X2Y113_SLICE_X0Y113_BO6;
  assign CLBLL_L_X2Y113_SLICE_X0Y113_C = CLBLL_L_X2Y113_SLICE_X0Y113_CO6;
  assign CLBLL_L_X2Y113_SLICE_X0Y113_D = CLBLL_L_X2Y113_SLICE_X0Y113_DO6;
  assign CLBLL_L_X2Y113_SLICE_X0Y113_AMUX = CLBLL_L_X2Y113_SLICE_X0Y113_AO5;
  assign CLBLL_L_X2Y113_SLICE_X1Y113_A = CLBLL_L_X2Y113_SLICE_X1Y113_AO6;
  assign CLBLL_L_X2Y113_SLICE_X1Y113_B = CLBLL_L_X2Y113_SLICE_X1Y113_BO6;
  assign CLBLL_L_X2Y113_SLICE_X1Y113_C = CLBLL_L_X2Y113_SLICE_X1Y113_CO6;
  assign CLBLL_L_X2Y113_SLICE_X1Y113_D = CLBLL_L_X2Y113_SLICE_X1Y113_DO6;
  assign CLBLL_L_X2Y113_SLICE_X1Y113_CMUX = CLBLL_L_X2Y113_SLICE_X1Y113_C5Q;
  assign CLBLL_L_X2Y114_SLICE_X0Y114_A = CLBLL_L_X2Y114_SLICE_X0Y114_AO6;
  assign CLBLL_L_X2Y114_SLICE_X0Y114_B = CLBLL_L_X2Y114_SLICE_X0Y114_BO6;
  assign CLBLL_L_X2Y114_SLICE_X0Y114_C = CLBLL_L_X2Y114_SLICE_X0Y114_CO6;
  assign CLBLL_L_X2Y114_SLICE_X0Y114_D = CLBLL_L_X2Y114_SLICE_X0Y114_DO6;
  assign CLBLL_L_X2Y114_SLICE_X1Y114_A = CLBLL_L_X2Y114_SLICE_X1Y114_AO6;
  assign CLBLL_L_X2Y114_SLICE_X1Y114_B = CLBLL_L_X2Y114_SLICE_X1Y114_BO6;
  assign CLBLL_L_X2Y114_SLICE_X1Y114_C = CLBLL_L_X2Y114_SLICE_X1Y114_CO6;
  assign CLBLL_L_X2Y114_SLICE_X1Y114_D = CLBLL_L_X2Y114_SLICE_X1Y114_DO6;
  assign CLBLL_L_X2Y114_SLICE_X1Y114_BMUX = CLBLL_L_X2Y114_SLICE_X1Y114_BO5;
  assign CLBLL_L_X2Y114_SLICE_X1Y114_CMUX = CLBLL_L_X2Y114_SLICE_X1Y114_CO5;
  assign CLBLL_L_X2Y115_SLICE_X0Y115_A = CLBLL_L_X2Y115_SLICE_X0Y115_AO6;
  assign CLBLL_L_X2Y115_SLICE_X0Y115_B = CLBLL_L_X2Y115_SLICE_X0Y115_BO6;
  assign CLBLL_L_X2Y115_SLICE_X0Y115_C = CLBLL_L_X2Y115_SLICE_X0Y115_CO6;
  assign CLBLL_L_X2Y115_SLICE_X0Y115_D = CLBLL_L_X2Y115_SLICE_X0Y115_DO6;
  assign CLBLL_L_X2Y115_SLICE_X1Y115_A = CLBLL_L_X2Y115_SLICE_X1Y115_AO6;
  assign CLBLL_L_X2Y115_SLICE_X1Y115_B = CLBLL_L_X2Y115_SLICE_X1Y115_BO6;
  assign CLBLL_L_X2Y115_SLICE_X1Y115_C = CLBLL_L_X2Y115_SLICE_X1Y115_CO6;
  assign CLBLL_L_X2Y115_SLICE_X1Y115_D = CLBLL_L_X2Y115_SLICE_X1Y115_DO6;
  assign CLBLL_L_X2Y116_SLICE_X0Y116_A = CLBLL_L_X2Y116_SLICE_X0Y116_AO6;
  assign CLBLL_L_X2Y116_SLICE_X0Y116_B = CLBLL_L_X2Y116_SLICE_X0Y116_BO6;
  assign CLBLL_L_X2Y116_SLICE_X0Y116_C = CLBLL_L_X2Y116_SLICE_X0Y116_CO6;
  assign CLBLL_L_X2Y116_SLICE_X0Y116_D = CLBLL_L_X2Y116_SLICE_X0Y116_DO6;
  assign CLBLL_L_X2Y116_SLICE_X1Y116_A = CLBLL_L_X2Y116_SLICE_X1Y116_AO6;
  assign CLBLL_L_X2Y116_SLICE_X1Y116_B = CLBLL_L_X2Y116_SLICE_X1Y116_BO6;
  assign CLBLL_L_X2Y116_SLICE_X1Y116_C = CLBLL_L_X2Y116_SLICE_X1Y116_CO6;
  assign CLBLL_L_X2Y116_SLICE_X1Y116_D = CLBLL_L_X2Y116_SLICE_X1Y116_DO6;
  assign CLBLL_L_X2Y117_SLICE_X0Y117_A = CLBLL_L_X2Y117_SLICE_X0Y117_AO6;
  assign CLBLL_L_X2Y117_SLICE_X0Y117_B = CLBLL_L_X2Y117_SLICE_X0Y117_BO6;
  assign CLBLL_L_X2Y117_SLICE_X0Y117_C = CLBLL_L_X2Y117_SLICE_X0Y117_CO6;
  assign CLBLL_L_X2Y117_SLICE_X0Y117_D = CLBLL_L_X2Y117_SLICE_X0Y117_DO6;
  assign CLBLL_L_X2Y117_SLICE_X0Y117_AMUX = CLBLL_L_X2Y117_SLICE_X0Y117_A5Q;
  assign CLBLL_L_X2Y117_SLICE_X0Y117_DMUX = CLBLL_L_X2Y117_SLICE_X0Y117_DO5;
  assign CLBLL_L_X2Y117_SLICE_X1Y117_A = CLBLL_L_X2Y117_SLICE_X1Y117_AO6;
  assign CLBLL_L_X2Y117_SLICE_X1Y117_B = CLBLL_L_X2Y117_SLICE_X1Y117_BO6;
  assign CLBLL_L_X2Y117_SLICE_X1Y117_C = CLBLL_L_X2Y117_SLICE_X1Y117_CO6;
  assign CLBLL_L_X2Y117_SLICE_X1Y117_D = CLBLL_L_X2Y117_SLICE_X1Y117_DO6;
  assign CLBLL_L_X2Y117_SLICE_X1Y117_CMUX = CLBLL_L_X2Y117_SLICE_X1Y117_CO6;
  assign CLBLL_L_X2Y118_SLICE_X0Y118_A = CLBLL_L_X2Y118_SLICE_X0Y118_AO6;
  assign CLBLL_L_X2Y118_SLICE_X0Y118_B = CLBLL_L_X2Y118_SLICE_X0Y118_BO6;
  assign CLBLL_L_X2Y118_SLICE_X0Y118_C = CLBLL_L_X2Y118_SLICE_X0Y118_CO6;
  assign CLBLL_L_X2Y118_SLICE_X0Y118_D = CLBLL_L_X2Y118_SLICE_X0Y118_DO6;
  assign CLBLL_L_X2Y118_SLICE_X1Y118_A = CLBLL_L_X2Y118_SLICE_X1Y118_AO6;
  assign CLBLL_L_X2Y118_SLICE_X1Y118_B = CLBLL_L_X2Y118_SLICE_X1Y118_BO6;
  assign CLBLL_L_X2Y118_SLICE_X1Y118_C = CLBLL_L_X2Y118_SLICE_X1Y118_CO6;
  assign CLBLL_L_X2Y118_SLICE_X1Y118_D = CLBLL_L_X2Y118_SLICE_X1Y118_DO6;
  assign CLBLL_L_X2Y119_SLICE_X0Y119_A = CLBLL_L_X2Y119_SLICE_X0Y119_AO6;
  assign CLBLL_L_X2Y119_SLICE_X0Y119_B = CLBLL_L_X2Y119_SLICE_X0Y119_BO6;
  assign CLBLL_L_X2Y119_SLICE_X0Y119_C = CLBLL_L_X2Y119_SLICE_X0Y119_CO6;
  assign CLBLL_L_X2Y119_SLICE_X0Y119_D = CLBLL_L_X2Y119_SLICE_X0Y119_DO6;
  assign CLBLL_L_X2Y119_SLICE_X1Y119_A = CLBLL_L_X2Y119_SLICE_X1Y119_AO6;
  assign CLBLL_L_X2Y119_SLICE_X1Y119_B = CLBLL_L_X2Y119_SLICE_X1Y119_BO6;
  assign CLBLL_L_X2Y119_SLICE_X1Y119_C = CLBLL_L_X2Y119_SLICE_X1Y119_CO6;
  assign CLBLL_L_X2Y119_SLICE_X1Y119_D = CLBLL_L_X2Y119_SLICE_X1Y119_DO6;
  assign CLBLL_L_X2Y119_SLICE_X1Y119_AMUX = CLBLL_L_X2Y119_SLICE_X1Y119_AO5;
  assign CLBLL_L_X2Y120_SLICE_X0Y120_A = CLBLL_L_X2Y120_SLICE_X0Y120_AO6;
  assign CLBLL_L_X2Y120_SLICE_X0Y120_B = CLBLL_L_X2Y120_SLICE_X0Y120_BO6;
  assign CLBLL_L_X2Y120_SLICE_X0Y120_C = CLBLL_L_X2Y120_SLICE_X0Y120_CO6;
  assign CLBLL_L_X2Y120_SLICE_X0Y120_D = CLBLL_L_X2Y120_SLICE_X0Y120_DO6;
  assign CLBLL_L_X2Y120_SLICE_X0Y120_AMUX = CLBLL_L_X2Y120_SLICE_X0Y120_AO5;
  assign CLBLL_L_X2Y120_SLICE_X1Y120_A = CLBLL_L_X2Y120_SLICE_X1Y120_AO6;
  assign CLBLL_L_X2Y120_SLICE_X1Y120_B = CLBLL_L_X2Y120_SLICE_X1Y120_BO6;
  assign CLBLL_L_X2Y120_SLICE_X1Y120_C = CLBLL_L_X2Y120_SLICE_X1Y120_CO6;
  assign CLBLL_L_X2Y120_SLICE_X1Y120_D = CLBLL_L_X2Y120_SLICE_X1Y120_DO6;
  assign CLBLL_L_X2Y120_SLICE_X1Y120_AMUX = CLBLL_L_X2Y120_SLICE_X1Y120_AO5;
  assign CLBLL_L_X2Y120_SLICE_X1Y120_CMUX = CLBLL_L_X2Y120_SLICE_X1Y120_CO6;
  assign CLBLL_L_X2Y121_SLICE_X0Y121_A = CLBLL_L_X2Y121_SLICE_X0Y121_AO6;
  assign CLBLL_L_X2Y121_SLICE_X0Y121_B = CLBLL_L_X2Y121_SLICE_X0Y121_BO6;
  assign CLBLL_L_X2Y121_SLICE_X0Y121_C = CLBLL_L_X2Y121_SLICE_X0Y121_CO6;
  assign CLBLL_L_X2Y121_SLICE_X0Y121_D = CLBLL_L_X2Y121_SLICE_X0Y121_DO6;
  assign CLBLL_L_X2Y121_SLICE_X0Y121_AMUX = CLBLL_L_X2Y121_SLICE_X0Y121_AO5;
  assign CLBLL_L_X2Y121_SLICE_X0Y121_BMUX = CLBLL_L_X2Y121_SLICE_X0Y121_BO5;
  assign CLBLL_L_X2Y121_SLICE_X1Y121_A = CLBLL_L_X2Y121_SLICE_X1Y121_AO6;
  assign CLBLL_L_X2Y121_SLICE_X1Y121_B = CLBLL_L_X2Y121_SLICE_X1Y121_BO6;
  assign CLBLL_L_X2Y121_SLICE_X1Y121_C = CLBLL_L_X2Y121_SLICE_X1Y121_CO6;
  assign CLBLL_L_X2Y121_SLICE_X1Y121_D = CLBLL_L_X2Y121_SLICE_X1Y121_DO6;
  assign CLBLL_L_X2Y121_SLICE_X1Y121_AMUX = CLBLL_L_X2Y121_SLICE_X1Y121_AO5;
  assign CLBLL_L_X2Y121_SLICE_X1Y121_BMUX = CLBLL_L_X2Y121_SLICE_X1Y121_BO5;
  assign CLBLL_L_X2Y122_SLICE_X0Y122_A = CLBLL_L_X2Y122_SLICE_X0Y122_AO6;
  assign CLBLL_L_X2Y122_SLICE_X0Y122_B = CLBLL_L_X2Y122_SLICE_X0Y122_BO6;
  assign CLBLL_L_X2Y122_SLICE_X0Y122_C = CLBLL_L_X2Y122_SLICE_X0Y122_CO6;
  assign CLBLL_L_X2Y122_SLICE_X0Y122_D = CLBLL_L_X2Y122_SLICE_X0Y122_DO6;
  assign CLBLL_L_X2Y122_SLICE_X0Y122_AMUX = CLBLL_L_X2Y122_SLICE_X0Y122_AO5;
  assign CLBLL_L_X2Y122_SLICE_X1Y122_A = CLBLL_L_X2Y122_SLICE_X1Y122_AO6;
  assign CLBLL_L_X2Y122_SLICE_X1Y122_B = CLBLL_L_X2Y122_SLICE_X1Y122_BO6;
  assign CLBLL_L_X2Y122_SLICE_X1Y122_C = CLBLL_L_X2Y122_SLICE_X1Y122_CO6;
  assign CLBLL_L_X2Y122_SLICE_X1Y122_D = CLBLL_L_X2Y122_SLICE_X1Y122_DO6;
  assign CLBLL_L_X2Y122_SLICE_X1Y122_BMUX = CLBLL_L_X2Y122_SLICE_X1Y122_BO6;
  assign CLBLL_L_X2Y123_SLICE_X0Y123_A = CLBLL_L_X2Y123_SLICE_X0Y123_AO6;
  assign CLBLL_L_X2Y123_SLICE_X0Y123_B = CLBLL_L_X2Y123_SLICE_X0Y123_BO6;
  assign CLBLL_L_X2Y123_SLICE_X0Y123_C = CLBLL_L_X2Y123_SLICE_X0Y123_CO6;
  assign CLBLL_L_X2Y123_SLICE_X0Y123_D = CLBLL_L_X2Y123_SLICE_X0Y123_DO6;
  assign CLBLL_L_X2Y123_SLICE_X1Y123_A = CLBLL_L_X2Y123_SLICE_X1Y123_AO6;
  assign CLBLL_L_X2Y123_SLICE_X1Y123_B = CLBLL_L_X2Y123_SLICE_X1Y123_BO6;
  assign CLBLL_L_X2Y123_SLICE_X1Y123_C = CLBLL_L_X2Y123_SLICE_X1Y123_CO6;
  assign CLBLL_L_X2Y123_SLICE_X1Y123_D = CLBLL_L_X2Y123_SLICE_X1Y123_DO6;
  assign CLBLL_L_X4Y110_SLICE_X4Y110_A = CLBLL_L_X4Y110_SLICE_X4Y110_AO6;
  assign CLBLL_L_X4Y110_SLICE_X4Y110_B = CLBLL_L_X4Y110_SLICE_X4Y110_BO6;
  assign CLBLL_L_X4Y110_SLICE_X4Y110_C = CLBLL_L_X4Y110_SLICE_X4Y110_CO6;
  assign CLBLL_L_X4Y110_SLICE_X4Y110_D = CLBLL_L_X4Y110_SLICE_X4Y110_DO6;
  assign CLBLL_L_X4Y110_SLICE_X4Y110_AMUX = CLBLL_L_X4Y110_SLICE_X4Y110_A5Q;
  assign CLBLL_L_X4Y110_SLICE_X4Y110_BMUX = CLBLL_L_X4Y110_SLICE_X4Y110_BO5;
  assign CLBLL_L_X4Y110_SLICE_X5Y110_A = CLBLL_L_X4Y110_SLICE_X5Y110_AO6;
  assign CLBLL_L_X4Y110_SLICE_X5Y110_B = CLBLL_L_X4Y110_SLICE_X5Y110_BO6;
  assign CLBLL_L_X4Y110_SLICE_X5Y110_C = CLBLL_L_X4Y110_SLICE_X5Y110_CO6;
  assign CLBLL_L_X4Y110_SLICE_X5Y110_D = CLBLL_L_X4Y110_SLICE_X5Y110_DO6;
  assign CLBLL_L_X4Y110_SLICE_X5Y110_CMUX = CLBLL_L_X4Y110_SLICE_X5Y110_CO5;
  assign CLBLL_L_X4Y111_SLICE_X4Y111_A = CLBLL_L_X4Y111_SLICE_X4Y111_AO6;
  assign CLBLL_L_X4Y111_SLICE_X4Y111_B = CLBLL_L_X4Y111_SLICE_X4Y111_BO6;
  assign CLBLL_L_X4Y111_SLICE_X4Y111_C = CLBLL_L_X4Y111_SLICE_X4Y111_CO6;
  assign CLBLL_L_X4Y111_SLICE_X4Y111_D = CLBLL_L_X4Y111_SLICE_X4Y111_DO6;
  assign CLBLL_L_X4Y111_SLICE_X4Y111_AMUX = CLBLL_L_X4Y111_SLICE_X4Y111_AO5;
  assign CLBLL_L_X4Y111_SLICE_X5Y111_A = CLBLL_L_X4Y111_SLICE_X5Y111_AO6;
  assign CLBLL_L_X4Y111_SLICE_X5Y111_B = CLBLL_L_X4Y111_SLICE_X5Y111_BO6;
  assign CLBLL_L_X4Y111_SLICE_X5Y111_C = CLBLL_L_X4Y111_SLICE_X5Y111_CO6;
  assign CLBLL_L_X4Y111_SLICE_X5Y111_D = CLBLL_L_X4Y111_SLICE_X5Y111_DO6;
  assign CLBLL_L_X4Y111_SLICE_X5Y111_AMUX = CLBLL_L_X4Y111_SLICE_X5Y111_A5Q;
  assign CLBLL_L_X4Y111_SLICE_X5Y111_DMUX = CLBLL_L_X4Y111_SLICE_X5Y111_DO6;
  assign CLBLL_L_X4Y112_SLICE_X4Y112_A = CLBLL_L_X4Y112_SLICE_X4Y112_AO6;
  assign CLBLL_L_X4Y112_SLICE_X4Y112_B = CLBLL_L_X4Y112_SLICE_X4Y112_BO6;
  assign CLBLL_L_X4Y112_SLICE_X4Y112_C = CLBLL_L_X4Y112_SLICE_X4Y112_CO6;
  assign CLBLL_L_X4Y112_SLICE_X4Y112_D = CLBLL_L_X4Y112_SLICE_X4Y112_DO6;
  assign CLBLL_L_X4Y112_SLICE_X5Y112_A = CLBLL_L_X4Y112_SLICE_X5Y112_AO6;
  assign CLBLL_L_X4Y112_SLICE_X5Y112_B = CLBLL_L_X4Y112_SLICE_X5Y112_BO6;
  assign CLBLL_L_X4Y112_SLICE_X5Y112_C = CLBLL_L_X4Y112_SLICE_X5Y112_CO6;
  assign CLBLL_L_X4Y112_SLICE_X5Y112_D = CLBLL_L_X4Y112_SLICE_X5Y112_DO6;
  assign CLBLL_L_X4Y112_SLICE_X5Y112_DMUX = CLBLL_L_X4Y112_SLICE_X5Y112_DO6;
  assign CLBLL_L_X4Y113_SLICE_X4Y113_A = CLBLL_L_X4Y113_SLICE_X4Y113_AO6;
  assign CLBLL_L_X4Y113_SLICE_X4Y113_B = CLBLL_L_X4Y113_SLICE_X4Y113_BO6;
  assign CLBLL_L_X4Y113_SLICE_X4Y113_C = CLBLL_L_X4Y113_SLICE_X4Y113_CO6;
  assign CLBLL_L_X4Y113_SLICE_X4Y113_D = CLBLL_L_X4Y113_SLICE_X4Y113_DO6;
  assign CLBLL_L_X4Y113_SLICE_X5Y113_A = CLBLL_L_X4Y113_SLICE_X5Y113_AO6;
  assign CLBLL_L_X4Y113_SLICE_X5Y113_B = CLBLL_L_X4Y113_SLICE_X5Y113_BO6;
  assign CLBLL_L_X4Y113_SLICE_X5Y113_C = CLBLL_L_X4Y113_SLICE_X5Y113_CO6;
  assign CLBLL_L_X4Y113_SLICE_X5Y113_D = CLBLL_L_X4Y113_SLICE_X5Y113_DO6;
  assign CLBLL_L_X4Y113_SLICE_X5Y113_DMUX = CLBLL_L_X4Y113_SLICE_X5Y113_DO5;
  assign CLBLL_L_X4Y114_SLICE_X4Y114_A = CLBLL_L_X4Y114_SLICE_X4Y114_AO6;
  assign CLBLL_L_X4Y114_SLICE_X4Y114_B = CLBLL_L_X4Y114_SLICE_X4Y114_BO6;
  assign CLBLL_L_X4Y114_SLICE_X4Y114_C = CLBLL_L_X4Y114_SLICE_X4Y114_CO6;
  assign CLBLL_L_X4Y114_SLICE_X4Y114_D = CLBLL_L_X4Y114_SLICE_X4Y114_DO6;
  assign CLBLL_L_X4Y114_SLICE_X5Y114_A = CLBLL_L_X4Y114_SLICE_X5Y114_AO6;
  assign CLBLL_L_X4Y114_SLICE_X5Y114_B = CLBLL_L_X4Y114_SLICE_X5Y114_BO6;
  assign CLBLL_L_X4Y114_SLICE_X5Y114_C = CLBLL_L_X4Y114_SLICE_X5Y114_CO6;
  assign CLBLL_L_X4Y114_SLICE_X5Y114_D = CLBLL_L_X4Y114_SLICE_X5Y114_DO6;
  assign CLBLL_L_X4Y114_SLICE_X5Y114_BMUX = CLBLL_L_X4Y114_SLICE_X5Y114_BO5;
  assign CLBLL_L_X4Y114_SLICE_X5Y114_CMUX = CLBLL_L_X4Y114_SLICE_X5Y114_CO6;
  assign CLBLL_L_X4Y115_SLICE_X4Y115_A = CLBLL_L_X4Y115_SLICE_X4Y115_AO6;
  assign CLBLL_L_X4Y115_SLICE_X4Y115_B = CLBLL_L_X4Y115_SLICE_X4Y115_BO6;
  assign CLBLL_L_X4Y115_SLICE_X4Y115_C = CLBLL_L_X4Y115_SLICE_X4Y115_CO6;
  assign CLBLL_L_X4Y115_SLICE_X4Y115_D = CLBLL_L_X4Y115_SLICE_X4Y115_DO6;
  assign CLBLL_L_X4Y115_SLICE_X4Y115_CMUX = CLBLL_L_X4Y115_SLICE_X4Y115_C5Q;
  assign CLBLL_L_X4Y115_SLICE_X5Y115_A = CLBLL_L_X4Y115_SLICE_X5Y115_AO6;
  assign CLBLL_L_X4Y115_SLICE_X5Y115_B = CLBLL_L_X4Y115_SLICE_X5Y115_BO6;
  assign CLBLL_L_X4Y115_SLICE_X5Y115_C = CLBLL_L_X4Y115_SLICE_X5Y115_CO6;
  assign CLBLL_L_X4Y115_SLICE_X5Y115_D = CLBLL_L_X4Y115_SLICE_X5Y115_DO6;
  assign CLBLL_L_X4Y116_SLICE_X4Y116_A = CLBLL_L_X4Y116_SLICE_X4Y116_AO6;
  assign CLBLL_L_X4Y116_SLICE_X4Y116_B = CLBLL_L_X4Y116_SLICE_X4Y116_BO6;
  assign CLBLL_L_X4Y116_SLICE_X4Y116_C = CLBLL_L_X4Y116_SLICE_X4Y116_CO6;
  assign CLBLL_L_X4Y116_SLICE_X4Y116_D = CLBLL_L_X4Y116_SLICE_X4Y116_DO6;
  assign CLBLL_L_X4Y116_SLICE_X4Y116_CMUX = CLBLL_L_X4Y116_SLICE_X4Y116_C5Q;
  assign CLBLL_L_X4Y116_SLICE_X5Y116_A = CLBLL_L_X4Y116_SLICE_X5Y116_AO6;
  assign CLBLL_L_X4Y116_SLICE_X5Y116_B = CLBLL_L_X4Y116_SLICE_X5Y116_BO6;
  assign CLBLL_L_X4Y116_SLICE_X5Y116_C = CLBLL_L_X4Y116_SLICE_X5Y116_CO6;
  assign CLBLL_L_X4Y116_SLICE_X5Y116_D = CLBLL_L_X4Y116_SLICE_X5Y116_DO6;
  assign CLBLL_L_X4Y116_SLICE_X5Y116_AMUX = CLBLL_L_X4Y116_SLICE_X5Y116_A5Q;
  assign CLBLL_L_X4Y116_SLICE_X5Y116_CMUX = CLBLL_L_X4Y116_SLICE_X5Y116_CO5;
  assign CLBLL_L_X4Y117_SLICE_X4Y117_A = CLBLL_L_X4Y117_SLICE_X4Y117_AO6;
  assign CLBLL_L_X4Y117_SLICE_X4Y117_B = CLBLL_L_X4Y117_SLICE_X4Y117_BO6;
  assign CLBLL_L_X4Y117_SLICE_X4Y117_C = CLBLL_L_X4Y117_SLICE_X4Y117_CO6;
  assign CLBLL_L_X4Y117_SLICE_X4Y117_D = CLBLL_L_X4Y117_SLICE_X4Y117_DO6;
  assign CLBLL_L_X4Y117_SLICE_X5Y117_A = CLBLL_L_X4Y117_SLICE_X5Y117_AO6;
  assign CLBLL_L_X4Y117_SLICE_X5Y117_B = CLBLL_L_X4Y117_SLICE_X5Y117_BO6;
  assign CLBLL_L_X4Y117_SLICE_X5Y117_C = CLBLL_L_X4Y117_SLICE_X5Y117_CO6;
  assign CLBLL_L_X4Y117_SLICE_X5Y117_D = CLBLL_L_X4Y117_SLICE_X5Y117_DO6;
  assign CLBLL_L_X4Y118_SLICE_X4Y118_A = CLBLL_L_X4Y118_SLICE_X4Y118_AO6;
  assign CLBLL_L_X4Y118_SLICE_X4Y118_B = CLBLL_L_X4Y118_SLICE_X4Y118_BO6;
  assign CLBLL_L_X4Y118_SLICE_X4Y118_C = CLBLL_L_X4Y118_SLICE_X4Y118_CO6;
  assign CLBLL_L_X4Y118_SLICE_X4Y118_D = CLBLL_L_X4Y118_SLICE_X4Y118_DO6;
  assign CLBLL_L_X4Y118_SLICE_X5Y118_A = CLBLL_L_X4Y118_SLICE_X5Y118_AO6;
  assign CLBLL_L_X4Y118_SLICE_X5Y118_B = CLBLL_L_X4Y118_SLICE_X5Y118_BO6;
  assign CLBLL_L_X4Y118_SLICE_X5Y118_C = CLBLL_L_X4Y118_SLICE_X5Y118_CO6;
  assign CLBLL_L_X4Y118_SLICE_X5Y118_D = CLBLL_L_X4Y118_SLICE_X5Y118_DO6;
  assign CLBLL_L_X4Y119_SLICE_X4Y119_A = CLBLL_L_X4Y119_SLICE_X4Y119_AO6;
  assign CLBLL_L_X4Y119_SLICE_X4Y119_B = CLBLL_L_X4Y119_SLICE_X4Y119_BO6;
  assign CLBLL_L_X4Y119_SLICE_X4Y119_C = CLBLL_L_X4Y119_SLICE_X4Y119_CO6;
  assign CLBLL_L_X4Y119_SLICE_X4Y119_D = CLBLL_L_X4Y119_SLICE_X4Y119_DO6;
  assign CLBLL_L_X4Y119_SLICE_X4Y119_BMUX = CLBLL_L_X4Y119_SLICE_X4Y119_B5Q;
  assign CLBLL_L_X4Y119_SLICE_X4Y119_CMUX = CLBLL_L_X4Y119_SLICE_X4Y119_C5Q;
  assign CLBLL_L_X4Y119_SLICE_X5Y119_A = CLBLL_L_X4Y119_SLICE_X5Y119_AO6;
  assign CLBLL_L_X4Y119_SLICE_X5Y119_B = CLBLL_L_X4Y119_SLICE_X5Y119_BO6;
  assign CLBLL_L_X4Y119_SLICE_X5Y119_C = CLBLL_L_X4Y119_SLICE_X5Y119_CO6;
  assign CLBLL_L_X4Y119_SLICE_X5Y119_D = CLBLL_L_X4Y119_SLICE_X5Y119_DO6;
  assign CLBLL_L_X4Y120_SLICE_X4Y120_A = CLBLL_L_X4Y120_SLICE_X4Y120_AO6;
  assign CLBLL_L_X4Y120_SLICE_X4Y120_B = CLBLL_L_X4Y120_SLICE_X4Y120_BO6;
  assign CLBLL_L_X4Y120_SLICE_X4Y120_C = CLBLL_L_X4Y120_SLICE_X4Y120_CO6;
  assign CLBLL_L_X4Y120_SLICE_X4Y120_D = CLBLL_L_X4Y120_SLICE_X4Y120_DO6;
  assign CLBLL_L_X4Y120_SLICE_X4Y120_DMUX = CLBLL_L_X4Y120_SLICE_X4Y120_DO6;
  assign CLBLL_L_X4Y120_SLICE_X5Y120_A = CLBLL_L_X4Y120_SLICE_X5Y120_AO6;
  assign CLBLL_L_X4Y120_SLICE_X5Y120_B = CLBLL_L_X4Y120_SLICE_X5Y120_BO6;
  assign CLBLL_L_X4Y120_SLICE_X5Y120_C = CLBLL_L_X4Y120_SLICE_X5Y120_CO6;
  assign CLBLL_L_X4Y120_SLICE_X5Y120_D = CLBLL_L_X4Y120_SLICE_X5Y120_DO6;
  assign CLBLL_L_X4Y120_SLICE_X5Y120_AMUX = CLBLL_L_X4Y120_SLICE_X5Y120_AO5;
  assign CLBLL_L_X4Y120_SLICE_X5Y120_BMUX = CLBLL_L_X4Y120_SLICE_X5Y120_BO5;
  assign CLBLL_L_X4Y121_SLICE_X4Y121_A = CLBLL_L_X4Y121_SLICE_X4Y121_AO6;
  assign CLBLL_L_X4Y121_SLICE_X4Y121_B = CLBLL_L_X4Y121_SLICE_X4Y121_BO6;
  assign CLBLL_L_X4Y121_SLICE_X4Y121_C = CLBLL_L_X4Y121_SLICE_X4Y121_CO6;
  assign CLBLL_L_X4Y121_SLICE_X4Y121_D = CLBLL_L_X4Y121_SLICE_X4Y121_DO6;
  assign CLBLL_L_X4Y121_SLICE_X4Y121_CMUX = CLBLL_L_X4Y121_SLICE_X4Y121_CO5;
  assign CLBLL_L_X4Y121_SLICE_X4Y121_DMUX = CLBLL_L_X4Y121_SLICE_X4Y121_DO5;
  assign CLBLL_L_X4Y121_SLICE_X5Y121_A = CLBLL_L_X4Y121_SLICE_X5Y121_AO6;
  assign CLBLL_L_X4Y121_SLICE_X5Y121_B = CLBLL_L_X4Y121_SLICE_X5Y121_BO6;
  assign CLBLL_L_X4Y121_SLICE_X5Y121_C = CLBLL_L_X4Y121_SLICE_X5Y121_CO6;
  assign CLBLL_L_X4Y121_SLICE_X5Y121_D = CLBLL_L_X4Y121_SLICE_X5Y121_DO6;
  assign CLBLL_L_X4Y121_SLICE_X5Y121_BMUX = CLBLL_L_X4Y121_SLICE_X5Y121_BO5;
  assign CLBLL_L_X4Y121_SLICE_X5Y121_CMUX = CLBLL_L_X4Y121_SLICE_X5Y121_CO5;
  assign CLBLL_L_X4Y122_SLICE_X4Y122_A = CLBLL_L_X4Y122_SLICE_X4Y122_AO6;
  assign CLBLL_L_X4Y122_SLICE_X4Y122_B = CLBLL_L_X4Y122_SLICE_X4Y122_BO6;
  assign CLBLL_L_X4Y122_SLICE_X4Y122_C = CLBLL_L_X4Y122_SLICE_X4Y122_CO6;
  assign CLBLL_L_X4Y122_SLICE_X4Y122_D = CLBLL_L_X4Y122_SLICE_X4Y122_DO6;
  assign CLBLL_L_X4Y122_SLICE_X4Y122_AMUX = CLBLL_L_X4Y122_SLICE_X4Y122_AO5;
  assign CLBLL_L_X4Y122_SLICE_X5Y122_A = CLBLL_L_X4Y122_SLICE_X5Y122_AO6;
  assign CLBLL_L_X4Y122_SLICE_X5Y122_B = CLBLL_L_X4Y122_SLICE_X5Y122_BO6;
  assign CLBLL_L_X4Y122_SLICE_X5Y122_C = CLBLL_L_X4Y122_SLICE_X5Y122_CO6;
  assign CLBLL_L_X4Y122_SLICE_X5Y122_D = CLBLL_L_X4Y122_SLICE_X5Y122_DO6;
  assign CLBLL_L_X4Y123_SLICE_X4Y123_A = CLBLL_L_X4Y123_SLICE_X4Y123_AO6;
  assign CLBLL_L_X4Y123_SLICE_X4Y123_B = CLBLL_L_X4Y123_SLICE_X4Y123_BO6;
  assign CLBLL_L_X4Y123_SLICE_X4Y123_C = CLBLL_L_X4Y123_SLICE_X4Y123_CO6;
  assign CLBLL_L_X4Y123_SLICE_X4Y123_D = CLBLL_L_X4Y123_SLICE_X4Y123_DO6;
  assign CLBLL_L_X4Y123_SLICE_X5Y123_A = CLBLL_L_X4Y123_SLICE_X5Y123_AO6;
  assign CLBLL_L_X4Y123_SLICE_X5Y123_B = CLBLL_L_X4Y123_SLICE_X5Y123_BO6;
  assign CLBLL_L_X4Y123_SLICE_X5Y123_C = CLBLL_L_X4Y123_SLICE_X5Y123_CO6;
  assign CLBLL_L_X4Y123_SLICE_X5Y123_D = CLBLL_L_X4Y123_SLICE_X5Y123_DO6;
  assign CLBLL_L_X4Y123_SLICE_X5Y123_AMUX = CLBLL_L_X4Y123_SLICE_X5Y123_AO5;
  assign CLBLL_L_X52Y126_SLICE_X78Y126_A = CLBLL_L_X52Y126_SLICE_X78Y126_AO6;
  assign CLBLL_L_X52Y126_SLICE_X78Y126_B = CLBLL_L_X52Y126_SLICE_X78Y126_BO6;
  assign CLBLL_L_X52Y126_SLICE_X78Y126_C = CLBLL_L_X52Y126_SLICE_X78Y126_CO6;
  assign CLBLL_L_X52Y126_SLICE_X78Y126_D = CLBLL_L_X52Y126_SLICE_X78Y126_DO6;
  assign CLBLL_L_X52Y126_SLICE_X79Y126_A = CLBLL_L_X52Y126_SLICE_X79Y126_AO6;
  assign CLBLL_L_X52Y126_SLICE_X79Y126_B = CLBLL_L_X52Y126_SLICE_X79Y126_BO6;
  assign CLBLL_L_X52Y126_SLICE_X79Y126_C = CLBLL_L_X52Y126_SLICE_X79Y126_CO6;
  assign CLBLL_L_X52Y126_SLICE_X79Y126_D = CLBLL_L_X52Y126_SLICE_X79Y126_DO6;
  assign CLBLM_L_X8Y110_SLICE_X10Y110_A = CLBLM_L_X8Y110_SLICE_X10Y110_AO6;
  assign CLBLM_L_X8Y110_SLICE_X10Y110_B = CLBLM_L_X8Y110_SLICE_X10Y110_BO6;
  assign CLBLM_L_X8Y110_SLICE_X10Y110_C = CLBLM_L_X8Y110_SLICE_X10Y110_CO6;
  assign CLBLM_L_X8Y110_SLICE_X10Y110_D = CLBLM_L_X8Y110_SLICE_X10Y110_DO6;
  assign CLBLM_L_X8Y110_SLICE_X11Y110_A = CLBLM_L_X8Y110_SLICE_X11Y110_AO6;
  assign CLBLM_L_X8Y110_SLICE_X11Y110_B = CLBLM_L_X8Y110_SLICE_X11Y110_BO6;
  assign CLBLM_L_X8Y110_SLICE_X11Y110_C = CLBLM_L_X8Y110_SLICE_X11Y110_CO6;
  assign CLBLM_L_X8Y110_SLICE_X11Y110_D = CLBLM_L_X8Y110_SLICE_X11Y110_DO6;
  assign CLBLM_L_X8Y111_SLICE_X10Y111_A = CLBLM_L_X8Y111_SLICE_X10Y111_AO6;
  assign CLBLM_L_X8Y111_SLICE_X10Y111_B = CLBLM_L_X8Y111_SLICE_X10Y111_BO6;
  assign CLBLM_L_X8Y111_SLICE_X10Y111_C = CLBLM_L_X8Y111_SLICE_X10Y111_CO6;
  assign CLBLM_L_X8Y111_SLICE_X10Y111_D = CLBLM_L_X8Y111_SLICE_X10Y111_DO6;
  assign CLBLM_L_X8Y111_SLICE_X11Y111_A = CLBLM_L_X8Y111_SLICE_X11Y111_AO6;
  assign CLBLM_L_X8Y111_SLICE_X11Y111_B = CLBLM_L_X8Y111_SLICE_X11Y111_BO6;
  assign CLBLM_L_X8Y111_SLICE_X11Y111_C = CLBLM_L_X8Y111_SLICE_X11Y111_CO6;
  assign CLBLM_L_X8Y111_SLICE_X11Y111_D = CLBLM_L_X8Y111_SLICE_X11Y111_DO6;
  assign CLBLM_L_X8Y112_SLICE_X10Y112_A = CLBLM_L_X8Y112_SLICE_X10Y112_AO6;
  assign CLBLM_L_X8Y112_SLICE_X10Y112_B = CLBLM_L_X8Y112_SLICE_X10Y112_BO6;
  assign CLBLM_L_X8Y112_SLICE_X10Y112_C = CLBLM_L_X8Y112_SLICE_X10Y112_CO6;
  assign CLBLM_L_X8Y112_SLICE_X10Y112_D = CLBLM_L_X8Y112_SLICE_X10Y112_DO6;
  assign CLBLM_L_X8Y112_SLICE_X11Y112_A = CLBLM_L_X8Y112_SLICE_X11Y112_AO6;
  assign CLBLM_L_X8Y112_SLICE_X11Y112_B = CLBLM_L_X8Y112_SLICE_X11Y112_BO6;
  assign CLBLM_L_X8Y112_SLICE_X11Y112_C = CLBLM_L_X8Y112_SLICE_X11Y112_CO6;
  assign CLBLM_L_X8Y112_SLICE_X11Y112_D = CLBLM_L_X8Y112_SLICE_X11Y112_DO6;
  assign CLBLM_L_X8Y112_SLICE_X11Y112_BMUX = CLBLM_L_X8Y112_SLICE_X11Y112_BO5;
  assign CLBLM_L_X8Y113_SLICE_X10Y113_A = CLBLM_L_X8Y113_SLICE_X10Y113_AO6;
  assign CLBLM_L_X8Y113_SLICE_X10Y113_B = CLBLM_L_X8Y113_SLICE_X10Y113_BO6;
  assign CLBLM_L_X8Y113_SLICE_X10Y113_C = CLBLM_L_X8Y113_SLICE_X10Y113_CO6;
  assign CLBLM_L_X8Y113_SLICE_X10Y113_D = CLBLM_L_X8Y113_SLICE_X10Y113_DO6;
  assign CLBLM_L_X8Y113_SLICE_X11Y113_A = CLBLM_L_X8Y113_SLICE_X11Y113_AO6;
  assign CLBLM_L_X8Y113_SLICE_X11Y113_B = CLBLM_L_X8Y113_SLICE_X11Y113_BO6;
  assign CLBLM_L_X8Y113_SLICE_X11Y113_C = CLBLM_L_X8Y113_SLICE_X11Y113_CO6;
  assign CLBLM_L_X8Y113_SLICE_X11Y113_D = CLBLM_L_X8Y113_SLICE_X11Y113_DO6;
  assign CLBLM_L_X8Y114_SLICE_X10Y114_A = CLBLM_L_X8Y114_SLICE_X10Y114_AO6;
  assign CLBLM_L_X8Y114_SLICE_X10Y114_B = CLBLM_L_X8Y114_SLICE_X10Y114_BO6;
  assign CLBLM_L_X8Y114_SLICE_X10Y114_C = CLBLM_L_X8Y114_SLICE_X10Y114_CO6;
  assign CLBLM_L_X8Y114_SLICE_X10Y114_D = CLBLM_L_X8Y114_SLICE_X10Y114_DO6;
  assign CLBLM_L_X8Y114_SLICE_X10Y114_BMUX = CLBLM_L_X8Y114_SLICE_X10Y114_B5Q;
  assign CLBLM_L_X8Y114_SLICE_X10Y114_CMUX = CLBLM_L_X8Y114_SLICE_X10Y114_C5Q;
  assign CLBLM_L_X8Y114_SLICE_X11Y114_A = CLBLM_L_X8Y114_SLICE_X11Y114_AO6;
  assign CLBLM_L_X8Y114_SLICE_X11Y114_B = CLBLM_L_X8Y114_SLICE_X11Y114_BO6;
  assign CLBLM_L_X8Y114_SLICE_X11Y114_C = CLBLM_L_X8Y114_SLICE_X11Y114_CO6;
  assign CLBLM_L_X8Y114_SLICE_X11Y114_D = CLBLM_L_X8Y114_SLICE_X11Y114_DO6;
  assign CLBLM_L_X8Y115_SLICE_X10Y115_A = CLBLM_L_X8Y115_SLICE_X10Y115_AO6;
  assign CLBLM_L_X8Y115_SLICE_X10Y115_B = CLBLM_L_X8Y115_SLICE_X10Y115_BO6;
  assign CLBLM_L_X8Y115_SLICE_X10Y115_C = CLBLM_L_X8Y115_SLICE_X10Y115_CO6;
  assign CLBLM_L_X8Y115_SLICE_X10Y115_D = CLBLM_L_X8Y115_SLICE_X10Y115_DO6;
  assign CLBLM_L_X8Y115_SLICE_X10Y115_BMUX = CLBLM_L_X8Y115_SLICE_X10Y115_BO5;
  assign CLBLM_L_X8Y115_SLICE_X10Y115_CMUX = CLBLM_L_X8Y115_SLICE_X10Y115_C5Q;
  assign CLBLM_L_X8Y115_SLICE_X11Y115_A = CLBLM_L_X8Y115_SLICE_X11Y115_AO6;
  assign CLBLM_L_X8Y115_SLICE_X11Y115_B = CLBLM_L_X8Y115_SLICE_X11Y115_BO6;
  assign CLBLM_L_X8Y115_SLICE_X11Y115_C = CLBLM_L_X8Y115_SLICE_X11Y115_CO6;
  assign CLBLM_L_X8Y115_SLICE_X11Y115_D = CLBLM_L_X8Y115_SLICE_X11Y115_DO6;
  assign CLBLM_L_X8Y115_SLICE_X11Y115_CMUX = CLBLM_L_X8Y115_SLICE_X11Y115_C5Q;
  assign CLBLM_L_X8Y116_SLICE_X10Y116_A = CLBLM_L_X8Y116_SLICE_X10Y116_AO6;
  assign CLBLM_L_X8Y116_SLICE_X10Y116_B = CLBLM_L_X8Y116_SLICE_X10Y116_BO6;
  assign CLBLM_L_X8Y116_SLICE_X10Y116_C = CLBLM_L_X8Y116_SLICE_X10Y116_CO6;
  assign CLBLM_L_X8Y116_SLICE_X10Y116_D = CLBLM_L_X8Y116_SLICE_X10Y116_DO6;
  assign CLBLM_L_X8Y116_SLICE_X11Y116_A = CLBLM_L_X8Y116_SLICE_X11Y116_AO6;
  assign CLBLM_L_X8Y116_SLICE_X11Y116_B = CLBLM_L_X8Y116_SLICE_X11Y116_BO6;
  assign CLBLM_L_X8Y116_SLICE_X11Y116_C = CLBLM_L_X8Y116_SLICE_X11Y116_CO6;
  assign CLBLM_L_X8Y116_SLICE_X11Y116_D = CLBLM_L_X8Y116_SLICE_X11Y116_DO6;
  assign CLBLM_L_X8Y116_SLICE_X11Y116_AMUX = CLBLM_L_X8Y116_SLICE_X11Y116_A5Q;
  assign CLBLM_L_X8Y116_SLICE_X11Y116_CMUX = CLBLM_L_X8Y116_SLICE_X11Y116_CO5;
  assign CLBLM_L_X8Y117_SLICE_X10Y117_A = CLBLM_L_X8Y117_SLICE_X10Y117_AO6;
  assign CLBLM_L_X8Y117_SLICE_X10Y117_B = CLBLM_L_X8Y117_SLICE_X10Y117_BO6;
  assign CLBLM_L_X8Y117_SLICE_X10Y117_C = CLBLM_L_X8Y117_SLICE_X10Y117_CO6;
  assign CLBLM_L_X8Y117_SLICE_X10Y117_D = CLBLM_L_X8Y117_SLICE_X10Y117_DO6;
  assign CLBLM_L_X8Y117_SLICE_X10Y117_DMUX = CLBLM_L_X8Y117_SLICE_X10Y117_DO5;
  assign CLBLM_L_X8Y117_SLICE_X11Y117_A = CLBLM_L_X8Y117_SLICE_X11Y117_AO6;
  assign CLBLM_L_X8Y117_SLICE_X11Y117_B = CLBLM_L_X8Y117_SLICE_X11Y117_BO6;
  assign CLBLM_L_X8Y117_SLICE_X11Y117_C = CLBLM_L_X8Y117_SLICE_X11Y117_CO6;
  assign CLBLM_L_X8Y117_SLICE_X11Y117_D = CLBLM_L_X8Y117_SLICE_X11Y117_DO6;
  assign CLBLM_L_X8Y118_SLICE_X10Y118_A = CLBLM_L_X8Y118_SLICE_X10Y118_AO6;
  assign CLBLM_L_X8Y118_SLICE_X10Y118_B = CLBLM_L_X8Y118_SLICE_X10Y118_BO6;
  assign CLBLM_L_X8Y118_SLICE_X10Y118_C = CLBLM_L_X8Y118_SLICE_X10Y118_CO6;
  assign CLBLM_L_X8Y118_SLICE_X10Y118_D = CLBLM_L_X8Y118_SLICE_X10Y118_DO6;
  assign CLBLM_L_X8Y118_SLICE_X10Y118_DMUX = CLBLM_L_X8Y118_SLICE_X10Y118_D5Q;
  assign CLBLM_L_X8Y118_SLICE_X11Y118_A = CLBLM_L_X8Y118_SLICE_X11Y118_AO6;
  assign CLBLM_L_X8Y118_SLICE_X11Y118_B = CLBLM_L_X8Y118_SLICE_X11Y118_BO6;
  assign CLBLM_L_X8Y118_SLICE_X11Y118_C = CLBLM_L_X8Y118_SLICE_X11Y118_CO6;
  assign CLBLM_L_X8Y118_SLICE_X11Y118_D = CLBLM_L_X8Y118_SLICE_X11Y118_DO6;
  assign CLBLM_L_X8Y118_SLICE_X11Y118_BMUX = CLBLM_L_X8Y118_SLICE_X11Y118_BO5;
  assign CLBLM_L_X8Y119_SLICE_X10Y119_A = CLBLM_L_X8Y119_SLICE_X10Y119_AO6;
  assign CLBLM_L_X8Y119_SLICE_X10Y119_B = CLBLM_L_X8Y119_SLICE_X10Y119_BO6;
  assign CLBLM_L_X8Y119_SLICE_X10Y119_C = CLBLM_L_X8Y119_SLICE_X10Y119_CO6;
  assign CLBLM_L_X8Y119_SLICE_X10Y119_D = CLBLM_L_X8Y119_SLICE_X10Y119_DO6;
  assign CLBLM_L_X8Y119_SLICE_X10Y119_AMUX = CLBLM_L_X8Y119_SLICE_X10Y119_A5Q;
  assign CLBLM_L_X8Y119_SLICE_X10Y119_DMUX = CLBLM_L_X8Y119_SLICE_X10Y119_DO5;
  assign CLBLM_L_X8Y119_SLICE_X11Y119_A = CLBLM_L_X8Y119_SLICE_X11Y119_AO6;
  assign CLBLM_L_X8Y119_SLICE_X11Y119_B = CLBLM_L_X8Y119_SLICE_X11Y119_BO6;
  assign CLBLM_L_X8Y119_SLICE_X11Y119_C = CLBLM_L_X8Y119_SLICE_X11Y119_CO6;
  assign CLBLM_L_X8Y119_SLICE_X11Y119_D = CLBLM_L_X8Y119_SLICE_X11Y119_DO6;
  assign CLBLM_L_X8Y119_SLICE_X11Y119_CMUX = CLBLM_L_X8Y119_SLICE_X11Y119_C5Q;
  assign CLBLM_L_X8Y120_SLICE_X10Y120_A = CLBLM_L_X8Y120_SLICE_X10Y120_AO6;
  assign CLBLM_L_X8Y120_SLICE_X10Y120_B = CLBLM_L_X8Y120_SLICE_X10Y120_BO6;
  assign CLBLM_L_X8Y120_SLICE_X10Y120_C = CLBLM_L_X8Y120_SLICE_X10Y120_CO6;
  assign CLBLM_L_X8Y120_SLICE_X10Y120_D = CLBLM_L_X8Y120_SLICE_X10Y120_DO6;
  assign CLBLM_L_X8Y120_SLICE_X10Y120_AMUX = CLBLM_L_X8Y120_SLICE_X10Y120_A5Q;
  assign CLBLM_L_X8Y120_SLICE_X10Y120_DMUX = CLBLM_L_X8Y120_SLICE_X10Y120_D5Q;
  assign CLBLM_L_X8Y120_SLICE_X11Y120_A = CLBLM_L_X8Y120_SLICE_X11Y120_AO6;
  assign CLBLM_L_X8Y120_SLICE_X11Y120_B = CLBLM_L_X8Y120_SLICE_X11Y120_BO6;
  assign CLBLM_L_X8Y120_SLICE_X11Y120_C = CLBLM_L_X8Y120_SLICE_X11Y120_CO6;
  assign CLBLM_L_X8Y120_SLICE_X11Y120_D = CLBLM_L_X8Y120_SLICE_X11Y120_DO6;
  assign CLBLM_L_X8Y120_SLICE_X11Y120_CMUX = CLBLM_L_X8Y120_SLICE_X11Y120_C5Q;
  assign CLBLM_L_X8Y121_SLICE_X10Y121_A = CLBLM_L_X8Y121_SLICE_X10Y121_AO6;
  assign CLBLM_L_X8Y121_SLICE_X10Y121_B = CLBLM_L_X8Y121_SLICE_X10Y121_BO6;
  assign CLBLM_L_X8Y121_SLICE_X10Y121_C = CLBLM_L_X8Y121_SLICE_X10Y121_CO6;
  assign CLBLM_L_X8Y121_SLICE_X10Y121_D = CLBLM_L_X8Y121_SLICE_X10Y121_DO6;
  assign CLBLM_L_X8Y121_SLICE_X11Y121_A = CLBLM_L_X8Y121_SLICE_X11Y121_AO6;
  assign CLBLM_L_X8Y121_SLICE_X11Y121_B = CLBLM_L_X8Y121_SLICE_X11Y121_BO6;
  assign CLBLM_L_X8Y121_SLICE_X11Y121_C = CLBLM_L_X8Y121_SLICE_X11Y121_CO6;
  assign CLBLM_L_X8Y121_SLICE_X11Y121_D = CLBLM_L_X8Y121_SLICE_X11Y121_DO6;
  assign CLBLM_L_X8Y122_SLICE_X10Y122_A = CLBLM_L_X8Y122_SLICE_X10Y122_AO6;
  assign CLBLM_L_X8Y122_SLICE_X10Y122_B = CLBLM_L_X8Y122_SLICE_X10Y122_BO6;
  assign CLBLM_L_X8Y122_SLICE_X10Y122_C = CLBLM_L_X8Y122_SLICE_X10Y122_CO6;
  assign CLBLM_L_X8Y122_SLICE_X10Y122_D = CLBLM_L_X8Y122_SLICE_X10Y122_DO6;
  assign CLBLM_L_X8Y122_SLICE_X10Y122_AMUX = CLBLM_L_X8Y122_SLICE_X10Y122_AO5;
  assign CLBLM_L_X8Y122_SLICE_X10Y122_BMUX = CLBLM_L_X8Y122_SLICE_X10Y122_BO5;
  assign CLBLM_L_X8Y122_SLICE_X11Y122_A = CLBLM_L_X8Y122_SLICE_X11Y122_AO6;
  assign CLBLM_L_X8Y122_SLICE_X11Y122_B = CLBLM_L_X8Y122_SLICE_X11Y122_BO6;
  assign CLBLM_L_X8Y122_SLICE_X11Y122_C = CLBLM_L_X8Y122_SLICE_X11Y122_CO6;
  assign CLBLM_L_X8Y122_SLICE_X11Y122_D = CLBLM_L_X8Y122_SLICE_X11Y122_DO6;
  assign CLBLM_L_X8Y122_SLICE_X11Y122_AMUX = CLBLM_L_X8Y122_SLICE_X11Y122_A5Q;
  assign CLBLM_L_X8Y123_SLICE_X10Y123_A = CLBLM_L_X8Y123_SLICE_X10Y123_AO6;
  assign CLBLM_L_X8Y123_SLICE_X10Y123_B = CLBLM_L_X8Y123_SLICE_X10Y123_BO6;
  assign CLBLM_L_X8Y123_SLICE_X10Y123_C = CLBLM_L_X8Y123_SLICE_X10Y123_CO6;
  assign CLBLM_L_X8Y123_SLICE_X10Y123_D = CLBLM_L_X8Y123_SLICE_X10Y123_DO6;
  assign CLBLM_L_X8Y123_SLICE_X10Y123_AMUX = CLBLM_L_X8Y123_SLICE_X10Y123_A5Q;
  assign CLBLM_L_X8Y123_SLICE_X10Y123_BMUX = CLBLM_L_X8Y123_SLICE_X10Y123_B5Q;
  assign CLBLM_L_X8Y123_SLICE_X11Y123_A = CLBLM_L_X8Y123_SLICE_X11Y123_AO6;
  assign CLBLM_L_X8Y123_SLICE_X11Y123_B = CLBLM_L_X8Y123_SLICE_X11Y123_BO6;
  assign CLBLM_L_X8Y123_SLICE_X11Y123_C = CLBLM_L_X8Y123_SLICE_X11Y123_CO6;
  assign CLBLM_L_X8Y123_SLICE_X11Y123_D = CLBLM_L_X8Y123_SLICE_X11Y123_DO6;
  assign CLBLM_L_X8Y123_SLICE_X11Y123_AMUX = CLBLM_L_X8Y123_SLICE_X11Y123_A5Q;
  assign CLBLM_L_X8Y128_SLICE_X10Y128_A = CLBLM_L_X8Y128_SLICE_X10Y128_AO6;
  assign CLBLM_L_X8Y128_SLICE_X10Y128_B = CLBLM_L_X8Y128_SLICE_X10Y128_BO6;
  assign CLBLM_L_X8Y128_SLICE_X10Y128_C = CLBLM_L_X8Y128_SLICE_X10Y128_CO6;
  assign CLBLM_L_X8Y128_SLICE_X10Y128_D = CLBLM_L_X8Y128_SLICE_X10Y128_DO6;
  assign CLBLM_L_X8Y128_SLICE_X10Y128_AMUX = CLBLM_L_X8Y128_SLICE_X10Y128_AO5;
  assign CLBLM_L_X8Y128_SLICE_X11Y128_A = CLBLM_L_X8Y128_SLICE_X11Y128_AO6;
  assign CLBLM_L_X8Y128_SLICE_X11Y128_B = CLBLM_L_X8Y128_SLICE_X11Y128_BO6;
  assign CLBLM_L_X8Y128_SLICE_X11Y128_C = CLBLM_L_X8Y128_SLICE_X11Y128_CO6;
  assign CLBLM_L_X8Y128_SLICE_X11Y128_D = CLBLM_L_X8Y128_SLICE_X11Y128_DO6;
  assign CLBLM_L_X8Y133_SLICE_X10Y133_A = CLBLM_L_X8Y133_SLICE_X10Y133_AO6;
  assign CLBLM_L_X8Y133_SLICE_X10Y133_B = CLBLM_L_X8Y133_SLICE_X10Y133_BO6;
  assign CLBLM_L_X8Y133_SLICE_X10Y133_C = CLBLM_L_X8Y133_SLICE_X10Y133_CO6;
  assign CLBLM_L_X8Y133_SLICE_X10Y133_D = CLBLM_L_X8Y133_SLICE_X10Y133_DO6;
  assign CLBLM_L_X8Y133_SLICE_X11Y133_A = CLBLM_L_X8Y133_SLICE_X11Y133_AO6;
  assign CLBLM_L_X8Y133_SLICE_X11Y133_B = CLBLM_L_X8Y133_SLICE_X11Y133_BO6;
  assign CLBLM_L_X8Y133_SLICE_X11Y133_C = CLBLM_L_X8Y133_SLICE_X11Y133_CO6;
  assign CLBLM_L_X8Y133_SLICE_X11Y133_D = CLBLM_L_X8Y133_SLICE_X11Y133_DO6;
  assign CLBLM_L_X8Y133_SLICE_X11Y133_AMUX = CLBLM_L_X8Y133_SLICE_X11Y133_AO5;
  assign CLBLM_L_X10Y110_SLICE_X12Y110_A = CLBLM_L_X10Y110_SLICE_X12Y110_AO6;
  assign CLBLM_L_X10Y110_SLICE_X12Y110_B = CLBLM_L_X10Y110_SLICE_X12Y110_BO6;
  assign CLBLM_L_X10Y110_SLICE_X12Y110_C = CLBLM_L_X10Y110_SLICE_X12Y110_CO6;
  assign CLBLM_L_X10Y110_SLICE_X12Y110_D = CLBLM_L_X10Y110_SLICE_X12Y110_DO6;
  assign CLBLM_L_X10Y110_SLICE_X13Y110_A = CLBLM_L_X10Y110_SLICE_X13Y110_AO6;
  assign CLBLM_L_X10Y110_SLICE_X13Y110_B = CLBLM_L_X10Y110_SLICE_X13Y110_BO6;
  assign CLBLM_L_X10Y110_SLICE_X13Y110_C = CLBLM_L_X10Y110_SLICE_X13Y110_CO6;
  assign CLBLM_L_X10Y110_SLICE_X13Y110_D = CLBLM_L_X10Y110_SLICE_X13Y110_DO6;
  assign CLBLM_L_X10Y110_SLICE_X13Y110_CMUX = CLBLM_L_X10Y110_SLICE_X13Y110_CO5;
  assign CLBLM_L_X10Y110_SLICE_X13Y110_DMUX = CLBLM_L_X10Y110_SLICE_X13Y110_DO5;
  assign CLBLM_L_X10Y111_SLICE_X12Y111_A = CLBLM_L_X10Y111_SLICE_X12Y111_AO6;
  assign CLBLM_L_X10Y111_SLICE_X12Y111_B = CLBLM_L_X10Y111_SLICE_X12Y111_BO6;
  assign CLBLM_L_X10Y111_SLICE_X12Y111_C = CLBLM_L_X10Y111_SLICE_X12Y111_CO6;
  assign CLBLM_L_X10Y111_SLICE_X12Y111_D = CLBLM_L_X10Y111_SLICE_X12Y111_DO6;
  assign CLBLM_L_X10Y111_SLICE_X12Y111_AMUX = CLBLM_L_X10Y111_SLICE_X12Y111_AO5;
  assign CLBLM_L_X10Y111_SLICE_X12Y111_BMUX = CLBLM_L_X10Y111_SLICE_X12Y111_BO5;
  assign CLBLM_L_X10Y111_SLICE_X13Y111_A = CLBLM_L_X10Y111_SLICE_X13Y111_AO6;
  assign CLBLM_L_X10Y111_SLICE_X13Y111_B = CLBLM_L_X10Y111_SLICE_X13Y111_BO6;
  assign CLBLM_L_X10Y111_SLICE_X13Y111_C = CLBLM_L_X10Y111_SLICE_X13Y111_CO6;
  assign CLBLM_L_X10Y111_SLICE_X13Y111_D = CLBLM_L_X10Y111_SLICE_X13Y111_DO6;
  assign CLBLM_L_X10Y111_SLICE_X13Y111_BMUX = CLBLM_L_X10Y111_SLICE_X13Y111_BO5;
  assign CLBLM_L_X10Y111_SLICE_X13Y111_CMUX = CLBLM_L_X10Y111_SLICE_X13Y111_CO5;
  assign CLBLM_L_X10Y112_SLICE_X12Y112_A = CLBLM_L_X10Y112_SLICE_X12Y112_AO6;
  assign CLBLM_L_X10Y112_SLICE_X12Y112_B = CLBLM_L_X10Y112_SLICE_X12Y112_BO6;
  assign CLBLM_L_X10Y112_SLICE_X12Y112_C = CLBLM_L_X10Y112_SLICE_X12Y112_CO6;
  assign CLBLM_L_X10Y112_SLICE_X12Y112_D = CLBLM_L_X10Y112_SLICE_X12Y112_DO6;
  assign CLBLM_L_X10Y112_SLICE_X12Y112_AMUX = CLBLM_L_X10Y112_SLICE_X12Y112_AO5;
  assign CLBLM_L_X10Y112_SLICE_X13Y112_A = CLBLM_L_X10Y112_SLICE_X13Y112_AO6;
  assign CLBLM_L_X10Y112_SLICE_X13Y112_B = CLBLM_L_X10Y112_SLICE_X13Y112_BO6;
  assign CLBLM_L_X10Y112_SLICE_X13Y112_C = CLBLM_L_X10Y112_SLICE_X13Y112_CO6;
  assign CLBLM_L_X10Y112_SLICE_X13Y112_D = CLBLM_L_X10Y112_SLICE_X13Y112_DO6;
  assign CLBLM_L_X10Y113_SLICE_X12Y113_A = CLBLM_L_X10Y113_SLICE_X12Y113_AO6;
  assign CLBLM_L_X10Y113_SLICE_X12Y113_B = CLBLM_L_X10Y113_SLICE_X12Y113_BO6;
  assign CLBLM_L_X10Y113_SLICE_X12Y113_C = CLBLM_L_X10Y113_SLICE_X12Y113_CO6;
  assign CLBLM_L_X10Y113_SLICE_X12Y113_D = CLBLM_L_X10Y113_SLICE_X12Y113_DO6;
  assign CLBLM_L_X10Y113_SLICE_X12Y113_AMUX = CLBLM_L_X10Y113_SLICE_X12Y113_AO5;
  assign CLBLM_L_X10Y113_SLICE_X13Y113_A = CLBLM_L_X10Y113_SLICE_X13Y113_AO6;
  assign CLBLM_L_X10Y113_SLICE_X13Y113_B = CLBLM_L_X10Y113_SLICE_X13Y113_BO6;
  assign CLBLM_L_X10Y113_SLICE_X13Y113_C = CLBLM_L_X10Y113_SLICE_X13Y113_CO6;
  assign CLBLM_L_X10Y113_SLICE_X13Y113_D = CLBLM_L_X10Y113_SLICE_X13Y113_DO6;
  assign CLBLM_L_X10Y113_SLICE_X13Y113_AMUX = CLBLM_L_X10Y113_SLICE_X13Y113_AO5;
  assign CLBLM_L_X10Y113_SLICE_X13Y113_CMUX = CLBLM_L_X10Y113_SLICE_X13Y113_CO6;
  assign CLBLM_L_X10Y114_SLICE_X12Y114_A = CLBLM_L_X10Y114_SLICE_X12Y114_AO6;
  assign CLBLM_L_X10Y114_SLICE_X12Y114_B = CLBLM_L_X10Y114_SLICE_X12Y114_BO6;
  assign CLBLM_L_X10Y114_SLICE_X12Y114_C = CLBLM_L_X10Y114_SLICE_X12Y114_CO6;
  assign CLBLM_L_X10Y114_SLICE_X12Y114_D = CLBLM_L_X10Y114_SLICE_X12Y114_DO6;
  assign CLBLM_L_X10Y114_SLICE_X12Y114_AMUX = CLBLM_L_X10Y114_SLICE_X12Y114_AO5;
  assign CLBLM_L_X10Y114_SLICE_X12Y114_BMUX = CLBLM_L_X10Y114_SLICE_X12Y114_BO5;
  assign CLBLM_L_X10Y114_SLICE_X13Y114_A = CLBLM_L_X10Y114_SLICE_X13Y114_AO6;
  assign CLBLM_L_X10Y114_SLICE_X13Y114_B = CLBLM_L_X10Y114_SLICE_X13Y114_BO6;
  assign CLBLM_L_X10Y114_SLICE_X13Y114_C = CLBLM_L_X10Y114_SLICE_X13Y114_CO6;
  assign CLBLM_L_X10Y114_SLICE_X13Y114_D = CLBLM_L_X10Y114_SLICE_X13Y114_DO6;
  assign CLBLM_L_X10Y114_SLICE_X13Y114_AMUX = CLBLM_L_X10Y114_SLICE_X13Y114_A5Q;
  assign CLBLM_L_X10Y114_SLICE_X13Y114_BMUX = CLBLM_L_X10Y114_SLICE_X13Y114_BO5;
  assign CLBLM_L_X10Y114_SLICE_X13Y114_DMUX = CLBLM_L_X10Y114_SLICE_X13Y114_D5Q;
  assign CLBLM_L_X10Y115_SLICE_X12Y115_A = CLBLM_L_X10Y115_SLICE_X12Y115_AO6;
  assign CLBLM_L_X10Y115_SLICE_X12Y115_B = CLBLM_L_X10Y115_SLICE_X12Y115_BO6;
  assign CLBLM_L_X10Y115_SLICE_X12Y115_C = CLBLM_L_X10Y115_SLICE_X12Y115_CO6;
  assign CLBLM_L_X10Y115_SLICE_X12Y115_D = CLBLM_L_X10Y115_SLICE_X12Y115_DO6;
  assign CLBLM_L_X10Y115_SLICE_X13Y115_A = CLBLM_L_X10Y115_SLICE_X13Y115_AO6;
  assign CLBLM_L_X10Y115_SLICE_X13Y115_B = CLBLM_L_X10Y115_SLICE_X13Y115_BO6;
  assign CLBLM_L_X10Y115_SLICE_X13Y115_C = CLBLM_L_X10Y115_SLICE_X13Y115_CO6;
  assign CLBLM_L_X10Y115_SLICE_X13Y115_D = CLBLM_L_X10Y115_SLICE_X13Y115_DO6;
  assign CLBLM_L_X10Y115_SLICE_X13Y115_AMUX = CLBLM_L_X10Y115_SLICE_X13Y115_AO6;
  assign CLBLM_L_X10Y116_SLICE_X12Y116_A = CLBLM_L_X10Y116_SLICE_X12Y116_AO6;
  assign CLBLM_L_X10Y116_SLICE_X12Y116_B = CLBLM_L_X10Y116_SLICE_X12Y116_BO6;
  assign CLBLM_L_X10Y116_SLICE_X12Y116_C = CLBLM_L_X10Y116_SLICE_X12Y116_CO6;
  assign CLBLM_L_X10Y116_SLICE_X12Y116_D = CLBLM_L_X10Y116_SLICE_X12Y116_DO6;
  assign CLBLM_L_X10Y116_SLICE_X12Y116_AMUX = CLBLM_L_X10Y116_SLICE_X12Y116_A5Q;
  assign CLBLM_L_X10Y116_SLICE_X12Y116_DMUX = CLBLM_L_X10Y116_SLICE_X12Y116_DO5;
  assign CLBLM_L_X10Y116_SLICE_X13Y116_A = CLBLM_L_X10Y116_SLICE_X13Y116_AO6;
  assign CLBLM_L_X10Y116_SLICE_X13Y116_B = CLBLM_L_X10Y116_SLICE_X13Y116_BO6;
  assign CLBLM_L_X10Y116_SLICE_X13Y116_C = CLBLM_L_X10Y116_SLICE_X13Y116_CO6;
  assign CLBLM_L_X10Y116_SLICE_X13Y116_D = CLBLM_L_X10Y116_SLICE_X13Y116_DO6;
  assign CLBLM_L_X10Y116_SLICE_X13Y116_AMUX = CLBLM_L_X10Y116_SLICE_X13Y116_AO5;
  assign CLBLM_L_X10Y116_SLICE_X13Y116_BMUX = CLBLM_L_X10Y116_SLICE_X13Y116_BO5;
  assign CLBLM_L_X10Y116_SLICE_X13Y116_CMUX = CLBLM_L_X10Y116_SLICE_X13Y116_CO5;
  assign CLBLM_L_X10Y117_SLICE_X12Y117_A = CLBLM_L_X10Y117_SLICE_X12Y117_AO6;
  assign CLBLM_L_X10Y117_SLICE_X12Y117_B = CLBLM_L_X10Y117_SLICE_X12Y117_BO6;
  assign CLBLM_L_X10Y117_SLICE_X12Y117_C = CLBLM_L_X10Y117_SLICE_X12Y117_CO6;
  assign CLBLM_L_X10Y117_SLICE_X12Y117_D = CLBLM_L_X10Y117_SLICE_X12Y117_DO6;
  assign CLBLM_L_X10Y117_SLICE_X13Y117_A = CLBLM_L_X10Y117_SLICE_X13Y117_AO6;
  assign CLBLM_L_X10Y117_SLICE_X13Y117_B = CLBLM_L_X10Y117_SLICE_X13Y117_BO6;
  assign CLBLM_L_X10Y117_SLICE_X13Y117_C = CLBLM_L_X10Y117_SLICE_X13Y117_CO6;
  assign CLBLM_L_X10Y117_SLICE_X13Y117_D = CLBLM_L_X10Y117_SLICE_X13Y117_DO6;
  assign CLBLM_L_X10Y118_SLICE_X12Y118_A = CLBLM_L_X10Y118_SLICE_X12Y118_AO6;
  assign CLBLM_L_X10Y118_SLICE_X12Y118_B = CLBLM_L_X10Y118_SLICE_X12Y118_BO6;
  assign CLBLM_L_X10Y118_SLICE_X12Y118_C = CLBLM_L_X10Y118_SLICE_X12Y118_CO6;
  assign CLBLM_L_X10Y118_SLICE_X12Y118_D = CLBLM_L_X10Y118_SLICE_X12Y118_DO6;
  assign CLBLM_L_X10Y118_SLICE_X12Y118_BMUX = CLBLM_L_X10Y118_SLICE_X12Y118_B5Q;
  assign CLBLM_L_X10Y118_SLICE_X13Y118_A = CLBLM_L_X10Y118_SLICE_X13Y118_AO6;
  assign CLBLM_L_X10Y118_SLICE_X13Y118_B = CLBLM_L_X10Y118_SLICE_X13Y118_BO6;
  assign CLBLM_L_X10Y118_SLICE_X13Y118_C = CLBLM_L_X10Y118_SLICE_X13Y118_CO6;
  assign CLBLM_L_X10Y118_SLICE_X13Y118_D = CLBLM_L_X10Y118_SLICE_X13Y118_DO6;
  assign CLBLM_L_X10Y119_SLICE_X12Y119_A = CLBLM_L_X10Y119_SLICE_X12Y119_AO6;
  assign CLBLM_L_X10Y119_SLICE_X12Y119_B = CLBLM_L_X10Y119_SLICE_X12Y119_BO6;
  assign CLBLM_L_X10Y119_SLICE_X12Y119_C = CLBLM_L_X10Y119_SLICE_X12Y119_CO6;
  assign CLBLM_L_X10Y119_SLICE_X12Y119_D = CLBLM_L_X10Y119_SLICE_X12Y119_DO6;
  assign CLBLM_L_X10Y119_SLICE_X13Y119_A = CLBLM_L_X10Y119_SLICE_X13Y119_AO6;
  assign CLBLM_L_X10Y119_SLICE_X13Y119_B = CLBLM_L_X10Y119_SLICE_X13Y119_BO6;
  assign CLBLM_L_X10Y119_SLICE_X13Y119_C = CLBLM_L_X10Y119_SLICE_X13Y119_CO6;
  assign CLBLM_L_X10Y119_SLICE_X13Y119_D = CLBLM_L_X10Y119_SLICE_X13Y119_DO6;
  assign CLBLM_L_X10Y120_SLICE_X12Y120_A = CLBLM_L_X10Y120_SLICE_X12Y120_AO6;
  assign CLBLM_L_X10Y120_SLICE_X12Y120_B = CLBLM_L_X10Y120_SLICE_X12Y120_BO6;
  assign CLBLM_L_X10Y120_SLICE_X12Y120_C = CLBLM_L_X10Y120_SLICE_X12Y120_CO6;
  assign CLBLM_L_X10Y120_SLICE_X12Y120_D = CLBLM_L_X10Y120_SLICE_X12Y120_DO6;
  assign CLBLM_L_X10Y120_SLICE_X13Y120_A = CLBLM_L_X10Y120_SLICE_X13Y120_AO6;
  assign CLBLM_L_X10Y120_SLICE_X13Y120_B = CLBLM_L_X10Y120_SLICE_X13Y120_BO6;
  assign CLBLM_L_X10Y120_SLICE_X13Y120_C = CLBLM_L_X10Y120_SLICE_X13Y120_CO6;
  assign CLBLM_L_X10Y120_SLICE_X13Y120_D = CLBLM_L_X10Y120_SLICE_X13Y120_DO6;
  assign CLBLM_L_X10Y120_SLICE_X13Y120_AMUX = CLBLM_L_X10Y120_SLICE_X13Y120_A5Q;
  assign CLBLM_L_X10Y121_SLICE_X12Y121_A = CLBLM_L_X10Y121_SLICE_X12Y121_AO6;
  assign CLBLM_L_X10Y121_SLICE_X12Y121_B = CLBLM_L_X10Y121_SLICE_X12Y121_BO6;
  assign CLBLM_L_X10Y121_SLICE_X12Y121_C = CLBLM_L_X10Y121_SLICE_X12Y121_CO6;
  assign CLBLM_L_X10Y121_SLICE_X12Y121_D = CLBLM_L_X10Y121_SLICE_X12Y121_DO6;
  assign CLBLM_L_X10Y121_SLICE_X13Y121_A = CLBLM_L_X10Y121_SLICE_X13Y121_AO6;
  assign CLBLM_L_X10Y121_SLICE_X13Y121_B = CLBLM_L_X10Y121_SLICE_X13Y121_BO6;
  assign CLBLM_L_X10Y121_SLICE_X13Y121_C = CLBLM_L_X10Y121_SLICE_X13Y121_CO6;
  assign CLBLM_L_X10Y121_SLICE_X13Y121_D = CLBLM_L_X10Y121_SLICE_X13Y121_DO6;
  assign CLBLM_L_X10Y122_SLICE_X12Y122_A = CLBLM_L_X10Y122_SLICE_X12Y122_AO6;
  assign CLBLM_L_X10Y122_SLICE_X12Y122_B = CLBLM_L_X10Y122_SLICE_X12Y122_BO6;
  assign CLBLM_L_X10Y122_SLICE_X12Y122_C = CLBLM_L_X10Y122_SLICE_X12Y122_CO6;
  assign CLBLM_L_X10Y122_SLICE_X12Y122_D = CLBLM_L_X10Y122_SLICE_X12Y122_DO6;
  assign CLBLM_L_X10Y122_SLICE_X12Y122_CMUX = CLBLM_L_X10Y122_SLICE_X12Y122_CO5;
  assign CLBLM_L_X10Y122_SLICE_X13Y122_A = CLBLM_L_X10Y122_SLICE_X13Y122_AO6;
  assign CLBLM_L_X10Y122_SLICE_X13Y122_B = CLBLM_L_X10Y122_SLICE_X13Y122_BO6;
  assign CLBLM_L_X10Y122_SLICE_X13Y122_C = CLBLM_L_X10Y122_SLICE_X13Y122_CO6;
  assign CLBLM_L_X10Y122_SLICE_X13Y122_D = CLBLM_L_X10Y122_SLICE_X13Y122_DO6;
  assign CLBLM_L_X10Y122_SLICE_X13Y122_AMUX = CLBLM_L_X10Y122_SLICE_X13Y122_A5Q;
  assign CLBLM_L_X10Y122_SLICE_X13Y122_DMUX = CLBLM_L_X10Y122_SLICE_X13Y122_DO6;
  assign CLBLM_L_X10Y123_SLICE_X12Y123_A = CLBLM_L_X10Y123_SLICE_X12Y123_AO6;
  assign CLBLM_L_X10Y123_SLICE_X12Y123_B = CLBLM_L_X10Y123_SLICE_X12Y123_BO6;
  assign CLBLM_L_X10Y123_SLICE_X12Y123_C = CLBLM_L_X10Y123_SLICE_X12Y123_CO6;
  assign CLBLM_L_X10Y123_SLICE_X12Y123_D = CLBLM_L_X10Y123_SLICE_X12Y123_DO6;
  assign CLBLM_L_X10Y123_SLICE_X12Y123_AMUX = CLBLM_L_X10Y123_SLICE_X12Y123_AO5;
  assign CLBLM_L_X10Y123_SLICE_X12Y123_CMUX = CLBLM_L_X10Y123_SLICE_X12Y123_CO6;
  assign CLBLM_L_X10Y123_SLICE_X13Y123_A = CLBLM_L_X10Y123_SLICE_X13Y123_AO6;
  assign CLBLM_L_X10Y123_SLICE_X13Y123_B = CLBLM_L_X10Y123_SLICE_X13Y123_BO6;
  assign CLBLM_L_X10Y123_SLICE_X13Y123_C = CLBLM_L_X10Y123_SLICE_X13Y123_CO6;
  assign CLBLM_L_X10Y123_SLICE_X13Y123_D = CLBLM_L_X10Y123_SLICE_X13Y123_DO6;
  assign CLBLM_L_X10Y124_SLICE_X12Y124_A = CLBLM_L_X10Y124_SLICE_X12Y124_AO6;
  assign CLBLM_L_X10Y124_SLICE_X12Y124_B = CLBLM_L_X10Y124_SLICE_X12Y124_BO6;
  assign CLBLM_L_X10Y124_SLICE_X12Y124_C = CLBLM_L_X10Y124_SLICE_X12Y124_CO6;
  assign CLBLM_L_X10Y124_SLICE_X12Y124_D = CLBLM_L_X10Y124_SLICE_X12Y124_DO6;
  assign CLBLM_L_X10Y124_SLICE_X13Y124_A = CLBLM_L_X10Y124_SLICE_X13Y124_AO6;
  assign CLBLM_L_X10Y124_SLICE_X13Y124_B = CLBLM_L_X10Y124_SLICE_X13Y124_BO6;
  assign CLBLM_L_X10Y124_SLICE_X13Y124_C = CLBLM_L_X10Y124_SLICE_X13Y124_CO6;
  assign CLBLM_L_X10Y124_SLICE_X13Y124_D = CLBLM_L_X10Y124_SLICE_X13Y124_DO6;
  assign CLBLM_L_X10Y124_SLICE_X13Y124_AMUX = CLBLM_L_X10Y124_SLICE_X13Y124_AO5;
  assign CLBLM_L_X10Y124_SLICE_X13Y124_BMUX = CLBLM_L_X10Y124_SLICE_X13Y124_BO5;
  assign CLBLM_L_X10Y124_SLICE_X13Y124_CMUX = CLBLM_L_X10Y124_SLICE_X13Y124_CO5;
  assign CLBLM_L_X10Y126_SLICE_X12Y126_A = CLBLM_L_X10Y126_SLICE_X12Y126_AO6;
  assign CLBLM_L_X10Y126_SLICE_X12Y126_B = CLBLM_L_X10Y126_SLICE_X12Y126_BO6;
  assign CLBLM_L_X10Y126_SLICE_X12Y126_C = CLBLM_L_X10Y126_SLICE_X12Y126_CO6;
  assign CLBLM_L_X10Y126_SLICE_X12Y126_D = CLBLM_L_X10Y126_SLICE_X12Y126_DO6;
  assign CLBLM_L_X10Y126_SLICE_X13Y126_A = CLBLM_L_X10Y126_SLICE_X13Y126_AO6;
  assign CLBLM_L_X10Y126_SLICE_X13Y126_B = CLBLM_L_X10Y126_SLICE_X13Y126_BO6;
  assign CLBLM_L_X10Y126_SLICE_X13Y126_C = CLBLM_L_X10Y126_SLICE_X13Y126_CO6;
  assign CLBLM_L_X10Y126_SLICE_X13Y126_D = CLBLM_L_X10Y126_SLICE_X13Y126_DO6;
  assign CLBLM_L_X10Y127_SLICE_X12Y127_A = CLBLM_L_X10Y127_SLICE_X12Y127_AO6;
  assign CLBLM_L_X10Y127_SLICE_X12Y127_B = CLBLM_L_X10Y127_SLICE_X12Y127_BO6;
  assign CLBLM_L_X10Y127_SLICE_X12Y127_C = CLBLM_L_X10Y127_SLICE_X12Y127_CO6;
  assign CLBLM_L_X10Y127_SLICE_X12Y127_D = CLBLM_L_X10Y127_SLICE_X12Y127_DO6;
  assign CLBLM_L_X10Y127_SLICE_X13Y127_A = CLBLM_L_X10Y127_SLICE_X13Y127_AO6;
  assign CLBLM_L_X10Y127_SLICE_X13Y127_B = CLBLM_L_X10Y127_SLICE_X13Y127_BO6;
  assign CLBLM_L_X10Y127_SLICE_X13Y127_C = CLBLM_L_X10Y127_SLICE_X13Y127_CO6;
  assign CLBLM_L_X10Y127_SLICE_X13Y127_D = CLBLM_L_X10Y127_SLICE_X13Y127_DO6;
  assign CLBLM_L_X10Y128_SLICE_X12Y128_A = CLBLM_L_X10Y128_SLICE_X12Y128_AO6;
  assign CLBLM_L_X10Y128_SLICE_X12Y128_B = CLBLM_L_X10Y128_SLICE_X12Y128_BO6;
  assign CLBLM_L_X10Y128_SLICE_X12Y128_C = CLBLM_L_X10Y128_SLICE_X12Y128_CO6;
  assign CLBLM_L_X10Y128_SLICE_X12Y128_D = CLBLM_L_X10Y128_SLICE_X12Y128_DO6;
  assign CLBLM_L_X10Y128_SLICE_X13Y128_A = CLBLM_L_X10Y128_SLICE_X13Y128_AO6;
  assign CLBLM_L_X10Y128_SLICE_X13Y128_B = CLBLM_L_X10Y128_SLICE_X13Y128_BO6;
  assign CLBLM_L_X10Y128_SLICE_X13Y128_C = CLBLM_L_X10Y128_SLICE_X13Y128_CO6;
  assign CLBLM_L_X10Y128_SLICE_X13Y128_D = CLBLM_L_X10Y128_SLICE_X13Y128_DO6;
  assign CLBLM_L_X10Y128_SLICE_X13Y128_AMUX = CLBLM_L_X10Y128_SLICE_X13Y128_AO5;
  assign CLBLM_L_X12Y115_SLICE_X16Y115_A = CLBLM_L_X12Y115_SLICE_X16Y115_AO6;
  assign CLBLM_L_X12Y115_SLICE_X16Y115_B = CLBLM_L_X12Y115_SLICE_X16Y115_BO6;
  assign CLBLM_L_X12Y115_SLICE_X16Y115_C = CLBLM_L_X12Y115_SLICE_X16Y115_CO6;
  assign CLBLM_L_X12Y115_SLICE_X16Y115_D = CLBLM_L_X12Y115_SLICE_X16Y115_DO6;
  assign CLBLM_L_X12Y115_SLICE_X17Y115_A = CLBLM_L_X12Y115_SLICE_X17Y115_AO6;
  assign CLBLM_L_X12Y115_SLICE_X17Y115_B = CLBLM_L_X12Y115_SLICE_X17Y115_BO6;
  assign CLBLM_L_X12Y115_SLICE_X17Y115_C = CLBLM_L_X12Y115_SLICE_X17Y115_CO6;
  assign CLBLM_L_X12Y115_SLICE_X17Y115_D = CLBLM_L_X12Y115_SLICE_X17Y115_DO6;
  assign CLBLM_L_X12Y118_SLICE_X16Y118_A = CLBLM_L_X12Y118_SLICE_X16Y118_AO6;
  assign CLBLM_L_X12Y118_SLICE_X16Y118_B = CLBLM_L_X12Y118_SLICE_X16Y118_BO6;
  assign CLBLM_L_X12Y118_SLICE_X16Y118_C = CLBLM_L_X12Y118_SLICE_X16Y118_CO6;
  assign CLBLM_L_X12Y118_SLICE_X16Y118_D = CLBLM_L_X12Y118_SLICE_X16Y118_DO6;
  assign CLBLM_L_X12Y118_SLICE_X17Y118_A = CLBLM_L_X12Y118_SLICE_X17Y118_AO6;
  assign CLBLM_L_X12Y118_SLICE_X17Y118_B = CLBLM_L_X12Y118_SLICE_X17Y118_BO6;
  assign CLBLM_L_X12Y118_SLICE_X17Y118_C = CLBLM_L_X12Y118_SLICE_X17Y118_CO6;
  assign CLBLM_L_X12Y118_SLICE_X17Y118_D = CLBLM_L_X12Y118_SLICE_X17Y118_DO6;
  assign CLBLM_L_X12Y119_SLICE_X16Y119_A = CLBLM_L_X12Y119_SLICE_X16Y119_AO6;
  assign CLBLM_L_X12Y119_SLICE_X16Y119_B = CLBLM_L_X12Y119_SLICE_X16Y119_BO6;
  assign CLBLM_L_X12Y119_SLICE_X16Y119_C = CLBLM_L_X12Y119_SLICE_X16Y119_CO6;
  assign CLBLM_L_X12Y119_SLICE_X16Y119_D = CLBLM_L_X12Y119_SLICE_X16Y119_DO6;
  assign CLBLM_L_X12Y119_SLICE_X17Y119_A = CLBLM_L_X12Y119_SLICE_X17Y119_AO6;
  assign CLBLM_L_X12Y119_SLICE_X17Y119_B = CLBLM_L_X12Y119_SLICE_X17Y119_BO6;
  assign CLBLM_L_X12Y119_SLICE_X17Y119_C = CLBLM_L_X12Y119_SLICE_X17Y119_CO6;
  assign CLBLM_L_X12Y119_SLICE_X17Y119_D = CLBLM_L_X12Y119_SLICE_X17Y119_DO6;
  assign CLBLM_L_X12Y119_SLICE_X17Y119_AMUX = CLBLM_L_X12Y119_SLICE_X17Y119_AO5;
  assign CLBLM_L_X12Y120_SLICE_X16Y120_A = CLBLM_L_X12Y120_SLICE_X16Y120_AO6;
  assign CLBLM_L_X12Y120_SLICE_X16Y120_B = CLBLM_L_X12Y120_SLICE_X16Y120_BO6;
  assign CLBLM_L_X12Y120_SLICE_X16Y120_C = CLBLM_L_X12Y120_SLICE_X16Y120_CO6;
  assign CLBLM_L_X12Y120_SLICE_X16Y120_D = CLBLM_L_X12Y120_SLICE_X16Y120_DO6;
  assign CLBLM_L_X12Y120_SLICE_X16Y120_AMUX = CLBLM_L_X12Y120_SLICE_X16Y120_AO5;
  assign CLBLM_L_X12Y120_SLICE_X17Y120_A = CLBLM_L_X12Y120_SLICE_X17Y120_AO6;
  assign CLBLM_L_X12Y120_SLICE_X17Y120_B = CLBLM_L_X12Y120_SLICE_X17Y120_BO6;
  assign CLBLM_L_X12Y120_SLICE_X17Y120_C = CLBLM_L_X12Y120_SLICE_X17Y120_CO6;
  assign CLBLM_L_X12Y120_SLICE_X17Y120_D = CLBLM_L_X12Y120_SLICE_X17Y120_DO6;
  assign CLBLM_L_X12Y120_SLICE_X17Y120_CMUX = CLBLM_L_X12Y120_SLICE_X17Y120_CO5;
  assign CLBLM_L_X12Y120_SLICE_X17Y120_DMUX = CLBLM_L_X12Y120_SLICE_X17Y120_DO5;
  assign CLBLM_L_X12Y121_SLICE_X16Y121_A = CLBLM_L_X12Y121_SLICE_X16Y121_AO6;
  assign CLBLM_L_X12Y121_SLICE_X16Y121_B = CLBLM_L_X12Y121_SLICE_X16Y121_BO6;
  assign CLBLM_L_X12Y121_SLICE_X16Y121_C = CLBLM_L_X12Y121_SLICE_X16Y121_CO6;
  assign CLBLM_L_X12Y121_SLICE_X16Y121_D = CLBLM_L_X12Y121_SLICE_X16Y121_DO6;
  assign CLBLM_L_X12Y121_SLICE_X17Y121_A = CLBLM_L_X12Y121_SLICE_X17Y121_AO6;
  assign CLBLM_L_X12Y121_SLICE_X17Y121_B = CLBLM_L_X12Y121_SLICE_X17Y121_BO6;
  assign CLBLM_L_X12Y121_SLICE_X17Y121_C = CLBLM_L_X12Y121_SLICE_X17Y121_CO6;
  assign CLBLM_L_X12Y121_SLICE_X17Y121_D = CLBLM_L_X12Y121_SLICE_X17Y121_DO6;
  assign CLBLM_R_X3Y110_SLICE_X2Y110_A = CLBLM_R_X3Y110_SLICE_X2Y110_AO6;
  assign CLBLM_R_X3Y110_SLICE_X2Y110_B = CLBLM_R_X3Y110_SLICE_X2Y110_BO6;
  assign CLBLM_R_X3Y110_SLICE_X2Y110_C = CLBLM_R_X3Y110_SLICE_X2Y110_CO6;
  assign CLBLM_R_X3Y110_SLICE_X2Y110_D = CLBLM_R_X3Y110_SLICE_X2Y110_DO6;
  assign CLBLM_R_X3Y110_SLICE_X3Y110_A = CLBLM_R_X3Y110_SLICE_X3Y110_AO6;
  assign CLBLM_R_X3Y110_SLICE_X3Y110_B = CLBLM_R_X3Y110_SLICE_X3Y110_BO6;
  assign CLBLM_R_X3Y110_SLICE_X3Y110_C = CLBLM_R_X3Y110_SLICE_X3Y110_CO6;
  assign CLBLM_R_X3Y110_SLICE_X3Y110_D = CLBLM_R_X3Y110_SLICE_X3Y110_DO6;
  assign CLBLM_R_X3Y111_SLICE_X2Y111_A = CLBLM_R_X3Y111_SLICE_X2Y111_AO6;
  assign CLBLM_R_X3Y111_SLICE_X2Y111_B = CLBLM_R_X3Y111_SLICE_X2Y111_BO6;
  assign CLBLM_R_X3Y111_SLICE_X2Y111_C = CLBLM_R_X3Y111_SLICE_X2Y111_CO6;
  assign CLBLM_R_X3Y111_SLICE_X2Y111_D = CLBLM_R_X3Y111_SLICE_X2Y111_DO6;
  assign CLBLM_R_X3Y111_SLICE_X2Y111_BMUX = CLBLM_R_X3Y111_SLICE_X2Y111_BO5;
  assign CLBLM_R_X3Y111_SLICE_X3Y111_A = CLBLM_R_X3Y111_SLICE_X3Y111_AO6;
  assign CLBLM_R_X3Y111_SLICE_X3Y111_B = CLBLM_R_X3Y111_SLICE_X3Y111_BO6;
  assign CLBLM_R_X3Y111_SLICE_X3Y111_C = CLBLM_R_X3Y111_SLICE_X3Y111_CO6;
  assign CLBLM_R_X3Y111_SLICE_X3Y111_D = CLBLM_R_X3Y111_SLICE_X3Y111_DO6;
  assign CLBLM_R_X3Y111_SLICE_X3Y111_AMUX = CLBLM_R_X3Y111_SLICE_X3Y111_AO5;
  assign CLBLM_R_X3Y111_SLICE_X3Y111_CMUX = CLBLM_R_X3Y111_SLICE_X3Y111_CO6;
  assign CLBLM_R_X3Y112_SLICE_X2Y112_A = CLBLM_R_X3Y112_SLICE_X2Y112_AO6;
  assign CLBLM_R_X3Y112_SLICE_X2Y112_B = CLBLM_R_X3Y112_SLICE_X2Y112_BO6;
  assign CLBLM_R_X3Y112_SLICE_X2Y112_C = CLBLM_R_X3Y112_SLICE_X2Y112_CO6;
  assign CLBLM_R_X3Y112_SLICE_X2Y112_D = CLBLM_R_X3Y112_SLICE_X2Y112_DO6;
  assign CLBLM_R_X3Y112_SLICE_X3Y112_A = CLBLM_R_X3Y112_SLICE_X3Y112_AO6;
  assign CLBLM_R_X3Y112_SLICE_X3Y112_B = CLBLM_R_X3Y112_SLICE_X3Y112_BO6;
  assign CLBLM_R_X3Y112_SLICE_X3Y112_C = CLBLM_R_X3Y112_SLICE_X3Y112_CO6;
  assign CLBLM_R_X3Y112_SLICE_X3Y112_D = CLBLM_R_X3Y112_SLICE_X3Y112_DO6;
  assign CLBLM_R_X3Y112_SLICE_X3Y112_BMUX = CLBLM_R_X3Y112_SLICE_X3Y112_B5Q;
  assign CLBLM_R_X3Y112_SLICE_X3Y112_CMUX = CLBLM_R_X3Y112_SLICE_X3Y112_C5Q;
  assign CLBLM_R_X3Y113_SLICE_X2Y113_A = CLBLM_R_X3Y113_SLICE_X2Y113_AO6;
  assign CLBLM_R_X3Y113_SLICE_X2Y113_B = CLBLM_R_X3Y113_SLICE_X2Y113_BO6;
  assign CLBLM_R_X3Y113_SLICE_X2Y113_C = CLBLM_R_X3Y113_SLICE_X2Y113_CO6;
  assign CLBLM_R_X3Y113_SLICE_X2Y113_D = CLBLM_R_X3Y113_SLICE_X2Y113_DO6;
  assign CLBLM_R_X3Y113_SLICE_X2Y113_CMUX = CLBLM_R_X3Y113_SLICE_X2Y113_CO5;
  assign CLBLM_R_X3Y113_SLICE_X2Y113_DMUX = CLBLM_R_X3Y113_SLICE_X2Y113_DO5;
  assign CLBLM_R_X3Y113_SLICE_X3Y113_A = CLBLM_R_X3Y113_SLICE_X3Y113_AO6;
  assign CLBLM_R_X3Y113_SLICE_X3Y113_B = CLBLM_R_X3Y113_SLICE_X3Y113_BO6;
  assign CLBLM_R_X3Y113_SLICE_X3Y113_C = CLBLM_R_X3Y113_SLICE_X3Y113_CO6;
  assign CLBLM_R_X3Y113_SLICE_X3Y113_D = CLBLM_R_X3Y113_SLICE_X3Y113_DO6;
  assign CLBLM_R_X3Y113_SLICE_X3Y113_BMUX = CLBLM_R_X3Y113_SLICE_X3Y113_BO5;
  assign CLBLM_R_X3Y114_SLICE_X2Y114_A = CLBLM_R_X3Y114_SLICE_X2Y114_AO6;
  assign CLBLM_R_X3Y114_SLICE_X2Y114_B = CLBLM_R_X3Y114_SLICE_X2Y114_BO6;
  assign CLBLM_R_X3Y114_SLICE_X2Y114_C = CLBLM_R_X3Y114_SLICE_X2Y114_CO6;
  assign CLBLM_R_X3Y114_SLICE_X2Y114_D = CLBLM_R_X3Y114_SLICE_X2Y114_DO6;
  assign CLBLM_R_X3Y114_SLICE_X2Y114_AMUX = CLBLM_R_X3Y114_SLICE_X2Y114_AO5;
  assign CLBLM_R_X3Y114_SLICE_X3Y114_A = CLBLM_R_X3Y114_SLICE_X3Y114_AO6;
  assign CLBLM_R_X3Y114_SLICE_X3Y114_B = CLBLM_R_X3Y114_SLICE_X3Y114_BO6;
  assign CLBLM_R_X3Y114_SLICE_X3Y114_C = CLBLM_R_X3Y114_SLICE_X3Y114_CO6;
  assign CLBLM_R_X3Y114_SLICE_X3Y114_D = CLBLM_R_X3Y114_SLICE_X3Y114_DO6;
  assign CLBLM_R_X3Y115_SLICE_X2Y115_A = CLBLM_R_X3Y115_SLICE_X2Y115_AO6;
  assign CLBLM_R_X3Y115_SLICE_X2Y115_B = CLBLM_R_X3Y115_SLICE_X2Y115_BO6;
  assign CLBLM_R_X3Y115_SLICE_X2Y115_C = CLBLM_R_X3Y115_SLICE_X2Y115_CO6;
  assign CLBLM_R_X3Y115_SLICE_X2Y115_D = CLBLM_R_X3Y115_SLICE_X2Y115_DO6;
  assign CLBLM_R_X3Y115_SLICE_X3Y115_A = CLBLM_R_X3Y115_SLICE_X3Y115_AO6;
  assign CLBLM_R_X3Y115_SLICE_X3Y115_B = CLBLM_R_X3Y115_SLICE_X3Y115_BO6;
  assign CLBLM_R_X3Y115_SLICE_X3Y115_C = CLBLM_R_X3Y115_SLICE_X3Y115_CO6;
  assign CLBLM_R_X3Y115_SLICE_X3Y115_D = CLBLM_R_X3Y115_SLICE_X3Y115_DO6;
  assign CLBLM_R_X3Y116_SLICE_X2Y116_A = CLBLM_R_X3Y116_SLICE_X2Y116_AO6;
  assign CLBLM_R_X3Y116_SLICE_X2Y116_B = CLBLM_R_X3Y116_SLICE_X2Y116_BO6;
  assign CLBLM_R_X3Y116_SLICE_X2Y116_C = CLBLM_R_X3Y116_SLICE_X2Y116_CO6;
  assign CLBLM_R_X3Y116_SLICE_X2Y116_D = CLBLM_R_X3Y116_SLICE_X2Y116_DO6;
  assign CLBLM_R_X3Y116_SLICE_X3Y116_A = CLBLM_R_X3Y116_SLICE_X3Y116_AO6;
  assign CLBLM_R_X3Y116_SLICE_X3Y116_B = CLBLM_R_X3Y116_SLICE_X3Y116_BO6;
  assign CLBLM_R_X3Y116_SLICE_X3Y116_C = CLBLM_R_X3Y116_SLICE_X3Y116_CO6;
  assign CLBLM_R_X3Y116_SLICE_X3Y116_D = CLBLM_R_X3Y116_SLICE_X3Y116_DO6;
  assign CLBLM_R_X3Y116_SLICE_X3Y116_AMUX = CLBLM_R_X3Y116_SLICE_X3Y116_A5Q;
  assign CLBLM_R_X3Y117_SLICE_X2Y117_A = CLBLM_R_X3Y117_SLICE_X2Y117_AO6;
  assign CLBLM_R_X3Y117_SLICE_X2Y117_B = CLBLM_R_X3Y117_SLICE_X2Y117_BO6;
  assign CLBLM_R_X3Y117_SLICE_X2Y117_C = CLBLM_R_X3Y117_SLICE_X2Y117_CO6;
  assign CLBLM_R_X3Y117_SLICE_X2Y117_D = CLBLM_R_X3Y117_SLICE_X2Y117_DO6;
  assign CLBLM_R_X3Y117_SLICE_X2Y117_BMUX = CLBLM_R_X3Y117_SLICE_X2Y117_BO5;
  assign CLBLM_R_X3Y117_SLICE_X3Y117_A = CLBLM_R_X3Y117_SLICE_X3Y117_AO6;
  assign CLBLM_R_X3Y117_SLICE_X3Y117_B = CLBLM_R_X3Y117_SLICE_X3Y117_BO6;
  assign CLBLM_R_X3Y117_SLICE_X3Y117_C = CLBLM_R_X3Y117_SLICE_X3Y117_CO6;
  assign CLBLM_R_X3Y117_SLICE_X3Y117_D = CLBLM_R_X3Y117_SLICE_X3Y117_DO6;
  assign CLBLM_R_X3Y117_SLICE_X3Y117_AMUX = CLBLM_R_X3Y117_SLICE_X3Y117_A5Q;
  assign CLBLM_R_X3Y117_SLICE_X3Y117_BMUX = CLBLM_R_X3Y117_SLICE_X3Y117_B5Q;
  assign CLBLM_R_X3Y117_SLICE_X3Y117_CMUX = CLBLM_R_X3Y117_SLICE_X3Y117_C5Q;
  assign CLBLM_R_X3Y118_SLICE_X2Y118_A = CLBLM_R_X3Y118_SLICE_X2Y118_AO6;
  assign CLBLM_R_X3Y118_SLICE_X2Y118_B = CLBLM_R_X3Y118_SLICE_X2Y118_BO6;
  assign CLBLM_R_X3Y118_SLICE_X2Y118_C = CLBLM_R_X3Y118_SLICE_X2Y118_CO6;
  assign CLBLM_R_X3Y118_SLICE_X2Y118_D = CLBLM_R_X3Y118_SLICE_X2Y118_DO6;
  assign CLBLM_R_X3Y118_SLICE_X3Y118_A = CLBLM_R_X3Y118_SLICE_X3Y118_AO6;
  assign CLBLM_R_X3Y118_SLICE_X3Y118_B = CLBLM_R_X3Y118_SLICE_X3Y118_BO6;
  assign CLBLM_R_X3Y118_SLICE_X3Y118_C = CLBLM_R_X3Y118_SLICE_X3Y118_CO6;
  assign CLBLM_R_X3Y118_SLICE_X3Y118_D = CLBLM_R_X3Y118_SLICE_X3Y118_DO6;
  assign CLBLM_R_X3Y119_SLICE_X2Y119_A = CLBLM_R_X3Y119_SLICE_X2Y119_AO6;
  assign CLBLM_R_X3Y119_SLICE_X2Y119_B = CLBLM_R_X3Y119_SLICE_X2Y119_BO6;
  assign CLBLM_R_X3Y119_SLICE_X2Y119_C = CLBLM_R_X3Y119_SLICE_X2Y119_CO6;
  assign CLBLM_R_X3Y119_SLICE_X2Y119_D = CLBLM_R_X3Y119_SLICE_X2Y119_DO6;
  assign CLBLM_R_X3Y119_SLICE_X3Y119_A = CLBLM_R_X3Y119_SLICE_X3Y119_AO6;
  assign CLBLM_R_X3Y119_SLICE_X3Y119_B = CLBLM_R_X3Y119_SLICE_X3Y119_BO6;
  assign CLBLM_R_X3Y119_SLICE_X3Y119_C = CLBLM_R_X3Y119_SLICE_X3Y119_CO6;
  assign CLBLM_R_X3Y119_SLICE_X3Y119_D = CLBLM_R_X3Y119_SLICE_X3Y119_DO6;
  assign CLBLM_R_X3Y120_SLICE_X2Y120_A = CLBLM_R_X3Y120_SLICE_X2Y120_AO6;
  assign CLBLM_R_X3Y120_SLICE_X2Y120_B = CLBLM_R_X3Y120_SLICE_X2Y120_BO6;
  assign CLBLM_R_X3Y120_SLICE_X2Y120_C = CLBLM_R_X3Y120_SLICE_X2Y120_CO6;
  assign CLBLM_R_X3Y120_SLICE_X2Y120_D = CLBLM_R_X3Y120_SLICE_X2Y120_DO6;
  assign CLBLM_R_X3Y120_SLICE_X3Y120_A = CLBLM_R_X3Y120_SLICE_X3Y120_AO6;
  assign CLBLM_R_X3Y120_SLICE_X3Y120_B = CLBLM_R_X3Y120_SLICE_X3Y120_BO6;
  assign CLBLM_R_X3Y120_SLICE_X3Y120_C = CLBLM_R_X3Y120_SLICE_X3Y120_CO6;
  assign CLBLM_R_X3Y120_SLICE_X3Y120_D = CLBLM_R_X3Y120_SLICE_X3Y120_DO6;
  assign CLBLM_R_X3Y120_SLICE_X3Y120_BMUX = CLBLM_R_X3Y120_SLICE_X3Y120_BO6;
  assign CLBLM_R_X3Y120_SLICE_X3Y120_DMUX = CLBLM_R_X3Y120_SLICE_X3Y120_DO6;
  assign CLBLM_R_X3Y121_SLICE_X2Y121_A = CLBLM_R_X3Y121_SLICE_X2Y121_AO6;
  assign CLBLM_R_X3Y121_SLICE_X2Y121_B = CLBLM_R_X3Y121_SLICE_X2Y121_BO6;
  assign CLBLM_R_X3Y121_SLICE_X2Y121_C = CLBLM_R_X3Y121_SLICE_X2Y121_CO6;
  assign CLBLM_R_X3Y121_SLICE_X2Y121_D = CLBLM_R_X3Y121_SLICE_X2Y121_DO6;
  assign CLBLM_R_X3Y121_SLICE_X2Y121_AMUX = CLBLM_R_X3Y121_SLICE_X2Y121_AO5;
  assign CLBLM_R_X3Y121_SLICE_X2Y121_CMUX = CLBLM_R_X3Y121_SLICE_X2Y121_CO6;
  assign CLBLM_R_X3Y121_SLICE_X3Y121_A = CLBLM_R_X3Y121_SLICE_X3Y121_AO6;
  assign CLBLM_R_X3Y121_SLICE_X3Y121_B = CLBLM_R_X3Y121_SLICE_X3Y121_BO6;
  assign CLBLM_R_X3Y121_SLICE_X3Y121_C = CLBLM_R_X3Y121_SLICE_X3Y121_CO6;
  assign CLBLM_R_X3Y121_SLICE_X3Y121_D = CLBLM_R_X3Y121_SLICE_X3Y121_DO6;
  assign CLBLM_R_X3Y121_SLICE_X3Y121_AMUX = CLBLM_R_X3Y121_SLICE_X3Y121_AO6;
  assign CLBLM_R_X3Y121_SLICE_X3Y121_DMUX = CLBLM_R_X3Y121_SLICE_X3Y121_DO6;
  assign CLBLM_R_X3Y122_SLICE_X2Y122_A = CLBLM_R_X3Y122_SLICE_X2Y122_AO6;
  assign CLBLM_R_X3Y122_SLICE_X2Y122_B = CLBLM_R_X3Y122_SLICE_X2Y122_BO6;
  assign CLBLM_R_X3Y122_SLICE_X2Y122_C = CLBLM_R_X3Y122_SLICE_X2Y122_CO6;
  assign CLBLM_R_X3Y122_SLICE_X2Y122_D = CLBLM_R_X3Y122_SLICE_X2Y122_DO6;
  assign CLBLM_R_X3Y122_SLICE_X2Y122_AMUX = CLBLM_R_X3Y122_SLICE_X2Y122_AO5;
  assign CLBLM_R_X3Y122_SLICE_X2Y122_BMUX = CLBLM_R_X3Y122_SLICE_X2Y122_BO5;
  assign CLBLM_R_X3Y122_SLICE_X2Y122_DMUX = CLBLM_R_X3Y122_SLICE_X2Y122_DO6;
  assign CLBLM_R_X3Y122_SLICE_X3Y122_A = CLBLM_R_X3Y122_SLICE_X3Y122_AO6;
  assign CLBLM_R_X3Y122_SLICE_X3Y122_B = CLBLM_R_X3Y122_SLICE_X3Y122_BO6;
  assign CLBLM_R_X3Y122_SLICE_X3Y122_C = CLBLM_R_X3Y122_SLICE_X3Y122_CO6;
  assign CLBLM_R_X3Y122_SLICE_X3Y122_D = CLBLM_R_X3Y122_SLICE_X3Y122_DO6;
  assign CLBLM_R_X3Y122_SLICE_X3Y122_AMUX = CLBLM_R_X3Y122_SLICE_X3Y122_AO5;
  assign CLBLM_R_X3Y123_SLICE_X2Y123_A = CLBLM_R_X3Y123_SLICE_X2Y123_AO6;
  assign CLBLM_R_X3Y123_SLICE_X2Y123_B = CLBLM_R_X3Y123_SLICE_X2Y123_BO6;
  assign CLBLM_R_X3Y123_SLICE_X2Y123_C = CLBLM_R_X3Y123_SLICE_X2Y123_CO6;
  assign CLBLM_R_X3Y123_SLICE_X2Y123_D = CLBLM_R_X3Y123_SLICE_X2Y123_DO6;
  assign CLBLM_R_X3Y123_SLICE_X3Y123_A = CLBLM_R_X3Y123_SLICE_X3Y123_AO6;
  assign CLBLM_R_X3Y123_SLICE_X3Y123_B = CLBLM_R_X3Y123_SLICE_X3Y123_BO6;
  assign CLBLM_R_X3Y123_SLICE_X3Y123_C = CLBLM_R_X3Y123_SLICE_X3Y123_CO6;
  assign CLBLM_R_X3Y123_SLICE_X3Y123_D = CLBLM_R_X3Y123_SLICE_X3Y123_DO6;
  assign CLBLM_R_X3Y123_SLICE_X3Y123_BMUX = CLBLM_R_X3Y123_SLICE_X3Y123_BO5;
  assign CLBLM_R_X3Y124_SLICE_X2Y124_A = CLBLM_R_X3Y124_SLICE_X2Y124_AO6;
  assign CLBLM_R_X3Y124_SLICE_X2Y124_B = CLBLM_R_X3Y124_SLICE_X2Y124_BO6;
  assign CLBLM_R_X3Y124_SLICE_X2Y124_C = CLBLM_R_X3Y124_SLICE_X2Y124_CO6;
  assign CLBLM_R_X3Y124_SLICE_X2Y124_D = CLBLM_R_X3Y124_SLICE_X2Y124_DO6;
  assign CLBLM_R_X3Y124_SLICE_X2Y124_AMUX = CLBLM_R_X3Y124_SLICE_X2Y124_AO5;
  assign CLBLM_R_X3Y124_SLICE_X2Y124_BMUX = CLBLM_R_X3Y124_SLICE_X2Y124_BO5;
  assign CLBLM_R_X3Y124_SLICE_X3Y124_A = CLBLM_R_X3Y124_SLICE_X3Y124_AO6;
  assign CLBLM_R_X3Y124_SLICE_X3Y124_B = CLBLM_R_X3Y124_SLICE_X3Y124_BO6;
  assign CLBLM_R_X3Y124_SLICE_X3Y124_C = CLBLM_R_X3Y124_SLICE_X3Y124_CO6;
  assign CLBLM_R_X3Y124_SLICE_X3Y124_D = CLBLM_R_X3Y124_SLICE_X3Y124_DO6;
  assign CLBLM_R_X5Y109_SLICE_X6Y109_A = CLBLM_R_X5Y109_SLICE_X6Y109_AO6;
  assign CLBLM_R_X5Y109_SLICE_X6Y109_B = CLBLM_R_X5Y109_SLICE_X6Y109_BO6;
  assign CLBLM_R_X5Y109_SLICE_X6Y109_C = CLBLM_R_X5Y109_SLICE_X6Y109_CO6;
  assign CLBLM_R_X5Y109_SLICE_X6Y109_D = CLBLM_R_X5Y109_SLICE_X6Y109_DO6;
  assign CLBLM_R_X5Y109_SLICE_X7Y109_A = CLBLM_R_X5Y109_SLICE_X7Y109_AO6;
  assign CLBLM_R_X5Y109_SLICE_X7Y109_B = CLBLM_R_X5Y109_SLICE_X7Y109_BO6;
  assign CLBLM_R_X5Y109_SLICE_X7Y109_C = CLBLM_R_X5Y109_SLICE_X7Y109_CO6;
  assign CLBLM_R_X5Y109_SLICE_X7Y109_D = CLBLM_R_X5Y109_SLICE_X7Y109_DO6;
  assign CLBLM_R_X5Y110_SLICE_X6Y110_A = CLBLM_R_X5Y110_SLICE_X6Y110_AO6;
  assign CLBLM_R_X5Y110_SLICE_X6Y110_B = CLBLM_R_X5Y110_SLICE_X6Y110_BO6;
  assign CLBLM_R_X5Y110_SLICE_X6Y110_C = CLBLM_R_X5Y110_SLICE_X6Y110_CO6;
  assign CLBLM_R_X5Y110_SLICE_X6Y110_D = CLBLM_R_X5Y110_SLICE_X6Y110_DO6;
  assign CLBLM_R_X5Y110_SLICE_X7Y110_A = CLBLM_R_X5Y110_SLICE_X7Y110_AO6;
  assign CLBLM_R_X5Y110_SLICE_X7Y110_B = CLBLM_R_X5Y110_SLICE_X7Y110_BO6;
  assign CLBLM_R_X5Y110_SLICE_X7Y110_C = CLBLM_R_X5Y110_SLICE_X7Y110_CO6;
  assign CLBLM_R_X5Y110_SLICE_X7Y110_D = CLBLM_R_X5Y110_SLICE_X7Y110_DO6;
  assign CLBLM_R_X5Y110_SLICE_X7Y110_AMUX = CLBLM_R_X5Y110_SLICE_X7Y110_AO5;
  assign CLBLM_R_X5Y110_SLICE_X7Y110_DMUX = CLBLM_R_X5Y110_SLICE_X7Y110_DO5;
  assign CLBLM_R_X5Y111_SLICE_X6Y111_A = CLBLM_R_X5Y111_SLICE_X6Y111_AO6;
  assign CLBLM_R_X5Y111_SLICE_X6Y111_B = CLBLM_R_X5Y111_SLICE_X6Y111_BO6;
  assign CLBLM_R_X5Y111_SLICE_X6Y111_C = CLBLM_R_X5Y111_SLICE_X6Y111_CO6;
  assign CLBLM_R_X5Y111_SLICE_X6Y111_D = CLBLM_R_X5Y111_SLICE_X6Y111_DO6;
  assign CLBLM_R_X5Y111_SLICE_X6Y111_CMUX = CLBLM_R_X5Y111_SLICE_X6Y111_C5Q;
  assign CLBLM_R_X5Y111_SLICE_X7Y111_A = CLBLM_R_X5Y111_SLICE_X7Y111_AO6;
  assign CLBLM_R_X5Y111_SLICE_X7Y111_B = CLBLM_R_X5Y111_SLICE_X7Y111_BO6;
  assign CLBLM_R_X5Y111_SLICE_X7Y111_C = CLBLM_R_X5Y111_SLICE_X7Y111_CO6;
  assign CLBLM_R_X5Y111_SLICE_X7Y111_D = CLBLM_R_X5Y111_SLICE_X7Y111_DO6;
  assign CLBLM_R_X5Y111_SLICE_X7Y111_CMUX = CLBLM_R_X5Y111_SLICE_X7Y111_CO5;
  assign CLBLM_R_X5Y112_SLICE_X6Y112_A = CLBLM_R_X5Y112_SLICE_X6Y112_AO6;
  assign CLBLM_R_X5Y112_SLICE_X6Y112_B = CLBLM_R_X5Y112_SLICE_X6Y112_BO6;
  assign CLBLM_R_X5Y112_SLICE_X6Y112_C = CLBLM_R_X5Y112_SLICE_X6Y112_CO6;
  assign CLBLM_R_X5Y112_SLICE_X6Y112_D = CLBLM_R_X5Y112_SLICE_X6Y112_DO6;
  assign CLBLM_R_X5Y112_SLICE_X6Y112_BMUX = CLBLM_R_X5Y112_SLICE_X6Y112_BO5;
  assign CLBLM_R_X5Y112_SLICE_X7Y112_A = CLBLM_R_X5Y112_SLICE_X7Y112_AO6;
  assign CLBLM_R_X5Y112_SLICE_X7Y112_B = CLBLM_R_X5Y112_SLICE_X7Y112_BO6;
  assign CLBLM_R_X5Y112_SLICE_X7Y112_C = CLBLM_R_X5Y112_SLICE_X7Y112_CO6;
  assign CLBLM_R_X5Y112_SLICE_X7Y112_D = CLBLM_R_X5Y112_SLICE_X7Y112_DO6;
  assign CLBLM_R_X5Y112_SLICE_X7Y112_AMUX = CLBLM_R_X5Y112_SLICE_X7Y112_AO5;
  assign CLBLM_R_X5Y113_SLICE_X6Y113_A = CLBLM_R_X5Y113_SLICE_X6Y113_AO6;
  assign CLBLM_R_X5Y113_SLICE_X6Y113_B = CLBLM_R_X5Y113_SLICE_X6Y113_BO6;
  assign CLBLM_R_X5Y113_SLICE_X6Y113_C = CLBLM_R_X5Y113_SLICE_X6Y113_CO6;
  assign CLBLM_R_X5Y113_SLICE_X6Y113_D = CLBLM_R_X5Y113_SLICE_X6Y113_DO6;
  assign CLBLM_R_X5Y113_SLICE_X6Y113_DMUX = CLBLM_R_X5Y113_SLICE_X6Y113_DO5;
  assign CLBLM_R_X5Y113_SLICE_X7Y113_A = CLBLM_R_X5Y113_SLICE_X7Y113_AO6;
  assign CLBLM_R_X5Y113_SLICE_X7Y113_B = CLBLM_R_X5Y113_SLICE_X7Y113_BO6;
  assign CLBLM_R_X5Y113_SLICE_X7Y113_C = CLBLM_R_X5Y113_SLICE_X7Y113_CO6;
  assign CLBLM_R_X5Y113_SLICE_X7Y113_D = CLBLM_R_X5Y113_SLICE_X7Y113_DO6;
  assign CLBLM_R_X5Y113_SLICE_X7Y113_AMUX = CLBLM_R_X5Y113_SLICE_X7Y113_A5Q;
  assign CLBLM_R_X5Y113_SLICE_X7Y113_BMUX = CLBLM_R_X5Y113_SLICE_X7Y113_BO6;
  assign CLBLM_R_X5Y114_SLICE_X6Y114_A = CLBLM_R_X5Y114_SLICE_X6Y114_AO6;
  assign CLBLM_R_X5Y114_SLICE_X6Y114_B = CLBLM_R_X5Y114_SLICE_X6Y114_BO6;
  assign CLBLM_R_X5Y114_SLICE_X6Y114_C = CLBLM_R_X5Y114_SLICE_X6Y114_CO6;
  assign CLBLM_R_X5Y114_SLICE_X6Y114_D = CLBLM_R_X5Y114_SLICE_X6Y114_DO6;
  assign CLBLM_R_X5Y114_SLICE_X7Y114_A = CLBLM_R_X5Y114_SLICE_X7Y114_AO6;
  assign CLBLM_R_X5Y114_SLICE_X7Y114_B = CLBLM_R_X5Y114_SLICE_X7Y114_BO6;
  assign CLBLM_R_X5Y114_SLICE_X7Y114_C = CLBLM_R_X5Y114_SLICE_X7Y114_CO6;
  assign CLBLM_R_X5Y114_SLICE_X7Y114_D = CLBLM_R_X5Y114_SLICE_X7Y114_DO6;
  assign CLBLM_R_X5Y114_SLICE_X7Y114_BMUX = CLBLM_R_X5Y114_SLICE_X7Y114_BO5;
  assign CLBLM_R_X5Y115_SLICE_X6Y115_A = CLBLM_R_X5Y115_SLICE_X6Y115_AO6;
  assign CLBLM_R_X5Y115_SLICE_X6Y115_B = CLBLM_R_X5Y115_SLICE_X6Y115_BO6;
  assign CLBLM_R_X5Y115_SLICE_X6Y115_C = CLBLM_R_X5Y115_SLICE_X6Y115_CO6;
  assign CLBLM_R_X5Y115_SLICE_X6Y115_D = CLBLM_R_X5Y115_SLICE_X6Y115_DO6;
  assign CLBLM_R_X5Y115_SLICE_X6Y115_CMUX = CLBLM_R_X5Y115_SLICE_X6Y115_CO5;
  assign CLBLM_R_X5Y115_SLICE_X7Y115_A = CLBLM_R_X5Y115_SLICE_X7Y115_AO6;
  assign CLBLM_R_X5Y115_SLICE_X7Y115_B = CLBLM_R_X5Y115_SLICE_X7Y115_BO6;
  assign CLBLM_R_X5Y115_SLICE_X7Y115_C = CLBLM_R_X5Y115_SLICE_X7Y115_CO6;
  assign CLBLM_R_X5Y115_SLICE_X7Y115_D = CLBLM_R_X5Y115_SLICE_X7Y115_DO6;
  assign CLBLM_R_X5Y115_SLICE_X7Y115_AMUX = CLBLM_R_X5Y115_SLICE_X7Y115_A5Q;
  assign CLBLM_R_X5Y115_SLICE_X7Y115_CMUX = CLBLM_R_X5Y115_SLICE_X7Y115_CO5;
  assign CLBLM_R_X5Y116_SLICE_X6Y116_A = CLBLM_R_X5Y116_SLICE_X6Y116_AO6;
  assign CLBLM_R_X5Y116_SLICE_X6Y116_B = CLBLM_R_X5Y116_SLICE_X6Y116_BO6;
  assign CLBLM_R_X5Y116_SLICE_X6Y116_C = CLBLM_R_X5Y116_SLICE_X6Y116_CO6;
  assign CLBLM_R_X5Y116_SLICE_X6Y116_D = CLBLM_R_X5Y116_SLICE_X6Y116_DO6;
  assign CLBLM_R_X5Y116_SLICE_X6Y116_AMUX = CLBLM_R_X5Y116_SLICE_X6Y116_A5Q;
  assign CLBLM_R_X5Y116_SLICE_X6Y116_CMUX = CLBLM_R_X5Y116_SLICE_X6Y116_CO5;
  assign CLBLM_R_X5Y116_SLICE_X7Y116_A = CLBLM_R_X5Y116_SLICE_X7Y116_AO6;
  assign CLBLM_R_X5Y116_SLICE_X7Y116_B = CLBLM_R_X5Y116_SLICE_X7Y116_BO6;
  assign CLBLM_R_X5Y116_SLICE_X7Y116_C = CLBLM_R_X5Y116_SLICE_X7Y116_CO6;
  assign CLBLM_R_X5Y116_SLICE_X7Y116_D = CLBLM_R_X5Y116_SLICE_X7Y116_DO6;
  assign CLBLM_R_X5Y116_SLICE_X7Y116_AMUX = CLBLM_R_X5Y116_SLICE_X7Y116_A5Q;
  assign CLBLM_R_X5Y116_SLICE_X7Y116_BMUX = CLBLM_R_X5Y116_SLICE_X7Y116_BO5;
  assign CLBLM_R_X5Y117_SLICE_X6Y117_A = CLBLM_R_X5Y117_SLICE_X6Y117_AO6;
  assign CLBLM_R_X5Y117_SLICE_X6Y117_B = CLBLM_R_X5Y117_SLICE_X6Y117_BO6;
  assign CLBLM_R_X5Y117_SLICE_X6Y117_C = CLBLM_R_X5Y117_SLICE_X6Y117_CO6;
  assign CLBLM_R_X5Y117_SLICE_X6Y117_D = CLBLM_R_X5Y117_SLICE_X6Y117_DO6;
  assign CLBLM_R_X5Y117_SLICE_X6Y117_DMUX = CLBLM_R_X5Y117_SLICE_X6Y117_D5Q;
  assign CLBLM_R_X5Y117_SLICE_X7Y117_A = CLBLM_R_X5Y117_SLICE_X7Y117_AO6;
  assign CLBLM_R_X5Y117_SLICE_X7Y117_B = CLBLM_R_X5Y117_SLICE_X7Y117_BO6;
  assign CLBLM_R_X5Y117_SLICE_X7Y117_C = CLBLM_R_X5Y117_SLICE_X7Y117_CO6;
  assign CLBLM_R_X5Y117_SLICE_X7Y117_D = CLBLM_R_X5Y117_SLICE_X7Y117_DO6;
  assign CLBLM_R_X5Y118_SLICE_X6Y118_A = CLBLM_R_X5Y118_SLICE_X6Y118_AO6;
  assign CLBLM_R_X5Y118_SLICE_X6Y118_B = CLBLM_R_X5Y118_SLICE_X6Y118_BO6;
  assign CLBLM_R_X5Y118_SLICE_X6Y118_C = CLBLM_R_X5Y118_SLICE_X6Y118_CO6;
  assign CLBLM_R_X5Y118_SLICE_X6Y118_D = CLBLM_R_X5Y118_SLICE_X6Y118_DO6;
  assign CLBLM_R_X5Y118_SLICE_X7Y118_A = CLBLM_R_X5Y118_SLICE_X7Y118_AO6;
  assign CLBLM_R_X5Y118_SLICE_X7Y118_B = CLBLM_R_X5Y118_SLICE_X7Y118_BO6;
  assign CLBLM_R_X5Y118_SLICE_X7Y118_C = CLBLM_R_X5Y118_SLICE_X7Y118_CO6;
  assign CLBLM_R_X5Y118_SLICE_X7Y118_D = CLBLM_R_X5Y118_SLICE_X7Y118_DO6;
  assign CLBLM_R_X5Y118_SLICE_X7Y118_BMUX = CLBLM_R_X5Y118_SLICE_X7Y118_BO5;
  assign CLBLM_R_X5Y119_SLICE_X6Y119_A = CLBLM_R_X5Y119_SLICE_X6Y119_AO6;
  assign CLBLM_R_X5Y119_SLICE_X6Y119_B = CLBLM_R_X5Y119_SLICE_X6Y119_BO6;
  assign CLBLM_R_X5Y119_SLICE_X6Y119_C = CLBLM_R_X5Y119_SLICE_X6Y119_CO6;
  assign CLBLM_R_X5Y119_SLICE_X6Y119_D = CLBLM_R_X5Y119_SLICE_X6Y119_DO6;
  assign CLBLM_R_X5Y119_SLICE_X6Y119_BMUX = CLBLM_R_X5Y119_SLICE_X6Y119_B5Q;
  assign CLBLM_R_X5Y119_SLICE_X7Y119_A = CLBLM_R_X5Y119_SLICE_X7Y119_AO6;
  assign CLBLM_R_X5Y119_SLICE_X7Y119_B = CLBLM_R_X5Y119_SLICE_X7Y119_BO6;
  assign CLBLM_R_X5Y119_SLICE_X7Y119_C = CLBLM_R_X5Y119_SLICE_X7Y119_CO6;
  assign CLBLM_R_X5Y119_SLICE_X7Y119_D = CLBLM_R_X5Y119_SLICE_X7Y119_DO6;
  assign CLBLM_R_X5Y120_SLICE_X6Y120_A = CLBLM_R_X5Y120_SLICE_X6Y120_AO6;
  assign CLBLM_R_X5Y120_SLICE_X6Y120_B = CLBLM_R_X5Y120_SLICE_X6Y120_BO6;
  assign CLBLM_R_X5Y120_SLICE_X6Y120_C = CLBLM_R_X5Y120_SLICE_X6Y120_CO6;
  assign CLBLM_R_X5Y120_SLICE_X6Y120_D = CLBLM_R_X5Y120_SLICE_X6Y120_DO6;
  assign CLBLM_R_X5Y120_SLICE_X6Y120_AMUX = CLBLM_R_X5Y120_SLICE_X6Y120_A5Q;
  assign CLBLM_R_X5Y120_SLICE_X6Y120_CMUX = CLBLM_R_X5Y120_SLICE_X6Y120_CO6;
  assign CLBLM_R_X5Y120_SLICE_X7Y120_A = CLBLM_R_X5Y120_SLICE_X7Y120_AO6;
  assign CLBLM_R_X5Y120_SLICE_X7Y120_B = CLBLM_R_X5Y120_SLICE_X7Y120_BO6;
  assign CLBLM_R_X5Y120_SLICE_X7Y120_C = CLBLM_R_X5Y120_SLICE_X7Y120_CO6;
  assign CLBLM_R_X5Y120_SLICE_X7Y120_D = CLBLM_R_X5Y120_SLICE_X7Y120_DO6;
  assign CLBLM_R_X5Y120_SLICE_X7Y120_DMUX = CLBLM_R_X5Y120_SLICE_X7Y120_DO5;
  assign CLBLM_R_X5Y121_SLICE_X6Y121_A = CLBLM_R_X5Y121_SLICE_X6Y121_AO6;
  assign CLBLM_R_X5Y121_SLICE_X6Y121_B = CLBLM_R_X5Y121_SLICE_X6Y121_BO6;
  assign CLBLM_R_X5Y121_SLICE_X6Y121_C = CLBLM_R_X5Y121_SLICE_X6Y121_CO6;
  assign CLBLM_R_X5Y121_SLICE_X6Y121_D = CLBLM_R_X5Y121_SLICE_X6Y121_DO6;
  assign CLBLM_R_X5Y121_SLICE_X6Y121_AMUX = CLBLM_R_X5Y121_SLICE_X6Y121_A5Q;
  assign CLBLM_R_X5Y121_SLICE_X6Y121_BMUX = CLBLM_R_X5Y121_SLICE_X6Y121_B5Q;
  assign CLBLM_R_X5Y121_SLICE_X6Y121_CMUX = CLBLM_R_X5Y121_SLICE_X6Y121_CO5;
  assign CLBLM_R_X5Y121_SLICE_X7Y121_A = CLBLM_R_X5Y121_SLICE_X7Y121_AO6;
  assign CLBLM_R_X5Y121_SLICE_X7Y121_B = CLBLM_R_X5Y121_SLICE_X7Y121_BO6;
  assign CLBLM_R_X5Y121_SLICE_X7Y121_C = CLBLM_R_X5Y121_SLICE_X7Y121_CO6;
  assign CLBLM_R_X5Y121_SLICE_X7Y121_D = CLBLM_R_X5Y121_SLICE_X7Y121_DO6;
  assign CLBLM_R_X5Y121_SLICE_X7Y121_AMUX = CLBLM_R_X5Y121_SLICE_X7Y121_A5Q;
  assign CLBLM_R_X5Y122_SLICE_X6Y122_A = CLBLM_R_X5Y122_SLICE_X6Y122_AO6;
  assign CLBLM_R_X5Y122_SLICE_X6Y122_B = CLBLM_R_X5Y122_SLICE_X6Y122_BO6;
  assign CLBLM_R_X5Y122_SLICE_X6Y122_C = CLBLM_R_X5Y122_SLICE_X6Y122_CO6;
  assign CLBLM_R_X5Y122_SLICE_X6Y122_D = CLBLM_R_X5Y122_SLICE_X6Y122_DO6;
  assign CLBLM_R_X5Y122_SLICE_X6Y122_AMUX = CLBLM_R_X5Y122_SLICE_X6Y122_AO5;
  assign CLBLM_R_X5Y122_SLICE_X6Y122_CMUX = CLBLM_R_X5Y122_SLICE_X6Y122_CO6;
  assign CLBLM_R_X5Y122_SLICE_X7Y122_A = CLBLM_R_X5Y122_SLICE_X7Y122_AO6;
  assign CLBLM_R_X5Y122_SLICE_X7Y122_B = CLBLM_R_X5Y122_SLICE_X7Y122_BO6;
  assign CLBLM_R_X5Y122_SLICE_X7Y122_C = CLBLM_R_X5Y122_SLICE_X7Y122_CO6;
  assign CLBLM_R_X5Y122_SLICE_X7Y122_D = CLBLM_R_X5Y122_SLICE_X7Y122_DO6;
  assign CLBLM_R_X5Y122_SLICE_X7Y122_AMUX = CLBLM_R_X5Y122_SLICE_X7Y122_A5Q;
  assign CLBLM_R_X5Y123_SLICE_X6Y123_A = CLBLM_R_X5Y123_SLICE_X6Y123_AO6;
  assign CLBLM_R_X5Y123_SLICE_X6Y123_B = CLBLM_R_X5Y123_SLICE_X6Y123_BO6;
  assign CLBLM_R_X5Y123_SLICE_X6Y123_C = CLBLM_R_X5Y123_SLICE_X6Y123_CO6;
  assign CLBLM_R_X5Y123_SLICE_X6Y123_D = CLBLM_R_X5Y123_SLICE_X6Y123_DO6;
  assign CLBLM_R_X5Y123_SLICE_X6Y123_DMUX = CLBLM_R_X5Y123_SLICE_X6Y123_DO5;
  assign CLBLM_R_X5Y123_SLICE_X7Y123_A = CLBLM_R_X5Y123_SLICE_X7Y123_AO6;
  assign CLBLM_R_X5Y123_SLICE_X7Y123_B = CLBLM_R_X5Y123_SLICE_X7Y123_BO6;
  assign CLBLM_R_X5Y123_SLICE_X7Y123_C = CLBLM_R_X5Y123_SLICE_X7Y123_CO6;
  assign CLBLM_R_X5Y123_SLICE_X7Y123_D = CLBLM_R_X5Y123_SLICE_X7Y123_DO6;
  assign CLBLM_R_X5Y124_SLICE_X6Y124_A = CLBLM_R_X5Y124_SLICE_X6Y124_AO6;
  assign CLBLM_R_X5Y124_SLICE_X6Y124_B = CLBLM_R_X5Y124_SLICE_X6Y124_BO6;
  assign CLBLM_R_X5Y124_SLICE_X6Y124_C = CLBLM_R_X5Y124_SLICE_X6Y124_CO6;
  assign CLBLM_R_X5Y124_SLICE_X6Y124_D = CLBLM_R_X5Y124_SLICE_X6Y124_DO6;
  assign CLBLM_R_X5Y124_SLICE_X7Y124_A = CLBLM_R_X5Y124_SLICE_X7Y124_AO6;
  assign CLBLM_R_X5Y124_SLICE_X7Y124_B = CLBLM_R_X5Y124_SLICE_X7Y124_BO6;
  assign CLBLM_R_X5Y124_SLICE_X7Y124_C = CLBLM_R_X5Y124_SLICE_X7Y124_CO6;
  assign CLBLM_R_X5Y124_SLICE_X7Y124_D = CLBLM_R_X5Y124_SLICE_X7Y124_DO6;
  assign CLBLM_R_X5Y125_SLICE_X6Y125_A = CLBLM_R_X5Y125_SLICE_X6Y125_AO6;
  assign CLBLM_R_X5Y125_SLICE_X6Y125_B = CLBLM_R_X5Y125_SLICE_X6Y125_BO6;
  assign CLBLM_R_X5Y125_SLICE_X6Y125_C = CLBLM_R_X5Y125_SLICE_X6Y125_CO6;
  assign CLBLM_R_X5Y125_SLICE_X6Y125_D = CLBLM_R_X5Y125_SLICE_X6Y125_DO6;
  assign CLBLM_R_X5Y125_SLICE_X6Y125_AMUX = CLBLM_R_X5Y125_SLICE_X6Y125_A5Q;
  assign CLBLM_R_X5Y125_SLICE_X6Y125_BMUX = CLBLM_R_X5Y125_SLICE_X6Y125_BO5;
  assign CLBLM_R_X5Y125_SLICE_X6Y125_CMUX = CLBLM_R_X5Y125_SLICE_X6Y125_CO5;
  assign CLBLM_R_X5Y125_SLICE_X7Y125_A = CLBLM_R_X5Y125_SLICE_X7Y125_AO6;
  assign CLBLM_R_X5Y125_SLICE_X7Y125_B = CLBLM_R_X5Y125_SLICE_X7Y125_BO6;
  assign CLBLM_R_X5Y125_SLICE_X7Y125_C = CLBLM_R_X5Y125_SLICE_X7Y125_CO6;
  assign CLBLM_R_X5Y125_SLICE_X7Y125_D = CLBLM_R_X5Y125_SLICE_X7Y125_DO6;
  assign CLBLM_R_X7Y109_SLICE_X8Y109_A = CLBLM_R_X7Y109_SLICE_X8Y109_AO6;
  assign CLBLM_R_X7Y109_SLICE_X8Y109_B = CLBLM_R_X7Y109_SLICE_X8Y109_BO6;
  assign CLBLM_R_X7Y109_SLICE_X8Y109_C = CLBLM_R_X7Y109_SLICE_X8Y109_CO6;
  assign CLBLM_R_X7Y109_SLICE_X8Y109_D = CLBLM_R_X7Y109_SLICE_X8Y109_DO6;
  assign CLBLM_R_X7Y109_SLICE_X9Y109_A = CLBLM_R_X7Y109_SLICE_X9Y109_AO6;
  assign CLBLM_R_X7Y109_SLICE_X9Y109_B = CLBLM_R_X7Y109_SLICE_X9Y109_BO6;
  assign CLBLM_R_X7Y109_SLICE_X9Y109_C = CLBLM_R_X7Y109_SLICE_X9Y109_CO6;
  assign CLBLM_R_X7Y109_SLICE_X9Y109_D = CLBLM_R_X7Y109_SLICE_X9Y109_DO6;
  assign CLBLM_R_X7Y110_SLICE_X8Y110_A = CLBLM_R_X7Y110_SLICE_X8Y110_AO6;
  assign CLBLM_R_X7Y110_SLICE_X8Y110_B = CLBLM_R_X7Y110_SLICE_X8Y110_BO6;
  assign CLBLM_R_X7Y110_SLICE_X8Y110_C = CLBLM_R_X7Y110_SLICE_X8Y110_CO6;
  assign CLBLM_R_X7Y110_SLICE_X8Y110_D = CLBLM_R_X7Y110_SLICE_X8Y110_DO6;
  assign CLBLM_R_X7Y110_SLICE_X8Y110_DMUX = CLBLM_R_X7Y110_SLICE_X8Y110_DO5;
  assign CLBLM_R_X7Y110_SLICE_X9Y110_A = CLBLM_R_X7Y110_SLICE_X9Y110_AO6;
  assign CLBLM_R_X7Y110_SLICE_X9Y110_B = CLBLM_R_X7Y110_SLICE_X9Y110_BO6;
  assign CLBLM_R_X7Y110_SLICE_X9Y110_C = CLBLM_R_X7Y110_SLICE_X9Y110_CO6;
  assign CLBLM_R_X7Y110_SLICE_X9Y110_D = CLBLM_R_X7Y110_SLICE_X9Y110_DO6;
  assign CLBLM_R_X7Y111_SLICE_X8Y111_A = CLBLM_R_X7Y111_SLICE_X8Y111_AO6;
  assign CLBLM_R_X7Y111_SLICE_X8Y111_B = CLBLM_R_X7Y111_SLICE_X8Y111_BO6;
  assign CLBLM_R_X7Y111_SLICE_X8Y111_C = CLBLM_R_X7Y111_SLICE_X8Y111_CO6;
  assign CLBLM_R_X7Y111_SLICE_X8Y111_D = CLBLM_R_X7Y111_SLICE_X8Y111_DO6;
  assign CLBLM_R_X7Y111_SLICE_X9Y111_A = CLBLM_R_X7Y111_SLICE_X9Y111_AO6;
  assign CLBLM_R_X7Y111_SLICE_X9Y111_B = CLBLM_R_X7Y111_SLICE_X9Y111_BO6;
  assign CLBLM_R_X7Y111_SLICE_X9Y111_C = CLBLM_R_X7Y111_SLICE_X9Y111_CO6;
  assign CLBLM_R_X7Y111_SLICE_X9Y111_D = CLBLM_R_X7Y111_SLICE_X9Y111_DO6;
  assign CLBLM_R_X7Y111_SLICE_X9Y111_AMUX = CLBLM_R_X7Y111_SLICE_X9Y111_AO5;
  assign CLBLM_R_X7Y111_SLICE_X9Y111_BMUX = CLBLM_R_X7Y111_SLICE_X9Y111_BO5;
  assign CLBLM_R_X7Y112_SLICE_X8Y112_A = CLBLM_R_X7Y112_SLICE_X8Y112_AO6;
  assign CLBLM_R_X7Y112_SLICE_X8Y112_B = CLBLM_R_X7Y112_SLICE_X8Y112_BO6;
  assign CLBLM_R_X7Y112_SLICE_X8Y112_C = CLBLM_R_X7Y112_SLICE_X8Y112_CO6;
  assign CLBLM_R_X7Y112_SLICE_X8Y112_D = CLBLM_R_X7Y112_SLICE_X8Y112_DO6;
  assign CLBLM_R_X7Y112_SLICE_X9Y112_A = CLBLM_R_X7Y112_SLICE_X9Y112_AO6;
  assign CLBLM_R_X7Y112_SLICE_X9Y112_B = CLBLM_R_X7Y112_SLICE_X9Y112_BO6;
  assign CLBLM_R_X7Y112_SLICE_X9Y112_C = CLBLM_R_X7Y112_SLICE_X9Y112_CO6;
  assign CLBLM_R_X7Y112_SLICE_X9Y112_D = CLBLM_R_X7Y112_SLICE_X9Y112_DO6;
  assign CLBLM_R_X7Y113_SLICE_X8Y113_A = CLBLM_R_X7Y113_SLICE_X8Y113_AO6;
  assign CLBLM_R_X7Y113_SLICE_X8Y113_B = CLBLM_R_X7Y113_SLICE_X8Y113_BO6;
  assign CLBLM_R_X7Y113_SLICE_X8Y113_C = CLBLM_R_X7Y113_SLICE_X8Y113_CO6;
  assign CLBLM_R_X7Y113_SLICE_X8Y113_D = CLBLM_R_X7Y113_SLICE_X8Y113_DO6;
  assign CLBLM_R_X7Y113_SLICE_X8Y113_BMUX = CLBLM_R_X7Y113_SLICE_X8Y113_BO5;
  assign CLBLM_R_X7Y113_SLICE_X9Y113_A = CLBLM_R_X7Y113_SLICE_X9Y113_AO6;
  assign CLBLM_R_X7Y113_SLICE_X9Y113_B = CLBLM_R_X7Y113_SLICE_X9Y113_BO6;
  assign CLBLM_R_X7Y113_SLICE_X9Y113_C = CLBLM_R_X7Y113_SLICE_X9Y113_CO6;
  assign CLBLM_R_X7Y113_SLICE_X9Y113_D = CLBLM_R_X7Y113_SLICE_X9Y113_DO6;
  assign CLBLM_R_X7Y113_SLICE_X9Y113_AMUX = CLBLM_R_X7Y113_SLICE_X9Y113_A5Q;
  assign CLBLM_R_X7Y114_SLICE_X8Y114_A = CLBLM_R_X7Y114_SLICE_X8Y114_AO6;
  assign CLBLM_R_X7Y114_SLICE_X8Y114_B = CLBLM_R_X7Y114_SLICE_X8Y114_BO6;
  assign CLBLM_R_X7Y114_SLICE_X8Y114_C = CLBLM_R_X7Y114_SLICE_X8Y114_CO6;
  assign CLBLM_R_X7Y114_SLICE_X8Y114_D = CLBLM_R_X7Y114_SLICE_X8Y114_DO6;
  assign CLBLM_R_X7Y114_SLICE_X9Y114_A = CLBLM_R_X7Y114_SLICE_X9Y114_AO6;
  assign CLBLM_R_X7Y114_SLICE_X9Y114_B = CLBLM_R_X7Y114_SLICE_X9Y114_BO6;
  assign CLBLM_R_X7Y114_SLICE_X9Y114_C = CLBLM_R_X7Y114_SLICE_X9Y114_CO6;
  assign CLBLM_R_X7Y114_SLICE_X9Y114_D = CLBLM_R_X7Y114_SLICE_X9Y114_DO6;
  assign CLBLM_R_X7Y115_SLICE_X8Y115_A = CLBLM_R_X7Y115_SLICE_X8Y115_AO6;
  assign CLBLM_R_X7Y115_SLICE_X8Y115_B = CLBLM_R_X7Y115_SLICE_X8Y115_BO6;
  assign CLBLM_R_X7Y115_SLICE_X8Y115_C = CLBLM_R_X7Y115_SLICE_X8Y115_CO6;
  assign CLBLM_R_X7Y115_SLICE_X8Y115_D = CLBLM_R_X7Y115_SLICE_X8Y115_DO6;
  assign CLBLM_R_X7Y115_SLICE_X8Y115_AMUX = CLBLM_R_X7Y115_SLICE_X8Y115_A5Q;
  assign CLBLM_R_X7Y115_SLICE_X8Y115_DMUX = CLBLM_R_X7Y115_SLICE_X8Y115_DO5;
  assign CLBLM_R_X7Y115_SLICE_X9Y115_A = CLBLM_R_X7Y115_SLICE_X9Y115_AO6;
  assign CLBLM_R_X7Y115_SLICE_X9Y115_B = CLBLM_R_X7Y115_SLICE_X9Y115_BO6;
  assign CLBLM_R_X7Y115_SLICE_X9Y115_C = CLBLM_R_X7Y115_SLICE_X9Y115_CO6;
  assign CLBLM_R_X7Y115_SLICE_X9Y115_D = CLBLM_R_X7Y115_SLICE_X9Y115_DO6;
  assign CLBLM_R_X7Y115_SLICE_X9Y115_BMUX = CLBLM_R_X7Y115_SLICE_X9Y115_B5Q;
  assign CLBLM_R_X7Y115_SLICE_X9Y115_CMUX = CLBLM_R_X7Y115_SLICE_X9Y115_C5Q;
  assign CLBLM_R_X7Y116_SLICE_X8Y116_A = CLBLM_R_X7Y116_SLICE_X8Y116_AO6;
  assign CLBLM_R_X7Y116_SLICE_X8Y116_B = CLBLM_R_X7Y116_SLICE_X8Y116_BO6;
  assign CLBLM_R_X7Y116_SLICE_X8Y116_C = CLBLM_R_X7Y116_SLICE_X8Y116_CO6;
  assign CLBLM_R_X7Y116_SLICE_X8Y116_D = CLBLM_R_X7Y116_SLICE_X8Y116_DO6;
  assign CLBLM_R_X7Y116_SLICE_X9Y116_A = CLBLM_R_X7Y116_SLICE_X9Y116_AO6;
  assign CLBLM_R_X7Y116_SLICE_X9Y116_B = CLBLM_R_X7Y116_SLICE_X9Y116_BO6;
  assign CLBLM_R_X7Y116_SLICE_X9Y116_C = CLBLM_R_X7Y116_SLICE_X9Y116_CO6;
  assign CLBLM_R_X7Y116_SLICE_X9Y116_D = CLBLM_R_X7Y116_SLICE_X9Y116_DO6;
  assign CLBLM_R_X7Y117_SLICE_X8Y117_A = CLBLM_R_X7Y117_SLICE_X8Y117_AO6;
  assign CLBLM_R_X7Y117_SLICE_X8Y117_B = CLBLM_R_X7Y117_SLICE_X8Y117_BO6;
  assign CLBLM_R_X7Y117_SLICE_X8Y117_C = CLBLM_R_X7Y117_SLICE_X8Y117_CO6;
  assign CLBLM_R_X7Y117_SLICE_X8Y117_D = CLBLM_R_X7Y117_SLICE_X8Y117_DO6;
  assign CLBLM_R_X7Y117_SLICE_X8Y117_AMUX = CLBLM_R_X7Y117_SLICE_X8Y117_A5Q;
  assign CLBLM_R_X7Y117_SLICE_X8Y117_DMUX = CLBLM_R_X7Y117_SLICE_X8Y117_DO5;
  assign CLBLM_R_X7Y117_SLICE_X9Y117_A = CLBLM_R_X7Y117_SLICE_X9Y117_AO6;
  assign CLBLM_R_X7Y117_SLICE_X9Y117_B = CLBLM_R_X7Y117_SLICE_X9Y117_BO6;
  assign CLBLM_R_X7Y117_SLICE_X9Y117_C = CLBLM_R_X7Y117_SLICE_X9Y117_CO6;
  assign CLBLM_R_X7Y117_SLICE_X9Y117_D = CLBLM_R_X7Y117_SLICE_X9Y117_DO6;
  assign CLBLM_R_X7Y118_SLICE_X8Y118_A = CLBLM_R_X7Y118_SLICE_X8Y118_AO6;
  assign CLBLM_R_X7Y118_SLICE_X8Y118_B = CLBLM_R_X7Y118_SLICE_X8Y118_BO6;
  assign CLBLM_R_X7Y118_SLICE_X8Y118_C = CLBLM_R_X7Y118_SLICE_X8Y118_CO6;
  assign CLBLM_R_X7Y118_SLICE_X8Y118_D = CLBLM_R_X7Y118_SLICE_X8Y118_DO6;
  assign CLBLM_R_X7Y118_SLICE_X9Y118_A = CLBLM_R_X7Y118_SLICE_X9Y118_AO6;
  assign CLBLM_R_X7Y118_SLICE_X9Y118_B = CLBLM_R_X7Y118_SLICE_X9Y118_BO6;
  assign CLBLM_R_X7Y118_SLICE_X9Y118_C = CLBLM_R_X7Y118_SLICE_X9Y118_CO6;
  assign CLBLM_R_X7Y118_SLICE_X9Y118_D = CLBLM_R_X7Y118_SLICE_X9Y118_DO6;
  assign CLBLM_R_X7Y119_SLICE_X8Y119_A = CLBLM_R_X7Y119_SLICE_X8Y119_AO6;
  assign CLBLM_R_X7Y119_SLICE_X8Y119_B = CLBLM_R_X7Y119_SLICE_X8Y119_BO6;
  assign CLBLM_R_X7Y119_SLICE_X8Y119_C = CLBLM_R_X7Y119_SLICE_X8Y119_CO6;
  assign CLBLM_R_X7Y119_SLICE_X8Y119_D = CLBLM_R_X7Y119_SLICE_X8Y119_DO6;
  assign CLBLM_R_X7Y119_SLICE_X8Y119_CMUX = CLBLM_R_X7Y119_SLICE_X8Y119_C5Q;
  assign CLBLM_R_X7Y119_SLICE_X8Y119_DMUX = CLBLM_R_X7Y119_SLICE_X8Y119_D5Q;
  assign CLBLM_R_X7Y119_SLICE_X9Y119_A = CLBLM_R_X7Y119_SLICE_X9Y119_AO6;
  assign CLBLM_R_X7Y119_SLICE_X9Y119_B = CLBLM_R_X7Y119_SLICE_X9Y119_BO6;
  assign CLBLM_R_X7Y119_SLICE_X9Y119_C = CLBLM_R_X7Y119_SLICE_X9Y119_CO6;
  assign CLBLM_R_X7Y119_SLICE_X9Y119_D = CLBLM_R_X7Y119_SLICE_X9Y119_DO6;
  assign CLBLM_R_X7Y119_SLICE_X9Y119_DMUX = CLBLM_R_X7Y119_SLICE_X9Y119_DO5;
  assign CLBLM_R_X7Y120_SLICE_X8Y120_A = CLBLM_R_X7Y120_SLICE_X8Y120_AO6;
  assign CLBLM_R_X7Y120_SLICE_X8Y120_B = CLBLM_R_X7Y120_SLICE_X8Y120_BO6;
  assign CLBLM_R_X7Y120_SLICE_X8Y120_C = CLBLM_R_X7Y120_SLICE_X8Y120_CO6;
  assign CLBLM_R_X7Y120_SLICE_X8Y120_D = CLBLM_R_X7Y120_SLICE_X8Y120_DO6;
  assign CLBLM_R_X7Y120_SLICE_X9Y120_A = CLBLM_R_X7Y120_SLICE_X9Y120_AO6;
  assign CLBLM_R_X7Y120_SLICE_X9Y120_B = CLBLM_R_X7Y120_SLICE_X9Y120_BO6;
  assign CLBLM_R_X7Y120_SLICE_X9Y120_C = CLBLM_R_X7Y120_SLICE_X9Y120_CO6;
  assign CLBLM_R_X7Y120_SLICE_X9Y120_D = CLBLM_R_X7Y120_SLICE_X9Y120_DO6;
  assign CLBLM_R_X7Y120_SLICE_X9Y120_AMUX = CLBLM_R_X7Y120_SLICE_X9Y120_A5Q;
  assign CLBLM_R_X7Y120_SLICE_X9Y120_DMUX = CLBLM_R_X7Y120_SLICE_X9Y120_D5Q;
  assign CLBLM_R_X7Y121_SLICE_X8Y121_A = CLBLM_R_X7Y121_SLICE_X8Y121_AO6;
  assign CLBLM_R_X7Y121_SLICE_X8Y121_B = CLBLM_R_X7Y121_SLICE_X8Y121_BO6;
  assign CLBLM_R_X7Y121_SLICE_X8Y121_C = CLBLM_R_X7Y121_SLICE_X8Y121_CO6;
  assign CLBLM_R_X7Y121_SLICE_X8Y121_D = CLBLM_R_X7Y121_SLICE_X8Y121_DO6;
  assign CLBLM_R_X7Y121_SLICE_X8Y121_CMUX = CLBLM_R_X7Y121_SLICE_X8Y121_C5Q;
  assign CLBLM_R_X7Y121_SLICE_X9Y121_A = CLBLM_R_X7Y121_SLICE_X9Y121_AO6;
  assign CLBLM_R_X7Y121_SLICE_X9Y121_B = CLBLM_R_X7Y121_SLICE_X9Y121_BO6;
  assign CLBLM_R_X7Y121_SLICE_X9Y121_C = CLBLM_R_X7Y121_SLICE_X9Y121_CO6;
  assign CLBLM_R_X7Y121_SLICE_X9Y121_D = CLBLM_R_X7Y121_SLICE_X9Y121_DO6;
  assign CLBLM_R_X7Y121_SLICE_X9Y121_AMUX = CLBLM_R_X7Y121_SLICE_X9Y121_A5Q;
  assign CLBLM_R_X7Y121_SLICE_X9Y121_CMUX = CLBLM_R_X7Y121_SLICE_X9Y121_CO5;
  assign CLBLM_R_X7Y121_SLICE_X9Y121_DMUX = CLBLM_R_X7Y121_SLICE_X9Y121_DO5;
  assign CLBLM_R_X7Y122_SLICE_X8Y122_A = CLBLM_R_X7Y122_SLICE_X8Y122_AO6;
  assign CLBLM_R_X7Y122_SLICE_X8Y122_B = CLBLM_R_X7Y122_SLICE_X8Y122_BO6;
  assign CLBLM_R_X7Y122_SLICE_X8Y122_C = CLBLM_R_X7Y122_SLICE_X8Y122_CO6;
  assign CLBLM_R_X7Y122_SLICE_X8Y122_D = CLBLM_R_X7Y122_SLICE_X8Y122_DO6;
  assign CLBLM_R_X7Y122_SLICE_X9Y122_A = CLBLM_R_X7Y122_SLICE_X9Y122_AO6;
  assign CLBLM_R_X7Y122_SLICE_X9Y122_B = CLBLM_R_X7Y122_SLICE_X9Y122_BO6;
  assign CLBLM_R_X7Y122_SLICE_X9Y122_C = CLBLM_R_X7Y122_SLICE_X9Y122_CO6;
  assign CLBLM_R_X7Y122_SLICE_X9Y122_D = CLBLM_R_X7Y122_SLICE_X9Y122_DO6;
  assign CLBLM_R_X7Y122_SLICE_X9Y122_AMUX = CLBLM_R_X7Y122_SLICE_X9Y122_A5Q;
  assign CLBLM_R_X7Y123_SLICE_X8Y123_A = CLBLM_R_X7Y123_SLICE_X8Y123_AO6;
  assign CLBLM_R_X7Y123_SLICE_X8Y123_B = CLBLM_R_X7Y123_SLICE_X8Y123_BO6;
  assign CLBLM_R_X7Y123_SLICE_X8Y123_C = CLBLM_R_X7Y123_SLICE_X8Y123_CO6;
  assign CLBLM_R_X7Y123_SLICE_X8Y123_D = CLBLM_R_X7Y123_SLICE_X8Y123_DO6;
  assign CLBLM_R_X7Y123_SLICE_X9Y123_A = CLBLM_R_X7Y123_SLICE_X9Y123_AO6;
  assign CLBLM_R_X7Y123_SLICE_X9Y123_B = CLBLM_R_X7Y123_SLICE_X9Y123_BO6;
  assign CLBLM_R_X7Y123_SLICE_X9Y123_C = CLBLM_R_X7Y123_SLICE_X9Y123_CO6;
  assign CLBLM_R_X7Y123_SLICE_X9Y123_D = CLBLM_R_X7Y123_SLICE_X9Y123_DO6;
  assign CLBLM_R_X7Y123_SLICE_X9Y123_BMUX = CLBLM_R_X7Y123_SLICE_X9Y123_BO5;
  assign CLBLM_R_X7Y124_SLICE_X8Y124_A = CLBLM_R_X7Y124_SLICE_X8Y124_AO6;
  assign CLBLM_R_X7Y124_SLICE_X8Y124_B = CLBLM_R_X7Y124_SLICE_X8Y124_BO6;
  assign CLBLM_R_X7Y124_SLICE_X8Y124_C = CLBLM_R_X7Y124_SLICE_X8Y124_CO6;
  assign CLBLM_R_X7Y124_SLICE_X8Y124_D = CLBLM_R_X7Y124_SLICE_X8Y124_DO6;
  assign CLBLM_R_X7Y124_SLICE_X8Y124_AMUX = CLBLM_R_X7Y124_SLICE_X8Y124_A5Q;
  assign CLBLM_R_X7Y124_SLICE_X8Y124_DMUX = CLBLM_R_X7Y124_SLICE_X8Y124_DO5;
  assign CLBLM_R_X7Y124_SLICE_X9Y124_A = CLBLM_R_X7Y124_SLICE_X9Y124_AO6;
  assign CLBLM_R_X7Y124_SLICE_X9Y124_B = CLBLM_R_X7Y124_SLICE_X9Y124_BO6;
  assign CLBLM_R_X7Y124_SLICE_X9Y124_C = CLBLM_R_X7Y124_SLICE_X9Y124_CO6;
  assign CLBLM_R_X7Y124_SLICE_X9Y124_D = CLBLM_R_X7Y124_SLICE_X9Y124_DO6;
  assign CLBLM_R_X7Y125_SLICE_X8Y125_A = CLBLM_R_X7Y125_SLICE_X8Y125_AO6;
  assign CLBLM_R_X7Y125_SLICE_X8Y125_B = CLBLM_R_X7Y125_SLICE_X8Y125_BO6;
  assign CLBLM_R_X7Y125_SLICE_X8Y125_C = CLBLM_R_X7Y125_SLICE_X8Y125_CO6;
  assign CLBLM_R_X7Y125_SLICE_X8Y125_D = CLBLM_R_X7Y125_SLICE_X8Y125_DO6;
  assign CLBLM_R_X7Y125_SLICE_X9Y125_A = CLBLM_R_X7Y125_SLICE_X9Y125_AO6;
  assign CLBLM_R_X7Y125_SLICE_X9Y125_B = CLBLM_R_X7Y125_SLICE_X9Y125_BO6;
  assign CLBLM_R_X7Y125_SLICE_X9Y125_C = CLBLM_R_X7Y125_SLICE_X9Y125_CO6;
  assign CLBLM_R_X7Y125_SLICE_X9Y125_D = CLBLM_R_X7Y125_SLICE_X9Y125_DO6;
  assign CLBLM_R_X7Y127_SLICE_X8Y127_A = CLBLM_R_X7Y127_SLICE_X8Y127_AO6;
  assign CLBLM_R_X7Y127_SLICE_X8Y127_B = CLBLM_R_X7Y127_SLICE_X8Y127_BO6;
  assign CLBLM_R_X7Y127_SLICE_X8Y127_C = CLBLM_R_X7Y127_SLICE_X8Y127_CO6;
  assign CLBLM_R_X7Y127_SLICE_X8Y127_D = CLBLM_R_X7Y127_SLICE_X8Y127_DO6;
  assign CLBLM_R_X7Y127_SLICE_X9Y127_A = CLBLM_R_X7Y127_SLICE_X9Y127_AO6;
  assign CLBLM_R_X7Y127_SLICE_X9Y127_B = CLBLM_R_X7Y127_SLICE_X9Y127_BO6;
  assign CLBLM_R_X7Y127_SLICE_X9Y127_C = CLBLM_R_X7Y127_SLICE_X9Y127_CO6;
  assign CLBLM_R_X7Y127_SLICE_X9Y127_D = CLBLM_R_X7Y127_SLICE_X9Y127_DO6;
  assign CLBLM_R_X7Y128_SLICE_X8Y128_A = CLBLM_R_X7Y128_SLICE_X8Y128_AO6;
  assign CLBLM_R_X7Y128_SLICE_X8Y128_B = CLBLM_R_X7Y128_SLICE_X8Y128_BO6;
  assign CLBLM_R_X7Y128_SLICE_X8Y128_C = CLBLM_R_X7Y128_SLICE_X8Y128_CO6;
  assign CLBLM_R_X7Y128_SLICE_X8Y128_D = CLBLM_R_X7Y128_SLICE_X8Y128_DO6;
  assign CLBLM_R_X7Y128_SLICE_X8Y128_AMUX = CLBLM_R_X7Y128_SLICE_X8Y128_AO5;
  assign CLBLM_R_X7Y128_SLICE_X9Y128_A = CLBLM_R_X7Y128_SLICE_X9Y128_AO6;
  assign CLBLM_R_X7Y128_SLICE_X9Y128_B = CLBLM_R_X7Y128_SLICE_X9Y128_BO6;
  assign CLBLM_R_X7Y128_SLICE_X9Y128_C = CLBLM_R_X7Y128_SLICE_X9Y128_CO6;
  assign CLBLM_R_X7Y128_SLICE_X9Y128_D = CLBLM_R_X7Y128_SLICE_X9Y128_DO6;
  assign CLBLM_R_X7Y151_SLICE_X8Y151_A = CLBLM_R_X7Y151_SLICE_X8Y151_AO6;
  assign CLBLM_R_X7Y151_SLICE_X8Y151_B = CLBLM_R_X7Y151_SLICE_X8Y151_BO6;
  assign CLBLM_R_X7Y151_SLICE_X8Y151_C = CLBLM_R_X7Y151_SLICE_X8Y151_CO6;
  assign CLBLM_R_X7Y151_SLICE_X8Y151_D = CLBLM_R_X7Y151_SLICE_X8Y151_DO6;
  assign CLBLM_R_X7Y151_SLICE_X9Y151_A = CLBLM_R_X7Y151_SLICE_X9Y151_AO6;
  assign CLBLM_R_X7Y151_SLICE_X9Y151_B = CLBLM_R_X7Y151_SLICE_X9Y151_BO6;
  assign CLBLM_R_X7Y151_SLICE_X9Y151_C = CLBLM_R_X7Y151_SLICE_X9Y151_CO6;
  assign CLBLM_R_X7Y151_SLICE_X9Y151_D = CLBLM_R_X7Y151_SLICE_X9Y151_DO6;
  assign CLBLM_R_X11Y113_SLICE_X14Y113_A = CLBLM_R_X11Y113_SLICE_X14Y113_AO6;
  assign CLBLM_R_X11Y113_SLICE_X14Y113_B = CLBLM_R_X11Y113_SLICE_X14Y113_BO6;
  assign CLBLM_R_X11Y113_SLICE_X14Y113_C = CLBLM_R_X11Y113_SLICE_X14Y113_CO6;
  assign CLBLM_R_X11Y113_SLICE_X14Y113_D = CLBLM_R_X11Y113_SLICE_X14Y113_DO6;
  assign CLBLM_R_X11Y113_SLICE_X15Y113_A = CLBLM_R_X11Y113_SLICE_X15Y113_AO6;
  assign CLBLM_R_X11Y113_SLICE_X15Y113_B = CLBLM_R_X11Y113_SLICE_X15Y113_BO6;
  assign CLBLM_R_X11Y113_SLICE_X15Y113_C = CLBLM_R_X11Y113_SLICE_X15Y113_CO6;
  assign CLBLM_R_X11Y113_SLICE_X15Y113_D = CLBLM_R_X11Y113_SLICE_X15Y113_DO6;
  assign CLBLM_R_X11Y114_SLICE_X14Y114_A = CLBLM_R_X11Y114_SLICE_X14Y114_AO6;
  assign CLBLM_R_X11Y114_SLICE_X14Y114_B = CLBLM_R_X11Y114_SLICE_X14Y114_BO6;
  assign CLBLM_R_X11Y114_SLICE_X14Y114_C = CLBLM_R_X11Y114_SLICE_X14Y114_CO6;
  assign CLBLM_R_X11Y114_SLICE_X14Y114_D = CLBLM_R_X11Y114_SLICE_X14Y114_DO6;
  assign CLBLM_R_X11Y114_SLICE_X14Y114_DMUX = CLBLM_R_X11Y114_SLICE_X14Y114_D5Q;
  assign CLBLM_R_X11Y114_SLICE_X15Y114_A = CLBLM_R_X11Y114_SLICE_X15Y114_AO6;
  assign CLBLM_R_X11Y114_SLICE_X15Y114_B = CLBLM_R_X11Y114_SLICE_X15Y114_BO6;
  assign CLBLM_R_X11Y114_SLICE_X15Y114_C = CLBLM_R_X11Y114_SLICE_X15Y114_CO6;
  assign CLBLM_R_X11Y114_SLICE_X15Y114_D = CLBLM_R_X11Y114_SLICE_X15Y114_DO6;
  assign CLBLM_R_X11Y115_SLICE_X14Y115_A = CLBLM_R_X11Y115_SLICE_X14Y115_AO6;
  assign CLBLM_R_X11Y115_SLICE_X14Y115_B = CLBLM_R_X11Y115_SLICE_X14Y115_BO6;
  assign CLBLM_R_X11Y115_SLICE_X14Y115_C = CLBLM_R_X11Y115_SLICE_X14Y115_CO6;
  assign CLBLM_R_X11Y115_SLICE_X14Y115_D = CLBLM_R_X11Y115_SLICE_X14Y115_DO6;
  assign CLBLM_R_X11Y115_SLICE_X15Y115_A = CLBLM_R_X11Y115_SLICE_X15Y115_AO6;
  assign CLBLM_R_X11Y115_SLICE_X15Y115_B = CLBLM_R_X11Y115_SLICE_X15Y115_BO6;
  assign CLBLM_R_X11Y115_SLICE_X15Y115_C = CLBLM_R_X11Y115_SLICE_X15Y115_CO6;
  assign CLBLM_R_X11Y115_SLICE_X15Y115_D = CLBLM_R_X11Y115_SLICE_X15Y115_DO6;
  assign CLBLM_R_X11Y116_SLICE_X14Y116_A = CLBLM_R_X11Y116_SLICE_X14Y116_AO6;
  assign CLBLM_R_X11Y116_SLICE_X14Y116_B = CLBLM_R_X11Y116_SLICE_X14Y116_BO6;
  assign CLBLM_R_X11Y116_SLICE_X14Y116_C = CLBLM_R_X11Y116_SLICE_X14Y116_CO6;
  assign CLBLM_R_X11Y116_SLICE_X14Y116_D = CLBLM_R_X11Y116_SLICE_X14Y116_DO6;
  assign CLBLM_R_X11Y116_SLICE_X14Y116_BMUX = CLBLM_R_X11Y116_SLICE_X14Y116_BO5;
  assign CLBLM_R_X11Y116_SLICE_X15Y116_A = CLBLM_R_X11Y116_SLICE_X15Y116_AO6;
  assign CLBLM_R_X11Y116_SLICE_X15Y116_B = CLBLM_R_X11Y116_SLICE_X15Y116_BO6;
  assign CLBLM_R_X11Y116_SLICE_X15Y116_C = CLBLM_R_X11Y116_SLICE_X15Y116_CO6;
  assign CLBLM_R_X11Y116_SLICE_X15Y116_D = CLBLM_R_X11Y116_SLICE_X15Y116_DO6;
  assign CLBLM_R_X11Y117_SLICE_X14Y117_A = CLBLM_R_X11Y117_SLICE_X14Y117_AO6;
  assign CLBLM_R_X11Y117_SLICE_X14Y117_B = CLBLM_R_X11Y117_SLICE_X14Y117_BO6;
  assign CLBLM_R_X11Y117_SLICE_X14Y117_C = CLBLM_R_X11Y117_SLICE_X14Y117_CO6;
  assign CLBLM_R_X11Y117_SLICE_X14Y117_D = CLBLM_R_X11Y117_SLICE_X14Y117_DO6;
  assign CLBLM_R_X11Y117_SLICE_X14Y117_DMUX = CLBLM_R_X11Y117_SLICE_X14Y117_DO5;
  assign CLBLM_R_X11Y117_SLICE_X15Y117_A = CLBLM_R_X11Y117_SLICE_X15Y117_AO6;
  assign CLBLM_R_X11Y117_SLICE_X15Y117_B = CLBLM_R_X11Y117_SLICE_X15Y117_BO6;
  assign CLBLM_R_X11Y117_SLICE_X15Y117_C = CLBLM_R_X11Y117_SLICE_X15Y117_CO6;
  assign CLBLM_R_X11Y117_SLICE_X15Y117_D = CLBLM_R_X11Y117_SLICE_X15Y117_DO6;
  assign CLBLM_R_X11Y118_SLICE_X14Y118_A = CLBLM_R_X11Y118_SLICE_X14Y118_AO6;
  assign CLBLM_R_X11Y118_SLICE_X14Y118_B = CLBLM_R_X11Y118_SLICE_X14Y118_BO6;
  assign CLBLM_R_X11Y118_SLICE_X14Y118_C = CLBLM_R_X11Y118_SLICE_X14Y118_CO6;
  assign CLBLM_R_X11Y118_SLICE_X14Y118_D = CLBLM_R_X11Y118_SLICE_X14Y118_DO6;
  assign CLBLM_R_X11Y118_SLICE_X14Y118_DMUX = CLBLM_R_X11Y118_SLICE_X14Y118_DO5;
  assign CLBLM_R_X11Y118_SLICE_X15Y118_A = CLBLM_R_X11Y118_SLICE_X15Y118_AO6;
  assign CLBLM_R_X11Y118_SLICE_X15Y118_B = CLBLM_R_X11Y118_SLICE_X15Y118_BO6;
  assign CLBLM_R_X11Y118_SLICE_X15Y118_C = CLBLM_R_X11Y118_SLICE_X15Y118_CO6;
  assign CLBLM_R_X11Y118_SLICE_X15Y118_D = CLBLM_R_X11Y118_SLICE_X15Y118_DO6;
  assign CLBLM_R_X11Y119_SLICE_X14Y119_A = CLBLM_R_X11Y119_SLICE_X14Y119_AO6;
  assign CLBLM_R_X11Y119_SLICE_X14Y119_B = CLBLM_R_X11Y119_SLICE_X14Y119_BO6;
  assign CLBLM_R_X11Y119_SLICE_X14Y119_C = CLBLM_R_X11Y119_SLICE_X14Y119_CO6;
  assign CLBLM_R_X11Y119_SLICE_X14Y119_D = CLBLM_R_X11Y119_SLICE_X14Y119_DO6;
  assign CLBLM_R_X11Y119_SLICE_X14Y119_AMUX = CLBLM_R_X11Y119_SLICE_X14Y119_AO5;
  assign CLBLM_R_X11Y119_SLICE_X14Y119_BMUX = CLBLM_R_X11Y119_SLICE_X14Y119_BO5;
  assign CLBLM_R_X11Y119_SLICE_X14Y119_CMUX = CLBLM_R_X11Y119_SLICE_X14Y119_CO5;
  assign CLBLM_R_X11Y119_SLICE_X15Y119_A = CLBLM_R_X11Y119_SLICE_X15Y119_AO6;
  assign CLBLM_R_X11Y119_SLICE_X15Y119_B = CLBLM_R_X11Y119_SLICE_X15Y119_BO6;
  assign CLBLM_R_X11Y119_SLICE_X15Y119_C = CLBLM_R_X11Y119_SLICE_X15Y119_CO6;
  assign CLBLM_R_X11Y119_SLICE_X15Y119_D = CLBLM_R_X11Y119_SLICE_X15Y119_DO6;
  assign CLBLM_R_X11Y120_SLICE_X14Y120_A = CLBLM_R_X11Y120_SLICE_X14Y120_AO6;
  assign CLBLM_R_X11Y120_SLICE_X14Y120_B = CLBLM_R_X11Y120_SLICE_X14Y120_BO6;
  assign CLBLM_R_X11Y120_SLICE_X14Y120_C = CLBLM_R_X11Y120_SLICE_X14Y120_CO6;
  assign CLBLM_R_X11Y120_SLICE_X14Y120_D = CLBLM_R_X11Y120_SLICE_X14Y120_DO6;
  assign CLBLM_R_X11Y120_SLICE_X14Y120_AMUX = CLBLM_R_X11Y120_SLICE_X14Y120_AO5;
  assign CLBLM_R_X11Y120_SLICE_X14Y120_BMUX = CLBLM_R_X11Y120_SLICE_X14Y120_BO5;
  assign CLBLM_R_X11Y120_SLICE_X15Y120_A = CLBLM_R_X11Y120_SLICE_X15Y120_AO6;
  assign CLBLM_R_X11Y120_SLICE_X15Y120_B = CLBLM_R_X11Y120_SLICE_X15Y120_BO6;
  assign CLBLM_R_X11Y120_SLICE_X15Y120_C = CLBLM_R_X11Y120_SLICE_X15Y120_CO6;
  assign CLBLM_R_X11Y120_SLICE_X15Y120_D = CLBLM_R_X11Y120_SLICE_X15Y120_DO6;
  assign CLBLM_R_X11Y121_SLICE_X14Y121_A = CLBLM_R_X11Y121_SLICE_X14Y121_AO6;
  assign CLBLM_R_X11Y121_SLICE_X14Y121_B = CLBLM_R_X11Y121_SLICE_X14Y121_BO6;
  assign CLBLM_R_X11Y121_SLICE_X14Y121_C = CLBLM_R_X11Y121_SLICE_X14Y121_CO6;
  assign CLBLM_R_X11Y121_SLICE_X14Y121_D = CLBLM_R_X11Y121_SLICE_X14Y121_DO6;
  assign CLBLM_R_X11Y121_SLICE_X14Y121_BMUX = CLBLM_R_X11Y121_SLICE_X14Y121_BO5;
  assign CLBLM_R_X11Y121_SLICE_X15Y121_A = CLBLM_R_X11Y121_SLICE_X15Y121_AO6;
  assign CLBLM_R_X11Y121_SLICE_X15Y121_B = CLBLM_R_X11Y121_SLICE_X15Y121_BO6;
  assign CLBLM_R_X11Y121_SLICE_X15Y121_C = CLBLM_R_X11Y121_SLICE_X15Y121_CO6;
  assign CLBLM_R_X11Y121_SLICE_X15Y121_D = CLBLM_R_X11Y121_SLICE_X15Y121_DO6;
  assign CLBLM_R_X11Y121_SLICE_X15Y121_AMUX = CLBLM_R_X11Y121_SLICE_X15Y121_AO6;
  assign CLBLM_R_X11Y122_SLICE_X14Y122_A = CLBLM_R_X11Y122_SLICE_X14Y122_AO6;
  assign CLBLM_R_X11Y122_SLICE_X14Y122_B = CLBLM_R_X11Y122_SLICE_X14Y122_BO6;
  assign CLBLM_R_X11Y122_SLICE_X14Y122_C = CLBLM_R_X11Y122_SLICE_X14Y122_CO6;
  assign CLBLM_R_X11Y122_SLICE_X14Y122_D = CLBLM_R_X11Y122_SLICE_X14Y122_DO6;
  assign CLBLM_R_X11Y122_SLICE_X15Y122_A = CLBLM_R_X11Y122_SLICE_X15Y122_AO6;
  assign CLBLM_R_X11Y122_SLICE_X15Y122_B = CLBLM_R_X11Y122_SLICE_X15Y122_BO6;
  assign CLBLM_R_X11Y122_SLICE_X15Y122_C = CLBLM_R_X11Y122_SLICE_X15Y122_CO6;
  assign CLBLM_R_X11Y122_SLICE_X15Y122_D = CLBLM_R_X11Y122_SLICE_X15Y122_DO6;
  assign CLBLM_R_X11Y123_SLICE_X14Y123_A = CLBLM_R_X11Y123_SLICE_X14Y123_AO6;
  assign CLBLM_R_X11Y123_SLICE_X14Y123_B = CLBLM_R_X11Y123_SLICE_X14Y123_BO6;
  assign CLBLM_R_X11Y123_SLICE_X14Y123_C = CLBLM_R_X11Y123_SLICE_X14Y123_CO6;
  assign CLBLM_R_X11Y123_SLICE_X14Y123_D = CLBLM_R_X11Y123_SLICE_X14Y123_DO6;
  assign CLBLM_R_X11Y123_SLICE_X14Y123_AMUX = CLBLM_R_X11Y123_SLICE_X14Y123_AO5;
  assign CLBLM_R_X11Y123_SLICE_X14Y123_BMUX = CLBLM_R_X11Y123_SLICE_X14Y123_BO5;
  assign CLBLM_R_X11Y123_SLICE_X15Y123_A = CLBLM_R_X11Y123_SLICE_X15Y123_AO6;
  assign CLBLM_R_X11Y123_SLICE_X15Y123_B = CLBLM_R_X11Y123_SLICE_X15Y123_BO6;
  assign CLBLM_R_X11Y123_SLICE_X15Y123_C = CLBLM_R_X11Y123_SLICE_X15Y123_CO6;
  assign CLBLM_R_X11Y123_SLICE_X15Y123_D = CLBLM_R_X11Y123_SLICE_X15Y123_DO6;
  assign CLBLM_R_X11Y128_SLICE_X14Y128_A = CLBLM_R_X11Y128_SLICE_X14Y128_AO6;
  assign CLBLM_R_X11Y128_SLICE_X14Y128_B = CLBLM_R_X11Y128_SLICE_X14Y128_BO6;
  assign CLBLM_R_X11Y128_SLICE_X14Y128_C = CLBLM_R_X11Y128_SLICE_X14Y128_CO6;
  assign CLBLM_R_X11Y128_SLICE_X14Y128_D = CLBLM_R_X11Y128_SLICE_X14Y128_DO6;
  assign CLBLM_R_X11Y128_SLICE_X14Y128_AMUX = CLBLM_R_X11Y128_SLICE_X14Y128_AO5;
  assign CLBLM_R_X11Y128_SLICE_X15Y128_A = CLBLM_R_X11Y128_SLICE_X15Y128_AO6;
  assign CLBLM_R_X11Y128_SLICE_X15Y128_B = CLBLM_R_X11Y128_SLICE_X15Y128_BO6;
  assign CLBLM_R_X11Y128_SLICE_X15Y128_C = CLBLM_R_X11Y128_SLICE_X15Y128_CO6;
  assign CLBLM_R_X11Y128_SLICE_X15Y128_D = CLBLM_R_X11Y128_SLICE_X15Y128_DO6;
  assign CLBLM_R_X13Y119_SLICE_X18Y119_A = CLBLM_R_X13Y119_SLICE_X18Y119_AO6;
  assign CLBLM_R_X13Y119_SLICE_X18Y119_B = CLBLM_R_X13Y119_SLICE_X18Y119_BO6;
  assign CLBLM_R_X13Y119_SLICE_X18Y119_C = CLBLM_R_X13Y119_SLICE_X18Y119_CO6;
  assign CLBLM_R_X13Y119_SLICE_X18Y119_D = CLBLM_R_X13Y119_SLICE_X18Y119_DO6;
  assign CLBLM_R_X13Y119_SLICE_X19Y119_A = CLBLM_R_X13Y119_SLICE_X19Y119_AO6;
  assign CLBLM_R_X13Y119_SLICE_X19Y119_B = CLBLM_R_X13Y119_SLICE_X19Y119_BO6;
  assign CLBLM_R_X13Y119_SLICE_X19Y119_C = CLBLM_R_X13Y119_SLICE_X19Y119_CO6;
  assign CLBLM_R_X13Y119_SLICE_X19Y119_D = CLBLM_R_X13Y119_SLICE_X19Y119_DO6;
  assign CLBLM_R_X13Y120_SLICE_X18Y120_A = CLBLM_R_X13Y120_SLICE_X18Y120_AO6;
  assign CLBLM_R_X13Y120_SLICE_X18Y120_B = CLBLM_R_X13Y120_SLICE_X18Y120_BO6;
  assign CLBLM_R_X13Y120_SLICE_X18Y120_C = CLBLM_R_X13Y120_SLICE_X18Y120_CO6;
  assign CLBLM_R_X13Y120_SLICE_X18Y120_D = CLBLM_R_X13Y120_SLICE_X18Y120_DO6;
  assign CLBLM_R_X13Y120_SLICE_X19Y120_A = CLBLM_R_X13Y120_SLICE_X19Y120_AO6;
  assign CLBLM_R_X13Y120_SLICE_X19Y120_B = CLBLM_R_X13Y120_SLICE_X19Y120_BO6;
  assign CLBLM_R_X13Y120_SLICE_X19Y120_C = CLBLM_R_X13Y120_SLICE_X19Y120_CO6;
  assign CLBLM_R_X13Y120_SLICE_X19Y120_D = CLBLM_R_X13Y120_SLICE_X19Y120_DO6;
  assign CLBLM_R_X37Y119_SLICE_X56Y119_A = CLBLM_R_X37Y119_SLICE_X56Y119_AO6;
  assign CLBLM_R_X37Y119_SLICE_X56Y119_B = CLBLM_R_X37Y119_SLICE_X56Y119_BO6;
  assign CLBLM_R_X37Y119_SLICE_X56Y119_C = CLBLM_R_X37Y119_SLICE_X56Y119_CO6;
  assign CLBLM_R_X37Y119_SLICE_X56Y119_D = CLBLM_R_X37Y119_SLICE_X56Y119_DO6;
  assign CLBLM_R_X37Y119_SLICE_X57Y119_A = CLBLM_R_X37Y119_SLICE_X57Y119_AO6;
  assign CLBLM_R_X37Y119_SLICE_X57Y119_B = CLBLM_R_X37Y119_SLICE_X57Y119_BO6;
  assign CLBLM_R_X37Y119_SLICE_X57Y119_C = CLBLM_R_X37Y119_SLICE_X57Y119_CO6;
  assign CLBLM_R_X37Y119_SLICE_X57Y119_D = CLBLM_R_X37Y119_SLICE_X57Y119_DO6;
  assign CLBLM_R_X103Y138_SLICE_X162Y138_A = CLBLM_R_X103Y138_SLICE_X162Y138_AO6;
  assign CLBLM_R_X103Y138_SLICE_X162Y138_B = CLBLM_R_X103Y138_SLICE_X162Y138_BO6;
  assign CLBLM_R_X103Y138_SLICE_X162Y138_C = CLBLM_R_X103Y138_SLICE_X162Y138_CO6;
  assign CLBLM_R_X103Y138_SLICE_X162Y138_D = CLBLM_R_X103Y138_SLICE_X162Y138_DO6;
  assign CLBLM_R_X103Y138_SLICE_X163Y138_A = CLBLM_R_X103Y138_SLICE_X163Y138_AO6;
  assign CLBLM_R_X103Y138_SLICE_X163Y138_B = CLBLM_R_X103Y138_SLICE_X163Y138_BO6;
  assign CLBLM_R_X103Y138_SLICE_X163Y138_C = CLBLM_R_X103Y138_SLICE_X163Y138_CO6;
  assign CLBLM_R_X103Y138_SLICE_X163Y138_D = CLBLM_R_X103Y138_SLICE_X163Y138_DO6;
  assign CLBLM_R_X103Y169_SLICE_X162Y169_A = CLBLM_R_X103Y169_SLICE_X162Y169_AO6;
  assign CLBLM_R_X103Y169_SLICE_X162Y169_B = CLBLM_R_X103Y169_SLICE_X162Y169_BO6;
  assign CLBLM_R_X103Y169_SLICE_X162Y169_C = CLBLM_R_X103Y169_SLICE_X162Y169_CO6;
  assign CLBLM_R_X103Y169_SLICE_X162Y169_D = CLBLM_R_X103Y169_SLICE_X162Y169_DO6;
  assign CLBLM_R_X103Y169_SLICE_X163Y169_A = CLBLM_R_X103Y169_SLICE_X163Y169_AO6;
  assign CLBLM_R_X103Y169_SLICE_X163Y169_B = CLBLM_R_X103Y169_SLICE_X163Y169_BO6;
  assign CLBLM_R_X103Y169_SLICE_X163Y169_C = CLBLM_R_X103Y169_SLICE_X163Y169_CO6;
  assign CLBLM_R_X103Y169_SLICE_X163Y169_D = CLBLM_R_X103Y169_SLICE_X163Y169_DO6;
  assign CLBLM_R_X103Y169_SLICE_X163Y169_AMUX = CLBLM_R_X103Y169_SLICE_X163Y169_AO5;
  assign CLBLM_R_X103Y172_SLICE_X162Y172_A = CLBLM_R_X103Y172_SLICE_X162Y172_AO6;
  assign CLBLM_R_X103Y172_SLICE_X162Y172_B = CLBLM_R_X103Y172_SLICE_X162Y172_BO6;
  assign CLBLM_R_X103Y172_SLICE_X162Y172_C = CLBLM_R_X103Y172_SLICE_X162Y172_CO6;
  assign CLBLM_R_X103Y172_SLICE_X162Y172_D = CLBLM_R_X103Y172_SLICE_X162Y172_DO6;
  assign CLBLM_R_X103Y172_SLICE_X163Y172_A = CLBLM_R_X103Y172_SLICE_X163Y172_AO6;
  assign CLBLM_R_X103Y172_SLICE_X163Y172_B = CLBLM_R_X103Y172_SLICE_X163Y172_BO6;
  assign CLBLM_R_X103Y172_SLICE_X163Y172_C = CLBLM_R_X103Y172_SLICE_X163Y172_CO6;
  assign CLBLM_R_X103Y172_SLICE_X163Y172_D = CLBLM_R_X103Y172_SLICE_X163Y172_DO6;
  assign CLBLM_R_X103Y172_SLICE_X163Y172_AMUX = CLBLM_R_X103Y172_SLICE_X163Y172_AO5;
  assign CLBLM_R_X103Y174_SLICE_X162Y174_A = CLBLM_R_X103Y174_SLICE_X162Y174_AO6;
  assign CLBLM_R_X103Y174_SLICE_X162Y174_B = CLBLM_R_X103Y174_SLICE_X162Y174_BO6;
  assign CLBLM_R_X103Y174_SLICE_X162Y174_C = CLBLM_R_X103Y174_SLICE_X162Y174_CO6;
  assign CLBLM_R_X103Y174_SLICE_X162Y174_D = CLBLM_R_X103Y174_SLICE_X162Y174_DO6;
  assign CLBLM_R_X103Y174_SLICE_X163Y174_A = CLBLM_R_X103Y174_SLICE_X163Y174_AO6;
  assign CLBLM_R_X103Y174_SLICE_X163Y174_B = CLBLM_R_X103Y174_SLICE_X163Y174_BO6;
  assign CLBLM_R_X103Y174_SLICE_X163Y174_C = CLBLM_R_X103Y174_SLICE_X163Y174_CO6;
  assign CLBLM_R_X103Y174_SLICE_X163Y174_D = CLBLM_R_X103Y174_SLICE_X163Y174_DO6;
  assign CLBLM_R_X103Y174_SLICE_X163Y174_AMUX = CLBLM_R_X103Y174_SLICE_X163Y174_AO5;
  assign CLBLM_R_X103Y177_SLICE_X162Y177_A = CLBLM_R_X103Y177_SLICE_X162Y177_AO6;
  assign CLBLM_R_X103Y177_SLICE_X162Y177_B = CLBLM_R_X103Y177_SLICE_X162Y177_BO6;
  assign CLBLM_R_X103Y177_SLICE_X162Y177_C = CLBLM_R_X103Y177_SLICE_X162Y177_CO6;
  assign CLBLM_R_X103Y177_SLICE_X162Y177_D = CLBLM_R_X103Y177_SLICE_X162Y177_DO6;
  assign CLBLM_R_X103Y177_SLICE_X163Y177_A = CLBLM_R_X103Y177_SLICE_X163Y177_AO6;
  assign CLBLM_R_X103Y177_SLICE_X163Y177_B = CLBLM_R_X103Y177_SLICE_X163Y177_BO6;
  assign CLBLM_R_X103Y177_SLICE_X163Y177_C = CLBLM_R_X103Y177_SLICE_X163Y177_CO6;
  assign CLBLM_R_X103Y177_SLICE_X163Y177_D = CLBLM_R_X103Y177_SLICE_X163Y177_DO6;
  assign CLBLM_R_X103Y177_SLICE_X163Y177_AMUX = CLBLM_R_X103Y177_SLICE_X163Y177_AO5;
  assign LIOI3_X0Y51_ILOGIC_X0Y52_O = LIOB33_X0Y51_IOB_X0Y52_I;
  assign LIOI3_X0Y51_ILOGIC_X0Y51_O = LIOB33_X0Y51_IOB_X0Y51_I;
  assign LIOI3_X0Y53_ILOGIC_X0Y54_O = LIOB33_X0Y53_IOB_X0Y54_I;
  assign LIOI3_X0Y53_ILOGIC_X0Y53_O = LIOB33_X0Y53_IOB_X0Y53_I;
  assign LIOI3_X0Y55_ILOGIC_X0Y56_O = LIOB33_X0Y55_IOB_X0Y56_I;
  assign LIOI3_X0Y55_ILOGIC_X0Y55_O = LIOB33_X0Y55_IOB_X0Y55_I;
  assign LIOI3_X0Y59_ILOGIC_X0Y60_O = LIOB33_X0Y59_IOB_X0Y60_I;
  assign LIOI3_X0Y59_ILOGIC_X0Y59_O = LIOB33_X0Y59_IOB_X0Y59_I;
  assign LIOI3_X0Y61_ILOGIC_X0Y62_O = LIOB33_X0Y61_IOB_X0Y62_I;
  assign LIOI3_X0Y61_ILOGIC_X0Y61_O = LIOB33_X0Y61_IOB_X0Y61_I;
  assign LIOI3_X0Y65_ILOGIC_X0Y66_O = LIOB33_X0Y65_IOB_X0Y66_I;
  assign LIOI3_X0Y65_ILOGIC_X0Y65_O = LIOB33_X0Y65_IOB_X0Y65_I;
  assign LIOI3_X0Y67_ILOGIC_X0Y68_O = LIOB33_X0Y67_IOB_X0Y68_I;
  assign LIOI3_X0Y67_ILOGIC_X0Y67_O = LIOB33_X0Y67_IOB_X0Y67_I;
  assign LIOI3_X0Y71_ILOGIC_X0Y72_O = LIOB33_X0Y71_IOB_X0Y72_I;
  assign LIOI3_X0Y71_ILOGIC_X0Y71_O = LIOB33_X0Y71_IOB_X0Y71_I;
  assign LIOI3_X0Y73_ILOGIC_X0Y74_O = LIOB33_X0Y73_IOB_X0Y74_I;
  assign LIOI3_X0Y73_ILOGIC_X0Y73_O = LIOB33_X0Y73_IOB_X0Y73_I;
  assign LIOI3_X0Y75_ILOGIC_X0Y76_O = LIOB33_X0Y75_IOB_X0Y76_I;
  assign LIOI3_X0Y75_ILOGIC_X0Y75_O = LIOB33_X0Y75_IOB_X0Y75_I;
  assign LIOI3_X0Y77_ILOGIC_X0Y78_O = LIOB33_X0Y77_IOB_X0Y78_I;
  assign LIOI3_X0Y77_ILOGIC_X0Y77_O = LIOB33_X0Y77_IOB_X0Y77_I;
  assign LIOI3_X0Y79_ILOGIC_X0Y79_O = LIOB33_X0Y79_IOB_X0Y79_I;
  assign LIOI3_X0Y79_OLOGIC_X0Y80_OQ = CLBLL_L_X2Y111_SLICE_X0Y111_AO6;
  assign LIOI3_X0Y79_OLOGIC_X0Y80_TQ = 1'b1;
  assign LIOI3_X0Y101_OLOGIC_X0Y102_OQ = CLBLL_L_X2Y111_SLICE_X0Y111_AO5;
  assign LIOI3_X0Y101_OLOGIC_X0Y102_TQ = 1'b1;
  assign LIOI3_X0Y101_OLOGIC_X0Y101_OQ = CLBLL_L_X2Y111_SLICE_X0Y111_CO6;
  assign LIOI3_X0Y101_OLOGIC_X0Y101_TQ = 1'b1;
  assign LIOI3_X0Y103_OLOGIC_X0Y104_OQ = CLBLL_L_X2Y111_SLICE_X0Y111_CO5;
  assign LIOI3_X0Y103_OLOGIC_X0Y104_TQ = 1'b1;
  assign LIOI3_X0Y103_OLOGIC_X0Y103_OQ = CLBLL_L_X2Y113_SLICE_X0Y113_AO6;
  assign LIOI3_X0Y103_OLOGIC_X0Y103_TQ = 1'b1;
  assign LIOI3_X0Y105_OLOGIC_X0Y106_OQ = CLBLL_L_X2Y111_SLICE_X0Y111_DO5;
  assign LIOI3_X0Y105_OLOGIC_X0Y106_TQ = 1'b1;
  assign LIOI3_X0Y105_OLOGIC_X0Y105_OQ = CLBLL_L_X2Y111_SLICE_X0Y111_DO6;
  assign LIOI3_X0Y105_OLOGIC_X0Y105_TQ = 1'b1;
  assign LIOI3_X0Y109_OLOGIC_X0Y110_OQ = CLBLL_L_X2Y110_SLICE_X0Y110_AO5;
  assign LIOI3_X0Y109_OLOGIC_X0Y110_TQ = 1'b1;
  assign LIOI3_X0Y109_OLOGIC_X0Y109_OQ = CLBLL_L_X2Y110_SLICE_X0Y110_AO6;
  assign LIOI3_X0Y109_OLOGIC_X0Y109_TQ = 1'b1;
  assign LIOI3_X0Y111_OLOGIC_X0Y112_OQ = CLBLM_R_X11Y114_SLICE_X14Y114_D5Q;
  assign LIOI3_X0Y111_OLOGIC_X0Y112_TQ = 1'b1;
  assign LIOI3_X0Y111_OLOGIC_X0Y111_OQ = 1'b0;
  assign LIOI3_X0Y111_OLOGIC_X0Y111_TQ = 1'b1;
  assign LIOI3_X0Y115_OLOGIC_X0Y116_OQ = CLBLM_L_X8Y123_SLICE_X11Y123_AQ;
  assign LIOI3_X0Y115_OLOGIC_X0Y116_TQ = 1'b1;
  assign LIOI3_X0Y115_OLOGIC_X0Y115_OQ = CLBLM_R_X11Y114_SLICE_X14Y114_DQ;
  assign LIOI3_X0Y115_OLOGIC_X0Y115_TQ = 1'b1;
  assign LIOI3_X0Y117_OLOGIC_X0Y118_OQ = CLBLL_L_X4Y116_SLICE_X4Y116_CQ;
  assign LIOI3_X0Y117_OLOGIC_X0Y118_TQ = 1'b1;
  assign LIOI3_X0Y117_OLOGIC_X0Y117_OQ = CLBLL_L_X4Y119_SLICE_X4Y119_BQ;
  assign LIOI3_X0Y117_OLOGIC_X0Y117_TQ = 1'b1;
  assign LIOI3_X0Y121_OLOGIC_X0Y122_OQ = CLBLM_R_X5Y121_SLICE_X6Y121_A5Q;
  assign LIOI3_X0Y121_OLOGIC_X0Y122_TQ = 1'b1;
  assign LIOI3_X0Y121_OLOGIC_X0Y121_OQ = CLBLM_L_X8Y123_SLICE_X11Y123_A5Q;
  assign LIOI3_X0Y121_OLOGIC_X0Y121_TQ = 1'b1;
  assign LIOI3_X0Y123_OLOGIC_X0Y124_OQ = CLBLL_L_X4Y116_SLICE_X4Y116_C5Q;
  assign LIOI3_X0Y123_OLOGIC_X0Y124_TQ = 1'b1;
  assign LIOI3_X0Y123_OLOGIC_X0Y123_OQ = CLBLM_R_X5Y117_SLICE_X6Y117_D5Q;
  assign LIOI3_X0Y123_OLOGIC_X0Y123_TQ = 1'b1;
  assign LIOI3_X0Y125_OLOGIC_X0Y126_OQ = CLBLM_R_X5Y124_SLICE_X6Y124_CQ;
  assign LIOI3_X0Y125_OLOGIC_X0Y126_TQ = 1'b1;
  assign LIOI3_X0Y125_OLOGIC_X0Y125_OQ = CLBLM_R_X7Y115_SLICE_X9Y115_CQ;
  assign LIOI3_X0Y125_OLOGIC_X0Y125_TQ = 1'b1;
  assign LIOI3_X0Y127_OLOGIC_X0Y128_OQ = CLBLL_L_X2Y117_SLICE_X0Y117_A5Q;
  assign LIOI3_X0Y127_OLOGIC_X0Y128_TQ = 1'b1;
  assign LIOI3_X0Y127_OLOGIC_X0Y127_OQ = CLBLL_L_X4Y121_SLICE_X4Y121_BQ;
  assign LIOI3_X0Y127_OLOGIC_X0Y127_TQ = 1'b1;
  assign LIOI3_X0Y129_OLOGIC_X0Y130_OQ = CLBLL_L_X52Y126_SLICE_X78Y126_AO6;
  assign LIOI3_X0Y129_OLOGIC_X0Y130_TQ = 1'b1;
  assign LIOI3_X0Y129_OLOGIC_X0Y129_OQ = CLBLM_R_X3Y115_SLICE_X3Y115_CQ;
  assign LIOI3_X0Y129_OLOGIC_X0Y129_TQ = 1'b1;
  assign LIOI3_X0Y133_OLOGIC_X0Y134_OQ = CLBLM_R_X7Y124_SLICE_X8Y124_BQ;
  assign LIOI3_X0Y133_OLOGIC_X0Y134_TQ = 1'b1;
  assign LIOI3_X0Y133_OLOGIC_X0Y133_OQ = CLBLM_R_X7Y124_SLICE_X8Y124_A5Q;
  assign LIOI3_X0Y133_OLOGIC_X0Y133_TQ = 1'b1;
  assign LIOI3_X0Y135_OLOGIC_X0Y136_OQ = CLBLM_R_X7Y124_SLICE_X8Y124_CQ;
  assign LIOI3_X0Y135_OLOGIC_X0Y136_TQ = 1'b1;
  assign LIOI3_X0Y135_OLOGIC_X0Y135_OQ = CLBLL_L_X4Y123_SLICE_X4Y123_AQ;
  assign LIOI3_X0Y135_OLOGIC_X0Y135_TQ = 1'b1;
  assign LIOI3_X0Y139_OLOGIC_X0Y140_OQ = CLBLL_L_X4Y123_SLICE_X4Y123_BQ;
  assign LIOI3_X0Y139_OLOGIC_X0Y140_TQ = 1'b1;
  assign LIOI3_X0Y139_OLOGIC_X0Y139_OQ = CLBLM_R_X5Y124_SLICE_X6Y124_AQ;
  assign LIOI3_X0Y139_OLOGIC_X0Y139_TQ = 1'b1;
  assign LIOI3_X0Y141_OLOGIC_X0Y142_OQ = LIOB33_X0Y53_IOB_X0Y54_I;
  assign LIOI3_X0Y141_OLOGIC_X0Y142_TQ = 1'b1;
  assign LIOI3_X0Y141_OLOGIC_X0Y141_OQ = CLBLM_R_X5Y123_SLICE_X6Y123_AQ;
  assign LIOI3_X0Y141_OLOGIC_X0Y141_TQ = 1'b1;
  assign LIOI3_X0Y145_OLOGIC_X0Y146_OQ = LIOB33_X0Y59_IOB_X0Y59_I;
  assign LIOI3_X0Y145_OLOGIC_X0Y146_TQ = 1'b1;
  assign LIOI3_X0Y145_OLOGIC_X0Y145_OQ = LIOB33_X0Y57_IOB_X0Y58_I;
  assign LIOI3_X0Y145_OLOGIC_X0Y145_TQ = 1'b1;
  assign LIOI3_X0Y147_OLOGIC_X0Y148_OQ = LIOB33_X0Y61_IOB_X0Y61_I;
  assign LIOI3_X0Y147_OLOGIC_X0Y148_TQ = 1'b1;
  assign LIOI3_X0Y147_OLOGIC_X0Y147_OQ = LIOB33_X0Y71_IOB_X0Y71_I;
  assign LIOI3_X0Y147_OLOGIC_X0Y147_TQ = 1'b1;
  assign LIOI3_X0Y151_OLOGIC_X0Y152_OQ = LIOB33_X0Y65_IOB_X0Y66_I;
  assign LIOI3_X0Y151_OLOGIC_X0Y152_TQ = 1'b1;
  assign LIOI3_X0Y151_OLOGIC_X0Y151_OQ = LIOB33_X0Y65_IOB_X0Y65_I;
  assign LIOI3_X0Y151_OLOGIC_X0Y151_TQ = 1'b1;
  assign LIOI3_X0Y153_OLOGIC_X0Y154_OQ = LIOB33_X0Y67_IOB_X0Y68_I;
  assign LIOI3_X0Y153_OLOGIC_X0Y154_TQ = 1'b1;
  assign LIOI3_X0Y153_OLOGIC_X0Y153_OQ = LIOB33_X0Y67_IOB_X0Y67_I;
  assign LIOI3_X0Y153_OLOGIC_X0Y153_TQ = 1'b1;
  assign LIOI3_X0Y155_OLOGIC_X0Y156_OQ = RIOB33_X105Y105_IOB_X1Y106_I;
  assign LIOI3_X0Y155_OLOGIC_X0Y156_TQ = 1'b1;
  assign LIOI3_X0Y155_OLOGIC_X0Y155_OQ = LIOB33_X0Y69_IOB_X0Y70_I;
  assign LIOI3_X0Y155_OLOGIC_X0Y155_TQ = 1'b1;
  assign LIOI3_X0Y159_OLOGIC_X0Y160_OQ = RIOB33_X105Y107_IOB_X1Y107_I;
  assign LIOI3_X0Y159_OLOGIC_X0Y160_TQ = 1'b1;
  assign LIOI3_X0Y159_OLOGIC_X0Y159_OQ = RIOB33_X105Y117_IOB_X1Y117_I;
  assign LIOI3_X0Y159_OLOGIC_X0Y159_TQ = 1'b1;
  assign LIOI3_X0Y161_OLOGIC_X0Y162_OQ = RIOB33_X105Y109_IOB_X1Y109_I;
  assign LIOI3_X0Y161_OLOGIC_X0Y162_TQ = 1'b1;
  assign LIOI3_X0Y161_OLOGIC_X0Y161_OQ = RIOB33_X105Y107_IOB_X1Y108_I;
  assign LIOI3_X0Y161_OLOGIC_X0Y161_TQ = 1'b1;
  assign LIOI3_X0Y165_OLOGIC_X0Y166_OQ = RIOB33_X105Y113_IOB_X1Y113_I;
  assign LIOI3_X0Y165_OLOGIC_X0Y166_TQ = 1'b1;
  assign LIOI3_X0Y165_OLOGIC_X0Y165_OQ = RIOB33_X105Y111_IOB_X1Y112_I;
  assign LIOI3_X0Y165_OLOGIC_X0Y165_TQ = 1'b1;
  assign LIOI3_X0Y167_OLOGIC_X0Y168_OQ = RIOB33_X105Y123_IOB_X1Y123_I;
  assign LIOI3_X0Y167_OLOGIC_X0Y168_TQ = 1'b1;
  assign LIOI3_X0Y167_OLOGIC_X0Y167_OQ = RIOB33_X105Y113_IOB_X1Y114_I;
  assign LIOI3_X0Y167_OLOGIC_X0Y167_TQ = 1'b1;
  assign LIOI3_X0Y171_OLOGIC_X0Y172_OQ = CLBLM_R_X103Y138_SLICE_X163Y138_AO6;
  assign LIOI3_X0Y171_OLOGIC_X0Y172_TQ = 1'b1;
  assign LIOI3_X0Y171_OLOGIC_X0Y171_OQ = LIOB33_SING_X0Y50_IOB_X0Y50_I;
  assign LIOI3_X0Y171_OLOGIC_X0Y171_TQ = 1'b1;
  assign LIOI3_X0Y173_OLOGIC_X0Y174_OQ = CLBLM_R_X7Y151_SLICE_X8Y151_AO6;
  assign LIOI3_X0Y173_OLOGIC_X0Y174_TQ = 1'b1;
  assign LIOI3_X0Y173_OLOGIC_X0Y173_OQ = CLBLM_L_X8Y133_SLICE_X11Y133_AO5;
  assign LIOI3_X0Y173_OLOGIC_X0Y173_TQ = 1'b1;
  assign LIOI3_X0Y175_OLOGIC_X0Y176_OQ = RIOB33_X105Y127_IOB_X1Y128_I;
  assign LIOI3_X0Y175_OLOGIC_X0Y176_TQ = 1'b1;
  assign LIOI3_X0Y175_OLOGIC_X0Y175_OQ = RIOB33_X105Y127_IOB_X1Y127_I;
  assign LIOI3_X0Y175_OLOGIC_X0Y175_TQ = 1'b1;
  assign LIOI3_X0Y177_OLOGIC_X0Y178_OQ = RIOB33_X105Y129_IOB_X1Y130_I;
  assign LIOI3_X0Y177_OLOGIC_X0Y178_TQ = 1'b1;
  assign LIOI3_X0Y177_OLOGIC_X0Y177_OQ = RIOB33_X105Y129_IOB_X1Y129_I;
  assign LIOI3_X0Y177_OLOGIC_X0Y177_TQ = 1'b1;
  assign LIOI3_X0Y179_OLOGIC_X0Y180_OQ = RIOB33_X105Y131_IOB_X1Y132_I;
  assign LIOI3_X0Y179_OLOGIC_X0Y180_TQ = 1'b1;
  assign LIOI3_X0Y179_OLOGIC_X0Y179_OQ = RIOB33_X105Y131_IOB_X1Y131_I;
  assign LIOI3_X0Y179_OLOGIC_X0Y179_TQ = 1'b1;
  assign LIOI3_X0Y183_OLOGIC_X0Y184_OQ = RIOB33_X105Y135_IOB_X1Y136_I;
  assign LIOI3_X0Y183_OLOGIC_X0Y184_TQ = 1'b1;
  assign LIOI3_X0Y183_OLOGIC_X0Y183_OQ = RIOB33_X105Y135_IOB_X1Y135_I;
  assign LIOI3_X0Y183_OLOGIC_X0Y183_TQ = 1'b1;
  assign LIOI3_X0Y185_OLOGIC_X0Y186_OQ = RIOB33_X105Y143_IOB_X1Y143_I;
  assign LIOI3_X0Y185_OLOGIC_X0Y186_TQ = 1'b1;
  assign LIOI3_X0Y185_OLOGIC_X0Y185_OQ = RIOB33_X105Y137_IOB_X1Y137_I;
  assign LIOI3_X0Y185_OLOGIC_X0Y185_TQ = 1'b1;
  assign LIOI3_X0Y189_OLOGIC_X0Y190_OQ = RIOB33_X105Y147_IOB_X1Y147_I;
  assign LIOI3_X0Y189_OLOGIC_X0Y190_TQ = 1'b1;
  assign LIOI3_X0Y189_OLOGIC_X0Y189_OQ = RIOB33_X105Y145_IOB_X1Y146_I;
  assign LIOI3_X0Y189_OLOGIC_X0Y189_TQ = 1'b1;
  assign LIOI3_X0Y191_OLOGIC_X0Y192_OQ = LIOB33_X0Y51_IOB_X0Y52_I;
  assign LIOI3_X0Y191_OLOGIC_X0Y192_TQ = 1'b1;
  assign LIOI3_X0Y191_OLOGIC_X0Y191_OQ = RIOB33_X105Y147_IOB_X1Y148_I;
  assign LIOI3_X0Y191_OLOGIC_X0Y191_TQ = 1'b1;
  assign LIOI3_X0Y195_OLOGIC_X0Y196_OQ = LIOB33_X0Y69_IOB_X0Y69_I;
  assign LIOI3_X0Y195_OLOGIC_X0Y196_TQ = 1'b1;
  assign LIOI3_X0Y195_OLOGIC_X0Y195_OQ = LIOB33_X0Y63_IOB_X0Y64_I;
  assign LIOI3_X0Y195_OLOGIC_X0Y195_TQ = 1'b1;
  assign LIOI3_X0Y197_OLOGIC_X0Y198_OQ = LIOB33_X0Y73_IOB_X0Y73_I;
  assign LIOI3_X0Y197_OLOGIC_X0Y198_TQ = 1'b1;
  assign LIOI3_X0Y197_OLOGIC_X0Y197_OQ = LIOB33_X0Y71_IOB_X0Y72_I;
  assign LIOI3_X0Y197_OLOGIC_X0Y197_TQ = 1'b1;
  assign LIOI3_SING_X0Y50_ILOGIC_X0Y50_O = LIOB33_SING_X0Y50_IOB_X0Y50_I;
  assign LIOI3_SING_X0Y100_OLOGIC_X0Y100_OQ = CLBLL_L_X2Y111_SLICE_X0Y111_BO6;
  assign LIOI3_SING_X0Y100_OLOGIC_X0Y100_TQ = 1'b1;
  assign LIOI3_SING_X0Y149_OLOGIC_X0Y149_OQ = LIOB33_X0Y61_IOB_X0Y62_I;
  assign LIOI3_SING_X0Y149_OLOGIC_X0Y149_TQ = 1'b1;
  assign LIOI3_SING_X0Y150_OLOGIC_X0Y150_OQ = LIOB33_X0Y63_IOB_X0Y63_I;
  assign LIOI3_SING_X0Y150_OLOGIC_X0Y150_TQ = 1'b1;
  assign LIOI3_SING_X0Y199_OLOGIC_X0Y199_OQ = LIOB33_X0Y73_IOB_X0Y74_I;
  assign LIOI3_SING_X0Y199_OLOGIC_X0Y199_TQ = 1'b1;
  assign LIOI3_TBYTESRC_X0Y57_ILOGIC_X0Y58_O = LIOB33_X0Y57_IOB_X0Y58_I;
  assign LIOI3_TBYTESRC_X0Y57_ILOGIC_X0Y57_O = LIOB33_X0Y57_IOB_X0Y57_I;
  assign LIOI3_TBYTESRC_X0Y69_ILOGIC_X0Y70_O = LIOB33_X0Y69_IOB_X0Y70_I;
  assign LIOI3_TBYTESRC_X0Y69_ILOGIC_X0Y69_O = LIOB33_X0Y69_IOB_X0Y69_I;
  assign LIOI3_TBYTESRC_X0Y107_OLOGIC_X0Y108_OQ = CLBLL_L_X2Y111_SLICE_X0Y111_BO5;
  assign LIOI3_TBYTESRC_X0Y107_OLOGIC_X0Y108_TQ = 1'b1;
  assign LIOI3_TBYTESRC_X0Y107_OLOGIC_X0Y107_OQ = CLBLL_L_X2Y109_SLICE_X0Y109_AO6;
  assign LIOI3_TBYTESRC_X0Y107_OLOGIC_X0Y107_TQ = 1'b1;
  assign LIOI3_TBYTESRC_X0Y119_OLOGIC_X0Y120_OQ = CLBLM_R_X3Y116_SLICE_X3Y116_A5Q;
  assign LIOI3_TBYTESRC_X0Y119_OLOGIC_X0Y120_TQ = 1'b1;
  assign LIOI3_TBYTESRC_X0Y119_OLOGIC_X0Y119_OQ = CLBLM_L_X8Y114_SLICE_X10Y114_CQ;
  assign LIOI3_TBYTESRC_X0Y119_OLOGIC_X0Y119_TQ = 1'b1;
  assign LIOI3_TBYTESRC_X0Y131_OLOGIC_X0Y132_OQ = CLBLM_R_X7Y128_SLICE_X8Y128_AQ;
  assign LIOI3_TBYTESRC_X0Y131_OLOGIC_X0Y132_TQ = 1'b1;
  assign LIOI3_TBYTESRC_X0Y131_OLOGIC_X0Y131_OQ = CLBLM_R_X7Y128_SLICE_X8Y128_AO5;
  assign LIOI3_TBYTESRC_X0Y131_OLOGIC_X0Y131_TQ = 1'b1;
  assign LIOI3_TBYTESRC_X0Y143_OLOGIC_X0Y144_OQ = LIOB33_X0Y57_IOB_X0Y57_I;
  assign LIOI3_TBYTESRC_X0Y143_OLOGIC_X0Y144_TQ = 1'b1;
  assign LIOI3_TBYTESRC_X0Y143_OLOGIC_X0Y143_OQ = LIOB33_X0Y55_IOB_X0Y55_I;
  assign LIOI3_TBYTESRC_X0Y143_OLOGIC_X0Y143_TQ = 1'b1;
  assign LIOI3_TBYTESRC_X0Y157_OLOGIC_X0Y158_OQ = RIOB33_X105Y115_IOB_X1Y116_I;
  assign LIOI3_TBYTESRC_X0Y157_OLOGIC_X0Y158_TQ = 1'b1;
  assign LIOI3_TBYTESRC_X0Y157_OLOGIC_X0Y157_OQ = RIOB33_X105Y115_IOB_X1Y115_I;
  assign LIOI3_TBYTESRC_X0Y157_OLOGIC_X0Y157_TQ = 1'b1;
  assign LIOI3_TBYTESRC_X0Y169_OLOGIC_X0Y170_OQ = RIOB33_SING_X105Y149_IOB_X1Y149_I;
  assign LIOI3_TBYTESRC_X0Y169_OLOGIC_X0Y170_TQ = 1'b1;
  assign LIOI3_TBYTESRC_X0Y169_OLOGIC_X0Y169_OQ = RIOB33_X105Y121_IOB_X1Y122_I;
  assign LIOI3_TBYTESRC_X0Y169_OLOGIC_X0Y169_TQ = 1'b1;
  assign LIOI3_TBYTESRC_X0Y181_OLOGIC_X0Y182_OQ = RIOB33_X105Y133_IOB_X1Y134_I;
  assign LIOI3_TBYTESRC_X0Y181_OLOGIC_X0Y182_TQ = 1'b1;
  assign LIOI3_TBYTESRC_X0Y181_OLOGIC_X0Y181_OQ = RIOB33_X105Y133_IOB_X1Y133_I;
  assign LIOI3_TBYTESRC_X0Y181_OLOGIC_X0Y181_TQ = 1'b1;
  assign LIOI3_TBYTESRC_X0Y193_OLOGIC_X0Y194_OQ = LIOB33_X0Y59_IOB_X0Y60_I;
  assign LIOI3_TBYTESRC_X0Y193_OLOGIC_X0Y194_TQ = 1'b1;
  assign LIOI3_TBYTESRC_X0Y193_OLOGIC_X0Y193_OQ = LIOB33_X0Y55_IOB_X0Y56_I;
  assign LIOI3_TBYTESRC_X0Y193_OLOGIC_X0Y193_TQ = 1'b1;
  assign LIOI3_TBYTETERM_X0Y63_ILOGIC_X0Y64_O = LIOB33_X0Y63_IOB_X0Y64_I;
  assign LIOI3_TBYTETERM_X0Y63_ILOGIC_X0Y63_O = LIOB33_X0Y63_IOB_X0Y63_I;
  assign LIOI3_TBYTETERM_X0Y113_OLOGIC_X0Y114_OQ = CLBLM_R_X5Y117_SLICE_X6Y117_DQ;
  assign LIOI3_TBYTETERM_X0Y113_OLOGIC_X0Y114_TQ = 1'b1;
  assign LIOI3_TBYTETERM_X0Y113_OLOGIC_X0Y113_OQ = RIOB33_X105Y121_IOB_X1Y121_I;
  assign LIOI3_TBYTETERM_X0Y113_OLOGIC_X0Y113_TQ = 1'b1;
  assign LIOI3_TBYTETERM_X0Y137_OLOGIC_X0Y138_OQ = CLBLM_R_X5Y125_SLICE_X6Y125_AQ;
  assign LIOI3_TBYTETERM_X0Y137_OLOGIC_X0Y138_TQ = 1'b1;
  assign LIOI3_TBYTETERM_X0Y137_OLOGIC_X0Y137_OQ = CLBLM_R_X5Y124_SLICE_X6Y124_BQ;
  assign LIOI3_TBYTETERM_X0Y137_OLOGIC_X0Y137_TQ = 1'b1;
  assign LIOI3_TBYTETERM_X0Y163_OLOGIC_X0Y164_OQ = RIOB33_X105Y111_IOB_X1Y111_I;
  assign LIOI3_TBYTETERM_X0Y163_OLOGIC_X0Y164_TQ = 1'b1;
  assign LIOI3_TBYTETERM_X0Y163_OLOGIC_X0Y163_OQ = RIOB33_X105Y109_IOB_X1Y110_I;
  assign LIOI3_TBYTETERM_X0Y163_OLOGIC_X0Y163_TQ = 1'b1;
  assign LIOI3_TBYTETERM_X0Y187_OLOGIC_X0Y188_OQ = RIOB33_X105Y145_IOB_X1Y145_I;
  assign LIOI3_TBYTETERM_X0Y187_OLOGIC_X0Y188_TQ = 1'b1;
  assign LIOI3_TBYTETERM_X0Y187_OLOGIC_X0Y187_OQ = RIOB33_X105Y143_IOB_X1Y144_I;
  assign LIOI3_TBYTETERM_X0Y187_OLOGIC_X0Y187_TQ = 1'b1;
  assign RIOI3_X105Y101_ILOGIC_X1Y102_O = RIOB33_X105Y101_IOB_X1Y102_I;
  assign RIOI3_X105Y101_ILOGIC_X1Y101_O = RIOB33_X105Y101_IOB_X1Y101_I;
  assign RIOI3_X105Y103_ILOGIC_X1Y104_O = RIOB33_X105Y103_IOB_X1Y104_I;
  assign RIOI3_X105Y103_ILOGIC_X1Y103_O = RIOB33_X105Y103_IOB_X1Y103_I;
  assign RIOI3_X105Y105_ILOGIC_X1Y106_O = RIOB33_X105Y105_IOB_X1Y106_I;
  assign RIOI3_X105Y105_ILOGIC_X1Y105_O = RIOB33_X105Y105_IOB_X1Y105_I;
  assign RIOI3_X105Y109_ILOGIC_X1Y110_O = RIOB33_X105Y109_IOB_X1Y110_I;
  assign RIOI3_X105Y109_ILOGIC_X1Y109_O = RIOB33_X105Y109_IOB_X1Y109_I;
  assign RIOI3_X105Y111_ILOGIC_X1Y112_O = RIOB33_X105Y111_IOB_X1Y112_I;
  assign RIOI3_X105Y111_ILOGIC_X1Y111_O = RIOB33_X105Y111_IOB_X1Y111_I;
  assign RIOI3_X105Y115_ILOGIC_X1Y116_O = RIOB33_X105Y115_IOB_X1Y116_I;
  assign RIOI3_X105Y115_ILOGIC_X1Y115_O = RIOB33_X105Y115_IOB_X1Y115_I;
  assign RIOI3_X105Y117_ILOGIC_X1Y118_O = RIOB33_X105Y117_IOB_X1Y118_I;
  assign RIOI3_X105Y117_ILOGIC_X1Y117_O = RIOB33_X105Y117_IOB_X1Y117_I;
  assign RIOI3_X105Y121_ILOGIC_X1Y122_O = RIOB33_X105Y121_IOB_X1Y122_I;
  assign RIOI3_X105Y121_ILOGIC_X1Y121_O = RIOB33_X105Y121_IOB_X1Y121_I;
  assign RIOI3_X105Y123_ILOGIC_X1Y124_O = RIOB33_X105Y123_IOB_X1Y124_I;
  assign RIOI3_X105Y123_ILOGIC_X1Y123_O = RIOB33_X105Y123_IOB_X1Y123_I;
  assign RIOI3_X105Y125_ILOGIC_X1Y126_O = RIOB33_X105Y125_IOB_X1Y126_I;
  assign RIOI3_X105Y125_ILOGIC_X1Y125_O = RIOB33_X105Y125_IOB_X1Y125_I;
  assign RIOI3_X105Y127_ILOGIC_X1Y128_O = RIOB33_X105Y127_IOB_X1Y128_I;
  assign RIOI3_X105Y127_ILOGIC_X1Y127_O = RIOB33_X105Y127_IOB_X1Y127_I;
  assign RIOI3_X105Y129_ILOGIC_X1Y130_O = RIOB33_X105Y129_IOB_X1Y130_I;
  assign RIOI3_X105Y129_ILOGIC_X1Y129_O = RIOB33_X105Y129_IOB_X1Y129_I;
  assign RIOI3_X105Y133_ILOGIC_X1Y134_O = RIOB33_X105Y133_IOB_X1Y134_I;
  assign RIOI3_X105Y133_ILOGIC_X1Y133_O = RIOB33_X105Y133_IOB_X1Y133_I;
  assign RIOI3_X105Y135_ILOGIC_X1Y136_O = RIOB33_X105Y135_IOB_X1Y136_I;
  assign RIOI3_X105Y135_ILOGIC_X1Y135_O = RIOB33_X105Y135_IOB_X1Y135_I;
  assign RIOI3_X105Y139_ILOGIC_X1Y140_O = RIOB33_X105Y139_IOB_X1Y140_I;
  assign RIOI3_X105Y139_ILOGIC_X1Y139_O = RIOB33_X105Y139_IOB_X1Y139_I;
  assign RIOI3_X105Y141_ILOGIC_X1Y142_O = RIOB33_X105Y141_IOB_X1Y142_I;
  assign RIOI3_X105Y141_ILOGIC_X1Y141_O = RIOB33_X105Y141_IOB_X1Y141_I;
  assign RIOI3_X105Y145_ILOGIC_X1Y146_O = RIOB33_X105Y145_IOB_X1Y146_I;
  assign RIOI3_X105Y145_ILOGIC_X1Y145_O = RIOB33_X105Y145_IOB_X1Y145_I;
  assign RIOI3_X105Y147_ILOGIC_X1Y148_O = RIOB33_X105Y147_IOB_X1Y148_I;
  assign RIOI3_X105Y147_ILOGIC_X1Y147_O = RIOB33_X105Y147_IOB_X1Y147_I;
  assign RIOI3_X105Y151_OLOGIC_X1Y152_OQ = RIOB33_SING_X105Y100_IOB_X1Y100_I;
  assign RIOI3_X105Y151_OLOGIC_X1Y152_TQ = 1'b1;
  assign RIOI3_X105Y151_OLOGIC_X1Y151_OQ = LIOB33_X0Y75_IOB_X0Y76_I;
  assign RIOI3_X105Y151_OLOGIC_X1Y151_TQ = 1'b1;
  assign RIOI3_X105Y153_OLOGIC_X1Y154_OQ = RIOB33_X105Y101_IOB_X1Y102_I;
  assign RIOI3_X105Y153_OLOGIC_X1Y154_TQ = 1'b1;
  assign RIOI3_X105Y153_OLOGIC_X1Y153_OQ = RIOB33_X105Y101_IOB_X1Y101_I;
  assign RIOI3_X105Y153_OLOGIC_X1Y153_TQ = 1'b1;
  assign RIOI3_X105Y155_OLOGIC_X1Y156_OQ = RIOB33_X105Y103_IOB_X1Y104_I;
  assign RIOI3_X105Y155_OLOGIC_X1Y156_TQ = 1'b1;
  assign RIOI3_X105Y155_OLOGIC_X1Y155_OQ = RIOB33_X105Y103_IOB_X1Y103_I;
  assign RIOI3_X105Y155_OLOGIC_X1Y155_TQ = 1'b1;
  assign RIOI3_X105Y159_OLOGIC_X1Y160_OQ = CLBLM_R_X11Y119_SLICE_X14Y119_CO6;
  assign RIOI3_X105Y159_OLOGIC_X1Y160_TQ = 1'b1;
  assign RIOI3_X105Y159_OLOGIC_X1Y159_OQ = CLBLM_R_X11Y113_SLICE_X15Y113_DO6;
  assign RIOI3_X105Y159_OLOGIC_X1Y159_TQ = 1'b1;
  assign RIOI3_X105Y161_OLOGIC_X1Y162_OQ = CLBLM_R_X11Y117_SLICE_X14Y117_DO6;
  assign RIOI3_X105Y161_OLOGIC_X1Y162_TQ = 1'b1;
  assign RIOI3_X105Y161_OLOGIC_X1Y161_OQ = CLBLM_R_X11Y119_SLICE_X14Y119_CO5;
  assign RIOI3_X105Y161_OLOGIC_X1Y161_TQ = 1'b1;
  assign RIOI3_X105Y165_OLOGIC_X1Y166_OQ = RIOB33_SING_X105Y149_IOB_X1Y149_I;
  assign RIOI3_X105Y165_OLOGIC_X1Y166_TQ = 1'b1;
  assign RIOI3_X105Y165_OLOGIC_X1Y165_OQ = RIOB33_X105Y125_IOB_X1Y125_I;
  assign RIOI3_X105Y165_OLOGIC_X1Y165_TQ = 1'b1;
  assign RIOI3_X105Y167_OLOGIC_X1Y168_OQ = CLBLM_R_X7Y151_SLICE_X8Y151_AO6;
  assign RIOI3_X105Y167_OLOGIC_X1Y168_TQ = 1'b1;
  assign RIOI3_X105Y167_OLOGIC_X1Y167_OQ = LIOB33_SING_X0Y50_IOB_X0Y50_I;
  assign RIOI3_X105Y167_OLOGIC_X1Y167_TQ = 1'b1;
  assign RIOI3_X105Y171_OLOGIC_X1Y172_OQ = CLBLM_R_X103Y172_SLICE_X163Y172_AO6;
  assign RIOI3_X105Y171_OLOGIC_X1Y172_TQ = 1'b1;
  assign RIOI3_X105Y171_OLOGIC_X1Y171_OQ = CLBLM_L_X8Y128_SLICE_X10Y128_AO5;
  assign RIOI3_X105Y171_OLOGIC_X1Y171_TQ = 1'b1;
  assign RIOI3_X105Y173_OLOGIC_X1Y174_OQ = CLBLM_R_X103Y174_SLICE_X163Y174_AO6;
  assign RIOI3_X105Y173_OLOGIC_X1Y174_TQ = 1'b1;
  assign RIOI3_X105Y173_OLOGIC_X1Y173_OQ = CLBLM_R_X103Y172_SLICE_X163Y172_AO5;
  assign RIOI3_X105Y173_OLOGIC_X1Y173_TQ = 1'b1;
  assign RIOI3_X105Y175_OLOGIC_X1Y176_OQ = CLBLM_R_X103Y174_SLICE_X163Y174_AO5;
  assign RIOI3_X105Y175_OLOGIC_X1Y176_TQ = 1'b1;
  assign RIOI3_X105Y175_OLOGIC_X1Y175_OQ = CLBLM_L_X10Y128_SLICE_X13Y128_AO6;
  assign RIOI3_X105Y175_OLOGIC_X1Y175_TQ = 1'b1;
  assign RIOI3_X105Y177_OLOGIC_X1Y178_OQ = CLBLM_R_X103Y177_SLICE_X163Y177_AO5;
  assign RIOI3_X105Y177_OLOGIC_X1Y178_TQ = 1'b1;
  assign RIOI3_X105Y177_OLOGIC_X1Y177_OQ = CLBLM_R_X103Y177_SLICE_X163Y177_AO6;
  assign RIOI3_X105Y177_OLOGIC_X1Y177_TQ = 1'b1;
  assign RIOI3_X105Y179_OLOGIC_X1Y180_OQ = CLBLM_R_X11Y113_SLICE_X15Y113_DO6;
  assign RIOI3_X105Y179_OLOGIC_X1Y180_TQ = 1'b1;
  assign RIOI3_X105Y179_OLOGIC_X1Y179_OQ = CLBLM_R_X11Y128_SLICE_X14Y128_AO5;
  assign RIOI3_X105Y179_OLOGIC_X1Y179_TQ = 1'b1;
  assign RIOI3_X105Y183_OLOGIC_X1Y184_OQ = CLBLM_R_X11Y117_SLICE_X14Y117_DO5;
  assign RIOI3_X105Y183_OLOGIC_X1Y184_TQ = 1'b1;
  assign RIOI3_X105Y183_OLOGIC_X1Y183_OQ = CLBLM_R_X11Y117_SLICE_X14Y117_DO6;
  assign RIOI3_X105Y183_OLOGIC_X1Y183_TQ = 1'b1;
  assign RIOI3_X105Y185_OLOGIC_X1Y186_OQ = CLBLM_L_X12Y115_SLICE_X16Y115_BQ;
  assign RIOI3_X105Y185_OLOGIC_X1Y186_TQ = 1'b1;
  assign RIOI3_X105Y185_OLOGIC_X1Y185_OQ = CLBLM_R_X7Y119_SLICE_X9Y119_DO5;
  assign RIOI3_X105Y185_OLOGIC_X1Y185_TQ = 1'b1;
  assign RIOI3_X105Y189_OLOGIC_X1Y190_OQ = CLBLM_R_X13Y119_SLICE_X18Y119_AQ;
  assign RIOI3_X105Y189_OLOGIC_X1Y190_TQ = 1'b1;
  assign RIOI3_X105Y189_OLOGIC_X1Y189_OQ = CLBLM_L_X8Y122_SLICE_X10Y122_AQ;
  assign RIOI3_X105Y189_OLOGIC_X1Y189_TQ = 1'b1;
  assign RIOI3_X105Y191_OLOGIC_X1Y192_OQ = CLBLM_L_X12Y115_SLICE_X16Y115_AQ;
  assign RIOI3_X105Y191_OLOGIC_X1Y192_TQ = 1'b1;
  assign RIOI3_X105Y191_OLOGIC_X1Y191_OQ = CLBLM_L_X8Y116_SLICE_X10Y116_AQ;
  assign RIOI3_X105Y191_OLOGIC_X1Y191_TQ = 1'b1;
  assign RIOI3_X105Y195_OLOGIC_X1Y196_OQ = CLBLM_R_X11Y120_SLICE_X14Y120_AQ;
  assign RIOI3_X105Y195_OLOGIC_X1Y196_TQ = 1'b1;
  assign RIOI3_X105Y195_OLOGIC_X1Y195_OQ = CLBLM_R_X11Y119_SLICE_X14Y119_AQ;
  assign RIOI3_X105Y195_OLOGIC_X1Y195_TQ = 1'b1;
  assign RIOI3_X105Y197_OLOGIC_X1Y198_OQ = CLBLM_L_X8Y122_SLICE_X10Y122_BO5;
  assign RIOI3_X105Y197_OLOGIC_X1Y198_TQ = 1'b1;
  assign RIOI3_X105Y197_OLOGIC_X1Y197_OQ = CLBLM_L_X8Y122_SLICE_X10Y122_BO5;
  assign RIOI3_X105Y197_OLOGIC_X1Y197_TQ = 1'b1;
  assign RIOI3_SING_X105Y100_ILOGIC_X1Y100_O = RIOB33_SING_X105Y100_IOB_X1Y100_I;
  assign RIOI3_SING_X105Y149_ILOGIC_X1Y149_O = RIOB33_SING_X105Y149_IOB_X1Y149_I;
  assign RIOI3_SING_X105Y150_OLOGIC_X1Y150_OQ = LIOB33_X0Y75_IOB_X0Y75_I;
  assign RIOI3_SING_X105Y150_OLOGIC_X1Y150_TQ = 1'b1;
  assign RIOI3_SING_X105Y199_OLOGIC_X1Y199_OQ = CLBLM_R_X11Y128_SLICE_X15Y128_AQ;
  assign RIOI3_SING_X105Y199_OLOGIC_X1Y199_TQ = 1'b1;
  assign RIOI3_TBYTESRC_X105Y107_ILOGIC_X1Y108_O = RIOB33_X105Y107_IOB_X1Y108_I;
  assign RIOI3_TBYTESRC_X105Y107_ILOGIC_X1Y107_O = RIOB33_X105Y107_IOB_X1Y107_I;
  assign RIOI3_TBYTESRC_X105Y119_ILOGIC_X1Y119_O = RIOB33_X105Y119_IOB_X1Y119_I;
  assign RIOI3_TBYTESRC_X105Y131_ILOGIC_X1Y132_O = RIOB33_X105Y131_IOB_X1Y132_I;
  assign RIOI3_TBYTESRC_X105Y131_ILOGIC_X1Y131_O = RIOB33_X105Y131_IOB_X1Y131_I;
  assign RIOI3_TBYTESRC_X105Y143_ILOGIC_X1Y144_O = RIOB33_X105Y143_IOB_X1Y144_I;
  assign RIOI3_TBYTESRC_X105Y143_ILOGIC_X1Y143_O = RIOB33_X105Y143_IOB_X1Y143_I;
  assign RIOI3_TBYTESRC_X105Y157_OLOGIC_X1Y158_OQ = CLBLM_R_X37Y119_SLICE_X56Y119_AO6;
  assign RIOI3_TBYTESRC_X105Y157_OLOGIC_X1Y158_TQ = 1'b1;
  assign RIOI3_TBYTESRC_X105Y157_OLOGIC_X1Y157_OQ = RIOB33_X105Y125_IOB_X1Y126_I;
  assign RIOI3_TBYTESRC_X105Y157_OLOGIC_X1Y157_TQ = 1'b1;
  assign RIOI3_TBYTESRC_X105Y169_OLOGIC_X1Y170_OQ = CLBLM_R_X103Y169_SLICE_X163Y169_AO5;
  assign RIOI3_TBYTESRC_X105Y169_OLOGIC_X1Y170_TQ = 1'b1;
  assign RIOI3_TBYTESRC_X105Y169_OLOGIC_X1Y169_OQ = CLBLM_R_X103Y169_SLICE_X163Y169_AO6;
  assign RIOI3_TBYTESRC_X105Y169_OLOGIC_X1Y169_TQ = 1'b1;
  assign RIOI3_TBYTESRC_X105Y181_OLOGIC_X1Y182_OQ = CLBLM_R_X11Y119_SLICE_X14Y119_CO5;
  assign RIOI3_TBYTESRC_X105Y181_OLOGIC_X1Y182_TQ = 1'b1;
  assign RIOI3_TBYTESRC_X105Y181_OLOGIC_X1Y181_OQ = CLBLM_R_X11Y119_SLICE_X14Y119_CO6;
  assign RIOI3_TBYTESRC_X105Y181_OLOGIC_X1Y181_TQ = 1'b1;
  assign RIOI3_TBYTESRC_X105Y193_OLOGIC_X1Y194_OQ = CLBLM_R_X11Y128_SLICE_X15Y128_AQ;
  assign RIOI3_TBYTESRC_X105Y193_OLOGIC_X1Y194_TQ = 1'b1;
  assign RIOI3_TBYTESRC_X105Y193_OLOGIC_X1Y193_OQ = CLBLM_L_X10Y124_SLICE_X13Y124_AQ;
  assign RIOI3_TBYTESRC_X105Y193_OLOGIC_X1Y193_TQ = 1'b1;
  assign RIOI3_TBYTETERM_X105Y113_ILOGIC_X1Y114_O = RIOB33_X105Y113_IOB_X1Y114_I;
  assign RIOI3_TBYTETERM_X105Y113_ILOGIC_X1Y113_O = RIOB33_X105Y113_IOB_X1Y113_I;
  assign RIOI3_TBYTETERM_X105Y137_ILOGIC_X1Y138_O = RIOB33_X105Y137_IOB_X1Y138_I;
  assign RIOI3_TBYTETERM_X105Y137_ILOGIC_X1Y137_O = RIOB33_X105Y137_IOB_X1Y137_I;
  assign RIOI3_TBYTETERM_X105Y163_OLOGIC_X1Y164_OQ = CLBLM_R_X7Y119_SLICE_X9Y119_DO5;
  assign RIOI3_TBYTETERM_X105Y163_OLOGIC_X1Y164_TQ = 1'b1;
  assign RIOI3_TBYTETERM_X105Y163_OLOGIC_X1Y163_OQ = CLBLM_R_X11Y117_SLICE_X14Y117_DO5;
  assign RIOI3_TBYTETERM_X105Y163_OLOGIC_X1Y163_TQ = 1'b1;
  assign RIOI3_TBYTETERM_X105Y187_OLOGIC_X1Y188_OQ = CLBLM_R_X11Y122_SLICE_X14Y122_AQ;
  assign RIOI3_TBYTETERM_X105Y187_OLOGIC_X1Y188_TQ = 1'b1;
  assign RIOI3_TBYTETERM_X105Y187_OLOGIC_X1Y187_OQ = CLBLM_L_X10Y114_SLICE_X12Y114_AQ;
  assign RIOI3_TBYTETERM_X105Y187_OLOGIC_X1Y187_TQ = 1'b1;
  assign CLBLM_R_X5Y121_SLICE_X6Y121_C4 = CLBLM_R_X5Y120_SLICE_X6Y120_AQ;
  assign CLBLM_R_X5Y121_SLICE_X6Y121_C5 = CLBLM_R_X5Y121_SLICE_X6Y121_B5Q;
  assign LIOB33_X0Y79_IOB_X0Y80_O = CLBLL_L_X2Y111_SLICE_X0Y111_AO6;
  assign CLBLM_R_X5Y121_SLICE_X6Y121_C6 = 1'b1;
  assign LIOB33_X0Y147_IOB_X0Y147_O = LIOB33_X0Y71_IOB_X0Y71_I;
  assign LIOB33_X0Y147_IOB_X0Y148_O = LIOB33_X0Y61_IOB_X0Y61_I;
  assign LIOI3_TBYTESRC_X0Y143_OLOGIC_X0Y143_T1 = 1'b1;
  assign CLBLM_R_X5Y121_SLICE_X6Y121_D2 = CLBLM_R_X5Y121_SLICE_X7Y121_CO6;
  assign CLBLM_R_X5Y121_SLICE_X6Y121_D3 = CLBLM_R_X5Y111_SLICE_X6Y111_AQ;
  assign LIOI3_X0Y155_OLOGIC_X0Y156_D1 = RIOB33_X105Y105_IOB_X1Y106_I;
  assign CLBLM_R_X5Y121_SLICE_X6Y121_D5 = CLBLM_R_X5Y121_SLICE_X7Y121_BO6;
  assign LIOI3_X0Y155_OLOGIC_X0Y156_T1 = 1'b1;
  assign LIOI3_X0Y155_OLOGIC_X0Y155_D1 = LIOB33_X0Y69_IOB_X0Y70_I;
  assign LIOI3_X0Y155_OLOGIC_X0Y155_T1 = 1'b1;
  assign CLBLM_R_X3Y119_SLICE_X3Y119_A1 = CLBLL_L_X4Y113_SLICE_X5Y113_CQ;
  assign CLBLM_R_X3Y119_SLICE_X3Y119_A2 = 1'b1;
  assign CLBLM_R_X3Y119_SLICE_X3Y119_A3 = CLBLM_R_X3Y119_SLICE_X3Y119_AQ;
  assign CLBLM_R_X3Y119_SLICE_X3Y119_A4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X3Y119_SLICE_X3Y119_A5 = CLBLM_R_X5Y115_SLICE_X6Y115_CO6;
  assign CLBLM_R_X3Y119_SLICE_X3Y119_A6 = CLBLL_L_X4Y123_SLICE_X4Y123_BQ;
  assign CLBLM_R_X3Y119_SLICE_X3Y119_B1 = CLBLL_L_X2Y122_SLICE_X1Y122_DO6;
  assign CLBLM_R_X3Y119_SLICE_X3Y119_B2 = RIOB33_X105Y131_IOB_X1Y131_I;
  assign CLBLM_R_X3Y119_SLICE_X3Y119_B3 = CLBLM_R_X3Y122_SLICE_X3Y122_AO6;
  assign CLBLM_R_X3Y119_SLICE_X3Y119_B4 = RIOB33_X105Y131_IOB_X1Y132_I;
  assign CLBLM_R_X3Y119_SLICE_X3Y119_B5 = CLBLM_R_X5Y122_SLICE_X7Y122_BQ;
  assign CLBLM_R_X3Y119_SLICE_X3Y119_B6 = CLBLM_L_X8Y119_SLICE_X11Y119_AQ;
  assign CLBLM_R_X3Y119_SLICE_X3Y119_C1 = CLBLL_L_X4Y120_SLICE_X5Y120_BO5;
  assign CLBLM_R_X3Y119_SLICE_X3Y119_C2 = CLBLM_L_X8Y119_SLICE_X11Y119_AQ;
  assign CLBLM_R_X3Y119_SLICE_X3Y119_C3 = CLBLL_L_X2Y120_SLICE_X0Y120_AO5;
  assign CLBLM_R_X3Y119_SLICE_X3Y119_C4 = CLBLM_R_X3Y121_SLICE_X2Y121_AO5;
  assign CLBLM_R_X3Y119_SLICE_X3Y119_C5 = CLBLM_R_X3Y113_SLICE_X3Y113_AQ;
  assign CLBLM_R_X3Y119_SLICE_X3Y119_C6 = CLBLM_R_X5Y122_SLICE_X7Y122_BQ;
  assign CLBLM_R_X3Y119_SLICE_X3Y119_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign RIOB33_SING_X105Y150_IOB_X1Y150_O = LIOB33_X0Y75_IOB_X0Y75_I;
  assign RIOI3_TBYTESRC_X105Y181_OLOGIC_X1Y182_D1 = CLBLM_R_X11Y119_SLICE_X14Y119_CO5;
  assign CLBLM_R_X3Y119_SLICE_X3Y119_D1 = 1'b1;
  assign CLBLM_R_X3Y119_SLICE_X3Y119_D2 = CLBLM_R_X3Y112_SLICE_X3Y112_C5Q;
  assign CLBLM_R_X3Y119_SLICE_X3Y119_D3 = RIOB33_X105Y109_IOB_X1Y109_I;
  assign CLBLM_R_X3Y119_SLICE_X3Y119_D4 = CLBLL_L_X2Y120_SLICE_X1Y120_AO6;
  assign CLBLM_R_X3Y119_SLICE_X3Y119_D5 = CLBLM_R_X3Y124_SLICE_X2Y124_AO6;
  assign CLBLM_R_X3Y119_SLICE_X3Y119_D6 = CLBLL_L_X2Y121_SLICE_X1Y121_BO6;
  assign RIOI3_TBYTESRC_X105Y181_OLOGIC_X1Y182_T1 = 1'b1;
  assign CLBLM_R_X3Y119_SLICE_X2Y119_A1 = CLBLL_L_X2Y119_SLICE_X1Y119_AO6;
  assign CLBLM_R_X3Y119_SLICE_X2Y119_A2 = CLBLL_L_X2Y120_SLICE_X1Y120_CO6;
  assign CLBLM_R_X3Y119_SLICE_X2Y119_A3 = CLBLM_R_X5Y118_SLICE_X6Y118_DO6;
  assign CLBLM_R_X3Y119_SLICE_X2Y119_A4 = CLBLM_R_X3Y119_SLICE_X2Y119_BO6;
  assign CLBLM_R_X3Y119_SLICE_X2Y119_A5 = CLBLM_R_X3Y118_SLICE_X2Y118_BO6;
  assign CLBLM_R_X3Y119_SLICE_X2Y119_A6 = CLBLM_R_X3Y119_SLICE_X2Y119_CO6;
  assign RIOI3_TBYTESRC_X105Y181_OLOGIC_X1Y181_D1 = CLBLM_R_X11Y119_SLICE_X14Y119_CO6;
  assign CLBLM_R_X3Y119_SLICE_X2Y119_B1 = CLBLL_L_X2Y121_SLICE_X1Y121_AO6;
  assign CLBLM_R_X3Y119_SLICE_X2Y119_B2 = CLBLL_L_X2Y122_SLICE_X0Y122_AO6;
  assign CLBLM_R_X3Y119_SLICE_X2Y119_B3 = CLBLL_L_X2Y120_SLICE_X0Y120_AO6;
  assign CLBLM_R_X3Y119_SLICE_X2Y119_B4 = RIOB33_X105Y111_IOB_X1Y112_I;
  assign CLBLM_R_X3Y119_SLICE_X2Y119_B5 = CLBLM_R_X3Y119_SLICE_X3Y119_AQ;
  assign CLBLM_R_X3Y119_SLICE_X2Y119_B6 = CLBLL_L_X4Y115_SLICE_X5Y115_DQ;
  assign CLBLM_R_X3Y119_SLICE_X2Y119_C1 = LIOB33_X0Y67_IOB_X0Y67_I;
  assign CLBLM_R_X3Y119_SLICE_X2Y119_C2 = CLBLM_R_X3Y112_SLICE_X3Y112_CQ;
  assign CLBLM_R_X3Y119_SLICE_X2Y119_C3 = CLBLL_L_X4Y122_SLICE_X4Y122_DO6;
  assign CLBLM_R_X3Y119_SLICE_X2Y119_C4 = RIOB33_X105Y137_IOB_X1Y137_I;
  assign CLBLM_R_X3Y119_SLICE_X2Y119_C5 = RIOB33_X105Y129_IOB_X1Y129_I;
  assign CLBLM_R_X3Y119_SLICE_X2Y119_C6 = CLBLL_L_X2Y121_SLICE_X0Y121_AO6;
  assign RIOI3_TBYTESRC_X105Y181_OLOGIC_X1Y181_T1 = 1'b1;
  assign CLBLM_R_X11Y123_SLICE_X15Y123_B1 = 1'b1;
  assign CLBLL_L_X4Y119_SLICE_X4Y119_A4 = CLBLL_L_X4Y115_SLICE_X4Y115_BQ;
  assign CLBLM_R_X3Y119_SLICE_X2Y119_D1 = CLBLM_R_X3Y115_SLICE_X2Y115_AQ;
  assign CLBLM_R_X3Y119_SLICE_X2Y119_D2 = RIOB33_X105Y135_IOB_X1Y136_I;
  assign CLBLM_R_X3Y119_SLICE_X2Y119_D3 = RIOB33_X105Y135_IOB_X1Y135_I;
  assign CLBLM_R_X3Y119_SLICE_X2Y119_D4 = CLBLM_R_X3Y122_SLICE_X3Y122_AO5;
  assign CLBLM_R_X3Y119_SLICE_X2Y119_D5 = RIOB33_X105Y111_IOB_X1Y111_I;
  assign CLBLM_R_X3Y119_SLICE_X2Y119_D6 = CLBLL_L_X2Y121_SLICE_X1Y121_BO6;
  assign CLBLL_L_X4Y119_SLICE_X4Y119_A5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLL_L_X4Y119_SLICE_X4Y119_A6 = CLBLM_R_X5Y115_SLICE_X6Y115_CO5;
  assign RIOB33_X105Y157_IOB_X1Y158_O = CLBLM_R_X37Y119_SLICE_X56Y119_AO6;
  assign RIOB33_X105Y157_IOB_X1Y157_O = RIOB33_X105Y125_IOB_X1Y126_I;
  assign CLBLL_L_X4Y119_SLICE_X4Y119_B1 = CLBLM_R_X7Y121_SLICE_X9Y121_AQ;
  assign CLBLL_L_X4Y119_SLICE_X4Y119_B3 = CLBLL_L_X2Y116_SLICE_X1Y116_AQ;
  assign CLBLL_L_X4Y119_SLICE_X4Y119_B4 = RIOB33_X105Y127_IOB_X1Y127_I;
  assign LIOI3_SING_X0Y199_OLOGIC_X0Y199_D1 = LIOB33_X0Y73_IOB_X0Y74_I;
  assign LIOB33_X0Y151_IOB_X0Y152_O = LIOB33_X0Y65_IOB_X0Y66_I;
  assign LIOB33_X0Y151_IOB_X0Y151_O = LIOB33_X0Y65_IOB_X0Y65_I;
  assign CLBLL_L_X4Y119_SLICE_X4Y119_C2 = CLBLM_R_X5Y110_SLICE_X7Y110_BQ;
  assign RIOB33_SING_X105Y199_IOB_X1Y199_O = CLBLM_R_X11Y128_SLICE_X15Y128_AQ;
  assign CLBLL_L_X4Y119_SLICE_X4Y119_C3 = CLBLM_R_X3Y119_SLICE_X3Y119_AQ;
  assign LIOI3_SING_X0Y199_OLOGIC_X0Y199_T1 = 1'b1;
  assign CLBLL_L_X4Y119_SLICE_X4Y119_C4 = CLBLL_L_X4Y116_SLICE_X5Y116_A5Q;
  assign RIOI3_X105Y139_ILOGIC_X1Y140_D = RIOB33_X105Y139_IOB_X1Y140_I;
  assign RIOI3_X105Y139_ILOGIC_X1Y139_D = RIOB33_X105Y139_IOB_X1Y139_I;
  assign RIOI3_X105Y109_ILOGIC_X1Y110_D = RIOB33_X105Y109_IOB_X1Y110_I;
  assign RIOI3_X105Y109_ILOGIC_X1Y109_D = RIOB33_X105Y109_IOB_X1Y109_I;
  assign CLBLM_R_X11Y128_SLICE_X15Y128_B5 = 1'b1;
  assign CLBLM_R_X11Y128_SLICE_X15Y128_B6 = 1'b1;
  assign CLBLM_L_X8Y117_SLICE_X11Y117_A1 = CLBLM_L_X8Y121_SLICE_X10Y121_DO6;
  assign CLBLM_R_X3Y120_SLICE_X3Y120_A1 = CLBLM_R_X3Y122_SLICE_X3Y122_AO5;
  assign CLBLM_R_X3Y120_SLICE_X3Y120_A2 = CLBLL_L_X2Y121_SLICE_X1Y121_BO6;
  assign CLBLM_R_X3Y120_SLICE_X3Y120_A3 = RIOB33_X105Y135_IOB_X1Y136_I;
  assign CLBLM_R_X3Y120_SLICE_X3Y120_A4 = RIOB33_X105Y111_IOB_X1Y112_I;
  assign CLBLM_R_X3Y120_SLICE_X3Y120_A5 = CLBLM_R_X3Y119_SLICE_X3Y119_AQ;
  assign CLBLM_R_X3Y120_SLICE_X3Y120_A6 = RIOB33_X105Y135_IOB_X1Y135_I;
  assign CLBLM_R_X3Y120_SLICE_X3Y120_B1 = CLBLM_R_X3Y118_SLICE_X3Y118_DO6;
  assign CLBLM_R_X3Y120_SLICE_X3Y120_B2 = CLBLL_L_X4Y120_SLICE_X5Y120_CO6;
  assign CLBLM_R_X3Y120_SLICE_X3Y120_B3 = CLBLL_L_X2Y121_SLICE_X1Y121_CO6;
  assign CLBLM_R_X3Y120_SLICE_X3Y120_B4 = CLBLM_R_X3Y120_SLICE_X3Y120_DO6;
  assign CLBLM_R_X3Y120_SLICE_X3Y120_B5 = CLBLM_R_X3Y122_SLICE_X2Y122_DO6;
  assign CLBLM_R_X3Y120_SLICE_X3Y120_B6 = CLBLM_R_X3Y118_SLICE_X3Y118_CO6;
  assign CLBLM_R_X11Y128_SLICE_X15Y128_C4 = 1'b1;
  assign CLBLM_R_X11Y128_SLICE_X15Y128_C5 = 1'b1;
  assign CLBLM_R_X3Y120_SLICE_X3Y120_C1 = CLBLM_R_X3Y112_SLICE_X2Y112_BQ;
  assign CLBLM_R_X3Y120_SLICE_X3Y120_C2 = CLBLL_L_X4Y122_SLICE_X4Y122_AO6;
  assign CLBLM_R_X3Y120_SLICE_X3Y120_C3 = CLBLM_R_X3Y124_SLICE_X2Y124_AO6;
  assign CLBLM_R_X3Y120_SLICE_X3Y120_C4 = 1'b1;
  assign CLBLM_R_X3Y120_SLICE_X3Y120_C5 = CLBLL_L_X4Y114_SLICE_X4Y114_CQ;
  assign CLBLM_R_X3Y120_SLICE_X3Y120_C6 = RIOB33_X105Y131_IOB_X1Y131_I;
  assign CLBLM_R_X11Y128_SLICE_X15Y128_C6 = 1'b1;
  assign CLBLM_R_X3Y120_SLICE_X3Y120_D1 = CLBLL_L_X2Y121_SLICE_X1Y121_AO6;
  assign CLBLM_R_X3Y120_SLICE_X3Y120_D2 = CLBLM_R_X3Y119_SLICE_X3Y119_DO6;
  assign CLBLM_R_X3Y120_SLICE_X3Y120_D3 = CLBLM_R_X3Y115_SLICE_X2Y115_DQ;
  assign CLBLM_R_X3Y120_SLICE_X3Y120_D4 = 1'b1;
  assign CLBLM_R_X3Y120_SLICE_X3Y120_D5 = CLBLM_R_X5Y120_SLICE_X7Y120_BQ;
  assign CLBLM_R_X3Y120_SLICE_X3Y120_D6 = CLBLL_L_X2Y120_SLICE_X0Y120_AO6;
  assign CLBLM_L_X12Y120_SLICE_X17Y120_C1 = CLBLM_R_X11Y118_SLICE_X14Y118_BQ;
  assign CLBLM_L_X12Y120_SLICE_X17Y120_C2 = CLBLM_L_X12Y120_SLICE_X16Y120_AO5;
  assign CLBLM_R_X3Y120_SLICE_X2Y120_A1 = CLBLL_L_X4Y122_SLICE_X4Y122_DO6;
  assign CLBLM_R_X3Y120_SLICE_X2Y120_A2 = CLBLL_L_X4Y115_SLICE_X5Y115_DQ;
  assign CLBLM_R_X3Y120_SLICE_X2Y120_A3 = CLBLM_R_X3Y120_SLICE_X3Y120_AO6;
  assign CLBLM_R_X3Y120_SLICE_X2Y120_A4 = CLBLM_R_X3Y120_SLICE_X2Y120_BO6;
  assign CLBLM_R_X3Y120_SLICE_X2Y120_A5 = CLBLL_L_X2Y121_SLICE_X1Y121_AO6;
  assign CLBLM_R_X3Y120_SLICE_X2Y120_A6 = CLBLM_R_X3Y118_SLICE_X2Y118_BO6;
  assign CLBLM_R_X3Y120_SLICE_X2Y120_B1 = CLBLM_R_X3Y124_SLICE_X2Y124_AO5;
  assign CLBLM_R_X3Y120_SLICE_X2Y120_B2 = RIOB33_X105Y129_IOB_X1Y129_I;
  assign CLBLM_R_X3Y120_SLICE_X2Y120_B3 = RIOB33_X105Y137_IOB_X1Y137_I;
  assign CLBLM_R_X3Y120_SLICE_X2Y120_B4 = CLBLL_L_X2Y121_SLICE_X1Y121_BO6;
  assign CLBLM_R_X3Y120_SLICE_X2Y120_B5 = CLBLM_R_X3Y112_SLICE_X3Y112_CQ;
  assign CLBLM_R_X3Y120_SLICE_X2Y120_B6 = LIOB33_X0Y67_IOB_X0Y67_I;
  assign CLBLM_R_X3Y120_SLICE_X2Y120_C1 = CLBLM_R_X3Y111_SLICE_X2Y111_AQ;
  assign CLBLM_R_X3Y120_SLICE_X2Y120_C2 = CLBLL_L_X2Y120_SLICE_X1Y120_AO6;
  assign CLBLM_R_X3Y120_SLICE_X2Y120_C3 = CLBLL_L_X2Y121_SLICE_X0Y121_BO6;
  assign CLBLM_R_X3Y120_SLICE_X2Y120_C4 = CLBLM_R_X3Y122_SLICE_X3Y122_AO6;
  assign CLBLM_R_X3Y120_SLICE_X2Y120_C5 = 1'b1;
  assign CLBLM_R_X3Y120_SLICE_X2Y120_C6 = CLBLM_R_X3Y116_SLICE_X2Y116_BQ;
  assign CLBLM_L_X12Y120_SLICE_X17Y120_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X11Y128_SLICE_X15Y128_D2 = 1'b1;
  assign CLBLM_L_X8Y117_SLICE_X11Y117_A5 = RIOB33_X105Y135_IOB_X1Y136_I;
  assign CLBLM_L_X10Y126_SLICE_X12Y126_C1 = 1'b1;
  assign CLBLM_R_X3Y120_SLICE_X2Y120_D1 = CLBLM_R_X3Y111_SLICE_X2Y111_AQ;
  assign CLBLM_R_X3Y120_SLICE_X2Y120_D2 = 1'b1;
  assign CLBLM_R_X3Y120_SLICE_X2Y120_D3 = CLBLM_R_X3Y119_SLICE_X2Y119_DO6;
  assign CLBLM_R_X3Y120_SLICE_X2Y120_D4 = CLBLL_L_X4Y120_SLICE_X5Y120_BO6;
  assign CLBLM_R_X3Y120_SLICE_X2Y120_D5 = CLBLM_R_X3Y122_SLICE_X2Y122_BO5;
  assign CLBLM_R_X3Y120_SLICE_X2Y120_D6 = CLBLM_R_X3Y116_SLICE_X2Y116_BQ;
  assign CLBLM_R_X11Y123_SLICE_X15Y123_C4 = 1'b1;
  assign CLBLM_L_X12Y115_SLICE_X17Y115_A1 = 1'b1;
  assign CLBLM_L_X12Y115_SLICE_X17Y115_A2 = 1'b1;
  assign CLBLM_L_X12Y115_SLICE_X17Y115_A3 = 1'b1;
  assign CLBLM_L_X12Y115_SLICE_X17Y115_A4 = 1'b1;
  assign CLBLM_L_X12Y115_SLICE_X17Y115_A5 = 1'b1;
  assign CLBLM_L_X12Y115_SLICE_X17Y115_A6 = 1'b1;
  assign CLBLM_R_X11Y128_SLICE_X15Y128_D6 = 1'b1;
  assign CLBLM_L_X12Y115_SLICE_X17Y115_B1 = 1'b1;
  assign CLBLM_L_X12Y115_SLICE_X17Y115_B2 = 1'b1;
  assign CLBLM_L_X12Y115_SLICE_X17Y115_B3 = 1'b1;
  assign CLBLM_L_X12Y115_SLICE_X17Y115_B4 = 1'b1;
  assign CLBLM_L_X12Y115_SLICE_X17Y115_B5 = 1'b1;
  assign CLBLM_L_X12Y115_SLICE_X17Y115_B6 = 1'b1;
  assign CLBLL_L_X4Y119_SLICE_X5Y119_A2 = CLBLM_R_X5Y115_SLICE_X6Y115_CO5;
  assign CLBLM_L_X12Y115_SLICE_X17Y115_C1 = 1'b1;
  assign CLBLM_L_X12Y115_SLICE_X17Y115_C2 = 1'b1;
  assign CLBLM_L_X12Y115_SLICE_X17Y115_C3 = 1'b1;
  assign CLBLM_L_X12Y115_SLICE_X17Y115_C4 = 1'b1;
  assign CLBLM_L_X12Y115_SLICE_X17Y115_C5 = 1'b1;
  assign CLBLM_L_X12Y115_SLICE_X17Y115_C6 = 1'b1;
  assign CLBLM_R_X11Y123_SLICE_X15Y123_C5 = 1'b1;
  assign CLBLM_R_X37Y119_SLICE_X57Y119_A1 = 1'b1;
  assign CLBLM_L_X12Y120_SLICE_X17Y120_D3 = 1'b1;
  assign CLBLM_R_X37Y119_SLICE_X57Y119_A2 = 1'b1;
  assign CLBLM_R_X37Y119_SLICE_X57Y119_A3 = 1'b1;
  assign CLBLM_R_X37Y119_SLICE_X57Y119_A4 = 1'b1;
  assign CLBLM_R_X37Y119_SLICE_X57Y119_A5 = 1'b1;
  assign CLBLM_R_X37Y119_SLICE_X57Y119_A6 = 1'b1;
  assign CLBLM_L_X12Y115_SLICE_X17Y115_D1 = 1'b1;
  assign CLBLM_L_X12Y115_SLICE_X17Y115_D2 = 1'b1;
  assign CLBLM_L_X12Y115_SLICE_X17Y115_D3 = 1'b1;
  assign CLBLM_L_X12Y115_SLICE_X17Y115_D4 = 1'b1;
  assign CLBLM_L_X12Y115_SLICE_X17Y115_D5 = 1'b1;
  assign CLBLM_L_X12Y115_SLICE_X17Y115_D6 = 1'b1;
  assign CLBLM_L_X12Y120_SLICE_X17Y120_D5 = CLBLM_L_X10Y119_SLICE_X13Y119_AQ;
  assign CLBLL_L_X4Y119_SLICE_X5Y119_A6 = CLBLM_R_X7Y117_SLICE_X8Y117_CQ;
  assign CLBLM_L_X12Y120_SLICE_X17Y120_D6 = 1'b1;
  assign CLBLM_R_X13Y119_SLICE_X19Y119_D1 = 1'b1;
  assign CLBLM_R_X37Y119_SLICE_X57Y119_B2 = 1'b1;
  assign CLBLM_R_X11Y123_SLICE_X15Y123_C6 = 1'b1;
  assign CLBLM_L_X12Y115_SLICE_X16Y115_A1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X12Y115_SLICE_X16Y115_A2 = 1'b1;
  assign CLBLM_L_X12Y115_SLICE_X16Y115_A3 = CLBLM_L_X12Y115_SLICE_X16Y115_AQ;
  assign CLBLM_L_X12Y115_SLICE_X16Y115_A4 = CLBLM_R_X7Y128_SLICE_X8Y128_AQ;
  assign CLBLM_L_X12Y115_SLICE_X16Y115_A5 = RIOB33_X105Y141_IOB_X1Y142_I;
  assign CLBLM_L_X12Y115_SLICE_X16Y115_A6 = CLBLM_R_X7Y115_SLICE_X9Y115_B5Q;
  assign CLBLM_R_X37Y119_SLICE_X57Y119_C1 = 1'b1;
  assign CLBLM_R_X37Y119_SLICE_X57Y119_C2 = 1'b1;
  assign CLBLM_R_X37Y119_SLICE_X57Y119_C3 = 1'b1;
  assign CLBLM_L_X12Y115_SLICE_X16Y115_B1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X12Y115_SLICE_X16Y115_B2 = CLBLM_L_X12Y115_SLICE_X16Y115_BQ;
  assign CLBLM_L_X12Y115_SLICE_X16Y115_B3 = CLBLM_R_X7Y114_SLICE_X8Y114_AQ;
  assign CLBLM_L_X12Y115_SLICE_X16Y115_B4 = CLBLM_R_X7Y128_SLICE_X8Y128_AQ;
  assign CLBLM_L_X12Y115_SLICE_X16Y115_B5 = RIOB33_X105Y141_IOB_X1Y142_I;
  assign CLBLM_L_X12Y115_SLICE_X16Y115_B6 = 1'b1;
  assign CLBLM_R_X13Y119_SLICE_X19Y119_D2 = 1'b1;
  assign CLBLM_R_X37Y119_SLICE_X57Y119_D1 = 1'b1;
  assign CLBLM_R_X37Y119_SLICE_X57Y119_D2 = 1'b1;
  assign CLBLM_L_X12Y115_SLICE_X16Y115_C1 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_L_X12Y115_SLICE_X16Y115_C2 = CLBLM_L_X12Y115_SLICE_X16Y115_CQ;
  assign CLBLM_L_X12Y115_SLICE_X16Y115_C3 = CLBLM_L_X12Y115_SLICE_X16Y115_DQ;
  assign CLBLM_L_X12Y115_SLICE_X16Y115_C4 = CLBLM_L_X12Y115_SLICE_X16Y115_BQ;
  assign CLBLM_L_X12Y115_SLICE_X16Y115_C5 = CLBLM_R_X3Y118_SLICE_X2Y118_AQ;
  assign CLBLM_L_X12Y115_SLICE_X16Y115_C6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLL_L_X4Y119_SLICE_X5Y119_B4 = CLBLL_L_X2Y120_SLICE_X0Y120_AO6;
  assign CLBLM_R_X37Y119_SLICE_X56Y119_A1 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_R_X37Y119_SLICE_X56Y119_A2 = CLBLM_R_X3Y117_SLICE_X3Y117_CQ;
  assign CLBLM_L_X12Y115_SLICE_X16Y115_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X37Y119_SLICE_X56Y119_A3 = 1'b1;
  assign CLBLM_R_X37Y119_SLICE_X56Y119_A4 = RIOB33_X105Y119_IOB_X1Y119_I;
  assign CLBLM_R_X37Y119_SLICE_X56Y119_A5 = 1'b1;
  assign CLBLM_R_X37Y119_SLICE_X56Y119_A6 = 1'b1;
  assign CLBLM_L_X12Y115_SLICE_X16Y115_D1 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_L_X12Y115_SLICE_X16Y115_D2 = CLBLM_L_X10Y114_SLICE_X13Y114_AQ;
  assign CLBLM_L_X12Y115_SLICE_X16Y115_D3 = CLBLM_L_X12Y115_SLICE_X16Y115_DQ;
  assign CLBLM_L_X12Y115_SLICE_X16Y115_D4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X12Y115_SLICE_X16Y115_D5 = CLBLM_R_X3Y118_SLICE_X2Y118_AQ;
  assign CLBLM_L_X12Y115_SLICE_X16Y115_D6 = CLBLM_L_X10Y114_SLICE_X13Y114_CQ;
  assign CLBLM_R_X13Y119_SLICE_X19Y119_D3 = 1'b1;
  assign CLBLM_R_X37Y119_SLICE_X56Y119_B1 = 1'b1;
  assign CLBLM_R_X37Y119_SLICE_X56Y119_B2 = 1'b1;
  assign CLBLM_R_X37Y119_SLICE_X56Y119_B3 = 1'b1;
  assign CLBLM_R_X37Y119_SLICE_X56Y119_B4 = 1'b1;
  assign CLBLM_R_X37Y119_SLICE_X56Y119_B5 = 1'b1;
  assign CLBLM_R_X37Y119_SLICE_X56Y119_B6 = 1'b1;
  assign CLBLM_R_X37Y119_SLICE_X56Y119_C1 = 1'b1;
  assign CLBLM_L_X12Y120_SLICE_X16Y120_A5 = CLBLM_L_X12Y121_SLICE_X16Y121_AQ;
  assign CLBLM_R_X37Y119_SLICE_X56Y119_C2 = 1'b1;
  assign CLBLM_R_X37Y119_SLICE_X56Y119_C3 = 1'b1;
  assign CLBLM_R_X37Y119_SLICE_X56Y119_C4 = 1'b1;
  assign CLBLM_R_X37Y119_SLICE_X56Y119_C5 = 1'b1;
  assign CLBLM_L_X12Y120_SLICE_X16Y120_A6 = 1'b1;
  assign CLBLM_R_X37Y119_SLICE_X56Y119_C6 = 1'b1;
  assign CLBLM_R_X13Y119_SLICE_X19Y119_D4 = 1'b1;
  assign CLBLM_R_X37Y119_SLICE_X56Y119_D1 = 1'b1;
  assign CLBLM_R_X37Y119_SLICE_X56Y119_D2 = 1'b1;
  assign CLBLM_R_X37Y119_SLICE_X56Y119_D3 = 1'b1;
  assign CLBLM_R_X37Y119_SLICE_X56Y119_D4 = 1'b1;
  assign CLBLM_R_X37Y119_SLICE_X56Y119_D5 = 1'b1;
  assign CLBLL_L_X4Y119_SLICE_X5Y119_C2 = RIOB33_X105Y133_IOB_X1Y133_I;
  assign CLBLM_L_X10Y122_SLICE_X13Y122_C1 = CLBLM_R_X11Y122_SLICE_X14Y122_BO6;
  assign CLBLM_R_X11Y128_SLICE_X14Y128_B5 = 1'b1;
  assign CLBLM_R_X37Y119_SLICE_X56Y119_D6 = 1'b1;
  assign CLBLL_L_X4Y119_SLICE_X5Y119_C3 = RIOB33_X105Y131_IOB_X1Y132_I;
  assign CLBLM_R_X11Y128_SLICE_X14Y128_B6 = 1'b1;
  assign RIOB33_X105Y169_IOB_X1Y170_O = CLBLM_R_X103Y169_SLICE_X163Y169_AO5;
  assign CLBLM_R_X13Y119_SLICE_X19Y119_D5 = 1'b1;
  assign RIOB33_X105Y169_IOB_X1Y169_O = CLBLM_R_X103Y169_SLICE_X163Y169_AO6;
  assign RIOI3_X105Y195_OLOGIC_X1Y196_D1 = CLBLM_R_X11Y120_SLICE_X14Y120_AQ;
  assign CLBLM_R_X13Y119_SLICE_X19Y119_D6 = 1'b1;
  assign CLBLM_R_X11Y128_SLICE_X14Y128_C3 = 1'b1;
  assign CLBLM_R_X11Y128_SLICE_X14Y128_C4 = 1'b1;
  assign CLBLM_R_X11Y128_SLICE_X14Y128_C5 = 1'b1;
  assign CLBLM_R_X11Y128_SLICE_X14Y128_C6 = 1'b1;
  assign RIOI3_X105Y195_OLOGIC_X1Y196_T1 = 1'b1;
  assign CLBLM_R_X3Y121_SLICE_X3Y121_A1 = CLBLM_R_X3Y117_SLICE_X3Y117_DO6;
  assign CLBLM_R_X3Y121_SLICE_X3Y121_A2 = CLBLM_R_X3Y122_SLICE_X3Y122_BO6;
  assign CLBLM_R_X3Y121_SLICE_X3Y121_A3 = CLBLM_R_X3Y119_SLICE_X3Y119_BO6;
  assign CLBLM_R_X3Y121_SLICE_X3Y121_A4 = CLBLM_R_X3Y121_SLICE_X3Y121_BO6;
  assign CLBLM_R_X3Y121_SLICE_X3Y121_A5 = CLBLM_R_X3Y120_SLICE_X2Y120_CO6;
  assign CLBLM_R_X3Y121_SLICE_X3Y121_A6 = CLBLM_R_X3Y119_SLICE_X2Y119_DO6;
  assign CLBLM_R_X11Y121_SLICE_X15Y121_B2 = 1'b1;
  assign CLBLM_R_X3Y121_SLICE_X3Y121_B1 = CLBLM_R_X3Y124_SLICE_X2Y124_AO5;
  assign CLBLM_R_X3Y121_SLICE_X3Y121_B2 = CLBLM_R_X5Y120_SLICE_X7Y120_CQ;
  assign CLBLM_R_X3Y121_SLICE_X3Y121_B3 = CLBLL_L_X2Y121_SLICE_X1Y121_BO5;
  assign CLBLM_R_X3Y121_SLICE_X3Y121_B4 = LIOB33_X0Y65_IOB_X0Y66_I;
  assign CLBLM_R_X3Y121_SLICE_X3Y121_B5 = CLBLM_L_X8Y122_SLICE_X10Y122_BO6;
  assign CLBLM_R_X3Y121_SLICE_X3Y121_B6 = CLBLL_L_X2Y121_SLICE_X1Y121_BO6;
  assign CLBLM_R_X3Y121_SLICE_X3Y121_C1 = RIOB33_X105Y131_IOB_X1Y132_I;
  assign CLBLM_R_X3Y121_SLICE_X3Y121_C2 = RIOB33_X105Y129_IOB_X1Y129_I;
  assign CLBLM_R_X3Y121_SLICE_X3Y121_C3 = RIOB33_X105Y135_IOB_X1Y136_I;
  assign CLBLM_R_X3Y121_SLICE_X3Y121_C4 = RIOB33_X105Y137_IOB_X1Y137_I;
  assign CLBLM_R_X3Y121_SLICE_X3Y121_C5 = RIOB33_X105Y129_IOB_X1Y130_I;
  assign CLBLM_R_X3Y121_SLICE_X3Y121_C6 = RIOB33_X105Y135_IOB_X1Y135_I;
  assign CLBLM_R_X11Y121_SLICE_X15Y121_B3 = CLBLM_R_X11Y118_SLICE_X14Y118_BQ;
  assign CLBLM_R_X3Y121_SLICE_X3Y121_D1 = CLBLM_L_X8Y122_SLICE_X10Y122_BO6;
  assign CLBLM_R_X3Y121_SLICE_X3Y121_D2 = CLBLM_R_X5Y120_SLICE_X7Y120_CQ;
  assign CLBLM_R_X3Y121_SLICE_X3Y121_D3 = CLBLM_R_X3Y123_SLICE_X3Y123_BO5;
  assign CLBLM_R_X3Y121_SLICE_X3Y121_D4 = CLBLM_R_X3Y117_SLICE_X3Y117_DO6;
  assign CLBLM_R_X3Y121_SLICE_X3Y121_D5 = LIOB33_X0Y65_IOB_X0Y66_I;
  assign CLBLM_R_X3Y121_SLICE_X3Y121_D6 = CLBLL_L_X2Y121_SLICE_X0Y121_AO6;
  assign CLBLM_R_X3Y121_SLICE_X2Y121_A1 = CLBLM_R_X3Y124_SLICE_X2Y124_AO6;
  assign CLBLM_R_X3Y121_SLICE_X2Y121_A2 = RIOB33_X105Y131_IOB_X1Y132_I;
  assign CLBLM_R_X3Y121_SLICE_X2Y121_A3 = RIOB33_X105Y133_IOB_X1Y134_I;
  assign CLBLM_R_X3Y121_SLICE_X2Y121_A4 = RIOB33_X105Y133_IOB_X1Y133_I;
  assign CLBLM_R_X3Y121_SLICE_X2Y121_A5 = RIOB33_X105Y131_IOB_X1Y131_I;
  assign CLBLM_R_X3Y121_SLICE_X2Y121_A6 = 1'b1;
  assign CLBLM_R_X11Y121_SLICE_X15Y121_B4 = 1'b1;
  assign CLBLM_R_X3Y121_SLICE_X2Y121_B1 = CLBLM_R_X3Y122_SLICE_X2Y122_CO6;
  assign CLBLM_R_X3Y121_SLICE_X2Y121_B2 = CLBLL_L_X4Y121_SLICE_X4Y121_DO6;
  assign CLBLM_R_X3Y121_SLICE_X2Y121_B3 = CLBLM_R_X3Y122_SLICE_X2Y122_AO6;
  assign CLBLM_R_X3Y121_SLICE_X2Y121_B4 = CLBLL_L_X2Y121_SLICE_X1Y121_AO6;
  assign CLBLM_R_X3Y121_SLICE_X2Y121_B5 = CLBLL_L_X2Y119_SLICE_X1Y119_AO6;
  assign CLBLM_R_X3Y121_SLICE_X2Y121_B6 = CLBLM_R_X3Y121_SLICE_X2Y121_AO5;
  assign LIOI3_X0Y159_OLOGIC_X0Y160_D1 = RIOB33_X105Y107_IOB_X1Y107_I;
  assign CLBLM_R_X3Y121_SLICE_X2Y121_C1 = CLBLM_R_X5Y118_SLICE_X6Y118_DO6;
  assign CLBLM_R_X3Y121_SLICE_X2Y121_C2 = CLBLM_R_X3Y121_SLICE_X3Y121_AO6;
  assign CLBLM_R_X3Y121_SLICE_X2Y121_C3 = CLBLM_R_X3Y120_SLICE_X2Y120_AO6;
  assign CLBLM_R_X3Y121_SLICE_X2Y121_C4 = CLBLL_L_X2Y121_SLICE_X1Y121_DO6;
  assign CLBLM_R_X3Y121_SLICE_X2Y121_C5 = CLBLL_L_X4Y122_SLICE_X5Y122_DO6;
  assign CLBLM_R_X3Y121_SLICE_X2Y121_C6 = CLBLM_R_X3Y121_SLICE_X2Y121_BO6;
  assign LIOI3_X0Y159_OLOGIC_X0Y160_T1 = 1'b1;
  assign CLBLM_R_X11Y121_SLICE_X15Y121_B5 = 1'b1;
  assign CLBLM_R_X3Y121_SLICE_X2Y121_D1 = CLBLM_R_X3Y122_SLICE_X2Y122_AO6;
  assign CLBLM_R_X3Y121_SLICE_X2Y121_D2 = CLBLL_L_X4Y121_SLICE_X4Y121_CO5;
  assign CLBLM_R_X3Y121_SLICE_X2Y121_D3 = CLBLM_R_X3Y122_SLICE_X2Y122_BO6;
  assign CLBLM_R_X3Y121_SLICE_X2Y121_D4 = CLBLL_L_X4Y121_SLICE_X5Y121_BO6;
  assign CLBLM_R_X3Y121_SLICE_X2Y121_D5 = CLBLL_L_X2Y120_SLICE_X0Y120_AO6;
  assign CLBLM_R_X3Y121_SLICE_X2Y121_D6 = CLBLM_R_X3Y123_SLICE_X3Y123_BO6;
  assign LIOI3_X0Y159_OLOGIC_X0Y159_D1 = RIOB33_X105Y117_IOB_X1Y117_I;
  assign LIOI3_X0Y159_OLOGIC_X0Y159_T1 = 1'b1;
  assign LIOB33_X0Y155_IOB_X0Y156_O = RIOB33_X105Y105_IOB_X1Y106_I;
  assign CLBLM_R_X11Y121_SLICE_X15Y121_B6 = CLBLM_R_X13Y119_SLICE_X18Y119_CQ;
  assign LIOB33_X0Y155_IOB_X0Y155_O = LIOB33_X0Y69_IOB_X0Y70_I;
  assign LIOB33_X0Y153_IOB_X0Y154_O = LIOB33_X0Y67_IOB_X0Y68_I;
  assign LIOB33_X0Y153_IOB_X0Y153_O = LIOB33_X0Y67_IOB_X0Y67_I;
  assign CLBLM_R_X13Y119_SLICE_X18Y119_A1 = CLBLM_L_X12Y118_SLICE_X16Y118_AQ;
  assign CLBLM_L_X10Y122_SLICE_X12Y122_C1 = CLBLM_L_X10Y124_SLICE_X12Y124_AQ;
  assign RIOI3_TBYTESRC_X105Y193_OLOGIC_X1Y194_D1 = CLBLM_R_X11Y128_SLICE_X15Y128_AQ;
  assign RIOI3_TBYTESRC_X105Y193_OLOGIC_X1Y194_T1 = 1'b1;
  assign CLBLM_L_X10Y122_SLICE_X12Y122_C5 = CLBLM_R_X7Y120_SLICE_X9Y120_A5Q;
  assign CLBLM_R_X13Y119_SLICE_X18Y119_A2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y122_SLICE_X12Y122_C6 = 1'b1;
  assign RIOI3_TBYTESRC_X105Y193_OLOGIC_X1Y193_D1 = CLBLM_L_X10Y124_SLICE_X13Y124_AQ;
  assign RIOI3_TBYTESRC_X105Y193_OLOGIC_X1Y193_T1 = 1'b1;
  assign RIOI3_TBYTETERM_X105Y113_ILOGIC_X1Y114_D = RIOB33_X105Y113_IOB_X1Y114_I;
  assign CLBLM_L_X10Y122_SLICE_X12Y122_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X13Y119_SLICE_X18Y119_A3 = CLBLM_R_X13Y119_SLICE_X18Y119_AQ;
  assign CLBLM_R_X13Y119_SLICE_X18Y119_A4 = RIOB33_X105Y141_IOB_X1Y142_I;
  assign CLBLM_R_X13Y119_SLICE_X18Y119_A5 = CLBLM_R_X7Y128_SLICE_X8Y128_AQ;
  assign RIOB33_X105Y167_IOB_X1Y168_O = CLBLM_R_X7Y151_SLICE_X8Y151_AO6;
  assign RIOI3_X105Y141_ILOGIC_X1Y142_D = RIOB33_X105Y141_IOB_X1Y142_I;
  assign RIOI3_X105Y141_ILOGIC_X1Y141_D = RIOB33_X105Y141_IOB_X1Y141_I;
  assign CLBLM_R_X3Y122_SLICE_X3Y122_A1 = RIOB33_X105Y129_IOB_X1Y129_I;
  assign CLBLM_R_X3Y122_SLICE_X3Y122_A2 = RIOB33_X105Y135_IOB_X1Y135_I;
  assign CLBLM_R_X3Y122_SLICE_X3Y122_A3 = RIOB33_X105Y129_IOB_X1Y130_I;
  assign CLBLM_R_X3Y122_SLICE_X3Y122_A4 = RIOB33_X105Y137_IOB_X1Y137_I;
  assign CLBLM_R_X3Y122_SLICE_X3Y122_A5 = RIOB33_X105Y135_IOB_X1Y136_I;
  assign CLBLM_R_X3Y122_SLICE_X3Y122_A6 = 1'b1;
  assign CLBLM_R_X3Y122_SLICE_X3Y122_B1 = CLBLM_R_X3Y113_SLICE_X3Y113_AQ;
  assign CLBLM_R_X3Y122_SLICE_X3Y122_B2 = RIOB33_X105Y131_IOB_X1Y131_I;
  assign CLBLM_R_X3Y122_SLICE_X3Y122_B3 = RIOB33_X105Y133_IOB_X1Y134_I;
  assign CLBLM_R_X3Y122_SLICE_X3Y122_B4 = CLBLM_R_X3Y124_SLICE_X2Y124_AO6;
  assign CLBLM_R_X3Y122_SLICE_X3Y122_B5 = RIOB33_X105Y133_IOB_X1Y133_I;
  assign CLBLM_R_X3Y122_SLICE_X3Y122_B6 = RIOB33_X105Y131_IOB_X1Y132_I;
  assign CLBLM_R_X3Y122_SLICE_X3Y122_C1 = RIOB33_X105Y137_IOB_X1Y137_I;
  assign CLBLM_R_X3Y122_SLICE_X3Y122_C2 = CLBLL_L_X2Y121_SLICE_X1Y121_BO6;
  assign CLBLM_R_X3Y122_SLICE_X3Y122_C3 = CLBLM_R_X3Y124_SLICE_X2Y124_AO5;
  assign CLBLM_R_X3Y122_SLICE_X3Y122_C4 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X3Y122_SLICE_X3Y122_C5 = RIOB33_X105Y129_IOB_X1Y129_I;
  assign CLBLM_R_X3Y122_SLICE_X3Y122_C6 = CLBLM_R_X5Y120_SLICE_X6Y120_AQ;
  assign CLBLM_R_X3Y122_SLICE_X3Y122_D1 = CLBLM_R_X5Y122_SLICE_X7Y122_AQ;
  assign CLBLM_R_X3Y122_SLICE_X3Y122_D2 = RIOB33_X105Y137_IOB_X1Y137_I;
  assign CLBLM_R_X3Y122_SLICE_X3Y122_D3 = CLBLL_L_X2Y121_SLICE_X0Y121_BO6;
  assign CLBLM_R_X3Y122_SLICE_X3Y122_D4 = RIOB33_X105Y117_IOB_X1Y117_I;
  assign CLBLM_R_X3Y122_SLICE_X3Y122_D5 = RIOB33_X105Y129_IOB_X1Y129_I;
  assign CLBLM_R_X3Y122_SLICE_X3Y122_D6 = CLBLM_R_X3Y124_SLICE_X2Y124_AO6;
  assign CLBLM_R_X3Y122_SLICE_X2Y122_A1 = CLBLM_R_X3Y124_SLICE_X2Y124_AO5;
  assign CLBLM_R_X3Y122_SLICE_X2Y122_A2 = RIOB33_X105Y133_IOB_X1Y134_I;
  assign CLBLM_R_X3Y122_SLICE_X2Y122_A3 = RIOB33_X105Y133_IOB_X1Y133_I;
  assign CLBLM_R_X3Y122_SLICE_X2Y122_A4 = RIOB33_X105Y131_IOB_X1Y131_I;
  assign CLBLM_R_X3Y122_SLICE_X2Y122_A5 = RIOB33_X105Y131_IOB_X1Y132_I;
  assign CLBLM_R_X3Y122_SLICE_X2Y122_A6 = 1'b1;
  assign CLBLM_R_X3Y122_SLICE_X2Y122_B1 = RIOB33_X105Y131_IOB_X1Y131_I;
  assign CLBLM_R_X3Y122_SLICE_X2Y122_B2 = RIOB33_X105Y133_IOB_X1Y133_I;
  assign CLBLM_R_X3Y122_SLICE_X2Y122_B3 = CLBLM_R_X3Y122_SLICE_X3Y122_AO6;
  assign CLBLM_R_X3Y122_SLICE_X2Y122_B4 = RIOB33_X105Y131_IOB_X1Y132_I;
  assign CLBLM_R_X3Y122_SLICE_X2Y122_B5 = RIOB33_X105Y133_IOB_X1Y134_I;
  assign CLBLM_R_X3Y122_SLICE_X2Y122_B6 = 1'b1;
  assign LIOI3_X0Y183_OLOGIC_X0Y184_T1 = 1'b1;
  assign RIOB33_X105Y167_IOB_X1Y167_O = LIOB33_SING_X0Y50_IOB_X0Y50_I;
  assign CLBLM_R_X3Y122_SLICE_X2Y122_C1 = CLBLL_L_X2Y121_SLICE_X0Y121_BO6;
  assign CLBLM_R_X3Y122_SLICE_X2Y122_C2 = CLBLM_R_X3Y122_SLICE_X3Y122_AO6;
  assign CLBLM_R_X3Y122_SLICE_X2Y122_C3 = CLBLL_L_X4Y121_SLICE_X5Y121_BO6;
  assign CLBLM_R_X3Y122_SLICE_X2Y122_C4 = CLBLM_R_X3Y124_SLICE_X2Y124_AO5;
  assign CLBLM_R_X3Y122_SLICE_X2Y122_C5 = CLBLL_L_X4Y122_SLICE_X4Y122_AO6;
  assign CLBLM_R_X3Y122_SLICE_X2Y122_C6 = RIOB33_X105Y131_IOB_X1Y131_I;
  assign LIOB33_X0Y157_IOB_X0Y158_O = RIOB33_X105Y115_IOB_X1Y116_I;
  assign LIOB33_X0Y157_IOB_X0Y157_O = RIOB33_X105Y115_IOB_X1Y115_I;
  assign CLBLM_R_X3Y122_SLICE_X2Y122_D1 = CLBLL_L_X2Y121_SLICE_X0Y121_DO6;
  assign CLBLM_R_X3Y122_SLICE_X2Y122_D2 = CLBLL_L_X2Y122_SLICE_X1Y122_CO6;
  assign CLBLM_R_X3Y122_SLICE_X2Y122_D3 = CLBLM_R_X3Y122_SLICE_X3Y122_DO6;
  assign CLBLM_R_X3Y122_SLICE_X2Y122_D4 = CLBLM_R_X3Y122_SLICE_X2Y122_AO5;
  assign CLBLM_R_X3Y122_SLICE_X2Y122_D5 = CLBLM_R_X5Y122_SLICE_X6Y122_DO6;
  assign CLBLM_R_X3Y122_SLICE_X2Y122_D6 = LIOB33_X0Y57_IOB_X0Y58_I;
  assign CLBLM_R_X7Y120_SLICE_X9Y120_C4 = CLBLL_L_X4Y115_SLICE_X4Y115_CQ;
  assign CLBLM_R_X7Y120_SLICE_X9Y120_C5 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X7Y120_SLICE_X9Y120_C6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign RIOI3_X105Y159_OLOGIC_X1Y160_D1 = CLBLM_R_X11Y119_SLICE_X14Y119_CO6;
  assign CLBLM_R_X7Y120_SLICE_X9Y120_D2 = CLBLM_L_X10Y124_SLICE_X12Y124_AQ;
  assign RIOI3_X105Y159_OLOGIC_X1Y160_T1 = 1'b1;
  assign CLBLM_R_X7Y120_SLICE_X9Y120_D5 = CLBLM_L_X8Y119_SLICE_X10Y119_AQ;
  assign CLBLM_R_X7Y120_SLICE_X9Y120_D6 = 1'b1;
  assign CLBLM_L_X10Y117_SLICE_X12Y117_D1 = 1'b1;
  assign CLBLM_L_X8Y114_SLICE_X11Y114_A1 = CLBLM_L_X10Y113_SLICE_X12Y113_DO6;
  assign CLBLM_L_X8Y114_SLICE_X11Y114_A2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y114_SLICE_X11Y114_A3 = CLBLM_L_X8Y114_SLICE_X11Y114_AQ;
  assign CLBLM_L_X10Y117_SLICE_X12Y117_D2 = 1'b1;
  assign CLBLM_L_X8Y114_SLICE_X11Y114_A5 = CLBLM_L_X8Y118_SLICE_X10Y118_AQ;
  assign CLBLM_L_X8Y114_SLICE_X11Y114_A6 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign RIOI3_X105Y159_OLOGIC_X1Y159_D1 = CLBLM_R_X11Y113_SLICE_X15Y113_DO6;
  assign CLBLM_L_X8Y114_SLICE_X11Y114_B1 = CLBLM_R_X7Y115_SLICE_X8Y115_CQ;
  assign CLBLM_L_X8Y114_SLICE_X11Y114_B2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y114_SLICE_X11Y114_B4 = 1'b1;
  assign CLBLM_R_X5Y122_SLICE_X7Y122_C2 = CLBLM_R_X5Y122_SLICE_X7Y122_CQ;
  assign CLBLM_R_X5Y122_SLICE_X7Y122_C3 = CLBLM_R_X3Y116_SLICE_X2Y116_DO6;
  assign CLBLM_L_X8Y114_SLICE_X11Y114_B6 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X5Y122_SLICE_X7Y122_C4 = CLBLM_R_X5Y122_SLICE_X7Y122_A5Q;
  assign CLBLM_R_X5Y122_SLICE_X7Y122_C5 = CLBLM_L_X10Y122_SLICE_X12Y122_BQ;
  assign CLBLM_R_X5Y122_SLICE_X7Y122_C6 = 1'b1;
  assign RIOI3_X105Y159_OLOGIC_X1Y159_T1 = 1'b1;
  assign CLBLM_L_X8Y114_SLICE_X11Y114_C1 = CLBLM_L_X8Y110_SLICE_X10Y110_BQ;
  assign CLBLM_R_X7Y120_SLICE_X8Y120_B5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y114_SLICE_X11Y114_C2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y120_SLICE_X8Y120_B6 = CLBLM_L_X8Y117_SLICE_X10Y117_CQ;
  assign CLBLM_L_X8Y114_SLICE_X11Y114_C3 = 1'b1;
  assign CLBLM_L_X8Y114_SLICE_X11Y114_C4 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X8Y114_SLICE_X11Y114_C5 = 1'b1;
  assign CLBLM_R_X3Y123_SLICE_X3Y123_A1 = 1'b1;
  assign CLBLM_R_X3Y123_SLICE_X3Y123_A2 = CLBLM_R_X3Y117_SLICE_X3Y117_AQ;
  assign CLBLM_R_X3Y123_SLICE_X3Y123_A3 = CLBLM_R_X3Y123_SLICE_X3Y123_AQ;
  assign CLBLM_R_X3Y123_SLICE_X3Y123_A4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X3Y123_SLICE_X3Y123_A5 = CLBLM_R_X7Y124_SLICE_X8Y124_BQ;
  assign CLBLM_R_X3Y123_SLICE_X3Y123_A6 = CLBLM_R_X3Y116_SLICE_X2Y116_DO6;
  assign CLBLM_R_X3Y123_SLICE_X3Y123_B1 = RIOB33_X105Y131_IOB_X1Y131_I;
  assign CLBLM_R_X3Y123_SLICE_X3Y123_B2 = RIOB33_X105Y133_IOB_X1Y133_I;
  assign CLBLM_R_X3Y123_SLICE_X3Y123_B3 = CLBLM_R_X3Y124_SLICE_X2Y124_AO5;
  assign CLBLM_R_X3Y123_SLICE_X3Y123_B4 = RIOB33_X105Y133_IOB_X1Y134_I;
  assign CLBLM_R_X3Y123_SLICE_X3Y123_B5 = RIOB33_X105Y131_IOB_X1Y132_I;
  assign CLBLM_R_X3Y123_SLICE_X3Y123_B6 = 1'b1;
  assign CLBLM_R_X5Y122_SLICE_X7Y122_D2 = CLBLM_L_X10Y126_SLICE_X12Y126_AQ;
  assign CLBLM_R_X3Y123_SLICE_X3Y123_C1 = RIOB33_X105Y133_IOB_X1Y134_I;
  assign CLBLM_R_X3Y123_SLICE_X3Y123_C2 = CLBLM_R_X3Y124_SLICE_X2Y124_AO5;
  assign CLBLM_R_X3Y123_SLICE_X3Y123_C3 = CLBLM_R_X7Y120_SLICE_X8Y120_CQ;
  assign CLBLM_R_X3Y123_SLICE_X3Y123_C4 = RIOB33_X105Y133_IOB_X1Y133_I;
  assign CLBLM_R_X3Y123_SLICE_X3Y123_C5 = RIOB33_X105Y131_IOB_X1Y131_I;
  assign CLBLM_R_X3Y123_SLICE_X3Y123_C6 = RIOB33_X105Y131_IOB_X1Y132_I;
  assign CLBLM_R_X7Y120_SLICE_X8Y120_C4 = CLBLM_R_X3Y116_SLICE_X2Y116_CO6;
  assign CLBLM_R_X3Y123_SLICE_X3Y123_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X5Y122_SLICE_X7Y122_D5 = 1'b1;
  assign CLBLM_R_X7Y120_SLICE_X8Y120_C5 = 1'b1;
  assign CLBLM_R_X3Y123_SLICE_X3Y123_D1 = CLBLM_R_X3Y124_SLICE_X3Y124_AO6;
  assign CLBLM_R_X3Y123_SLICE_X3Y123_D2 = CLBLL_L_X4Y123_SLICE_X4Y123_DO6;
  assign CLBLM_R_X3Y123_SLICE_X3Y123_D3 = CLBLM_R_X3Y123_SLICE_X2Y123_DO6;
  assign CLBLM_R_X3Y123_SLICE_X3Y123_D4 = CLBLM_R_X3Y122_SLICE_X3Y122_CO6;
  assign CLBLM_R_X3Y123_SLICE_X3Y123_D5 = CLBLL_L_X2Y117_SLICE_X1Y117_BQ;
  assign CLBLM_R_X3Y123_SLICE_X3Y123_D6 = CLBLM_R_X3Y123_SLICE_X3Y123_BO6;
  assign CLBLM_R_X5Y122_SLICE_X7Y122_D6 = CLBLM_R_X7Y120_SLICE_X9Y120_D5Q;
  assign CLBLM_R_X7Y120_SLICE_X8Y120_C6 = CLBLM_R_X7Y120_SLICE_X9Y120_BQ;
  assign LIOB33_X0Y159_IOB_X0Y160_O = RIOB33_X105Y107_IOB_X1Y107_I;
  assign LIOB33_X0Y159_IOB_X0Y159_O = RIOB33_X105Y117_IOB_X1Y117_I;
  assign CLBLM_R_X3Y123_SLICE_X2Y123_A1 = RIOB33_X105Y115_IOB_X1Y115_I;
  assign CLBLM_R_X3Y123_SLICE_X2Y123_A2 = CLBLL_L_X2Y121_SLICE_X0Y121_BO6;
  assign CLBLM_R_X3Y123_SLICE_X2Y123_A3 = CLBLM_R_X7Y119_SLICE_X8Y119_C5Q;
  assign CLBLM_R_X3Y123_SLICE_X2Y123_A4 = RIOB33_X105Y129_IOB_X1Y129_I;
  assign CLBLM_R_X3Y123_SLICE_X2Y123_A5 = RIOB33_X105Y137_IOB_X1Y137_I;
  assign CLBLM_R_X3Y123_SLICE_X2Y123_A6 = CLBLM_R_X3Y124_SLICE_X2Y124_AO6;
  assign CLBLM_L_X8Y114_SLICE_X11Y114_D1 = CLBLM_L_X8Y115_SLICE_X11Y115_C5Q;
  assign LIOI3_X0Y183_OLOGIC_X0Y183_D1 = RIOB33_X105Y135_IOB_X1Y135_I;
  assign CLBLM_R_X3Y123_SLICE_X2Y123_B1 = CLBLL_L_X2Y117_SLICE_X0Y117_AQ;
  assign CLBLM_R_X3Y123_SLICE_X2Y123_B2 = CLBLM_R_X3Y123_SLICE_X3Y123_BO6;
  assign CLBLM_R_X3Y123_SLICE_X2Y123_B3 = CLBLL_L_X2Y122_SLICE_X1Y122_AO6;
  assign CLBLM_R_X3Y123_SLICE_X2Y123_B4 = CLBLM_R_X3Y123_SLICE_X3Y123_CO6;
  assign CLBLM_R_X3Y123_SLICE_X2Y123_B5 = CLBLM_R_X3Y123_SLICE_X2Y123_AO6;
  assign CLBLM_R_X3Y123_SLICE_X2Y123_B6 = CLBLM_R_X3Y123_SLICE_X2Y123_CO6;
  assign CLBLM_R_X3Y123_SLICE_X2Y123_C1 = RIOB33_X105Y131_IOB_X1Y132_I;
  assign CLBLM_R_X3Y123_SLICE_X2Y123_C2 = RIOB33_X105Y131_IOB_X1Y131_I;
  assign CLBLM_R_X3Y123_SLICE_X2Y123_C3 = CLBLM_R_X3Y124_SLICE_X2Y124_BO5;
  assign CLBLM_R_X3Y123_SLICE_X2Y123_C4 = CLBLM_R_X3Y124_SLICE_X2Y124_AO5;
  assign CLBLM_R_X3Y123_SLICE_X2Y123_C5 = LIOB33_X0Y55_IOB_X0Y55_I;
  assign CLBLM_R_X3Y123_SLICE_X2Y123_C6 = CLBLL_L_X4Y119_SLICE_X4Y119_DQ;
  assign CLBLM_R_X5Y122_SLICE_X6Y122_A2 = CLBLM_L_X8Y121_SLICE_X11Y121_AQ;
  assign CLBLM_R_X3Y123_SLICE_X2Y123_D1 = CLBLM_R_X3Y123_SLICE_X3Y123_AQ;
  assign CLBLM_R_X3Y123_SLICE_X2Y123_D2 = CLBLM_R_X3Y124_SLICE_X2Y124_AO5;
  assign CLBLM_R_X3Y123_SLICE_X2Y123_D3 = RIOB33_X105Y131_IOB_X1Y131_I;
  assign CLBLM_R_X3Y123_SLICE_X2Y123_D4 = LIOB33_X0Y57_IOB_X0Y57_I;
  assign CLBLM_R_X3Y123_SLICE_X2Y123_D5 = CLBLM_R_X3Y124_SLICE_X2Y124_BO5;
  assign CLBLM_R_X3Y123_SLICE_X2Y123_D6 = RIOB33_X105Y131_IOB_X1Y132_I;
  assign LIOI3_TBYTESRC_X0Y157_OLOGIC_X0Y158_D1 = RIOB33_X105Y115_IOB_X1Y116_I;
  assign CLBLM_L_X12Y118_SLICE_X17Y118_A1 = CLBLM_R_X11Y119_SLICE_X15Y119_AQ;
  assign CLBLM_L_X12Y118_SLICE_X17Y118_A2 = 1'b1;
  assign CLBLM_L_X12Y118_SLICE_X17Y118_A3 = CLBLM_R_X11Y119_SLICE_X15Y119_BQ;
  assign CLBLM_L_X12Y118_SLICE_X17Y118_A4 = CLBLM_L_X12Y118_SLICE_X16Y118_BQ;
  assign CLBLM_L_X12Y118_SLICE_X17Y118_A5 = CLBLM_R_X13Y119_SLICE_X18Y119_DO6;
  assign CLBLM_L_X12Y118_SLICE_X17Y118_A6 = CLBLM_L_X12Y120_SLICE_X17Y120_BQ;
  assign CLBLM_L_X12Y118_SLICE_X17Y118_B1 = 1'b1;
  assign CLBLM_L_X12Y118_SLICE_X17Y118_B2 = 1'b1;
  assign CLBLM_L_X12Y118_SLICE_X17Y118_B3 = 1'b1;
  assign CLBLM_L_X12Y118_SLICE_X17Y118_B4 = 1'b1;
  assign CLBLM_L_X12Y118_SLICE_X17Y118_B5 = 1'b1;
  assign CLBLM_L_X12Y118_SLICE_X17Y118_B6 = 1'b1;
  assign CLBLM_L_X12Y118_SLICE_X17Y118_C1 = 1'b1;
  assign CLBLM_L_X12Y118_SLICE_X17Y118_C2 = 1'b1;
  assign CLBLM_L_X12Y118_SLICE_X17Y118_C3 = 1'b1;
  assign CLBLM_L_X12Y118_SLICE_X17Y118_C4 = 1'b1;
  assign CLBLM_L_X12Y118_SLICE_X17Y118_C5 = 1'b1;
  assign CLBLM_L_X12Y118_SLICE_X17Y118_C6 = 1'b1;
  assign CLBLM_L_X12Y118_SLICE_X17Y118_D1 = 1'b1;
  assign CLBLM_L_X12Y118_SLICE_X17Y118_D2 = 1'b1;
  assign CLBLM_L_X12Y118_SLICE_X17Y118_D3 = 1'b1;
  assign CLBLM_L_X12Y118_SLICE_X17Y118_D4 = 1'b1;
  assign CLBLM_L_X12Y118_SLICE_X17Y118_D5 = 1'b1;
  assign CLBLM_L_X12Y118_SLICE_X17Y118_D6 = 1'b1;
  assign CLBLM_L_X12Y118_SLICE_X16Y118_A1 = CLBLM_R_X11Y120_SLICE_X14Y120_AO5;
  assign CLBLM_L_X12Y118_SLICE_X16Y118_A2 = CLBLM_R_X11Y118_SLICE_X14Y118_CQ;
  assign CLBLM_L_X12Y118_SLICE_X16Y118_A3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X12Y118_SLICE_X16Y118_A4 = CLBLM_L_X12Y120_SLICE_X17Y120_CO5;
  assign CLBLM_L_X12Y118_SLICE_X16Y118_A5 = 1'b1;
  assign CLBLM_L_X12Y118_SLICE_X16Y118_A6 = CLBLM_L_X12Y118_SLICE_X16Y118_CO6;
  assign CLBLM_L_X12Y118_SLICE_X16Y118_B1 = CLBLM_R_X11Y120_SLICE_X14Y120_AO5;
  assign CLBLM_L_X12Y118_SLICE_X16Y118_B2 = CLBLM_L_X12Y120_SLICE_X17Y120_CO5;
  assign CLBLM_L_X12Y118_SLICE_X16Y118_B3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X12Y118_SLICE_X16Y118_B4 = CLBLM_L_X12Y119_SLICE_X16Y119_BO6;
  assign CLBLM_L_X12Y118_SLICE_X16Y118_B5 = CLBLM_L_X12Y118_SLICE_X16Y118_BQ;
  assign CLBLM_L_X12Y118_SLICE_X16Y118_B6 = CLBLM_R_X7Y118_SLICE_X9Y118_CQ;
  assign CLBLM_R_X5Y122_SLICE_X6Y122_B6 = CLBLM_R_X5Y125_SLICE_X6Y125_A5Q;
  assign CLBLM_L_X12Y118_SLICE_X16Y118_C1 = CLBLM_R_X11Y118_SLICE_X14Y118_DO5;
  assign CLBLM_L_X12Y118_SLICE_X16Y118_C2 = CLBLM_L_X12Y118_SLICE_X16Y118_AQ;
  assign CLBLM_L_X12Y118_SLICE_X16Y118_C3 = CLBLM_R_X11Y118_SLICE_X15Y118_CQ;
  assign CLBLM_L_X12Y118_SLICE_X16Y118_C4 = CLBLM_L_X12Y119_SLICE_X17Y119_DO6;
  assign CLBLM_L_X12Y118_SLICE_X16Y118_C5 = CLBLM_L_X12Y119_SLICE_X16Y119_DO6;
  assign CLBLM_L_X12Y118_SLICE_X16Y118_C6 = CLBLM_L_X12Y118_SLICE_X17Y118_AO6;
  assign CLBLM_L_X12Y118_SLICE_X16Y118_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X12Y118_SLICE_X16Y118_D1 = 1'b1;
  assign CLBLM_L_X12Y118_SLICE_X16Y118_D2 = 1'b1;
  assign CLBLM_L_X12Y118_SLICE_X16Y118_D3 = 1'b1;
  assign CLBLM_L_X12Y118_SLICE_X16Y118_D4 = 1'b1;
  assign CLBLM_L_X12Y118_SLICE_X16Y118_D5 = 1'b1;
  assign CLBLM_L_X12Y118_SLICE_X16Y118_D6 = 1'b1;
  assign LIOI3_X0Y161_OLOGIC_X0Y162_D1 = RIOB33_X105Y109_IOB_X1Y109_I;
  assign CLBLM_L_X8Y114_SLICE_X10Y114_B5 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign LIOI3_X0Y161_OLOGIC_X0Y162_T1 = 1'b1;
  assign CLBLM_L_X8Y114_SLICE_X10Y114_B6 = 1'b1;
  assign LIOI3_X0Y101_OLOGIC_X0Y102_D1 = CLBLL_L_X2Y111_SLICE_X0Y111_AO5;
  assign CLBLM_R_X5Y122_SLICE_X6Y122_C4 = CLBLM_R_X13Y119_SLICE_X18Y119_BQ;
  assign CLBLM_R_X5Y122_SLICE_X6Y122_C5 = CLBLM_R_X7Y123_SLICE_X8Y123_CQ;
  assign LIOI3_X0Y161_OLOGIC_X0Y161_D1 = RIOB33_X105Y107_IOB_X1Y108_I;
  assign CLBLM_R_X5Y122_SLICE_X6Y122_C6 = CLBLM_R_X3Y124_SLICE_X2Y124_BO6;
  assign LIOI3_X0Y101_OLOGIC_X0Y102_T1 = 1'b1;
  assign LIOI3_X0Y161_OLOGIC_X0Y161_T1 = 1'b1;
  assign LIOI3_X0Y101_OLOGIC_X0Y101_D1 = CLBLL_L_X2Y111_SLICE_X0Y111_CO6;
  assign CLBLM_L_X8Y114_SLICE_X10Y114_C1 = RIOB33_X105Y103_IOB_X1Y103_I;
  assign CLBLM_L_X8Y114_SLICE_X10Y114_C2 = CLBLM_R_X5Y113_SLICE_X6Y113_BQ;
  assign LIOI3_X0Y101_OLOGIC_X0Y101_T1 = 1'b1;
  assign CLBLM_L_X8Y114_SLICE_X10Y114_C5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y117_SLICE_X10Y117_A1 = 1'b1;
  assign RIOB33_X105Y159_IOB_X1Y160_O = CLBLM_R_X11Y119_SLICE_X14Y119_CO6;
  assign RIOB33_X105Y159_IOB_X1Y159_O = CLBLM_R_X11Y113_SLICE_X15Y113_DO6;
  assign CLBLM_L_X8Y117_SLICE_X10Y117_A3 = CLBLM_L_X8Y117_SLICE_X10Y117_AQ;
  assign CLBLL_L_X4Y123_SLICE_X4Y123_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X3Y124_SLICE_X3Y124_A1 = RIOB33_X105Y115_IOB_X1Y116_I;
  assign CLBLM_R_X3Y124_SLICE_X3Y124_A2 = RIOB33_X105Y133_IOB_X1Y133_I;
  assign CLBLM_R_X3Y124_SLICE_X3Y124_A3 = CLBLM_R_X3Y124_SLICE_X2Y124_AO6;
  assign CLBLM_R_X3Y124_SLICE_X3Y124_A4 = RIOB33_X105Y133_IOB_X1Y134_I;
  assign CLBLM_R_X3Y124_SLICE_X3Y124_A5 = RIOB33_X105Y131_IOB_X1Y132_I;
  assign CLBLM_R_X3Y124_SLICE_X3Y124_A6 = RIOB33_X105Y131_IOB_X1Y131_I;
  assign CLBLM_R_X3Y124_SLICE_X3Y124_B1 = 1'b1;
  assign CLBLM_R_X3Y124_SLICE_X3Y124_B2 = 1'b1;
  assign CLBLM_R_X3Y124_SLICE_X3Y124_B3 = 1'b1;
  assign CLBLM_R_X3Y124_SLICE_X3Y124_B4 = 1'b1;
  assign CLBLM_R_X3Y124_SLICE_X3Y124_B5 = 1'b1;
  assign CLBLM_R_X3Y124_SLICE_X3Y124_B6 = 1'b1;
  assign LIOB33_X0Y161_IOB_X0Y161_O = RIOB33_X105Y107_IOB_X1Y108_I;
  assign LIOB33_X0Y161_IOB_X0Y162_O = RIOB33_X105Y109_IOB_X1Y109_I;
  assign CLBLM_R_X3Y124_SLICE_X3Y124_C1 = 1'b1;
  assign CLBLM_R_X3Y124_SLICE_X3Y124_C2 = 1'b1;
  assign CLBLM_R_X3Y124_SLICE_X3Y124_C3 = 1'b1;
  assign CLBLM_R_X3Y124_SLICE_X3Y124_C4 = 1'b1;
  assign CLBLM_R_X3Y124_SLICE_X3Y124_C5 = 1'b1;
  assign CLBLM_R_X3Y124_SLICE_X3Y124_C6 = 1'b1;
  assign CLBLM_L_X8Y117_SLICE_X10Y117_A5 = CLBLM_L_X8Y115_SLICE_X11Y115_AQ;
  assign CLBLM_R_X3Y124_SLICE_X3Y124_D1 = 1'b1;
  assign CLBLM_R_X3Y124_SLICE_X3Y124_D2 = 1'b1;
  assign CLBLM_R_X3Y124_SLICE_X3Y124_D3 = 1'b1;
  assign CLBLM_R_X3Y124_SLICE_X3Y124_D4 = 1'b1;
  assign CLBLM_R_X3Y124_SLICE_X3Y124_D5 = 1'b1;
  assign CLBLM_R_X3Y124_SLICE_X3Y124_D6 = 1'b1;
  assign CLBLM_R_X3Y124_SLICE_X2Y124_A1 = RIOB33_X105Y129_IOB_X1Y129_I;
  assign CLBLM_R_X3Y124_SLICE_X2Y124_A2 = RIOB33_X105Y137_IOB_X1Y137_I;
  assign CLBLM_R_X3Y124_SLICE_X2Y124_A3 = RIOB33_X105Y135_IOB_X1Y136_I;
  assign CLBLM_R_X3Y124_SLICE_X2Y124_A4 = RIOB33_X105Y135_IOB_X1Y135_I;
  assign CLBLM_R_X3Y124_SLICE_X2Y124_A5 = RIOB33_X105Y129_IOB_X1Y130_I;
  assign CLBLM_R_X3Y124_SLICE_X2Y124_A6 = 1'b1;
  assign CLBLM_L_X8Y117_SLICE_X10Y117_A6 = CLBLM_R_X5Y119_SLICE_X7Y119_AO6;
  assign CLBLM_R_X3Y124_SLICE_X2Y124_B1 = 1'b1;
  assign CLBLM_R_X3Y124_SLICE_X2Y124_B2 = RIOB33_X105Y133_IOB_X1Y133_I;
  assign CLBLM_R_X3Y124_SLICE_X2Y124_B3 = 1'b1;
  assign CLBLM_R_X3Y124_SLICE_X2Y124_B4 = RIOB33_X105Y133_IOB_X1Y134_I;
  assign CLBLM_R_X3Y124_SLICE_X2Y124_B5 = RIOB33_X105Y131_IOB_X1Y132_I;
  assign CLBLM_R_X3Y124_SLICE_X2Y124_B6 = 1'b1;
  assign CLBLL_L_X4Y120_SLICE_X4Y120_A4 = CLBLL_L_X2Y121_SLICE_X1Y121_CO6;
  assign CLBLM_R_X3Y124_SLICE_X2Y124_C1 = 1'b1;
  assign CLBLM_R_X3Y124_SLICE_X2Y124_C2 = 1'b1;
  assign CLBLM_R_X3Y124_SLICE_X2Y124_C3 = 1'b1;
  assign CLBLM_R_X3Y124_SLICE_X2Y124_C4 = 1'b1;
  assign CLBLM_R_X3Y124_SLICE_X2Y124_C5 = 1'b1;
  assign CLBLM_R_X3Y124_SLICE_X2Y124_C6 = 1'b1;
  assign LIOI3_TBYTESRC_X0Y157_OLOGIC_X0Y158_T1 = 1'b1;
  assign CLBLM_R_X3Y124_SLICE_X2Y124_D1 = 1'b1;
  assign CLBLM_R_X3Y124_SLICE_X2Y124_D2 = 1'b1;
  assign CLBLM_R_X3Y124_SLICE_X2Y124_D3 = 1'b1;
  assign CLBLM_R_X3Y124_SLICE_X2Y124_D4 = 1'b1;
  assign CLBLM_R_X3Y124_SLICE_X2Y124_D5 = 1'b1;
  assign CLBLM_R_X3Y124_SLICE_X2Y124_D6 = 1'b1;
  assign CLBLM_L_X12Y119_SLICE_X17Y119_A1 = CLBLM_R_X7Y120_SLICE_X9Y120_AQ;
  assign CLBLM_L_X12Y119_SLICE_X17Y119_A2 = CLBLM_R_X13Y119_SLICE_X18Y119_CQ;
  assign CLBLM_L_X12Y119_SLICE_X17Y119_A3 = CLBLM_L_X10Y116_SLICE_X12Y116_DO5;
  assign CLBLM_L_X12Y119_SLICE_X17Y119_A4 = CLBLM_R_X11Y119_SLICE_X15Y119_CQ;
  assign CLBLM_L_X12Y119_SLICE_X17Y119_A5 = CLBLM_L_X12Y120_SLICE_X16Y120_AO5;
  assign CLBLM_L_X12Y119_SLICE_X17Y119_A6 = 1'b1;
  assign CLBLL_L_X4Y120_SLICE_X4Y120_B1 = CLBLL_L_X4Y118_SLICE_X4Y118_DO6;
  assign CLBLM_L_X12Y119_SLICE_X17Y119_B1 = CLBLM_R_X13Y120_SLICE_X18Y120_CO6;
  assign CLBLM_L_X12Y119_SLICE_X17Y119_B2 = CLBLM_R_X11Y118_SLICE_X14Y118_DO5;
  assign CLBLM_L_X12Y119_SLICE_X17Y119_B3 = CLBLM_R_X13Y119_SLICE_X18Y119_DO6;
  assign CLBLM_L_X12Y119_SLICE_X17Y119_B4 = CLBLM_L_X12Y119_SLICE_X17Y119_DO6;
  assign CLBLM_L_X12Y119_SLICE_X17Y119_B5 = CLBLM_R_X11Y117_SLICE_X15Y117_AQ;
  assign CLBLM_L_X12Y119_SLICE_X17Y119_B6 = CLBLM_R_X11Y119_SLICE_X15Y119_AQ;
  assign CLBLL_L_X4Y120_SLICE_X4Y120_B2 = CLBLL_L_X2Y121_SLICE_X1Y121_CO6;
  assign RIOI3_X105Y145_ILOGIC_X1Y146_D = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLL_L_X4Y120_SLICE_X4Y120_B3 = CLBLM_R_X3Y123_SLICE_X3Y123_DO6;
  assign CLBLM_L_X12Y119_SLICE_X17Y119_C1 = CLBLM_L_X12Y118_SLICE_X16Y118_AQ;
  assign CLBLM_L_X12Y119_SLICE_X17Y119_C2 = CLBLM_R_X11Y119_SLICE_X15Y119_AQ;
  assign CLBLM_L_X12Y119_SLICE_X17Y119_C3 = CLBLM_L_X12Y118_SLICE_X16Y118_BQ;
  assign CLBLM_L_X12Y119_SLICE_X17Y119_C4 = CLBLM_R_X13Y119_SLICE_X18Y119_DO6;
  assign CLBLM_L_X12Y119_SLICE_X17Y119_C5 = CLBLM_L_X12Y120_SLICE_X17Y120_BQ;
  assign CLBLM_L_X12Y119_SLICE_X17Y119_C6 = CLBLM_R_X11Y119_SLICE_X15Y119_BQ;
  assign CLBLL_L_X4Y120_SLICE_X4Y120_B4 = CLBLL_L_X4Y120_SLICE_X4Y120_DO6;
  assign LIOI3_TBYTETERM_X0Y63_ILOGIC_X0Y64_D = LIOB33_X0Y63_IOB_X0Y64_I;
  assign CLBLL_L_X4Y120_SLICE_X4Y120_B5 = CLBLL_L_X4Y119_SLICE_X5Y119_BO6;
  assign LIOI3_TBYTETERM_X0Y63_ILOGIC_X0Y63_D = LIOB33_X0Y63_IOB_X0Y63_I;
  assign CLBLM_L_X12Y119_SLICE_X17Y119_D1 = CLBLM_L_X10Y116_SLICE_X12Y116_DO5;
  assign CLBLM_L_X12Y119_SLICE_X17Y119_D2 = CLBLM_L_X10Y119_SLICE_X13Y119_AQ;
  assign CLBLM_L_X12Y119_SLICE_X17Y119_D3 = CLBLM_R_X11Y118_SLICE_X14Y118_BQ;
  assign CLBLM_L_X12Y119_SLICE_X17Y119_D4 = CLBLM_R_X7Y120_SLICE_X9Y120_AQ;
  assign CLBLM_L_X12Y119_SLICE_X17Y119_D5 = CLBLM_R_X13Y119_SLICE_X18Y119_CQ;
  assign CLBLM_L_X12Y119_SLICE_X17Y119_D6 = CLBLM_R_X11Y119_SLICE_X15Y119_CQ;
  assign CLBLM_L_X12Y119_SLICE_X16Y119_A1 = CLBLM_R_X13Y120_SLICE_X18Y120_AO6;
  assign CLBLM_L_X12Y119_SLICE_X16Y119_A2 = CLBLM_L_X10Y117_SLICE_X12Y117_BQ;
  assign CLBLM_L_X12Y119_SLICE_X16Y119_A3 = CLBLM_L_X12Y119_SLICE_X17Y119_DO6;
  assign CLBLM_L_X12Y119_SLICE_X16Y119_A4 = CLBLM_R_X13Y120_SLICE_X18Y120_BO6;
  assign CLBLM_L_X12Y119_SLICE_X16Y119_A5 = CLBLM_R_X11Y119_SLICE_X15Y119_BQ;
  assign CLBLM_L_X12Y119_SLICE_X16Y119_A6 = CLBLM_R_X11Y118_SLICE_X14Y118_DO5;
  assign CLBLM_L_X12Y119_SLICE_X16Y119_B1 = CLBLM_R_X13Y120_SLICE_X18Y120_AO6;
  assign CLBLM_L_X12Y119_SLICE_X16Y119_B2 = CLBLM_R_X11Y118_SLICE_X14Y118_DO5;
  assign CLBLM_L_X12Y119_SLICE_X16Y119_B3 = CLBLM_L_X12Y119_SLICE_X17Y119_DO6;
  assign CLBLM_L_X12Y119_SLICE_X16Y119_B4 = CLBLM_R_X13Y120_SLICE_X18Y120_BO6;
  assign CLBLM_L_X12Y119_SLICE_X16Y119_B5 = CLBLM_R_X11Y119_SLICE_X15Y119_BQ;
  assign CLBLL_L_X4Y120_SLICE_X4Y120_C2 = CLBLL_L_X4Y117_SLICE_X4Y117_CO6;
  assign CLBLM_L_X12Y119_SLICE_X16Y119_B6 = CLBLM_L_X10Y118_SLICE_X13Y118_BQ;
  assign CLBLL_L_X4Y120_SLICE_X4Y120_C3 = CLBLL_L_X2Y122_SLICE_X0Y122_AO6;
  assign CLBLM_L_X12Y119_SLICE_X16Y119_C1 = CLBLM_L_X12Y118_SLICE_X16Y118_AQ;
  assign CLBLM_L_X12Y119_SLICE_X16Y119_C2 = CLBLM_R_X13Y120_SLICE_X18Y120_CO6;
  assign CLBLM_L_X12Y119_SLICE_X16Y119_C3 = CLBLM_L_X12Y120_SLICE_X17Y120_BQ;
  assign CLBLM_L_X12Y119_SLICE_X16Y119_C4 = CLBLM_R_X11Y119_SLICE_X15Y119_AQ;
  assign CLBLM_L_X12Y119_SLICE_X16Y119_C5 = CLBLM_R_X11Y119_SLICE_X15Y119_BQ;
  assign CLBLM_L_X12Y119_SLICE_X16Y119_C6 = CLBLM_L_X12Y118_SLICE_X16Y118_BQ;
  assign CLBLM_R_X7Y123_SLICE_X9Y123_C4 = CLBLM_L_X10Y118_SLICE_X12Y118_B5Q;
  assign CLBLL_L_X4Y120_SLICE_X4Y120_C5 = 1'b1;
  assign CLBLM_L_X12Y119_SLICE_X16Y119_D1 = CLBLM_R_X11Y119_SLICE_X15Y119_BQ;
  assign CLBLM_L_X12Y119_SLICE_X16Y119_D2 = CLBLM_L_X12Y120_SLICE_X17Y120_BQ;
  assign CLBLM_L_X12Y119_SLICE_X16Y119_D3 = CLBLM_R_X11Y119_SLICE_X15Y119_AQ;
  assign CLBLM_L_X12Y119_SLICE_X16Y119_D4 = CLBLM_R_X13Y120_SLICE_X18Y120_CO6;
  assign CLBLM_L_X12Y119_SLICE_X16Y119_D5 = 1'b1;
  assign CLBLM_L_X12Y119_SLICE_X16Y119_D6 = CLBLM_L_X12Y118_SLICE_X16Y118_BQ;
  assign CLBLL_L_X4Y123_SLICE_X4Y123_D2 = RIOB33_X105Y131_IOB_X1Y131_I;
  assign LIOI3_X0Y125_OLOGIC_X0Y125_T1 = 1'b1;
  assign CLBLM_R_X103Y138_SLICE_X163Y138_A1 = RIOB33_X105Y139_IOB_X1Y139_I;
  assign CLBLM_L_X8Y117_SLICE_X10Y117_B1 = CLBLM_R_X3Y118_SLICE_X2Y118_AQ;
  assign CLBLM_R_X103Y138_SLICE_X163Y138_A2 = 1'b1;
  assign CLBLM_R_X103Y138_SLICE_X163Y138_A3 = 1'b1;
  assign CLBLM_R_X103Y138_SLICE_X163Y138_A4 = RIOB33_X105Y137_IOB_X1Y138_I;
  assign CLBLM_R_X103Y138_SLICE_X163Y138_A5 = 1'b1;
  assign CLBLM_R_X103Y138_SLICE_X163Y138_A6 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X103Y138_SLICE_X163Y138_B1 = 1'b1;
  assign CLBLL_L_X4Y123_SLICE_X4Y123_D3 = CLBLM_R_X3Y124_SLICE_X2Y124_AO5;
  assign CLBLM_R_X103Y138_SLICE_X163Y138_B3 = 1'b1;
  assign CLBLM_R_X103Y138_SLICE_X163Y138_B4 = 1'b1;
  assign CLBLM_R_X103Y138_SLICE_X163Y138_B5 = 1'b1;
  assign CLBLM_R_X103Y138_SLICE_X163Y138_B6 = 1'b1;
  assign CLBLM_R_X103Y138_SLICE_X163Y138_B2 = 1'b1;
  assign CLBLM_R_X103Y138_SLICE_X163Y138_C1 = 1'b1;
  assign CLBLM_R_X103Y138_SLICE_X163Y138_C2 = 1'b1;
  assign CLBLM_R_X103Y138_SLICE_X163Y138_C3 = 1'b1;
  assign CLBLM_R_X103Y138_SLICE_X163Y138_C4 = 1'b1;
  assign CLBLM_R_X103Y138_SLICE_X163Y138_C5 = 1'b1;
  assign CLBLM_R_X103Y138_SLICE_X163Y138_C6 = 1'b1;
  assign CLBLM_L_X8Y117_SLICE_X10Y117_B2 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign RIOB33_X105Y171_IOB_X1Y172_O = CLBLM_R_X103Y172_SLICE_X163Y172_AO6;
  assign CLBLL_L_X4Y120_SLICE_X4Y120_D3 = CLBLM_R_X3Y120_SLICE_X3Y120_CO6;
  assign CLBLM_R_X103Y138_SLICE_X163Y138_D1 = 1'b1;
  assign CLBLL_L_X4Y123_SLICE_X4Y123_D4 = RIOB33_X105Y133_IOB_X1Y134_I;
  assign CLBLL_L_X4Y120_SLICE_X4Y120_D4 = CLBLM_R_X7Y120_SLICE_X8Y120_BQ;
  assign CLBLM_R_X103Y138_SLICE_X163Y138_D2 = 1'b1;
  assign CLBLM_R_X103Y138_SLICE_X163Y138_D3 = 1'b1;
  assign CLBLM_R_X103Y138_SLICE_X163Y138_D4 = 1'b1;
  assign CLBLM_R_X103Y138_SLICE_X163Y138_D5 = 1'b1;
  assign CLBLL_L_X4Y120_SLICE_X4Y120_D5 = 1'b1;
  assign CLBLM_R_X103Y138_SLICE_X163Y138_D6 = 1'b1;
  assign CLBLL_L_X4Y120_SLICE_X4Y120_D6 = CLBLM_R_X3Y122_SLICE_X2Y122_BO5;
  assign CLBLM_R_X103Y138_SLICE_X162Y138_A1 = 1'b1;
  assign CLBLM_R_X103Y138_SLICE_X162Y138_A2 = 1'b1;
  assign CLBLM_R_X103Y138_SLICE_X162Y138_A3 = 1'b1;
  assign CLBLM_L_X8Y117_SLICE_X10Y117_B3 = CLBLM_R_X3Y116_SLICE_X3Y116_AQ;
  assign CLBLM_R_X103Y138_SLICE_X162Y138_A4 = 1'b1;
  assign CLBLM_R_X103Y138_SLICE_X162Y138_A5 = 1'b1;
  assign CLBLM_R_X103Y138_SLICE_X162Y138_A6 = 1'b1;
  assign LIOI3_TBYTETERM_X0Y137_OLOGIC_X0Y138_D1 = CLBLM_R_X5Y125_SLICE_X6Y125_AQ;
  assign CLBLM_R_X103Y138_SLICE_X162Y138_B1 = 1'b1;
  assign CLBLM_R_X103Y138_SLICE_X162Y138_B2 = 1'b1;
  assign CLBLL_L_X4Y123_SLICE_X4Y123_D5 = CLBLM_R_X5Y122_SLICE_X6Y122_AQ;
  assign CLBLM_R_X103Y138_SLICE_X162Y138_B3 = 1'b1;
  assign CLBLM_R_X103Y138_SLICE_X162Y138_B4 = 1'b1;
  assign CLBLM_R_X103Y138_SLICE_X162Y138_B5 = 1'b1;
  assign CLBLM_R_X103Y138_SLICE_X162Y138_B6 = 1'b1;
  assign CLBLM_R_X7Y124_SLICE_X9Y124_D5 = 1'b1;
  assign CLBLM_R_X103Y138_SLICE_X162Y138_C1 = 1'b1;
  assign CLBLM_R_X103Y138_SLICE_X162Y138_C2 = 1'b1;
  assign CLBLM_R_X103Y138_SLICE_X162Y138_C3 = 1'b1;
  assign CLBLM_R_X103Y138_SLICE_X162Y138_C4 = 1'b1;
  assign CLBLM_R_X103Y138_SLICE_X162Y138_C5 = 1'b1;
  assign CLBLM_R_X103Y138_SLICE_X162Y138_C6 = 1'b1;
  assign CLBLM_L_X8Y117_SLICE_X10Y117_B4 = CLBLM_L_X8Y119_SLICE_X10Y119_BQ;
  assign CLBLL_L_X4Y123_SLICE_X4Y123_D6 = RIOB33_X105Y133_IOB_X1Y133_I;
  assign CLBLM_R_X103Y138_SLICE_X162Y138_D1 = 1'b1;
  assign CLBLM_R_X103Y138_SLICE_X162Y138_D2 = 1'b1;
  assign CLBLM_R_X103Y138_SLICE_X162Y138_D3 = 1'b1;
  assign CLBLM_R_X103Y138_SLICE_X162Y138_D4 = 1'b1;
  assign CLBLM_R_X103Y138_SLICE_X162Y138_D5 = 1'b1;
  assign CLBLM_R_X103Y138_SLICE_X162Y138_D6 = 1'b1;
  assign LIOB33_X0Y163_IOB_X0Y163_O = RIOB33_X105Y109_IOB_X1Y110_I;
  assign LIOB33_X0Y163_IOB_X0Y164_O = RIOB33_X105Y111_IOB_X1Y111_I;
  assign CLBLM_L_X8Y117_SLICE_X10Y117_B5 = CLBLM_L_X8Y117_SLICE_X10Y117_BQ;
  assign LIOI3_TBYTETERM_X0Y137_OLOGIC_X0Y138_T1 = 1'b1;
  assign CLBLM_L_X8Y117_SLICE_X10Y117_B6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X11Y121_SLICE_X14Y121_B4 = CLBLM_L_X10Y121_SLICE_X13Y121_AQ;
  assign CLBLM_R_X11Y121_SLICE_X14Y121_B5 = CLBLM_L_X10Y120_SLICE_X13Y120_AQ;
  assign LIOI3_TBYTETERM_X0Y137_OLOGIC_X0Y137_D1 = CLBLM_R_X5Y124_SLICE_X6Y124_BQ;
  assign CLBLM_R_X11Y121_SLICE_X14Y121_B6 = 1'b1;
  assign CLBLM_R_X7Y124_SLICE_X9Y124_D6 = 1'b1;
  assign CLBLM_L_X12Y120_SLICE_X17Y120_A1 = CLBLM_L_X12Y120_SLICE_X16Y120_CO6;
  assign CLBLM_L_X12Y120_SLICE_X17Y120_A2 = 1'b1;
  assign CLBLM_L_X12Y120_SLICE_X17Y120_A3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X12Y120_SLICE_X17Y120_A4 = CLBLM_R_X11Y120_SLICE_X14Y120_AO5;
  assign CLBLM_L_X12Y120_SLICE_X17Y120_A5 = CLBLM_L_X12Y120_SLICE_X17Y120_CO5;
  assign CLBLM_L_X12Y120_SLICE_X17Y120_A6 = CLBLM_R_X13Y119_SLICE_X18Y119_BQ;
  assign CLBLL_L_X4Y120_SLICE_X5Y120_A2 = CLBLL_L_X4Y120_SLICE_X4Y120_BO6;
  assign CLBLM_L_X12Y120_SLICE_X17Y120_B1 = CLBLM_L_X12Y119_SLICE_X17Y119_BO6;
  assign CLBLM_L_X12Y120_SLICE_X17Y120_B2 = CLBLM_L_X12Y120_SLICE_X17Y120_BQ;
  assign CLBLM_L_X12Y120_SLICE_X17Y120_B3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X12Y120_SLICE_X17Y120_B4 = CLBLM_R_X11Y120_SLICE_X14Y120_AO5;
  assign CLBLM_L_X12Y120_SLICE_X17Y120_B5 = CLBLM_L_X12Y120_SLICE_X17Y120_CO5;
  assign CLBLM_L_X12Y120_SLICE_X17Y120_B6 = CLBLM_R_X5Y120_SLICE_X6Y120_BQ;
  assign CLBLM_L_X10Y110_SLICE_X13Y110_A1 = CLBLM_R_X7Y120_SLICE_X9Y120_DQ;
  assign CLBLM_L_X10Y110_SLICE_X13Y110_A2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X12Y120_SLICE_X17Y120_C3 = CLBLM_R_X11Y119_SLICE_X15Y119_CQ;
  assign CLBLM_L_X12Y120_SLICE_X17Y120_C4 = CLBLM_R_X13Y119_SLICE_X18Y119_CQ;
  assign CLBLM_L_X12Y120_SLICE_X17Y120_C5 = CLBLM_L_X10Y119_SLICE_X13Y119_AQ;
  assign CLBLM_L_X12Y120_SLICE_X17Y120_C6 = 1'b1;
  assign CLBLM_L_X10Y110_SLICE_X13Y110_A3 = CLBLM_L_X10Y110_SLICE_X13Y110_AQ;
  assign CLBLM_L_X10Y110_SLICE_X13Y110_A4 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X10Y110_SLICE_X13Y110_A5 = CLBLM_L_X10Y112_SLICE_X12Y112_DQ;
  assign CLBLM_L_X10Y110_SLICE_X13Y110_A6 = CLBLM_L_X10Y110_SLICE_X13Y110_CO6;
  assign CLBLM_L_X10Y110_SLICE_X13Y110_B1 = CLBLM_L_X10Y110_SLICE_X13Y110_DO6;
  assign CLBLM_L_X10Y110_SLICE_X13Y110_B2 = CLBLM_L_X10Y110_SLICE_X13Y110_BQ;
  assign CLBLM_L_X10Y110_SLICE_X13Y110_B3 = CLBLM_L_X10Y116_SLICE_X13Y116_AQ;
  assign CLBLM_L_X10Y110_SLICE_X13Y110_B4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y110_SLICE_X13Y110_B5 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X12Y120_SLICE_X17Y120_D2 = 1'b1;
  assign CLBLM_L_X10Y110_SLICE_X13Y110_B6 = CLBLM_R_X7Y120_SLICE_X9Y120_DQ;
  assign CLBLM_L_X12Y120_SLICE_X17Y120_D1 = CLBLM_R_X11Y118_SLICE_X14Y118_BQ;
  assign CLBLM_L_X10Y110_SLICE_X13Y110_C1 = CLBLM_L_X10Y110_SLICE_X12Y110_AQ;
  assign CLBLM_L_X10Y110_SLICE_X13Y110_C2 = CLBLM_L_X10Y113_SLICE_X12Y113_DO6;
  assign CLBLM_L_X10Y110_SLICE_X13Y110_C3 = CLBLM_L_X10Y110_SLICE_X13Y110_BQ;
  assign CLBLM_L_X10Y110_SLICE_X13Y110_C4 = CLBLM_R_X11Y115_SLICE_X14Y115_AQ;
  assign CLBLM_L_X10Y110_SLICE_X13Y110_C5 = CLBLM_L_X10Y110_SLICE_X13Y110_AQ;
  assign CLBLM_L_X10Y110_SLICE_X13Y110_C6 = 1'b1;
  assign CLBLM_L_X12Y120_SLICE_X17Y120_D4 = CLBLM_R_X11Y119_SLICE_X15Y119_CQ;
  assign CLBLM_L_X10Y110_SLICE_X13Y110_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X12Y120_SLICE_X16Y120_A1 = CLBLM_L_X12Y119_SLICE_X16Y119_CO6;
  assign CLBLM_L_X12Y120_SLICE_X16Y120_A2 = CLBLM_R_X11Y118_SLICE_X14Y118_DO5;
  assign CLBLM_L_X12Y120_SLICE_X16Y120_A3 = CLBLM_L_X12Y119_SLICE_X17Y119_CO6;
  assign CLBLM_L_X12Y120_SLICE_X16Y120_A4 = 1'b1;
  assign CLBLM_L_X12Y121_SLICE_X17Y121_D5 = 1'b1;
  assign CLBLM_L_X10Y110_SLICE_X13Y110_D1 = CLBLM_L_X10Y110_SLICE_X12Y110_AQ;
  assign CLBLM_L_X10Y110_SLICE_X13Y110_D2 = CLBLM_R_X11Y115_SLICE_X14Y115_AQ;
  assign CLBLM_L_X10Y110_SLICE_X13Y110_D3 = CLBLM_L_X10Y110_SLICE_X13Y110_BQ;
  assign CLBLM_L_X12Y120_SLICE_X16Y120_B1 = CLBLM_R_X11Y118_SLICE_X14Y118_DO5;
  assign CLBLM_L_X12Y120_SLICE_X16Y120_B2 = CLBLM_L_X12Y120_SLICE_X17Y120_DO6;
  assign CLBLM_L_X12Y120_SLICE_X16Y120_B3 = CLBLM_R_X11Y118_SLICE_X15Y118_AQ;
  assign CLBLM_L_X12Y120_SLICE_X16Y120_B4 = CLBLM_L_X12Y120_SLICE_X17Y120_AQ;
  assign CLBLM_L_X12Y120_SLICE_X16Y120_B5 = CLBLM_R_X11Y117_SLICE_X14Y117_AQ;
  assign CLBLM_L_X12Y120_SLICE_X16Y120_B6 = CLBLM_L_X12Y119_SLICE_X17Y119_DO6;
  assign CLBLM_L_X10Y110_SLICE_X13Y110_D4 = CLBLM_L_X10Y110_SLICE_X13Y110_AQ;
  assign CLBLM_L_X10Y110_SLICE_X13Y110_D5 = CLBLM_L_X10Y113_SLICE_X12Y113_DO6;
  assign CLBLM_L_X10Y110_SLICE_X12Y110_A1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y110_SLICE_X12Y110_A2 = CLBLM_L_X10Y110_SLICE_X13Y110_DO5;
  assign CLBLM_L_X12Y120_SLICE_X16Y120_C1 = CLBLM_R_X11Y118_SLICE_X15Y118_AQ;
  assign CLBLM_L_X12Y120_SLICE_X16Y120_C2 = CLBLM_L_X12Y120_SLICE_X17Y120_AQ;
  assign CLBLM_L_X12Y120_SLICE_X16Y120_C3 = CLBLM_L_X12Y120_SLICE_X17Y120_DO6;
  assign CLBLM_L_X12Y120_SLICE_X16Y120_C4 = CLBLM_R_X11Y118_SLICE_X14Y118_DO5;
  assign CLBLM_L_X12Y120_SLICE_X16Y120_C5 = CLBLM_L_X12Y119_SLICE_X17Y119_DO6;
  assign CLBLM_L_X12Y120_SLICE_X16Y120_C6 = CLBLM_L_X10Y118_SLICE_X13Y118_AQ;
  assign CLBLM_L_X10Y110_SLICE_X12Y110_A3 = CLBLM_L_X10Y110_SLICE_X12Y110_AQ;
  assign CLBLM_L_X10Y110_SLICE_X12Y110_A4 = CLBLM_R_X7Y120_SLICE_X9Y120_DQ;
  assign CLBLM_L_X10Y110_SLICE_X12Y110_A5 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X10Y110_SLICE_X12Y110_A6 = CLBLM_R_X5Y114_SLICE_X7Y114_AQ;
  assign CLBLM_L_X10Y110_SLICE_X12Y110_B1 = CLBLM_R_X5Y111_SLICE_X7Y111_DO6;
  assign CLBLM_L_X10Y110_SLICE_X12Y110_B2 = CLBLM_L_X10Y110_SLICE_X12Y110_BQ;
  assign CLBLM_L_X10Y110_SLICE_X12Y110_B3 = CLBLM_L_X10Y110_SLICE_X12Y110_AQ;
  assign CLBLM_L_X10Y110_SLICE_X12Y110_B4 = CLBLM_L_X8Y116_SLICE_X11Y116_BQ;
  assign CLBLM_L_X12Y120_SLICE_X16Y120_D1 = CLBLM_L_X12Y121_SLICE_X16Y121_AQ;
  assign CLBLM_L_X12Y120_SLICE_X16Y120_D2 = CLBLM_L_X12Y119_SLICE_X16Y119_CO6;
  assign CLBLM_L_X12Y120_SLICE_X16Y120_D3 = CLBLM_R_X11Y118_SLICE_X14Y118_DO5;
  assign CLBLM_L_X12Y120_SLICE_X16Y120_D4 = CLBLM_L_X12Y119_SLICE_X17Y119_CO6;
  assign CLBLM_L_X12Y120_SLICE_X16Y120_D5 = CLBLM_L_X10Y120_SLICE_X12Y120_DQ;
  assign CLBLM_L_X12Y120_SLICE_X16Y120_D6 = CLBLM_L_X12Y119_SLICE_X17Y119_DO6;
  assign CLBLM_L_X10Y110_SLICE_X12Y110_C1 = 1'b1;
  assign CLBLM_L_X10Y110_SLICE_X12Y110_C2 = 1'b1;
  assign CLBLM_L_X10Y110_SLICE_X12Y110_C3 = 1'b1;
  assign CLBLM_L_X10Y110_SLICE_X12Y110_C4 = 1'b1;
  assign CLBLM_L_X10Y110_SLICE_X12Y110_C5 = 1'b1;
  assign CLBLM_L_X10Y110_SLICE_X12Y110_C6 = 1'b1;
  assign CLBLM_L_X10Y110_SLICE_X12Y110_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X12Y121_SLICE_X16Y121_A2 = 1'b1;
  assign CLBLL_L_X4Y120_SLICE_X5Y120_C1 = CLBLM_R_X5Y120_SLICE_X6Y120_BQ;
  assign CLBLM_L_X12Y121_SLICE_X16Y121_A3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign RIOI3_TBYTETERM_X105Y163_OLOGIC_X1Y164_D1 = CLBLM_R_X7Y119_SLICE_X9Y119_DO5;
  assign CLBLM_L_X10Y110_SLICE_X12Y110_D1 = 1'b1;
  assign CLBLM_L_X10Y110_SLICE_X12Y110_D2 = 1'b1;
  assign CLBLM_L_X10Y110_SLICE_X12Y110_D3 = 1'b1;
  assign CLBLM_L_X10Y110_SLICE_X12Y110_D4 = 1'b1;
  assign CLBLM_L_X10Y110_SLICE_X12Y110_D5 = 1'b1;
  assign CLBLM_L_X10Y110_SLICE_X12Y110_D6 = 1'b1;
  assign CLBLL_L_X4Y120_SLICE_X5Y120_C4 = CLBLM_R_X7Y117_SLICE_X9Y117_DQ;
  assign CLBLL_L_X4Y120_SLICE_X5Y120_C3 = CLBLL_L_X4Y121_SLICE_X4Y121_DO5;
  assign CLBLL_L_X4Y120_SLICE_X5Y120_C5 = CLBLL_L_X4Y121_SLICE_X5Y121_AQ;
  assign CLBLM_R_X11Y122_SLICE_X14Y122_C4 = 1'b1;
  assign CLBLM_R_X7Y123_SLICE_X9Y123_D5 = 1'b1;
  assign CLBLM_R_X11Y121_SLICE_X14Y121_C2 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign LIOB33_X0Y165_IOB_X0Y166_O = RIOB33_X105Y113_IOB_X1Y113_I;
  assign LIOB33_X0Y165_IOB_X0Y165_O = RIOB33_X105Y111_IOB_X1Y112_I;
  assign CLBLM_R_X7Y123_SLICE_X9Y123_D6 = CLBLM_R_X7Y123_SLICE_X9Y123_AQ;
  assign CLBLM_R_X11Y121_SLICE_X14Y121_C3 = CLBLM_R_X13Y119_SLICE_X18Y119_BQ;
  assign LIOI3_X0Y165_OLOGIC_X0Y166_D1 = RIOB33_X105Y113_IOB_X1Y113_I;
  assign CLBLM_R_X11Y121_SLICE_X14Y121_C4 = RIOB33_X105Y121_IOB_X1Y121_I;
  assign LIOI3_X0Y165_OLOGIC_X0Y166_T1 = 1'b1;
  assign LIOI3_X0Y103_OLOGIC_X0Y104_D1 = CLBLL_L_X2Y111_SLICE_X0Y111_CO5;
  assign LIOI3_X0Y165_OLOGIC_X0Y165_D1 = RIOB33_X105Y111_IOB_X1Y112_I;
  assign LIOI3_X0Y103_OLOGIC_X0Y104_T1 = 1'b1;
  assign CLBLM_R_X11Y121_SLICE_X14Y121_C5 = CLBLM_R_X7Y114_SLICE_X8Y114_BQ;
  assign LIOI3_X0Y165_OLOGIC_X0Y165_T1 = 1'b1;
  assign LIOI3_X0Y103_OLOGIC_X0Y103_D1 = CLBLL_L_X2Y113_SLICE_X0Y113_AO6;
  assign LIOI3_X0Y103_OLOGIC_X0Y103_T1 = 1'b1;
  assign CLBLM_R_X11Y121_SLICE_X14Y121_C6 = 1'b1;
  assign RIOI3_TBYTETERM_X105Y163_OLOGIC_X1Y163_T1 = 1'b1;
  assign CLBLM_L_X12Y121_SLICE_X17Y121_A1 = 1'b1;
  assign CLBLM_L_X12Y121_SLICE_X17Y121_A2 = 1'b1;
  assign CLBLM_L_X12Y121_SLICE_X17Y121_A3 = 1'b1;
  assign CLBLM_L_X12Y121_SLICE_X17Y121_A4 = 1'b1;
  assign CLBLM_L_X12Y121_SLICE_X17Y121_A5 = 1'b1;
  assign CLBLM_L_X12Y121_SLICE_X17Y121_A6 = 1'b1;
  assign CLBLM_L_X12Y121_SLICE_X17Y121_B1 = 1'b1;
  assign CLBLM_L_X12Y121_SLICE_X17Y121_B2 = 1'b1;
  assign CLBLM_L_X12Y121_SLICE_X17Y121_B3 = 1'b1;
  assign CLBLM_L_X12Y121_SLICE_X17Y121_B4 = 1'b1;
  assign CLBLM_L_X12Y121_SLICE_X17Y121_B5 = 1'b1;
  assign CLBLM_L_X12Y121_SLICE_X17Y121_B6 = 1'b1;
  assign CLBLM_L_X12Y121_SLICE_X17Y121_C1 = 1'b1;
  assign CLBLM_L_X12Y121_SLICE_X17Y121_C2 = 1'b1;
  assign CLBLM_L_X12Y121_SLICE_X17Y121_C3 = 1'b1;
  assign CLBLM_L_X12Y121_SLICE_X17Y121_C4 = 1'b1;
  assign CLBLM_L_X12Y121_SLICE_X17Y121_C5 = 1'b1;
  assign CLBLM_L_X12Y121_SLICE_X17Y121_C6 = 1'b1;
  assign CLBLM_L_X10Y111_SLICE_X13Y111_A1 = CLBLM_L_X10Y111_SLICE_X12Y111_CO6;
  assign CLBLM_L_X10Y111_SLICE_X13Y111_A2 = CLBLM_R_X7Y128_SLICE_X8Y128_AQ;
  assign CLBLM_L_X10Y111_SLICE_X13Y111_A3 = CLBLM_R_X7Y119_SLICE_X8Y119_D5Q;
  assign CLBLM_L_X10Y111_SLICE_X13Y111_A4 = 1'b1;
  assign CLBLM_L_X10Y111_SLICE_X13Y111_A5 = RIOB33_X105Y141_IOB_X1Y142_I;
  assign CLBLM_L_X10Y111_SLICE_X13Y111_A6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y111_SLICE_X13Y111_B1 = CLBLM_R_X5Y111_SLICE_X7Y111_DO6;
  assign CLBLM_L_X10Y111_SLICE_X13Y111_B2 = CLBLM_L_X10Y112_SLICE_X13Y112_CQ;
  assign CLBLM_L_X10Y111_SLICE_X13Y111_B3 = CLBLM_R_X7Y110_SLICE_X8Y110_CQ;
  assign CLBLM_L_X10Y111_SLICE_X13Y111_B4 = CLBLL_L_X4Y110_SLICE_X5Y110_AQ;
  assign CLBLM_L_X10Y111_SLICE_X13Y111_B5 = CLBLM_L_X8Y110_SLICE_X10Y110_BQ;
  assign CLBLM_L_X10Y111_SLICE_X13Y111_B6 = 1'b1;
  assign CLBLM_L_X12Y121_SLICE_X17Y121_D1 = 1'b1;
  assign CLBLM_L_X10Y111_SLICE_X13Y111_C1 = CLBLM_L_X10Y112_SLICE_X13Y112_CQ;
  assign CLBLM_L_X10Y111_SLICE_X13Y111_C2 = CLBLM_L_X10Y117_SLICE_X12Y117_AQ;
  assign CLBLM_L_X10Y111_SLICE_X13Y111_C3 = CLBLL_L_X4Y110_SLICE_X5Y110_AQ;
  assign CLBLM_L_X10Y111_SLICE_X13Y111_C4 = CLBLM_R_X7Y110_SLICE_X8Y110_CQ;
  assign CLBLM_L_X10Y111_SLICE_X13Y111_C5 = CLBLM_L_X8Y110_SLICE_X10Y110_BQ;
  assign CLBLM_L_X10Y111_SLICE_X13Y111_C6 = 1'b1;
  assign CLBLM_L_X10Y111_SLICE_X13Y111_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X12Y121_SLICE_X16Y121_A1 = CLBLM_L_X12Y120_SLICE_X16Y120_DO6;
  assign CLBLM_L_X12Y121_SLICE_X16Y121_A4 = CLBLM_R_X11Y119_SLICE_X15Y119_CQ;
  assign CLBLM_L_X12Y121_SLICE_X16Y121_A5 = CLBLM_L_X12Y120_SLICE_X17Y120_CO5;
  assign CLBLM_L_X12Y121_SLICE_X16Y121_A6 = CLBLM_R_X11Y120_SLICE_X14Y120_AO5;
  assign CLBLM_L_X10Y111_SLICE_X13Y111_D1 = 1'b1;
  assign CLBLM_L_X10Y111_SLICE_X13Y111_D2 = 1'b1;
  assign CLBLM_L_X10Y111_SLICE_X13Y111_D3 = 1'b1;
  assign CLBLM_L_X10Y111_SLICE_X13Y111_D4 = 1'b1;
  assign CLBLM_L_X10Y111_SLICE_X13Y111_D5 = 1'b1;
  assign CLBLM_L_X10Y111_SLICE_X13Y111_D6 = 1'b1;
  assign CLBLM_L_X12Y121_SLICE_X16Y121_B1 = 1'b1;
  assign CLBLM_L_X12Y121_SLICE_X16Y121_B2 = 1'b1;
  assign CLBLM_L_X12Y121_SLICE_X16Y121_B3 = 1'b1;
  assign CLBLM_L_X12Y121_SLICE_X16Y121_B4 = 1'b1;
  assign CLBLM_L_X12Y121_SLICE_X16Y121_B5 = 1'b1;
  assign CLBLM_L_X12Y121_SLICE_X16Y121_B6 = 1'b1;
  assign CLBLM_L_X10Y111_SLICE_X12Y111_A1 = CLBLM_L_X10Y112_SLICE_X13Y112_CQ;
  assign CLBLM_L_X12Y121_SLICE_X16Y121_C1 = 1'b1;
  assign CLBLM_L_X12Y121_SLICE_X16Y121_C2 = 1'b1;
  assign CLBLM_L_X12Y121_SLICE_X16Y121_C3 = 1'b1;
  assign CLBLM_L_X12Y121_SLICE_X16Y121_C4 = 1'b1;
  assign CLBLM_L_X12Y121_SLICE_X16Y121_C5 = 1'b1;
  assign CLBLM_L_X12Y121_SLICE_X16Y121_C6 = 1'b1;
  assign CLBLM_L_X10Y111_SLICE_X12Y111_A2 = CLBLM_R_X7Y110_SLICE_X8Y110_CQ;
  assign CLBLM_L_X10Y111_SLICE_X12Y111_A3 = CLBLM_L_X10Y115_SLICE_X12Y115_AQ;
  assign CLBLM_L_X10Y111_SLICE_X12Y111_A4 = CLBLL_L_X4Y110_SLICE_X5Y110_AQ;
  assign CLBLM_L_X12Y121_SLICE_X16Y121_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X10Y111_SLICE_X12Y111_A5 = CLBLM_L_X8Y110_SLICE_X10Y110_BQ;
  assign CLBLM_L_X10Y111_SLICE_X12Y111_A6 = 1'b1;
  assign CLBLM_L_X10Y111_SLICE_X12Y111_B1 = CLBLM_L_X10Y112_SLICE_X13Y112_CQ;
  assign CLBLM_L_X10Y111_SLICE_X12Y111_B2 = CLBLL_L_X4Y110_SLICE_X5Y110_AQ;
  assign CLBLM_L_X12Y121_SLICE_X16Y121_D1 = 1'b1;
  assign CLBLM_L_X12Y121_SLICE_X16Y121_D2 = 1'b1;
  assign CLBLM_L_X12Y121_SLICE_X16Y121_D3 = 1'b1;
  assign CLBLM_L_X12Y121_SLICE_X16Y121_D4 = 1'b1;
  assign CLBLM_L_X12Y121_SLICE_X16Y121_D5 = 1'b1;
  assign CLBLM_L_X12Y121_SLICE_X16Y121_D6 = 1'b1;
  assign CLBLM_L_X10Y111_SLICE_X12Y111_B6 = 1'b1;
  assign CLBLM_L_X10Y111_SLICE_X12Y111_C1 = CLBLM_L_X10Y111_SLICE_X13Y111_AQ;
  assign CLBLM_L_X10Y111_SLICE_X12Y111_C2 = CLBLM_R_X7Y115_SLICE_X9Y115_BQ;
  assign CLBLM_L_X10Y111_SLICE_X12Y111_C3 = CLBLM_R_X5Y111_SLICE_X7Y111_DO6;
  assign CLBLM_L_X10Y111_SLICE_X12Y111_C4 = CLBLM_L_X10Y111_SLICE_X12Y111_AO5;
  assign CLBLM_L_X10Y111_SLICE_X12Y111_C5 = CLBLM_L_X10Y111_SLICE_X12Y111_BO5;
  assign CLBLM_L_X10Y111_SLICE_X12Y111_C6 = CLBLM_L_X10Y117_SLICE_X12Y117_AQ;
  assign CLBLM_L_X10Y111_SLICE_X12Y111_D1 = CLBLM_L_X10Y112_SLICE_X12Y112_AO6;
  assign CLBLM_L_X10Y111_SLICE_X12Y111_D2 = CLBLM_L_X10Y122_SLICE_X13Y122_A5Q;
  assign CLBLM_L_X10Y111_SLICE_X12Y111_D3 = CLBLM_R_X5Y119_SLICE_X7Y119_CO6;
  assign CLBLM_L_X10Y111_SLICE_X12Y111_D4 = CLBLM_L_X10Y116_SLICE_X13Y116_CQ;
  assign CLBLM_L_X10Y111_SLICE_X12Y111_D5 = CLBLL_L_X2Y119_SLICE_X1Y119_BO6;
  assign CLBLM_L_X10Y111_SLICE_X12Y111_D6 = CLBLM_L_X10Y111_SLICE_X12Y111_BO6;
  assign RIOI3_X105Y147_ILOGIC_X1Y148_D = RIOB33_X105Y147_IOB_X1Y148_I;
  assign RIOI3_X105Y147_ILOGIC_X1Y147_D = RIOB33_X105Y147_IOB_X1Y147_I;
  assign RIOB33_X105Y171_IOB_X1Y171_O = CLBLM_L_X8Y128_SLICE_X10Y128_AO5;
  assign LIOB33_X0Y167_IOB_X0Y168_O = RIOB33_X105Y123_IOB_X1Y123_I;
  assign CLBLM_L_X10Y123_SLICE_X12Y123_D1 = CLBLM_L_X8Y123_SLICE_X10Y123_AQ;
  assign LIOB33_X0Y167_IOB_X0Y167_O = RIOB33_X105Y113_IOB_X1Y114_I;
  assign CLBLM_R_X11Y119_SLICE_X15Y119_C4 = CLBLM_R_X11Y119_SLICE_X14Y119_BO6;
  assign CLBLM_R_X11Y119_SLICE_X15Y119_C5 = CLBLM_L_X8Y120_SLICE_X11Y120_AQ;
  assign CLBLM_R_X11Y119_SLICE_X15Y119_C6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X11Y119_SLICE_X15Y119_D1 = CLBLM_R_X11Y118_SLICE_X14Y118_DO5;
  assign CLBLM_R_X11Y119_SLICE_X15Y119_D2 = CLBLM_R_X11Y120_SLICE_X14Y120_AO5;
  assign CLBLM_R_X11Y119_SLICE_X15Y119_D3 = CLBLM_R_X11Y119_SLICE_X14Y119_DO6;
  assign CLBLM_R_X11Y119_SLICE_X15Y119_D4 = CLBLM_L_X12Y119_SLICE_X17Y119_DO6;
  assign CLBLM_R_X7Y121_SLICE_X9Y121_C4 = CLBLM_L_X8Y118_SLICE_X10Y118_CQ;
  assign CLBLM_R_X7Y121_SLICE_X9Y121_C5 = CLBLM_L_X8Y120_SLICE_X10Y120_CQ;
  assign CLBLM_R_X7Y121_SLICE_X9Y121_C6 = 1'b1;
  assign CLBLM_L_X10Y112_SLICE_X13Y112_A1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y112_SLICE_X13Y112_A2 = CLBLM_R_X3Y118_SLICE_X2Y118_AQ;
  assign CLBLM_L_X10Y112_SLICE_X13Y112_A3 = CLBLM_L_X10Y112_SLICE_X13Y112_AQ;
  assign CLBLM_L_X10Y112_SLICE_X13Y112_A4 = CLBLM_R_X5Y114_SLICE_X6Y114_DQ;
  assign CLBLM_L_X10Y112_SLICE_X13Y112_A5 = CLBLM_R_X7Y112_SLICE_X8Y112_DO6;
  assign CLBLM_L_X10Y112_SLICE_X13Y112_A6 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_L_X10Y112_SLICE_X13Y112_B1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y112_SLICE_X13Y112_B2 = CLBLM_L_X10Y112_SLICE_X13Y112_BQ;
  assign CLBLM_L_X10Y112_SLICE_X13Y112_B3 = CLBLM_L_X10Y113_SLICE_X12Y113_DO6;
  assign CLBLM_L_X10Y112_SLICE_X13Y112_B4 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X10Y112_SLICE_X13Y112_B5 = CLBLM_R_X11Y113_SLICE_X14Y113_AQ;
  assign CLBLM_L_X10Y112_SLICE_X13Y112_B6 = CLBLM_L_X8Y118_SLICE_X10Y118_DQ;
  assign CLBLM_R_X11Y119_SLICE_X14Y119_B6 = 1'b1;
  assign CLBLM_L_X10Y112_SLICE_X13Y112_C1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y112_SLICE_X13Y112_C2 = CLBLM_L_X10Y111_SLICE_X13Y111_BO5;
  assign CLBLM_L_X10Y112_SLICE_X13Y112_C3 = CLBLM_L_X8Y118_SLICE_X10Y118_DQ;
  assign CLBLM_L_X10Y112_SLICE_X13Y112_C4 = CLBLM_L_X12Y120_SLICE_X17Y120_BQ;
  assign CLBLM_L_X10Y112_SLICE_X13Y112_C5 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X10Y112_SLICE_X13Y112_C6 = CLBLM_L_X10Y112_SLICE_X13Y112_CQ;
  assign CLBLM_L_X10Y112_SLICE_X13Y112_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X10Y112_SLICE_X13Y112_D1 = CLBLM_L_X8Y111_SLICE_X10Y111_AQ;
  assign CLBLM_L_X10Y112_SLICE_X13Y112_D2 = CLBLM_L_X8Y111_SLICE_X10Y111_DO6;
  assign CLBLM_L_X10Y112_SLICE_X13Y112_D3 = CLBLM_L_X10Y120_SLICE_X12Y120_BQ;
  assign CLBLM_L_X10Y112_SLICE_X13Y112_D4 = CLBLM_L_X10Y112_SLICE_X13Y112_BQ;
  assign CLBLM_L_X10Y112_SLICE_X13Y112_D5 = 1'b1;
  assign CLBLM_L_X10Y112_SLICE_X13Y112_D6 = CLBLM_L_X12Y115_SLICE_X16Y115_CQ;
  assign CLBLM_L_X10Y112_SLICE_X12Y112_A1 = CLBLL_L_X4Y110_SLICE_X5Y110_AQ;
  assign CLBLM_L_X10Y112_SLICE_X12Y112_A2 = CLBLM_R_X7Y110_SLICE_X8Y110_CQ;
  assign CLBLM_L_X10Y112_SLICE_X12Y112_A3 = CLBLM_L_X8Y110_SLICE_X10Y110_BQ;
  assign CLBLM_L_X10Y112_SLICE_X12Y112_A4 = CLBLM_R_X11Y117_SLICE_X14Y117_BQ;
  assign CLBLM_L_X10Y112_SLICE_X12Y112_A5 = CLBLM_L_X10Y112_SLICE_X13Y112_CQ;
  assign CLBLM_L_X10Y112_SLICE_X12Y112_A6 = 1'b1;
  assign CLBLM_R_X7Y121_SLICE_X9Y121_D2 = CLBLM_R_X7Y121_SLICE_X8Y121_BQ;
  assign CLBLM_L_X10Y112_SLICE_X12Y112_B1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y112_SLICE_X12Y112_B2 = CLBLM_R_X3Y118_SLICE_X2Y118_AQ;
  assign CLBLM_L_X10Y112_SLICE_X12Y112_B3 = CLBLM_R_X7Y112_SLICE_X8Y112_DO6;
  assign CLBLM_L_X10Y112_SLICE_X12Y112_B4 = CLBLM_R_X3Y112_SLICE_X3Y112_B5Q;
  assign CLBLM_L_X10Y112_SLICE_X12Y112_B5 = CLBLM_L_X10Y112_SLICE_X12Y112_BQ;
  assign CLBLM_L_X10Y112_SLICE_X12Y112_B6 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_R_X11Y119_SLICE_X14Y119_C4 = CLBLM_R_X11Y118_SLICE_X14Y118_CQ;
  assign CLBLM_R_X7Y121_SLICE_X9Y121_D5 = CLBLM_R_X7Y121_SLICE_X9Y121_AQ;
  assign CLBLM_R_X11Y119_SLICE_X14Y119_C5 = CLBLM_R_X3Y117_SLICE_X3Y117_BQ;
  assign CLBLM_L_X10Y112_SLICE_X12Y112_C1 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X10Y112_SLICE_X12Y112_C2 = CLBLM_L_X10Y112_SLICE_X12Y112_CQ;
  assign CLBLM_L_X10Y112_SLICE_X12Y112_C3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y112_SLICE_X12Y112_C4 = CLBLM_L_X10Y113_SLICE_X12Y113_DO6;
  assign CLBLM_L_X10Y112_SLICE_X12Y112_C5 = CLBLM_R_X11Y114_SLICE_X14Y114_AQ;
  assign CLBLM_L_X10Y112_SLICE_X12Y112_C6 = CLBLM_R_X5Y112_SLICE_X6Y112_AQ;
  assign CLBLM_R_X7Y121_SLICE_X9Y121_D6 = 1'b1;
  assign CLBLM_R_X11Y119_SLICE_X14Y119_C6 = 1'b1;
  assign CLBLM_L_X10Y112_SLICE_X12Y112_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X11Y119_SLICE_X14Y119_CE = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y112_SLICE_X12Y112_D1 = CLBLM_L_X10Y112_SLICE_X12Y112_BQ;
  assign CLBLM_L_X10Y112_SLICE_X12Y112_D2 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_L_X10Y112_SLICE_X12Y112_D3 = CLBLM_L_X10Y112_SLICE_X12Y112_DQ;
  assign CLBLM_L_X10Y112_SLICE_X12Y112_D4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y112_SLICE_X12Y112_D5 = CLBLM_R_X3Y118_SLICE_X2Y118_AQ;
  assign CLBLM_L_X10Y112_SLICE_X12Y112_D6 = CLBLM_L_X10Y113_SLICE_X12Y113_BQ;
  assign LIOB33_X0Y169_IOB_X0Y169_O = RIOB33_X105Y121_IOB_X1Y122_I;
  assign LIOB33_X0Y169_IOB_X0Y170_O = RIOB33_SING_X105Y149_IOB_X1Y149_I;
  assign CLBLM_L_X8Y115_SLICE_X11Y115_B1 = CLBLM_L_X10Y111_SLICE_X13Y111_AQ;
  assign CLBLM_L_X8Y115_SLICE_X11Y115_B2 = CLBLM_L_X8Y115_SLICE_X11Y115_BQ;
  assign CLBLM_R_X5Y123_SLICE_X7Y123_C1 = 1'b1;
  assign CLBLM_L_X8Y115_SLICE_X11Y115_B3 = CLBLM_R_X3Y118_SLICE_X2Y118_AQ;
  assign CLBLM_R_X11Y119_SLICE_X14Y119_D5 = CLBLM_L_X12Y120_SLICE_X17Y120_AQ;
  assign CLBLM_R_X5Y123_SLICE_X7Y123_C2 = 1'b1;
  assign CLBLM_L_X8Y115_SLICE_X11Y115_B4 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_R_X5Y123_SLICE_X7Y123_C3 = 1'b1;
  assign CLBLM_R_X5Y123_SLICE_X7Y123_C4 = 1'b1;
  assign CLBLM_R_X5Y123_SLICE_X7Y123_C5 = 1'b1;
  assign CLBLM_R_X5Y123_SLICE_X7Y123_C6 = 1'b1;
  assign LIOI3_X0Y109_OLOGIC_X0Y109_D1 = CLBLL_L_X2Y110_SLICE_X0Y110_AO6;
  assign CLBLM_R_X7Y121_SLICE_X8Y121_B5 = CLBLM_R_X5Y117_SLICE_X7Y117_AQ;
  assign CLBLM_R_X7Y121_SLICE_X8Y121_B6 = CLBLM_L_X8Y120_SLICE_X10Y120_CQ;
  assign CLBLM_L_X8Y115_SLICE_X11Y115_C4 = CLBLM_L_X8Y119_SLICE_X10Y119_A5Q;
  assign CLBLM_L_X8Y115_SLICE_X11Y115_C5 = CLBLM_L_X8Y113_SLICE_X11Y113_AQ;
  assign CLBLM_R_X5Y123_SLICE_X7Y123_D1 = 1'b1;
  assign CLBLM_R_X5Y123_SLICE_X7Y123_D2 = 1'b1;
  assign CLBLM_R_X7Y121_SLICE_X8Y121_C4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X5Y123_SLICE_X7Y123_D5 = 1'b1;
  assign CLBLM_R_X7Y121_SLICE_X8Y121_C5 = CLBLM_R_X7Y122_SLICE_X9Y122_A5Q;
  assign CLBLM_R_X5Y123_SLICE_X7Y123_D6 = 1'b1;
  assign CLBLM_R_X7Y121_SLICE_X8Y121_C6 = 1'b1;
  assign LIOI3_X0Y109_OLOGIC_X0Y109_T1 = 1'b1;
  assign LIOI3_X0Y167_OLOGIC_X0Y168_D1 = RIOB33_X105Y123_IOB_X1Y123_I;
  assign CLBLM_R_X5Y123_SLICE_X6Y123_A5 = CLBLL_L_X4Y123_SLICE_X4Y123_BQ;
  assign LIOI3_X0Y167_OLOGIC_X0Y168_T1 = 1'b1;
  assign LIOI3_X0Y105_OLOGIC_X0Y106_D1 = CLBLL_L_X2Y111_SLICE_X0Y111_DO5;
  assign CLBLM_L_X10Y113_SLICE_X13Y113_A1 = CLBLM_R_X7Y111_SLICE_X9Y111_DO6;
  assign CLBLM_L_X10Y113_SLICE_X13Y113_A2 = CLBLM_L_X10Y114_SLICE_X13Y114_AQ;
  assign CLBLM_L_X10Y113_SLICE_X13Y113_A3 = CLBLM_L_X8Y114_SLICE_X11Y114_AQ;
  assign CLBLM_L_X10Y113_SLICE_X13Y113_A4 = CLBLM_L_X10Y110_SLICE_X13Y110_CO5;
  assign CLBLM_L_X10Y113_SLICE_X13Y113_A5 = CLBLM_L_X10Y113_SLICE_X13Y113_CO6;
  assign CLBLM_L_X10Y113_SLICE_X13Y113_A6 = 1'b1;
  assign LIOI3_X0Y167_OLOGIC_X0Y167_D1 = RIOB33_X105Y113_IOB_X1Y114_I;
  assign CLBLM_R_X7Y121_SLICE_X8Y121_D5 = CLBLM_R_X7Y121_SLICE_X8Y121_AQ;
  assign CLBLM_L_X10Y113_SLICE_X13Y113_B1 = CLBLM_L_X10Y112_SLICE_X13Y112_DO6;
  assign CLBLM_L_X10Y113_SLICE_X13Y113_B2 = CLBLM_R_X7Y111_SLICE_X9Y111_DO6;
  assign CLBLM_L_X10Y113_SLICE_X13Y113_B3 = CLBLM_L_X10Y110_SLICE_X13Y110_CO5;
  assign CLBLM_L_X10Y113_SLICE_X13Y113_B4 = CLBLM_L_X10Y113_SLICE_X12Y113_DO6;
  assign CLBLM_L_X10Y113_SLICE_X13Y113_B5 = CLBLM_L_X8Y113_SLICE_X10Y113_AO6;
  assign CLBLM_L_X10Y113_SLICE_X13Y113_B6 = CLBLM_L_X10Y113_SLICE_X13Y113_AO5;
  assign LIOI3_X0Y105_OLOGIC_X0Y106_T1 = 1'b1;
  assign RIOI3_X105Y151_OLOGIC_X1Y152_D1 = RIOB33_SING_X105Y100_IOB_X1Y100_I;
  assign LIOI3_X0Y167_OLOGIC_X0Y167_T1 = 1'b1;
  assign CLBLM_L_X10Y113_SLICE_X13Y113_C1 = CLBLM_L_X8Y114_SLICE_X11Y114_AQ;
  assign CLBLM_L_X10Y113_SLICE_X13Y113_C2 = CLBLM_L_X8Y113_SLICE_X11Y113_AQ;
  assign CLBLM_L_X10Y113_SLICE_X13Y113_C3 = CLBLM_R_X11Y113_SLICE_X15Y113_AQ;
  assign CLBLM_L_X10Y113_SLICE_X13Y113_C4 = CLBLM_R_X11Y113_SLICE_X14Y113_DO6;
  assign CLBLM_L_X10Y113_SLICE_X13Y113_C5 = CLBLM_L_X10Y113_SLICE_X13Y113_DO6;
  assign CLBLM_L_X10Y113_SLICE_X13Y113_C6 = CLBLM_L_X8Y112_SLICE_X10Y112_BQ;
  assign LIOI3_X0Y105_OLOGIC_X0Y105_D1 = CLBLL_L_X2Y111_SLICE_X0Y111_DO6;
  assign RIOI3_X105Y151_OLOGIC_X1Y152_T1 = 1'b1;
  assign LIOI3_TBYTETERM_X0Y113_OLOGIC_X0Y114_D1 = CLBLM_R_X5Y117_SLICE_X6Y117_DQ;
  assign CLBLM_L_X10Y113_SLICE_X13Y113_D1 = CLBLM_R_X11Y113_SLICE_X14Y113_AQ;
  assign CLBLM_L_X10Y113_SLICE_X13Y113_D2 = CLBLM_R_X11Y113_SLICE_X15Y113_BQ;
  assign CLBLM_L_X10Y113_SLICE_X13Y113_D3 = CLBLM_R_X11Y114_SLICE_X14Y114_AQ;
  assign CLBLM_L_X10Y113_SLICE_X13Y113_D4 = CLBLM_L_X8Y112_SLICE_X10Y112_AQ;
  assign CLBLM_L_X10Y113_SLICE_X13Y113_D5 = CLBLM_R_X11Y114_SLICE_X14Y114_BQ;
  assign CLBLM_L_X10Y113_SLICE_X13Y113_D6 = CLBLM_L_X10Y112_SLICE_X12Y112_CQ;
  assign CLBLM_R_X5Y123_SLICE_X6Y123_B3 = CLBLM_R_X7Y122_SLICE_X9Y122_BO6;
  assign LIOI3_X0Y105_OLOGIC_X0Y105_T1 = 1'b1;
  assign CLBLM_R_X5Y123_SLICE_X6Y123_B4 = CLBLL_L_X4Y115_SLICE_X5Y115_BQ;
  assign LIOI3_TBYTETERM_X0Y113_OLOGIC_X0Y114_T1 = 1'b1;
  assign RIOI3_X105Y151_OLOGIC_X1Y151_D1 = LIOB33_X0Y75_IOB_X0Y76_I;
  assign RIOI3_TBYTETERM_X105Y187_OLOGIC_X1Y188_T1 = 1'b1;
  assign CLBLM_L_X10Y113_SLICE_X12Y113_A1 = CLBLM_L_X10Y112_SLICE_X13Y112_CQ;
  assign CLBLM_L_X10Y113_SLICE_X12Y113_A2 = CLBLM_R_X7Y110_SLICE_X8Y110_CQ;
  assign CLBLM_L_X10Y113_SLICE_X12Y113_A3 = CLBLM_L_X8Y110_SLICE_X10Y110_BQ;
  assign CLBLM_L_X10Y113_SLICE_X12Y113_A4 = CLBLL_L_X4Y110_SLICE_X5Y110_AQ;
  assign CLBLM_L_X10Y113_SLICE_X12Y113_A5 = CLBLM_R_X7Y112_SLICE_X9Y112_CQ;
  assign CLBLM_L_X10Y113_SLICE_X12Y113_A6 = 1'b1;
  assign CLBLM_R_X5Y123_SLICE_X6Y123_B5 = CLBLM_R_X5Y123_SLICE_X7Y123_AQ;
  assign CLBLM_R_X5Y123_SLICE_X6Y123_B6 = CLBLM_R_X5Y123_SLICE_X6Y123_BQ;
  assign LIOI3_TBYTETERM_X0Y113_OLOGIC_X0Y113_D1 = RIOB33_X105Y121_IOB_X1Y121_I;
  assign RIOI3_X105Y151_OLOGIC_X1Y151_T1 = 1'b1;
  assign CLBLM_L_X10Y113_SLICE_X12Y113_B1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y113_SLICE_X12Y113_B2 = CLBLM_L_X10Y113_SLICE_X12Y113_BQ;
  assign CLBLM_L_X10Y113_SLICE_X12Y113_B3 = CLBLM_L_X10Y114_SLICE_X13Y114_DQ;
  assign CLBLM_L_X10Y113_SLICE_X12Y113_B4 = CLBLM_R_X11Y123_SLICE_X14Y123_CO6;
  assign CLBLM_L_X10Y113_SLICE_X12Y113_B5 = CLBLM_L_X8Y111_SLICE_X11Y111_AO6;
  assign CLBLM_L_X10Y113_SLICE_X12Y113_B6 = CLBLM_L_X10Y113_SLICE_X12Y113_CO6;
  assign LIOB33_X0Y171_IOB_X0Y171_O = LIOB33_SING_X0Y50_IOB_X0Y50_I;
  assign LIOB33_X0Y171_IOB_X0Y172_O = CLBLM_R_X103Y138_SLICE_X163Y138_AO6;
  assign LIOI3_TBYTETERM_X0Y113_OLOGIC_X0Y113_T1 = 1'b1;
  assign CLBLM_L_X10Y113_SLICE_X12Y113_C1 = CLBLM_L_X10Y114_SLICE_X13Y114_DQ;
  assign CLBLM_L_X10Y113_SLICE_X12Y113_C2 = CLBLM_L_X8Y110_SLICE_X10Y110_BQ;
  assign CLBLM_L_X10Y113_SLICE_X12Y113_C3 = CLBLM_R_X5Y111_SLICE_X7Y111_DO6;
  assign CLBLM_L_X10Y113_SLICE_X12Y113_C4 = CLBLL_L_X4Y110_SLICE_X5Y110_AQ;
  assign CLBLM_L_X10Y113_SLICE_X12Y113_C5 = CLBLM_L_X10Y116_SLICE_X13Y116_AO5;
  assign CLBLM_L_X10Y113_SLICE_X12Y113_C6 = CLBLM_L_X10Y111_SLICE_X12Y111_AO5;
  assign CLBLM_L_X10Y113_SLICE_X12Y113_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X10Y113_SLICE_X12Y113_D1 = 1'b1;
  assign CLBLM_L_X10Y113_SLICE_X12Y113_D2 = 1'b1;
  assign CLBLM_L_X10Y113_SLICE_X12Y113_D3 = CLBLL_L_X2Y113_SLICE_X1Y113_AQ;
  assign CLBLM_L_X10Y113_SLICE_X12Y113_D4 = CLBLM_R_X3Y118_SLICE_X2Y118_AQ;
  assign CLBLM_L_X10Y113_SLICE_X12Y113_D5 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_L_X10Y113_SLICE_X12Y113_D6 = CLBLM_R_X5Y110_SLICE_X7Y110_BQ;
  assign CLBLM_R_X5Y123_SLICE_X6Y123_C2 = CLBLM_R_X5Y123_SLICE_X6Y123_CQ;
  assign CLBLM_R_X5Y123_SLICE_X6Y123_C3 = CLBLM_R_X3Y115_SLICE_X2Y115_BQ;
  assign CLBLM_R_X5Y123_SLICE_X6Y123_C4 = 1'b1;
  assign CLBLM_R_X103Y169_SLICE_X162Y169_D3 = 1'b1;
  assign CLBLM_R_X7Y111_SLICE_X9Y111_A3 = CLBLL_L_X2Y120_SLICE_X1Y120_DO6;
  assign CLBLM_R_X5Y123_SLICE_X6Y123_C5 = CLBLM_R_X7Y122_SLICE_X9Y122_BO6;
  assign LIOI3_X0Y185_OLOGIC_X0Y185_D1 = RIOB33_X105Y137_IOB_X1Y137_I;
  assign CLBLM_R_X7Y111_SLICE_X9Y111_A4 = CLBLM_R_X5Y117_SLICE_X7Y117_DO6;
  assign CLBLM_R_X5Y123_SLICE_X6Y123_C6 = CLBLM_R_X5Y123_SLICE_X6Y123_DO5;
  assign CLBLM_L_X8Y115_SLICE_X10Y115_C2 = CLBLM_R_X7Y116_SLICE_X9Y116_AQ;
  assign CLBLM_L_X8Y115_SLICE_X10Y115_C3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y115_SLICE_X10Y115_C4 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X7Y111_SLICE_X9Y111_B3 = CLBLM_L_X10Y112_SLICE_X13Y112_CQ;
  assign CLBLM_R_X7Y111_SLICE_X9Y111_B4 = CLBLM_L_X8Y110_SLICE_X10Y110_BQ;
  assign CLBLM_R_X7Y111_SLICE_X9Y111_B5 = CLBLM_R_X7Y110_SLICE_X8Y110_CQ;
  assign CLBLM_R_X7Y111_SLICE_X9Y111_B6 = 1'b1;
  assign CLBLM_L_X8Y115_SLICE_X10Y115_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X5Y123_SLICE_X6Y123_D5 = RIOB33_X105Y127_IOB_X1Y127_I;
  assign CLBLM_R_X7Y111_SLICE_X9Y111_C5 = CLBLM_R_X5Y111_SLICE_X7Y111_DO6;
  assign CLBLM_R_X103Y169_SLICE_X162Y169_D4 = 1'b1;
  assign CLBLL_L_X4Y123_SLICE_X5Y123_C4 = 1'b1;
  assign CLBLL_L_X4Y123_SLICE_X5Y123_C6 = 1'b1;
  assign CLBLM_L_X10Y114_SLICE_X13Y114_A1 = CLBLM_L_X10Y113_SLICE_X12Y113_DO6;
  assign CLBLM_L_X10Y114_SLICE_X13Y114_A2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y114_SLICE_X13Y114_A3 = CLBLM_L_X10Y114_SLICE_X13Y114_AQ;
  assign CLBLM_L_X10Y114_SLICE_X13Y114_A4 = CLBLM_R_X7Y112_SLICE_X8Y112_BQ;
  assign CLBLM_L_X10Y114_SLICE_X13Y114_A5 = CLBLM_L_X8Y114_SLICE_X11Y114_AQ;
  assign CLBLM_L_X10Y114_SLICE_X13Y114_A6 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X10Y114_SLICE_X13Y114_AX = CLBLM_L_X10Y114_SLICE_X13Y114_BO6;
  assign CLBLM_L_X10Y114_SLICE_X13Y114_B1 = CLBLL_L_X4Y114_SLICE_X5Y114_AQ;
  assign CLBLM_L_X10Y114_SLICE_X13Y114_B2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y114_SLICE_X13Y114_B3 = CLBLM_L_X10Y112_SLICE_X13Y112_AQ;
  assign CLBLM_L_X10Y114_SLICE_X13Y114_B4 = RIOB33_X105Y121_IOB_X1Y121_I;
  assign CLBLM_L_X10Y114_SLICE_X13Y114_B5 = CLBLM_R_X11Y116_SLICE_X14Y116_DQ;
  assign CLBLM_L_X10Y114_SLICE_X13Y114_B6 = 1'b1;
  assign CLBLM_L_X10Y114_SLICE_X13Y114_C1 = CLBLM_R_X3Y113_SLICE_X3Y113_AQ;
  assign CLBLM_L_X10Y114_SLICE_X13Y114_C2 = CLBLM_L_X10Y114_SLICE_X12Y114_CO6;
  assign CLBLM_L_X10Y114_SLICE_X13Y114_C3 = 1'b1;
  assign CLBLM_L_X10Y114_SLICE_X13Y114_C4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y114_SLICE_X13Y114_C5 = CLBLM_R_X7Y128_SLICE_X8Y128_AQ;
  assign CLBLM_L_X10Y114_SLICE_X13Y114_C6 = RIOB33_X105Y141_IOB_X1Y142_I;
  assign CLBLM_L_X10Y114_SLICE_X13Y114_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign LIOB33_X0Y173_IOB_X0Y174_O = CLBLM_R_X7Y151_SLICE_X8Y151_AO6;
  assign LIOB33_X0Y173_IOB_X0Y173_O = CLBLM_L_X8Y133_SLICE_X11Y133_AO5;
  assign RIOI3_TBYTETERM_X105Y187_OLOGIC_X1Y187_D1 = CLBLM_L_X10Y114_SLICE_X12Y114_AQ;
  assign CLBLM_L_X10Y114_SLICE_X13Y114_D1 = CLBLM_R_X7Y110_SLICE_X8Y110_CQ;
  assign CLBLM_L_X10Y114_SLICE_X13Y114_D2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y114_SLICE_X13Y114_D3 = CLBLM_R_X11Y120_SLICE_X15Y120_CQ;
  assign CLBLM_L_X10Y114_SLICE_X13Y114_D4 = CLBLM_L_X10Y114_SLICE_X13Y114_A5Q;
  assign CLBLM_L_X10Y114_SLICE_X13Y114_D5 = CLBLM_L_X10Y113_SLICE_X12Y113_BQ;
  assign CLBLM_L_X10Y114_SLICE_X13Y114_D6 = 1'b1;
  assign CLBLM_L_X10Y114_SLICE_X12Y114_A1 = CLBLM_L_X8Y110_SLICE_X10Y110_AQ;
  assign CLBLM_L_X10Y114_SLICE_X12Y114_A2 = CLBLM_R_X7Y110_SLICE_X8Y110_CQ;
  assign CLBLM_L_X10Y114_SLICE_X12Y114_A3 = CLBLL_L_X4Y110_SLICE_X5Y110_AQ;
  assign CLBLM_L_X10Y114_SLICE_X12Y114_A4 = CLBLM_L_X10Y112_SLICE_X13Y112_CQ;
  assign CLBLM_L_X10Y114_SLICE_X12Y114_A5 = CLBLM_L_X8Y110_SLICE_X10Y110_BQ;
  assign CLBLM_L_X10Y114_SLICE_X12Y114_A6 = 1'b1;
  assign LIOI3_X0Y171_OLOGIC_X0Y171_T1 = 1'b1;
  assign CLBLM_L_X10Y114_SLICE_X12Y114_AX = CLBLM_R_X11Y114_SLICE_X14Y114_DQ;
  assign CLBLM_L_X10Y114_SLICE_X12Y114_B1 = CLBLM_L_X8Y114_SLICE_X10Y114_DQ;
  assign CLBLM_L_X10Y114_SLICE_X12Y114_B2 = CLBLM_L_X10Y115_SLICE_X12Y115_BQ;
  assign CLBLM_L_X10Y114_SLICE_X12Y114_B3 = CLBLM_L_X8Y115_SLICE_X11Y115_C5Q;
  assign CLBLM_L_X10Y114_SLICE_X12Y114_B4 = RIOB33_X105Y121_IOB_X1Y121_I;
  assign CLBLM_L_X10Y114_SLICE_X12Y114_B5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y114_SLICE_X12Y114_B6 = 1'b1;
  assign CLBLL_L_X4Y110_SLICE_X4Y110_A1 = CLBLM_R_X3Y112_SLICE_X3Y112_C5Q;
  assign CLBLL_L_X4Y110_SLICE_X4Y110_A2 = CLBLM_R_X3Y118_SLICE_X2Y118_AQ;
  assign CLBLL_L_X4Y110_SLICE_X4Y110_A3 = CLBLL_L_X4Y110_SLICE_X4Y110_AQ;
  assign CLBLL_L_X4Y110_SLICE_X4Y110_A4 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLL_L_X4Y110_SLICE_X4Y110_A5 = 1'b1;
  assign CLBLL_L_X4Y110_SLICE_X4Y110_A6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y114_SLICE_X12Y114_C1 = CLBLM_L_X10Y114_SLICE_X13Y114_CQ;
  assign CLBLL_L_X4Y110_SLICE_X4Y110_AX = CLBLL_L_X4Y110_SLICE_X4Y110_BO6;
  assign CLBLM_L_X10Y114_SLICE_X12Y114_C2 = CLBLM_L_X10Y115_SLICE_X12Y115_AQ;
  assign CLBLL_L_X4Y110_SLICE_X4Y110_B1 = CLBLM_L_X8Y120_SLICE_X11Y120_CQ;
  assign CLBLL_L_X4Y110_SLICE_X4Y110_B2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLL_L_X4Y110_SLICE_X4Y110_B3 = CLBLM_R_X5Y121_SLICE_X6Y121_B5Q;
  assign CLBLL_L_X4Y110_SLICE_X4Y110_B4 = CLBLL_L_X4Y110_SLICE_X4Y110_DQ;
  assign CLBLL_L_X4Y110_SLICE_X4Y110_B5 = RIOB33_X105Y121_IOB_X1Y121_I;
  assign CLBLL_L_X4Y110_SLICE_X4Y110_B6 = 1'b1;
  assign CLBLM_L_X10Y114_SLICE_X12Y114_C4 = CLBLM_L_X10Y114_SLICE_X12Y114_AO5;
  assign CLBLM_L_X10Y114_SLICE_X12Y114_C5 = CLBLM_R_X5Y111_SLICE_X7Y111_DO6;
  assign CLBLM_L_X10Y114_SLICE_X12Y114_CE = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLL_L_X4Y110_SLICE_X4Y110_C1 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLL_L_X4Y110_SLICE_X4Y110_C2 = CLBLL_L_X4Y110_SLICE_X4Y110_AQ;
  assign CLBLL_L_X4Y110_SLICE_X4Y110_C3 = CLBLM_L_X10Y116_SLICE_X12Y116_CQ;
  assign CLBLL_L_X4Y110_SLICE_X4Y110_C4 = 1'b1;
  assign CLBLL_L_X4Y110_SLICE_X4Y110_C5 = CLBLL_L_X4Y110_SLICE_X4Y110_BO5;
  assign CLBLL_L_X4Y110_SLICE_X4Y110_C6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y114_SLICE_X12Y114_D1 = CLBLM_L_X10Y117_SLICE_X12Y117_AQ;
  assign CLBLL_L_X4Y110_SLICE_X4Y110_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X10Y114_SLICE_X12Y114_D2 = CLBLM_L_X8Y110_SLICE_X10Y110_AQ;
  assign CLBLM_L_X10Y114_SLICE_X12Y114_D3 = CLBLM_R_X11Y117_SLICE_X14Y117_BQ;
  assign CLBLM_L_X10Y114_SLICE_X12Y114_D4 = CLBLL_L_X4Y110_SLICE_X5Y110_BQ;
  assign CLBLM_L_X10Y114_SLICE_X12Y114_D5 = CLBLM_R_X7Y112_SLICE_X9Y112_CQ;
  assign CLBLM_L_X10Y114_SLICE_X12Y114_D6 = CLBLM_R_X5Y114_SLICE_X6Y114_DQ;
  assign CLBLL_L_X4Y110_SLICE_X4Y110_D1 = CLBLM_R_X3Y118_SLICE_X2Y118_AQ;
  assign CLBLL_L_X4Y110_SLICE_X4Y110_D2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLL_L_X4Y110_SLICE_X4Y110_D3 = CLBLL_L_X4Y110_SLICE_X4Y110_DQ;
  assign CLBLL_L_X4Y110_SLICE_X4Y110_D4 = CLBLM_R_X5Y112_SLICE_X7Y112_AO6;
  assign CLBLL_L_X4Y110_SLICE_X4Y110_D5 = CLBLM_R_X3Y111_SLICE_X3Y111_BQ;
  assign CLBLL_L_X4Y110_SLICE_X4Y110_D6 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLL_L_X4Y110_SLICE_X5Y110_A1 = CLBLM_R_X3Y111_SLICE_X2Y111_AQ;
  assign CLBLL_L_X4Y110_SLICE_X5Y110_A2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLL_L_X4Y110_SLICE_X5Y110_A3 = CLBLL_L_X4Y110_SLICE_X5Y110_AQ;
  assign CLBLL_L_X4Y110_SLICE_X5Y110_A4 = CLBLM_L_X10Y111_SLICE_X13Y111_BO6;
  assign CLBLL_L_X4Y110_SLICE_X5Y110_A5 = CLBLM_R_X7Y110_SLICE_X8Y110_DO5;
  assign CLBLL_L_X4Y110_SLICE_X5Y110_A6 = CLBLL_L_X4Y110_SLICE_X5Y110_CO6;
  assign CLBLL_L_X4Y110_SLICE_X5Y110_B1 = CLBLM_R_X5Y111_SLICE_X7Y111_DO6;
  assign CLBLL_L_X4Y110_SLICE_X5Y110_B2 = CLBLL_L_X4Y110_SLICE_X5Y110_BQ;
  assign CLBLL_L_X4Y110_SLICE_X5Y110_B3 = CLBLM_R_X5Y114_SLICE_X6Y114_DQ;
  assign CLBLL_L_X4Y110_SLICE_X5Y110_B4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLL_L_X4Y110_SLICE_X5Y110_B5 = CLBLL_L_X4Y113_SLICE_X5Y113_AQ;
  assign CLBLL_L_X4Y110_SLICE_X5Y110_B6 = 1'b1;
  assign CLBLL_L_X4Y110_SLICE_X5Y110_C1 = CLBLM_L_X8Y118_SLICE_X10Y118_DQ;
  assign CLBLL_L_X4Y110_SLICE_X5Y110_C2 = CLBLM_R_X5Y114_SLICE_X6Y114_BQ;
  assign CLBLL_L_X4Y110_SLICE_X5Y110_C3 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLL_L_X4Y110_SLICE_X5Y110_C4 = CLBLM_R_X3Y110_SLICE_X3Y110_BQ;
  assign CLBLL_L_X4Y110_SLICE_X5Y110_C5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLL_L_X4Y110_SLICE_X5Y110_C6 = 1'b1;
  assign CLBLL_L_X4Y110_SLICE_X5Y110_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLL_L_X4Y110_SLICE_X5Y110_D1 = CLBLM_R_X5Y109_SLICE_X6Y109_BQ;
  assign CLBLL_L_X4Y110_SLICE_X5Y110_D2 = CLBLM_R_X3Y110_SLICE_X3Y110_BQ;
  assign CLBLL_L_X4Y110_SLICE_X5Y110_D3 = 1'b1;
  assign CLBLL_L_X4Y110_SLICE_X5Y110_D4 = CLBLM_R_X5Y109_SLICE_X6Y109_AQ;
  assign CLBLL_L_X4Y110_SLICE_X5Y110_D5 = CLBLL_L_X4Y110_SLICE_X4Y110_AQ;
  assign CLBLL_L_X4Y110_SLICE_X5Y110_D6 = 1'b1;
  assign LIOB33_X0Y109_IOB_X0Y110_O = CLBLL_L_X2Y110_SLICE_X0Y110_AO5;
  assign LIOB33_X0Y109_IOB_X0Y109_O = CLBLL_L_X2Y110_SLICE_X0Y110_AO6;
  assign LIOI3_TBYTESRC_X0Y107_OLOGIC_X0Y108_D1 = CLBLL_L_X2Y111_SLICE_X0Y111_BO5;
  assign CLBLM_R_X5Y125_SLICE_X6Y125_B5 = CLBLM_R_X5Y125_SLICE_X6Y125_CO6;
  assign CLBLM_R_X5Y125_SLICE_X6Y125_B6 = 1'b1;
  assign LIOI3_TBYTETERM_X0Y187_OLOGIC_X0Y188_D1 = RIOB33_X105Y145_IOB_X1Y145_I;
  assign LIOB33_X0Y175_IOB_X0Y176_O = RIOB33_X105Y127_IOB_X1Y128_I;
  assign CLBLM_L_X10Y115_SLICE_X13Y115_A1 = CLBLM_R_X5Y111_SLICE_X7Y111_DO6;
  assign CLBLM_L_X10Y115_SLICE_X13Y115_A2 = CLBLM_R_X11Y115_SLICE_X14Y115_CQ;
  assign CLBLM_L_X10Y115_SLICE_X13Y115_A3 = CLBLM_L_X10Y111_SLICE_X13Y111_CO6;
  assign CLBLM_L_X10Y115_SLICE_X13Y115_A4 = CLBLM_L_X10Y115_SLICE_X12Y115_BQ;
  assign CLBLM_L_X10Y115_SLICE_X13Y115_A5 = CLBLM_L_X10Y112_SLICE_X13Y112_CQ;
  assign CLBLM_L_X10Y115_SLICE_X13Y115_A6 = CLBLM_L_X10Y116_SLICE_X13Y116_CQ;
  assign LIOB33_X0Y175_IOB_X0Y175_O = RIOB33_X105Y127_IOB_X1Y127_I;
  assign CLBLM_L_X10Y115_SLICE_X13Y115_B1 = CLBLM_R_X11Y115_SLICE_X14Y115_BQ;
  assign CLBLM_L_X10Y115_SLICE_X13Y115_B2 = CLBLM_R_X5Y111_SLICE_X7Y111_DO6;
  assign CLBLM_L_X10Y115_SLICE_X13Y115_B3 = CLBLM_L_X10Y111_SLICE_X13Y111_CO6;
  assign CLBLM_L_X10Y115_SLICE_X13Y115_B4 = CLBLM_L_X10Y112_SLICE_X13Y112_CQ;
  assign CLBLM_L_X10Y115_SLICE_X13Y115_B5 = CLBLM_R_X7Y112_SLICE_X9Y112_CQ;
  assign CLBLM_L_X10Y115_SLICE_X13Y115_B6 = CLBLM_R_X7Y115_SLICE_X9Y115_B5Q;
  assign CLBLM_L_X10Y115_SLICE_X13Y115_C1 = CLBLM_L_X8Y117_SLICE_X11Y117_BQ;
  assign CLBLM_L_X10Y115_SLICE_X13Y115_C2 = CLBLM_L_X10Y117_SLICE_X13Y117_BQ;
  assign CLBLM_L_X10Y115_SLICE_X13Y115_C3 = CLBLM_L_X10Y114_SLICE_X12Y114_DO6;
  assign CLBLM_L_X10Y115_SLICE_X13Y115_C4 = 1'b1;
  assign CLBLM_L_X10Y115_SLICE_X13Y115_C5 = CLBLM_L_X10Y115_SLICE_X13Y115_DO6;
  assign CLBLM_L_X10Y115_SLICE_X13Y115_C6 = CLBLM_L_X10Y115_SLICE_X12Y115_BQ;
  assign CLBLM_L_X10Y115_SLICE_X13Y115_D1 = CLBLM_R_X11Y115_SLICE_X15Y115_BQ;
  assign CLBLM_L_X10Y115_SLICE_X13Y115_D2 = CLBLM_R_X11Y115_SLICE_X15Y115_DQ;
  assign CLBLM_L_X10Y115_SLICE_X13Y115_D3 = 1'b1;
  assign CLBLM_L_X10Y115_SLICE_X13Y115_D4 = 1'b1;
  assign CLBLM_L_X10Y115_SLICE_X13Y115_D5 = CLBLM_L_X10Y115_SLICE_X12Y115_AQ;
  assign CLBLM_L_X10Y115_SLICE_X13Y115_D6 = CLBLM_L_X10Y119_SLICE_X12Y119_BQ;
  assign LIOI3_X0Y133_OLOGIC_X0Y134_D1 = CLBLM_R_X7Y124_SLICE_X8Y124_BQ;
  assign CLBLM_L_X10Y115_SLICE_X12Y115_A1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y115_SLICE_X12Y115_A2 = CLBLM_L_X10Y115_SLICE_X12Y115_AQ;
  assign CLBLM_L_X10Y115_SLICE_X12Y115_A3 = CLBLM_L_X8Y117_SLICE_X11Y117_BQ;
  assign CLBLM_L_X10Y115_SLICE_X12Y115_A4 = 1'b1;
  assign CLBLM_L_X10Y115_SLICE_X12Y115_A5 = CLBLM_L_X8Y123_SLICE_X11Y123_AQ;
  assign CLBLM_L_X10Y115_SLICE_X12Y115_A6 = CLBLM_R_X5Y111_SLICE_X7Y111_DO6;
  assign CLBLM_L_X10Y115_SLICE_X12Y115_B1 = CLBLM_R_X5Y111_SLICE_X7Y111_DO6;
  assign CLBLM_L_X10Y115_SLICE_X12Y115_B2 = CLBLM_L_X10Y115_SLICE_X12Y115_BQ;
  assign CLBLL_L_X4Y111_SLICE_X4Y111_A1 = CLBLL_L_X2Y113_SLICE_X1Y113_BQ;
  assign CLBLL_L_X4Y111_SLICE_X4Y111_A2 = CLBLL_L_X4Y111_SLICE_X5Y111_DO6;
  assign CLBLL_L_X4Y111_SLICE_X4Y111_A3 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLL_L_X4Y111_SLICE_X4Y111_A4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLL_L_X4Y111_SLICE_X4Y111_A5 = CLBLM_R_X3Y118_SLICE_X2Y118_AQ;
  assign CLBLL_L_X4Y111_SLICE_X4Y111_A6 = 1'b1;
  assign CLBLM_L_X10Y115_SLICE_X12Y115_B3 = 1'b1;
  assign CLBLM_L_X10Y115_SLICE_X12Y115_C1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLL_L_X4Y111_SLICE_X4Y111_B1 = CLBLM_R_X5Y115_SLICE_X6Y115_CO6;
  assign CLBLL_L_X4Y111_SLICE_X4Y111_B2 = CLBLL_L_X4Y111_SLICE_X4Y111_BQ;
  assign CLBLL_L_X4Y111_SLICE_X4Y111_B3 = 1'b1;
  assign CLBLL_L_X4Y111_SLICE_X4Y111_B4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLL_L_X4Y111_SLICE_X4Y111_B5 = CLBLM_R_X5Y111_SLICE_X6Y111_BQ;
  assign CLBLL_L_X4Y111_SLICE_X4Y111_B6 = CLBLM_R_X7Y109_SLICE_X8Y109_BQ;
  assign CLBLM_L_X10Y115_SLICE_X12Y115_C2 = CLBLM_L_X10Y115_SLICE_X12Y115_CQ;
  assign CLBLM_L_X10Y115_SLICE_X12Y115_C3 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X10Y115_SLICE_X12Y115_C4 = CLBLM_R_X7Y115_SLICE_X9Y115_DQ;
  assign CLBLL_L_X4Y111_SLICE_X4Y111_C1 = CLBLL_L_X4Y112_SLICE_X5Y112_AQ;
  assign CLBLL_L_X4Y111_SLICE_X4Y111_C2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLL_L_X4Y111_SLICE_X4Y111_C3 = CLBLM_R_X7Y121_SLICE_X9Y121_AQ;
  assign CLBLL_L_X4Y111_SLICE_X4Y111_C4 = CLBLM_R_X5Y112_SLICE_X7Y112_CO6;
  assign CLBLM_L_X10Y115_SLICE_X12Y115_D1 = 1'b1;
  assign CLBLM_L_X10Y115_SLICE_X12Y115_D2 = CLBLM_R_X5Y111_SLICE_X7Y111_DO6;
  assign CLBLM_L_X10Y115_SLICE_X12Y115_D3 = CLBLM_L_X10Y115_SLICE_X12Y115_DQ;
  assign CLBLM_L_X10Y115_SLICE_X12Y115_D4 = CLBLM_L_X10Y110_SLICE_X12Y110_BQ;
  assign CLBLL_L_X4Y111_SLICE_X4Y111_C6 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLL_L_X4Y111_SLICE_X4Y111_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLL_L_X4Y111_SLICE_X4Y111_C5 = 1'b1;
  assign CLBLM_L_X10Y115_SLICE_X12Y115_D5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLL_L_X4Y111_SLICE_X4Y111_D1 = CLBLL_L_X4Y112_SLICE_X5Y112_AQ;
  assign CLBLL_L_X4Y111_SLICE_X4Y111_D2 = 1'b1;
  assign CLBLL_L_X4Y111_SLICE_X4Y111_D3 = CLBLL_L_X4Y111_SLICE_X4Y111_DQ;
  assign CLBLL_L_X4Y111_SLICE_X4Y111_D4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLL_L_X4Y111_SLICE_X4Y111_D5 = 1'b1;
  assign CLBLL_L_X4Y111_SLICE_X4Y111_D6 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign LIOI3_X0Y133_OLOGIC_X0Y134_T1 = 1'b1;
  assign LIOI3_X0Y171_OLOGIC_X0Y172_D1 = CLBLM_R_X103Y138_SLICE_X163Y138_AO6;
  assign RIOI3_SING_X105Y100_ILOGIC_X1Y100_D = RIOB33_SING_X105Y100_IOB_X1Y100_I;
  assign LIOI3_X0Y171_OLOGIC_X0Y172_T1 = 1'b1;
  assign LIOI3_X0Y109_OLOGIC_X0Y110_D1 = CLBLL_L_X2Y110_SLICE_X0Y110_AO5;
  assign LIOI3_X0Y171_OLOGIC_X0Y171_D1 = LIOB33_SING_X0Y50_IOB_X0Y50_I;
  assign LIOI3_X0Y109_OLOGIC_X0Y110_T1 = 1'b1;
  assign CLBLM_R_X13Y119_SLICE_X19Y119_A1 = 1'b1;
  assign CLBLM_R_X13Y119_SLICE_X19Y119_A2 = 1'b1;
  assign CLBLM_R_X13Y119_SLICE_X19Y119_A3 = 1'b1;
  assign CLBLM_R_X13Y119_SLICE_X19Y119_A4 = 1'b1;
  assign CLBLM_R_X13Y119_SLICE_X19Y119_A5 = 1'b1;
  assign CLBLL_L_X4Y111_SLICE_X5Y111_A1 = 1'b1;
  assign CLBLL_L_X4Y111_SLICE_X5Y111_A2 = CLBLL_L_X4Y111_SLICE_X5Y111_BQ;
  assign CLBLL_L_X4Y111_SLICE_X5Y111_A3 = CLBLL_L_X4Y111_SLICE_X5Y111_AQ;
  assign CLBLL_L_X4Y111_SLICE_X5Y111_A4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLL_L_X4Y111_SLICE_X5Y111_A5 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLL_L_X4Y111_SLICE_X5Y111_A6 = 1'b1;
  assign CLBLM_R_X13Y119_SLICE_X19Y119_B1 = 1'b1;
  assign CLBLM_R_X13Y119_SLICE_X19Y119_B2 = 1'b1;
  assign CLBLL_L_X4Y111_SLICE_X5Y111_AX = CLBLL_L_X4Y110_SLICE_X5Y110_CO5;
  assign CLBLM_R_X13Y119_SLICE_X19Y119_B3 = 1'b1;
  assign CLBLL_L_X4Y111_SLICE_X5Y111_B1 = 1'b1;
  assign CLBLL_L_X4Y111_SLICE_X5Y111_B2 = CLBLM_R_X5Y110_SLICE_X6Y110_BO6;
  assign CLBLL_L_X4Y111_SLICE_X5Y111_B3 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLL_L_X4Y111_SLICE_X5Y111_B4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLL_L_X4Y111_SLICE_X5Y111_B5 = CLBLM_R_X7Y120_SLICE_X8Y120_DQ;
  assign CLBLL_L_X4Y111_SLICE_X5Y111_B6 = CLBLL_L_X4Y112_SLICE_X5Y112_DO6;
  assign CLBLM_R_X13Y119_SLICE_X19Y119_B4 = 1'b1;
  assign CLBLM_R_X13Y119_SLICE_X19Y119_B5 = 1'b1;
  assign CLBLM_R_X13Y119_SLICE_X19Y119_B6 = 1'b1;
  assign CLBLL_L_X4Y111_SLICE_X5Y111_C1 = CLBLL_L_X4Y114_SLICE_X5Y114_DO6;
  assign CLBLL_L_X4Y111_SLICE_X5Y111_C2 = CLBLM_R_X5Y111_SLICE_X6Y111_CQ;
  assign CLBLL_L_X4Y111_SLICE_X5Y111_C3 = CLBLM_R_X7Y113_SLICE_X8Y113_AQ;
  assign CLBLL_L_X4Y111_SLICE_X5Y111_C4 = CLBLL_L_X4Y114_SLICE_X5Y114_BO6;
  assign CLBLL_L_X4Y111_SLICE_X5Y111_C5 = CLBLM_R_X3Y115_SLICE_X3Y115_DQ;
  assign CLBLL_L_X4Y111_SLICE_X5Y111_C6 = CLBLL_L_X4Y115_SLICE_X4Y115_BQ;
  assign CLBLM_R_X13Y119_SLICE_X19Y119_C3 = 1'b1;
  assign CLBLM_R_X13Y119_SLICE_X19Y119_C4 = 1'b1;
  assign CLBLL_L_X4Y111_SLICE_X5Y111_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X13Y119_SLICE_X19Y119_C6 = 1'b1;
  assign CLBLM_R_X7Y151_SLICE_X9Y151_A1 = 1'b1;
  assign CLBLM_R_X7Y151_SLICE_X9Y151_A2 = 1'b1;
  assign CLBLM_R_X7Y151_SLICE_X9Y151_A3 = 1'b1;
  assign CLBLL_L_X4Y111_SLICE_X5Y111_D1 = CLBLL_L_X4Y111_SLICE_X4Y111_AQ;
  assign CLBLL_L_X4Y111_SLICE_X5Y111_D2 = 1'b1;
  assign CLBLL_L_X4Y111_SLICE_X5Y111_D3 = CLBLL_L_X4Y120_SLICE_X4Y120_BO6;
  assign CLBLL_L_X4Y111_SLICE_X5Y111_D4 = CLBLM_R_X5Y116_SLICE_X7Y116_CQ;
  assign CLBLL_L_X4Y111_SLICE_X5Y111_D5 = CLBLM_R_X7Y109_SLICE_X8Y109_AQ;
  assign CLBLL_L_X4Y111_SLICE_X5Y111_D6 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X7Y151_SLICE_X9Y151_A4 = 1'b1;
  assign CLBLM_R_X7Y151_SLICE_X9Y151_A5 = 1'b1;
  assign CLBLM_R_X7Y151_SLICE_X9Y151_A6 = 1'b1;
  assign CLBLM_R_X7Y151_SLICE_X9Y151_B1 = 1'b1;
  assign CLBLM_R_X7Y151_SLICE_X9Y151_B2 = 1'b1;
  assign CLBLM_R_X7Y151_SLICE_X9Y151_B3 = 1'b1;
  assign CLBLM_R_X7Y151_SLICE_X9Y151_B4 = 1'b1;
  assign CLBLM_R_X7Y151_SLICE_X9Y151_B5 = 1'b1;
  assign CLBLM_R_X7Y151_SLICE_X9Y151_B6 = 1'b1;
  assign CLBLM_R_X7Y151_SLICE_X9Y151_C1 = 1'b1;
  assign CLBLM_R_X7Y151_SLICE_X9Y151_C2 = 1'b1;
  assign CLBLM_R_X7Y151_SLICE_X9Y151_C3 = 1'b1;
  assign CLBLM_R_X7Y151_SLICE_X9Y151_C4 = 1'b1;
  assign CLBLM_R_X7Y151_SLICE_X9Y151_C5 = 1'b1;
  assign CLBLM_R_X7Y151_SLICE_X9Y151_C6 = 1'b1;
  assign CLBLM_R_X13Y119_SLICE_X18Y119_B1 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X13Y119_SLICE_X18Y119_B2 = CLBLM_R_X13Y119_SLICE_X18Y119_BQ;
  assign CLBLM_R_X13Y119_SLICE_X18Y119_B3 = CLBLM_R_X11Y117_SLICE_X14Y117_BQ;
  assign CLBLM_R_X13Y119_SLICE_X18Y119_B4 = RIOB33_X105Y121_IOB_X1Y121_I;
  assign CLBLM_R_X13Y119_SLICE_X18Y119_B5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y151_SLICE_X9Y151_D1 = 1'b1;
  assign CLBLM_R_X7Y151_SLICE_X9Y151_D2 = 1'b1;
  assign CLBLM_R_X7Y151_SLICE_X9Y151_D3 = 1'b1;
  assign CLBLM_R_X7Y151_SLICE_X9Y151_D4 = 1'b1;
  assign CLBLM_R_X7Y151_SLICE_X9Y151_D5 = 1'b1;
  assign CLBLM_R_X7Y151_SLICE_X9Y151_D6 = 1'b1;
  assign CLBLM_R_X13Y119_SLICE_X18Y119_C1 = CLBLM_R_X11Y120_SLICE_X14Y120_BO6;
  assign CLBLM_R_X13Y119_SLICE_X18Y119_C2 = CLBLM_R_X13Y119_SLICE_X18Y119_CQ;
  assign CLBLM_R_X13Y119_SLICE_X18Y119_C3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X13Y119_SLICE_X18Y119_C4 = CLBLL_L_X4Y118_SLICE_X5Y118_CQ;
  assign CLBLM_R_X13Y119_SLICE_X18Y119_C5 = RIOB33_X105Y121_IOB_X1Y121_I;
  assign CLBLM_R_X7Y151_SLICE_X8Y151_A1 = 1'b1;
  assign CLBLM_R_X7Y151_SLICE_X8Y151_A2 = 1'b1;
  assign CLBLM_R_X7Y151_SLICE_X8Y151_A3 = 1'b1;
  assign CLBLM_R_X7Y151_SLICE_X8Y151_A4 = 1'b1;
  assign CLBLM_R_X7Y151_SLICE_X8Y151_A5 = 1'b1;
  assign CLBLM_R_X7Y151_SLICE_X8Y151_A6 = CLBLM_R_X5Y113_SLICE_X7Y113_A5Q;
  assign CLBLM_R_X13Y119_SLICE_X18Y119_D1 = CLBLM_R_X11Y118_SLICE_X15Y118_AQ;
  assign CLBLM_R_X13Y119_SLICE_X18Y119_D2 = CLBLM_L_X12Y120_SLICE_X17Y120_AQ;
  assign CLBLM_R_X13Y119_SLICE_X18Y119_D3 = CLBLM_L_X10Y119_SLICE_X13Y119_AQ;
  assign CLBLM_R_X7Y151_SLICE_X8Y151_B1 = 1'b1;
  assign CLBLM_R_X7Y151_SLICE_X8Y151_B2 = 1'b1;
  assign CLBLM_R_X7Y151_SLICE_X8Y151_B3 = 1'b1;
  assign CLBLM_R_X7Y151_SLICE_X8Y151_B4 = 1'b1;
  assign CLBLM_R_X7Y151_SLICE_X8Y151_B5 = 1'b1;
  assign CLBLM_R_X7Y151_SLICE_X8Y151_B6 = 1'b1;
  assign LIOI3_X0Y133_OLOGIC_X0Y133_T1 = 1'b1;
  assign LIOI3_TBYTESRC_X0Y119_OLOGIC_X0Y120_T1 = 1'b1;
  assign CLBLM_R_X7Y151_SLICE_X8Y151_C1 = 1'b1;
  assign CLBLM_R_X7Y151_SLICE_X8Y151_C2 = 1'b1;
  assign CLBLM_R_X7Y151_SLICE_X8Y151_C3 = 1'b1;
  assign CLBLM_R_X7Y151_SLICE_X8Y151_C4 = 1'b1;
  assign CLBLM_R_X7Y151_SLICE_X8Y151_C5 = 1'b1;
  assign CLBLM_R_X7Y151_SLICE_X8Y151_C6 = 1'b1;
  assign CLBLM_R_X7Y151_SLICE_X8Y151_D1 = 1'b1;
  assign CLBLM_R_X7Y151_SLICE_X8Y151_D2 = 1'b1;
  assign CLBLM_R_X7Y151_SLICE_X8Y151_D3 = 1'b1;
  assign CLBLM_R_X7Y151_SLICE_X8Y151_D4 = 1'b1;
  assign CLBLM_R_X7Y151_SLICE_X8Y151_D5 = 1'b1;
  assign CLBLM_R_X7Y151_SLICE_X8Y151_D6 = 1'b1;
  assign LIOB33_X0Y177_IOB_X0Y178_O = RIOB33_X105Y129_IOB_X1Y130_I;
  assign LIOB33_X0Y177_IOB_X0Y177_O = RIOB33_X105Y129_IOB_X1Y129_I;
  assign CLBLM_R_X103Y172_SLICE_X162Y172_D3 = 1'b1;
  assign CLBLM_L_X10Y124_SLICE_X12Y124_B1 = 1'b1;
  assign CLBLM_L_X10Y116_SLICE_X13Y116_A1 = RIOB33_X105Y103_IOB_X1Y104_I;
  assign CLBLM_L_X10Y116_SLICE_X13Y116_A2 = CLBLM_L_X10Y117_SLICE_X13Y117_AQ;
  assign CLBLM_L_X10Y116_SLICE_X13Y116_A3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y116_SLICE_X13Y116_A4 = CLBLM_L_X10Y115_SLICE_X13Y115_CO6;
  assign CLBLM_L_X10Y116_SLICE_X13Y116_A5 = CLBLM_L_X10Y116_SLICE_X13Y116_DQ;
  assign CLBLM_L_X10Y116_SLICE_X13Y116_A6 = 1'b1;
  assign CLBLM_L_X10Y116_SLICE_X13Y116_AX = CLBLM_R_X11Y116_SLICE_X14Y116_BO6;
  assign CLBLM_L_X10Y116_SLICE_X13Y116_B1 = CLBLM_L_X10Y117_SLICE_X13Y117_DQ;
  assign CLBLM_L_X10Y116_SLICE_X13Y116_B2 = CLBLM_L_X10Y112_SLICE_X13Y112_BQ;
  assign CLBLM_L_X10Y116_SLICE_X13Y116_B3 = CLBLM_R_X5Y119_SLICE_X6Y119_BQ;
  assign CLBLM_L_X10Y116_SLICE_X13Y116_B4 = RIOB33_X105Y121_IOB_X1Y121_I;
  assign CLBLM_L_X10Y116_SLICE_X13Y116_B5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y116_SLICE_X13Y116_B6 = 1'b1;
  assign CLBLM_R_X5Y121_SLICE_X7Y121_D1 = CLBLM_R_X5Y123_SLICE_X7Y123_AQ;
  assign CLBLM_L_X10Y116_SLICE_X13Y116_C1 = CLBLM_L_X10Y116_SLICE_X12Y116_AQ;
  assign CLBLM_L_X10Y116_SLICE_X13Y116_C2 = CLBLM_L_X8Y119_SLICE_X10Y119_BQ;
  assign CLBLM_L_X10Y116_SLICE_X13Y116_C3 = CLBLM_L_X10Y116_SLICE_X13Y116_BQ;
  assign CLBLM_L_X10Y116_SLICE_X13Y116_C4 = CLBLM_L_X8Y116_SLICE_X11Y116_A5Q;
  assign CLBLM_L_X10Y116_SLICE_X13Y116_C5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y116_SLICE_X13Y116_C6 = 1'b1;
  assign CLBLM_L_X10Y116_SLICE_X13Y116_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X10Y116_SLICE_X13Y116_D1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y116_SLICE_X13Y116_D2 = CLBLM_L_X10Y117_SLICE_X13Y117_AQ;
  assign CLBLM_L_X10Y116_SLICE_X13Y116_D3 = CLBLM_L_X10Y116_SLICE_X13Y116_DQ;
  assign CLBLM_L_X10Y116_SLICE_X13Y116_D4 = CLBLM_R_X7Y117_SLICE_X8Y117_A5Q;
  assign CLBLM_L_X10Y116_SLICE_X13Y116_D5 = CLBLM_R_X5Y111_SLICE_X7Y111_DO6;
  assign CLBLM_L_X10Y116_SLICE_X13Y116_D6 = 1'b1;
  assign CLBLM_R_X5Y121_SLICE_X7Y121_D2 = CLBLM_R_X7Y121_SLICE_X9Y121_BQ;
  assign CLBLM_L_X10Y116_SLICE_X12Y116_A1 = CLBLM_L_X10Y114_SLICE_X12Y114_AQ;
  assign CLBLM_L_X10Y116_SLICE_X12Y116_A2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y116_SLICE_X12Y116_A3 = CLBLM_L_X10Y116_SLICE_X12Y116_AQ;
  assign CLBLM_L_X10Y116_SLICE_X12Y116_A4 = CLBLM_L_X10Y116_SLICE_X12Y116_DO5;
  assign CLBLM_L_X10Y116_SLICE_X12Y116_A5 = CLBLM_L_X8Y116_SLICE_X11Y116_CO5;
  assign CLBLM_L_X10Y116_SLICE_X12Y116_A6 = CLBLM_R_X11Y119_SLICE_X14Y119_AO6;
  assign CLBLM_L_X10Y124_SLICE_X12Y124_C1 = 1'b1;
  assign CLBLL_L_X4Y112_SLICE_X4Y112_A1 = CLBLM_R_X5Y114_SLICE_X6Y114_AQ;
  assign CLBLL_L_X4Y112_SLICE_X4Y112_A2 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLL_L_X4Y112_SLICE_X4Y112_A3 = CLBLL_L_X4Y112_SLICE_X4Y112_AQ;
  assign CLBLL_L_X4Y112_SLICE_X4Y112_A4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLL_L_X4Y112_SLICE_X4Y112_A5 = CLBLM_R_X3Y118_SLICE_X2Y118_AQ;
  assign CLBLL_L_X4Y112_SLICE_X4Y112_A6 = CLBLM_R_X3Y115_SLICE_X2Y115_CQ;
  assign CLBLM_L_X10Y116_SLICE_X12Y116_AX = CLBLM_L_X10Y114_SLICE_X12Y114_BO6;
  assign CLBLM_L_X10Y116_SLICE_X12Y116_B1 = CLBLM_L_X10Y116_SLICE_X12Y116_DO6;
  assign CLBLM_L_X10Y116_SLICE_X12Y116_B2 = CLBLM_L_X10Y116_SLICE_X12Y116_BQ;
  assign CLBLL_L_X4Y112_SLICE_X4Y112_B1 = 1'b1;
  assign CLBLL_L_X4Y112_SLICE_X4Y112_B2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLL_L_X4Y112_SLICE_X4Y112_B3 = CLBLM_R_X5Y112_SLICE_X6Y112_BO6;
  assign CLBLL_L_X4Y112_SLICE_X4Y112_B4 = CLBLL_L_X4Y113_SLICE_X5Y113_CQ;
  assign CLBLL_L_X4Y112_SLICE_X4Y112_B5 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLL_L_X4Y112_SLICE_X4Y112_B6 = CLBLM_R_X3Y115_SLICE_X2Y115_CQ;
  assign CLBLM_L_X10Y116_SLICE_X12Y116_B5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y116_SLICE_X12Y116_B6 = CLBLM_R_X11Y119_SLICE_X14Y119_AO6;
  assign CLBLL_L_X4Y112_SLICE_X4Y112_C1 = 1'b1;
  assign CLBLL_L_X4Y112_SLICE_X4Y112_C2 = CLBLL_L_X4Y111_SLICE_X4Y111_CQ;
  assign CLBLL_L_X4Y112_SLICE_X4Y112_C3 = CLBLM_R_X7Y122_SLICE_X9Y122_BQ;
  assign CLBLL_L_X4Y112_SLICE_X4Y112_C4 = CLBLL_L_X4Y111_SLICE_X5Y111_A5Q;
  assign CLBLL_L_X4Y112_SLICE_X4Y112_C5 = 1'b1;
  assign CLBLL_L_X4Y112_SLICE_X4Y112_C6 = CLBLL_L_X4Y111_SLICE_X5Y111_BQ;
  assign CLBLM_L_X10Y116_SLICE_X12Y116_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X10Y116_SLICE_X12Y116_C5 = CLBLM_L_X10Y119_SLICE_X12Y119_CQ;
  assign CLBLL_L_X4Y112_SLICE_X4Y112_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X10Y116_SLICE_X12Y116_D1 = CLBLM_L_X10Y116_SLICE_X12Y116_BQ;
  assign CLBLM_L_X10Y116_SLICE_X12Y116_D2 = CLBLM_L_X8Y116_SLICE_X11Y116_A5Q;
  assign CLBLM_L_X10Y116_SLICE_X12Y116_D3 = CLBLM_R_X11Y116_SLICE_X14Y116_CQ;
  assign CLBLM_L_X10Y116_SLICE_X12Y116_D4 = CLBLM_L_X8Y119_SLICE_X10Y119_BQ;
  assign CLBLL_L_X4Y112_SLICE_X4Y112_D1 = 1'b1;
  assign CLBLL_L_X4Y112_SLICE_X4Y112_D2 = 1'b1;
  assign CLBLL_L_X4Y112_SLICE_X4Y112_D3 = 1'b1;
  assign CLBLL_L_X4Y112_SLICE_X4Y112_D4 = CLBLM_R_X7Y120_SLICE_X9Y120_CQ;
  assign CLBLL_L_X4Y112_SLICE_X4Y112_D5 = 1'b1;
  assign CLBLL_L_X4Y112_SLICE_X4Y112_D6 = CLBLM_R_X5Y114_SLICE_X7Y114_AQ;
  assign CLBLM_L_X10Y116_SLICE_X12Y116_D5 = CLBLM_L_X10Y116_SLICE_X12Y116_AQ;
  assign CLBLM_L_X10Y116_SLICE_X12Y116_D6 = 1'b1;
  assign CLBLM_L_X10Y124_SLICE_X12Y124_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLL_L_X4Y112_SLICE_X5Y112_A1 = CLBLM_R_X5Y114_SLICE_X7Y114_DO6;
  assign CLBLL_L_X4Y112_SLICE_X5Y112_A2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLL_L_X4Y112_SLICE_X5Y112_A3 = CLBLM_R_X5Y111_SLICE_X6Y111_BQ;
  assign CLBLL_L_X4Y112_SLICE_X5Y112_A4 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLL_L_X4Y112_SLICE_X5Y112_A5 = CLBLL_L_X4Y112_SLICE_X4Y112_AQ;
  assign CLBLL_L_X4Y112_SLICE_X5Y112_A6 = 1'b1;
  assign CLBLM_R_X11Y120_SLICE_X15Y120_C2 = 1'b1;
  assign CLBLM_R_X11Y120_SLICE_X15Y120_C3 = CLBLM_R_X7Y121_SLICE_X9Y121_DO6;
  assign CLBLM_R_X13Y120_SLICE_X19Y120_A1 = 1'b1;
  assign CLBLL_L_X4Y112_SLICE_X5Y112_B1 = CLBLM_L_X10Y116_SLICE_X13Y116_AQ;
  assign CLBLL_L_X4Y112_SLICE_X5Y112_B2 = 1'b1;
  assign CLBLL_L_X4Y112_SLICE_X5Y112_B3 = CLBLM_R_X3Y112_SLICE_X3Y112_BQ;
  assign CLBLL_L_X4Y112_SLICE_X5Y112_B4 = CLBLL_L_X4Y112_SLICE_X4Y112_CO6;
  assign CLBLL_L_X4Y112_SLICE_X5Y112_B5 = CLBLL_L_X4Y114_SLICE_X5Y114_CO6;
  assign CLBLL_L_X4Y112_SLICE_X5Y112_B6 = CLBLL_L_X4Y112_SLICE_X5Y112_CO6;
  assign CLBLM_R_X11Y120_SLICE_X15Y120_C4 = CLBLM_R_X11Y119_SLICE_X14Y119_AO6;
  assign CLBLM_R_X11Y120_SLICE_X15Y120_C5 = CLBLM_R_X11Y120_SLICE_X15Y120_DO6;
  assign CLBLM_R_X13Y120_SLICE_X19Y120_B1 = 1'b1;
  assign CLBLL_L_X4Y112_SLICE_X5Y112_C1 = CLBLL_L_X2Y113_SLICE_X1Y113_BQ;
  assign CLBLL_L_X4Y112_SLICE_X5Y112_C2 = CLBLM_R_X5Y114_SLICE_X6Y114_BQ;
  assign CLBLL_L_X4Y112_SLICE_X5Y112_C3 = 1'b1;
  assign CLBLL_L_X4Y112_SLICE_X5Y112_C4 = CLBLM_R_X5Y111_SLICE_X6Y111_BQ;
  assign CLBLL_L_X4Y112_SLICE_X5Y112_C5 = CLBLL_L_X4Y113_SLICE_X4Y113_BQ;
  assign CLBLL_L_X4Y112_SLICE_X5Y112_C6 = CLBLM_R_X7Y117_SLICE_X8Y117_CQ;
  assign CLBLM_R_X11Y120_SLICE_X15Y120_C6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLL_L_X4Y112_SLICE_X5Y112_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X13Y120_SLICE_X19Y120_C1 = 1'b1;
  assign CLBLM_R_X13Y120_SLICE_X19Y120_C2 = 1'b1;
  assign CLBLM_R_X13Y120_SLICE_X19Y120_C3 = 1'b1;
  assign CLBLM_R_X13Y120_SLICE_X19Y120_C4 = 1'b1;
  assign CLBLM_R_X13Y120_SLICE_X19Y120_C6 = 1'b1;
  assign CLBLL_L_X4Y112_SLICE_X5Y112_D1 = 1'b1;
  assign CLBLL_L_X4Y112_SLICE_X5Y112_D2 = 1'b1;
  assign CLBLL_L_X4Y112_SLICE_X5Y112_D3 = CLBLM_L_X8Y120_SLICE_X10Y120_BQ;
  assign CLBLL_L_X4Y112_SLICE_X5Y112_D4 = CLBLM_L_X10Y116_SLICE_X13Y116_AQ;
  assign CLBLL_L_X4Y112_SLICE_X5Y112_D5 = CLBLM_R_X7Y122_SLICE_X9Y122_BQ;
  assign CLBLL_L_X4Y112_SLICE_X5Y112_D6 = CLBLL_L_X4Y111_SLICE_X5Y111_BQ;
  assign CLBLM_R_X13Y120_SLICE_X19Y120_D1 = 1'b1;
  assign CLBLM_R_X13Y120_SLICE_X19Y120_D2 = 1'b1;
  assign CLBLM_R_X13Y120_SLICE_X19Y120_D3 = 1'b1;
  assign CLBLM_R_X13Y120_SLICE_X19Y120_D4 = 1'b1;
  assign CLBLM_R_X13Y120_SLICE_X19Y120_D5 = 1'b1;
  assign CLBLM_R_X13Y120_SLICE_X18Y120_A1 = CLBLM_L_X12Y120_SLICE_X17Y120_BQ;
  assign CLBLM_R_X13Y120_SLICE_X18Y120_A2 = CLBLM_R_X11Y119_SLICE_X15Y119_AQ;
  assign CLBLM_R_X13Y120_SLICE_X18Y120_A3 = CLBLM_R_X11Y118_SLICE_X15Y118_AQ;
  assign CLBLM_R_X13Y120_SLICE_X18Y120_A4 = CLBLM_L_X12Y120_SLICE_X17Y120_AQ;
  assign CLBLM_R_X13Y120_SLICE_X18Y120_A5 = CLBLM_R_X11Y120_SLICE_X15Y120_AQ;
  assign CLBLM_R_X13Y120_SLICE_X18Y120_A6 = CLBLM_L_X12Y120_SLICE_X17Y120_DO6;
  assign CLBLM_R_X13Y120_SLICE_X18Y120_B1 = CLBLM_L_X12Y120_SLICE_X17Y120_BQ;
  assign CLBLM_R_X13Y120_SLICE_X18Y120_B2 = CLBLM_R_X11Y119_SLICE_X15Y119_AQ;
  assign CLBLM_R_X13Y120_SLICE_X18Y120_B3 = CLBLM_R_X11Y118_SLICE_X15Y118_AQ;
  assign CLBLM_R_X13Y120_SLICE_X18Y120_B4 = CLBLM_L_X12Y120_SLICE_X17Y120_DO6;
  assign CLBLM_R_X13Y120_SLICE_X18Y120_B5 = CLBLM_R_X11Y120_SLICE_X15Y120_AQ;
  assign CLBLM_R_X13Y120_SLICE_X18Y120_B6 = CLBLM_L_X12Y120_SLICE_X17Y120_AQ;
  assign CLBLM_R_X13Y120_SLICE_X18Y120_C1 = CLBLM_R_X11Y118_SLICE_X15Y118_AQ;
  assign CLBLM_R_X11Y120_SLICE_X15Y120_D1 = CLBLM_R_X11Y120_SLICE_X15Y120_BQ;
  assign CLBLM_R_X13Y120_SLICE_X18Y120_C2 = CLBLM_R_X11Y120_SLICE_X15Y120_AQ;
  assign CLBLM_R_X13Y120_SLICE_X18Y120_C3 = CLBLM_L_X10Y119_SLICE_X13Y119_AQ;
  assign CLBLM_R_X13Y120_SLICE_X18Y120_C4 = CLBLM_R_X11Y119_SLICE_X15Y119_CQ;
  assign CLBLM_R_X13Y120_SLICE_X18Y120_C5 = CLBLM_R_X11Y118_SLICE_X14Y118_BQ;
  assign CLBLM_R_X11Y120_SLICE_X15Y120_D2 = CLBLM_R_X11Y120_SLICE_X15Y120_CQ;
  assign CLBLM_R_X13Y120_SLICE_X18Y120_C6 = CLBLM_L_X12Y120_SLICE_X17Y120_AQ;
  assign CLBLM_R_X13Y120_SLICE_X18Y120_D1 = 1'b1;
  assign CLBLM_R_X13Y120_SLICE_X18Y120_D2 = 1'b1;
  assign CLBLM_R_X13Y120_SLICE_X18Y120_D3 = 1'b1;
  assign CLBLM_R_X13Y120_SLICE_X18Y120_D4 = 1'b1;
  assign CLBLM_R_X13Y120_SLICE_X18Y120_D5 = 1'b1;
  assign CLBLM_R_X11Y120_SLICE_X15Y120_D5 = CLBLM_L_X8Y119_SLICE_X10Y119_CQ;
  assign CLBLM_R_X13Y120_SLICE_X18Y120_D6 = 1'b1;
  assign LIOI3_X0Y195_OLOGIC_X0Y196_T1 = 1'b1;
  assign CLBLM_R_X11Y120_SLICE_X15Y120_D6 = CLBLM_L_X12Y120_SLICE_X17Y120_CO6;
  assign LIOB33_X0Y179_IOB_X0Y180_O = RIOB33_X105Y131_IOB_X1Y132_I;
  assign LIOB33_X0Y179_IOB_X0Y179_O = RIOB33_X105Y131_IOB_X1Y131_I;
  assign CLBLL_L_X2Y109_SLICE_X0Y109_A4 = CLBLL_L_X2Y110_SLICE_X0Y110_BO6;
  assign LIOI3_X0Y195_OLOGIC_X0Y195_D1 = LIOB33_X0Y63_IOB_X0Y64_I;
  assign CLBLL_L_X2Y109_SLICE_X0Y109_A6 = 1'b1;
  assign CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_I0 = LIOB33_X0Y77_IOB_X0Y78_I;
  assign CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_I1 = 1'b1;
  assign CLBLM_R_X7Y122_SLICE_X9Y122_C4 = CLBLM_L_X10Y124_SLICE_X12Y124_AQ;
  assign CLBLM_L_X10Y117_SLICE_X13Y117_A1 = CLBLM_L_X10Y119_SLICE_X12Y119_CQ;
  assign CLBLM_L_X10Y117_SLICE_X13Y117_A2 = CLBLM_L_X10Y119_SLICE_X12Y119_BQ;
  assign CLBLM_L_X10Y117_SLICE_X13Y117_A3 = CLBLM_L_X10Y117_SLICE_X13Y117_AQ;
  assign CLBLM_L_X10Y117_SLICE_X13Y117_A4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y117_SLICE_X13Y117_A5 = CLBLM_R_X5Y119_SLICE_X7Y119_AO6;
  assign CLBLM_L_X10Y117_SLICE_X13Y117_A6 = 1'b1;
  assign CLBLL_L_X2Y109_SLICE_X0Y109_B4 = 1'b1;
  assign CLBLM_R_X7Y122_SLICE_X9Y122_C5 = CLBLM_R_X7Y123_SLICE_X9Y123_BO5;
  assign CLBLM_R_X7Y122_SLICE_X9Y122_C6 = CLBLM_R_X5Y120_SLICE_X6Y120_A5Q;
  assign CLBLM_L_X10Y117_SLICE_X13Y117_B1 = 1'b1;
  assign CLBLM_L_X10Y117_SLICE_X13Y117_B2 = CLBLM_L_X10Y117_SLICE_X13Y117_BQ;
  assign CLBLM_L_X10Y117_SLICE_X13Y117_B3 = CLBLM_R_X5Y119_SLICE_X7Y119_AO6;
  assign CLBLM_L_X10Y117_SLICE_X13Y117_B4 = CLBLM_R_X11Y118_SLICE_X15Y118_BQ;
  assign CLBLM_L_X10Y117_SLICE_X13Y117_B5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y117_SLICE_X13Y117_B6 = CLBLM_R_X11Y115_SLICE_X15Y115_BQ;
  assign CLBLL_L_X2Y109_SLICE_X0Y109_B5 = 1'b1;
  assign CLBLL_L_X2Y109_SLICE_X0Y109_B6 = 1'b1;
  assign CLBLM_R_X11Y120_SLICE_X14Y120_B4 = CLBLM_R_X11Y120_SLICE_X15Y120_BQ;
  assign CLBLM_L_X10Y117_SLICE_X13Y117_C1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y117_SLICE_X13Y117_C2 = CLBLM_L_X10Y117_SLICE_X13Y117_CQ;
  assign CLBLM_L_X10Y117_SLICE_X13Y117_C3 = CLBLM_L_X10Y116_SLICE_X13Y116_DQ;
  assign CLBLM_L_X10Y117_SLICE_X13Y117_C4 = CLBLM_R_X7Y119_SLICE_X8Y119_D5Q;
  assign CLBLM_L_X10Y117_SLICE_X13Y117_C5 = CLBLM_R_X3Y112_SLICE_X3Y112_AQ;
  assign CLBLM_L_X10Y117_SLICE_X13Y117_C6 = CLBLM_L_X10Y113_SLICE_X13Y113_BO6;
  assign CLBLM_R_X11Y120_SLICE_X14Y120_B5 = CLBLM_R_X11Y119_SLICE_X15Y119_CQ;
  assign LIOI3_X0Y195_OLOGIC_X0Y195_T1 = 1'b1;
  assign CLBLM_L_X10Y117_SLICE_X13Y117_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X11Y120_SLICE_X14Y120_B6 = 1'b1;
  assign CLBLM_L_X10Y117_SLICE_X13Y117_D1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y117_SLICE_X13Y117_D2 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_L_X10Y117_SLICE_X13Y117_D3 = CLBLM_L_X10Y117_SLICE_X13Y117_DQ;
  assign CLBLM_L_X10Y117_SLICE_X13Y117_D4 = CLBLM_R_X13Y119_SLICE_X18Y119_AQ;
  assign CLBLM_L_X10Y117_SLICE_X13Y117_D5 = CLBLM_R_X3Y118_SLICE_X2Y118_AQ;
  assign CLBLM_L_X10Y117_SLICE_X13Y117_D6 = CLBLM_R_X7Y113_SLICE_X8Y113_CO6;
  assign CLBLL_L_X2Y109_SLICE_X0Y109_C1 = 1'b1;
  assign CLBLL_L_X2Y109_SLICE_X0Y109_C2 = 1'b1;
  assign CLBLM_L_X10Y117_SLICE_X12Y117_A1 = 1'b1;
  assign CLBLM_L_X10Y117_SLICE_X12Y117_A2 = CLBLM_R_X11Y116_SLICE_X15Y116_AQ;
  assign CLBLM_L_X10Y117_SLICE_X12Y117_A3 = CLBLM_L_X10Y117_SLICE_X12Y117_AQ;
  assign CLBLM_L_X10Y117_SLICE_X12Y117_A4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y117_SLICE_X12Y117_A5 = CLBLM_R_X7Y112_SLICE_X9Y112_CQ;
  assign CLBLM_L_X10Y117_SLICE_X12Y117_A6 = CLBLM_R_X5Y111_SLICE_X7Y111_DO6;
  assign CLBLL_L_X4Y113_SLICE_X4Y113_A1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLL_L_X4Y113_SLICE_X4Y113_A2 = CLBLM_R_X5Y110_SLICE_X7Y110_BQ;
  assign CLBLL_L_X4Y113_SLICE_X4Y113_A3 = CLBLL_L_X4Y113_SLICE_X4Y113_AQ;
  assign CLBLL_L_X4Y113_SLICE_X4Y113_A4 = CLBLM_R_X11Y113_SLICE_X15Y113_AQ;
  assign CLBLM_L_X10Y117_SLICE_X12Y117_B1 = CLBLL_L_X2Y117_SLICE_X0Y117_AQ;
  assign CLBLM_L_X10Y117_SLICE_X12Y117_B2 = CLBLM_L_X10Y117_SLICE_X12Y117_BQ;
  assign CLBLM_L_X10Y117_SLICE_X12Y117_B3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y117_SLICE_X12Y117_B4 = CLBLM_R_X11Y117_SLICE_X15Y117_AQ;
  assign CLBLM_L_X10Y117_SLICE_X12Y117_B5 = CLBLM_R_X11Y119_SLICE_X14Y119_AO6;
  assign CLBLM_L_X10Y117_SLICE_X12Y117_B6 = CLBLM_L_X12Y119_SLICE_X17Y119_AO5;
  assign CLBLL_L_X4Y113_SLICE_X4Y113_A6 = CLBLL_L_X4Y113_SLICE_X4Y113_CO6;
  assign CLBLL_L_X4Y113_SLICE_X4Y113_B1 = CLBLL_L_X4Y113_SLICE_X4Y113_DO6;
  assign CLBLL_L_X4Y113_SLICE_X4Y113_B2 = CLBLM_R_X5Y115_SLICE_X6Y115_BQ;
  assign CLBLM_L_X10Y117_SLICE_X12Y117_C1 = CLBLM_L_X10Y112_SLICE_X13Y112_CQ;
  assign CLBLM_L_X10Y117_SLICE_X12Y117_C2 = CLBLM_L_X10Y118_SLICE_X12Y118_BQ;
  assign CLBLM_L_X10Y117_SLICE_X12Y117_C3 = CLBLL_L_X4Y110_SLICE_X5Y110_BQ;
  assign CLBLM_L_X10Y117_SLICE_X12Y117_C4 = CLBLM_L_X10Y113_SLICE_X12Y113_AO5;
  assign CLBLM_L_X10Y117_SLICE_X12Y117_C5 = CLBLM_R_X5Y111_SLICE_X7Y111_DO6;
  assign CLBLM_L_X10Y117_SLICE_X12Y117_C6 = CLBLM_L_X10Y118_SLICE_X12Y118_AQ;
  assign CLBLL_L_X4Y113_SLICE_X4Y113_C1 = CLBLM_R_X3Y111_SLICE_X3Y111_BQ;
  assign CLBLL_L_X4Y113_SLICE_X4Y113_C2 = CLBLL_L_X4Y118_SLICE_X5Y118_AQ;
  assign CLBLM_L_X10Y117_SLICE_X12Y117_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLL_L_X4Y113_SLICE_X4Y113_C3 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLL_L_X4Y113_SLICE_X4Y113_C4 = CLBLM_R_X3Y118_SLICE_X2Y118_AQ;
  assign CLBLL_L_X4Y113_SLICE_X4Y113_C5 = CLBLM_R_X3Y112_SLICE_X3Y112_AQ;
  assign CLBLL_L_X4Y113_SLICE_X4Y113_C6 = CLBLM_R_X5Y116_SLICE_X6Y116_BQ;
  assign CLBLL_L_X4Y113_SLICE_X4Y113_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLL_L_X4Y113_SLICE_X4Y113_D1 = CLBLM_L_X8Y120_SLICE_X11Y120_CQ;
  assign CLBLM_L_X10Y117_SLICE_X12Y117_D3 = 1'b1;
  assign CLBLL_L_X4Y113_SLICE_X4Y113_D2 = CLBLL_L_X4Y111_SLICE_X4Y111_DQ;
  assign CLBLM_L_X10Y117_SLICE_X12Y117_D5 = 1'b1;
  assign CLBLM_L_X10Y117_SLICE_X12Y117_D6 = 1'b1;
  assign CLBLL_L_X4Y113_SLICE_X4Y113_D3 = RIOB33_X105Y121_IOB_X1Y121_I;
  assign CLBLL_L_X4Y113_SLICE_X4Y113_D4 = CLBLL_L_X4Y112_SLICE_X4Y112_DO6;
  assign CLBLL_L_X4Y113_SLICE_X4Y113_D5 = CLBLL_L_X4Y121_SLICE_X4Y121_AQ;
  assign CLBLL_L_X4Y113_SLICE_X4Y113_D6 = CLBLL_L_X4Y114_SLICE_X4Y114_BQ;
  assign CLBLM_L_X10Y117_SLICE_X12Y117_D4 = 1'b1;
  assign CLBLM_L_X8Y116_SLICE_X11Y116_A1 = CLBLM_L_X8Y121_SLICE_X10Y121_CQ;
  assign CLBLM_R_X37Y119_SLICE_X57Y119_B5 = 1'b1;
  assign CLBLM_R_X37Y119_SLICE_X57Y119_B6 = 1'b1;
  assign RIOI3_SING_X105Y150_OLOGIC_X1Y150_T1 = 1'b1;
  assign CLBLM_L_X8Y116_SLICE_X11Y116_A5 = 1'b1;
  assign CLBLL_L_X4Y113_SLICE_X5Y113_A1 = CLBLM_R_X5Y117_SLICE_X6Y117_BQ;
  assign CLBLL_L_X4Y113_SLICE_X5Y113_A2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLL_L_X4Y113_SLICE_X5Y113_A3 = CLBLL_L_X4Y112_SLICE_X5Y112_BO6;
  assign CLBLL_L_X4Y113_SLICE_X5Y113_A4 = CLBLL_L_X4Y113_SLICE_X5Y113_AQ;
  assign CLBLL_L_X4Y113_SLICE_X5Y113_A5 = 1'b1;
  assign CLBLL_L_X4Y113_SLICE_X5Y113_A6 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLL_L_X4Y113_SLICE_X5Y113_B1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLL_L_X4Y113_SLICE_X5Y113_B2 = CLBLL_L_X4Y113_SLICE_X5Y113_BQ;
  assign CLBLL_L_X4Y113_SLICE_X5Y113_B3 = 1'b1;
  assign CLBLL_L_X4Y113_SLICE_X5Y113_B4 = CLBLL_L_X4Y113_SLICE_X4Y113_BQ;
  assign CLBLL_L_X4Y113_SLICE_X5Y113_B5 = CLBLM_R_X11Y114_SLICE_X14Y114_D5Q;
  assign CLBLL_L_X4Y113_SLICE_X5Y113_B6 = CLBLM_R_X5Y115_SLICE_X6Y115_CO6;
  assign CLBLM_L_X8Y116_SLICE_X11Y116_AX = CLBLM_L_X8Y116_SLICE_X11Y116_CO6;
  assign CLBLM_R_X37Y119_SLICE_X57Y119_C4 = 1'b1;
  assign CLBLL_L_X4Y113_SLICE_X5Y113_C1 = 1'b1;
  assign CLBLL_L_X4Y113_SLICE_X5Y113_C2 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLL_L_X4Y113_SLICE_X5Y113_C3 = CLBLM_R_X3Y117_SLICE_X3Y117_BQ;
  assign CLBLL_L_X4Y113_SLICE_X5Y113_C4 = CLBLM_R_X5Y114_SLICE_X6Y114_CQ;
  assign CLBLL_L_X4Y113_SLICE_X5Y113_C5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLL_L_X4Y113_SLICE_X5Y113_C6 = CLBLL_L_X4Y113_SLICE_X5Y113_DO5;
  assign CLBLM_L_X8Y116_SLICE_X11Y116_B1 = 1'b1;
  assign CLBLM_R_X37Y119_SLICE_X57Y119_C5 = 1'b1;
  assign CLBLL_L_X4Y113_SLICE_X5Y113_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X37Y119_SLICE_X57Y119_C6 = 1'b1;
  assign CLBLM_L_X8Y116_SLICE_X11Y116_B2 = CLBLM_L_X8Y116_SLICE_X11Y116_BQ;
  assign CLBLM_R_X11Y120_SLICE_X14Y120_D4 = CLBLM_L_X10Y119_SLICE_X13Y119_AQ;
  assign CLBLL_L_X4Y113_SLICE_X5Y113_D1 = CLBLM_R_X5Y113_SLICE_X6Y113_AQ;
  assign CLBLL_L_X4Y113_SLICE_X5Y113_D2 = CLBLM_L_X8Y115_SLICE_X11Y115_C5Q;
  assign CLBLL_L_X4Y113_SLICE_X5Y113_D3 = CLBLM_R_X3Y113_SLICE_X2Y113_AQ;
  assign CLBLL_L_X4Y113_SLICE_X5Y113_D4 = RIOB33_X105Y121_IOB_X1Y121_I;
  assign CLBLL_L_X4Y113_SLICE_X5Y113_D5 = CLBLM_R_X3Y116_SLICE_X3Y116_BQ;
  assign CLBLL_L_X4Y113_SLICE_X5Y113_D6 = 1'b1;
  assign CLBLM_L_X8Y116_SLICE_X11Y116_B4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X11Y120_SLICE_X14Y120_D5 = CLBLM_R_X11Y120_SLICE_X14Y120_BO5;
  assign CLBLM_R_X5Y124_SLICE_X7Y124_C4 = 1'b1;
  assign CLBLM_R_X5Y124_SLICE_X7Y124_C5 = 1'b1;
  assign CLBLM_R_X5Y124_SLICE_X7Y124_C6 = 1'b1;
  assign CLBLM_R_X7Y122_SLICE_X8Y122_B5 = CLBLM_R_X7Y112_SLICE_X9Y112_CQ;
  assign CLBLM_R_X7Y122_SLICE_X8Y122_B6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y116_SLICE_X11Y116_C3 = CLBLM_R_X7Y111_SLICE_X8Y111_AQ;
  assign CLBLM_R_X37Y119_SLICE_X57Y119_D3 = 1'b1;
  assign LIOI3_X0Y173_OLOGIC_X0Y174_D1 = CLBLM_R_X7Y151_SLICE_X8Y151_AO6;
  assign CLBLM_L_X8Y116_SLICE_X11Y116_C4 = CLBLM_L_X8Y116_SLICE_X11Y116_A5Q;
  assign CLBLM_R_X37Y119_SLICE_X57Y119_D4 = 1'b1;
  assign CLBLM_R_X37Y119_SLICE_X57Y119_D5 = 1'b1;
  assign LIOB33_X0Y181_IOB_X0Y182_O = RIOB33_X105Y133_IOB_X1Y134_I;
  assign LIOB33_X0Y181_IOB_X0Y181_O = RIOB33_X105Y133_IOB_X1Y133_I;
  assign LIOI3_X0Y173_OLOGIC_X0Y174_T1 = 1'b1;
  assign CLBLM_R_X37Y119_SLICE_X57Y119_D6 = 1'b1;
  assign LIOI3_X0Y111_OLOGIC_X0Y112_D1 = CLBLM_R_X11Y114_SLICE_X14Y114_D5Q;
  assign LIOI3_X0Y173_OLOGIC_X0Y173_D1 = CLBLM_L_X8Y133_SLICE_X11Y133_AO5;
  assign LIOI3_X0Y111_OLOGIC_X0Y112_T1 = 1'b1;
  assign RIOI3_X105Y155_OLOGIC_X1Y156_D1 = RIOB33_X105Y103_IOB_X1Y104_I;
  assign LIOI3_X0Y173_OLOGIC_X0Y173_T1 = 1'b1;
  assign CLBLM_R_X7Y122_SLICE_X8Y122_C4 = CLBLM_R_X7Y122_SLICE_X8Y122_BQ;
  assign LIOI3_X0Y111_OLOGIC_X0Y111_D1 = 1'b0;
  assign CLBLM_R_X5Y124_SLICE_X7Y124_D5 = 1'b1;
  assign CLBLM_R_X7Y122_SLICE_X8Y122_C5 = 1'b1;
  assign RIOI3_X105Y155_OLOGIC_X1Y156_T1 = 1'b1;
  assign CLBLM_R_X5Y124_SLICE_X7Y124_D6 = 1'b1;
  assign CLBLM_R_X7Y122_SLICE_X8Y122_C6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign LIOI3_TBYTETERM_X0Y163_OLOGIC_X0Y164_D1 = RIOB33_X105Y111_IOB_X1Y111_I;
  assign LIOI3_X0Y111_OLOGIC_X0Y111_T1 = 1'b1;
  assign RIOI3_X105Y155_OLOGIC_X1Y155_D1 = RIOB33_X105Y103_IOB_X1Y103_I;
  assign LIOI3_TBYTETERM_X0Y163_OLOGIC_X0Y164_T1 = 1'b1;
  assign RIOI3_X105Y155_OLOGIC_X1Y155_T1 = 1'b1;
  assign LIOI3_TBYTETERM_X0Y163_OLOGIC_X0Y163_D1 = RIOB33_X105Y109_IOB_X1Y110_I;
  assign CLBLM_L_X10Y114_SLICE_X12Y114_C3 = CLBLM_L_X10Y127_SLICE_X12Y127_AQ;
  assign LIOI3_TBYTETERM_X0Y163_OLOGIC_X0Y163_T1 = 1'b1;
  assign CLBLM_L_X10Y114_SLICE_X12Y114_C6 = CLBLM_L_X10Y112_SLICE_X12Y112_AO5;
  assign CLBLM_L_X10Y118_SLICE_X13Y118_A1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y118_SLICE_X13Y118_A2 = CLBLM_L_X12Y119_SLICE_X17Y119_AO5;
  assign CLBLM_L_X10Y118_SLICE_X13Y118_A3 = CLBLM_L_X10Y118_SLICE_X13Y118_AQ;
  assign CLBLM_L_X10Y118_SLICE_X13Y118_A4 = CLBLM_L_X8Y114_SLICE_X11Y114_BQ;
  assign CLBLM_L_X10Y114_SLICE_X12Y114_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X10Y118_SLICE_X13Y118_A5 = CLBLM_R_X11Y119_SLICE_X14Y119_AO6;
  assign CLBLM_L_X10Y118_SLICE_X13Y118_A6 = CLBLM_L_X10Y120_SLICE_X12Y120_CQ;
  assign CLBLM_R_X5Y124_SLICE_X6Y124_A6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y118_SLICE_X13Y118_B1 = CLBLM_L_X12Y119_SLICE_X17Y119_AO5;
  assign CLBLM_L_X10Y118_SLICE_X13Y118_B2 = CLBLM_L_X10Y118_SLICE_X13Y118_BQ;
  assign CLBLM_L_X10Y118_SLICE_X13Y118_B3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y118_SLICE_X13Y118_B4 = CLBLM_L_X10Y117_SLICE_X12Y117_BQ;
  assign CLBLM_L_X10Y118_SLICE_X13Y118_B5 = CLBLM_R_X11Y119_SLICE_X14Y119_AO6;
  assign CLBLM_L_X10Y118_SLICE_X13Y118_B6 = CLBLM_R_X7Y117_SLICE_X8Y117_CQ;
  assign CLBLM_L_X10Y118_SLICE_X13Y118_C1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y118_SLICE_X13Y118_C2 = CLBLL_L_X4Y110_SLICE_X4Y110_CQ;
  assign CLBLM_L_X10Y118_SLICE_X13Y118_C3 = CLBLM_L_X10Y116_SLICE_X13Y116_BO5;
  assign CLBLM_L_X10Y118_SLICE_X13Y118_C4 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X10Y118_SLICE_X13Y118_C5 = 1'b1;
  assign CLBLM_L_X10Y118_SLICE_X13Y118_C6 = CLBLM_L_X8Y122_SLICE_X11Y122_AQ;
  assign CLBLM_L_X10Y118_SLICE_X13Y118_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_CE0 = 1'b1;
  assign CLBLM_L_X10Y118_SLICE_X13Y118_D1 = CLBLM_L_X10Y115_SLICE_X13Y115_CO6;
  assign CLBLM_L_X10Y118_SLICE_X13Y118_D2 = CLBLM_R_X11Y113_SLICE_X15Y113_CO6;
  assign CLBLM_L_X10Y118_SLICE_X13Y118_D3 = CLBLM_R_X7Y118_SLICE_X8Y118_BQ;
  assign CLBLM_L_X10Y118_SLICE_X13Y118_D4 = CLBLM_R_X7Y123_SLICE_X9Y123_CO6;
  assign CLBLM_L_X10Y118_SLICE_X13Y118_D5 = CLBLM_R_X11Y119_SLICE_X14Y119_BO5;
  assign CLBLM_L_X10Y118_SLICE_X13Y118_D6 = CLBLM_L_X10Y113_SLICE_X13Y113_CO6;
  assign CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_CE1 = 1'b1;
  assign CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_IGNORE0 = 1'b1;
  assign CLBLM_L_X8Y116_SLICE_X10Y116_A5 = CLBLM_L_X10Y114_SLICE_X13Y114_DQ;
  assign CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_IGNORE1 = 1'b1;
  assign CLBLL_L_X4Y114_SLICE_X4Y114_A1 = CLBLM_R_X3Y115_SLICE_X3Y115_DQ;
  assign CLBLL_L_X4Y114_SLICE_X4Y114_A2 = CLBLM_R_X5Y115_SLICE_X6Y115_CO6;
  assign CLBLM_L_X10Y118_SLICE_X12Y118_A1 = 1'b1;
  assign CLBLM_L_X10Y118_SLICE_X12Y118_A2 = CLBLM_L_X10Y117_SLICE_X12Y117_CO6;
  assign CLBLM_L_X10Y118_SLICE_X12Y118_A3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y118_SLICE_X12Y118_A4 = RIOB33_X105Y141_IOB_X1Y142_I;
  assign CLBLM_L_X10Y118_SLICE_X12Y118_A5 = CLBLM_R_X7Y128_SLICE_X8Y128_AQ;
  assign CLBLM_L_X10Y118_SLICE_X12Y118_A6 = CLBLM_L_X8Y119_SLICE_X11Y119_CQ;
  assign CLBLL_L_X4Y114_SLICE_X4Y114_A3 = CLBLL_L_X4Y114_SLICE_X4Y114_AQ;
  assign CLBLL_L_X4Y114_SLICE_X4Y114_A4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLL_L_X4Y114_SLICE_X4Y114_A5 = CLBLL_L_X4Y111_SLICE_X4Y111_BQ;
  assign CLBLL_L_X4Y114_SLICE_X4Y114_A6 = 1'b1;
  assign CLBLM_L_X10Y118_SLICE_X12Y118_B1 = CLBLM_L_X10Y123_SLICE_X13Y123_BO6;
  assign CLBLM_L_X10Y118_SLICE_X12Y118_B2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y118_SLICE_X12Y118_B3 = CLBLM_R_X5Y110_SLICE_X7Y110_BQ;
  assign CLBLM_L_X10Y118_SLICE_X12Y118_B4 = 1'b1;
  assign CLBLM_L_X10Y118_SLICE_X12Y118_B5 = CLBLM_L_X10Y116_SLICE_X12Y116_A5Q;
  assign CLBLL_L_X4Y114_SLICE_X4Y114_B1 = CLBLL_L_X4Y115_SLICE_X4Y115_CQ;
  assign CLBLL_L_X4Y114_SLICE_X4Y114_B2 = CLBLL_L_X4Y114_SLICE_X4Y114_BQ;
  assign CLBLL_L_X4Y114_SLICE_X4Y114_B3 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLL_L_X4Y114_SLICE_X4Y114_B4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLL_L_X4Y114_SLICE_X4Y114_B5 = 1'b1;
  assign CLBLL_L_X4Y114_SLICE_X4Y114_B6 = CLBLL_L_X4Y113_SLICE_X5Y113_CQ;
  assign CLBLL_L_X4Y114_SLICE_X4Y114_C1 = CLBLM_L_X10Y113_SLICE_X13Y113_BO6;
  assign CLBLL_L_X4Y114_SLICE_X4Y114_C2 = CLBLL_L_X4Y114_SLICE_X4Y114_CQ;
  assign CLBLL_L_X4Y114_SLICE_X4Y114_C3 = CLBLL_L_X4Y113_SLICE_X4Y113_AQ;
  assign CLBLM_L_X10Y118_SLICE_X12Y118_C5 = CLBLM_L_X10Y118_SLICE_X12Y118_DO6;
  assign CLBLM_L_X10Y118_SLICE_X12Y118_C6 = CLBLM_R_X7Y119_SLICE_X9Y119_BQ;
  assign CLBLL_L_X4Y114_SLICE_X4Y114_C4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLL_L_X4Y114_SLICE_X4Y114_C5 = CLBLM_R_X7Y119_SLICE_X8Y119_D5Q;
  assign CLBLL_L_X4Y114_SLICE_X4Y114_C6 = CLBLL_L_X4Y116_SLICE_X4Y116_BQ;
  assign CLBLM_L_X10Y118_SLICE_X12Y118_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLL_L_X4Y114_SLICE_X4Y114_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X10Y118_SLICE_X12Y118_C3 = CLBLM_L_X10Y119_SLICE_X12Y119_DO6;
  assign CLBLL_L_X4Y114_SLICE_X4Y114_D1 = CLBLL_L_X4Y114_SLICE_X5Y114_AQ;
  assign CLBLL_L_X4Y114_SLICE_X4Y114_D2 = CLBLM_R_X5Y114_SLICE_X7Y114_AQ;
  assign CLBLL_L_X4Y114_SLICE_X4Y114_D3 = RIOB33_X105Y121_IOB_X1Y121_I;
  assign CLBLL_L_X4Y114_SLICE_X4Y114_D4 = CLBLM_R_X5Y114_SLICE_X7Y114_BO5;
  assign CLBLL_L_X4Y114_SLICE_X4Y114_D5 = CLBLL_L_X4Y116_SLICE_X4Y116_BQ;
  assign CLBLL_L_X4Y114_SLICE_X4Y114_D6 = CLBLM_R_X7Y120_SLICE_X9Y120_CQ;
  assign CLBLM_L_X10Y118_SLICE_X12Y118_D1 = 1'b1;
  assign CLBLM_L_X10Y114_SLICE_X12Y114_SR = CLBLM_R_X11Y123_SLICE_X14Y123_CO6;
  assign CLBLM_L_X10Y118_SLICE_X12Y118_D2 = 1'b1;
  assign CLBLM_L_X10Y118_SLICE_X12Y118_D3 = CLBLM_L_X8Y119_SLICE_X11Y119_BQ;
  assign CLBLM_L_X10Y118_SLICE_X12Y118_D4 = CLBLM_L_X10Y118_SLICE_X13Y118_CQ;
  assign CLBLM_L_X10Y118_SLICE_X12Y118_D5 = CLBLM_L_X10Y119_SLICE_X12Y119_CQ;
  assign CLBLM_L_X10Y118_SLICE_X12Y118_D6 = CLBLM_L_X10Y116_SLICE_X12Y116_CQ;
  assign CLBLM_R_X5Y124_SLICE_X6Y124_C4 = CLBLM_R_X5Y125_SLICE_X6Y125_BO5;
  assign CLBLM_R_X103Y172_SLICE_X162Y172_D5 = 1'b1;
  assign CLBLM_R_X5Y124_SLICE_X6Y124_C5 = CLBLM_R_X5Y116_SLICE_X6Y116_BQ;
  assign CLBLL_L_X4Y114_SLICE_X5Y114_A1 = CLBLL_L_X4Y115_SLICE_X5Y115_CQ;
  assign CLBLL_L_X4Y114_SLICE_X5Y114_A2 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLL_L_X4Y114_SLICE_X5Y114_A3 = 1'b1;
  assign CLBLL_L_X4Y114_SLICE_X5Y114_A4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLL_L_X4Y114_SLICE_X5Y114_A5 = 1'b1;
  assign CLBLL_L_X4Y114_SLICE_X5Y114_A6 = CLBLM_R_X3Y114_SLICE_X2Y114_DQ;
  assign CLBLM_R_X5Y124_SLICE_X6Y124_C6 = CLBLM_R_X5Y123_SLICE_X6Y123_AQ;
  assign CLBLM_R_X7Y112_SLICE_X9Y112_A5 = CLBLM_R_X7Y112_SLICE_X8Y112_AQ;
  assign CLBLL_L_X4Y114_SLICE_X5Y114_B1 = CLBLM_R_X5Y121_SLICE_X6Y121_AQ;
  assign CLBLL_L_X4Y114_SLICE_X5Y114_B2 = CLBLM_R_X5Y115_SLICE_X6Y115_BQ;
  assign CLBLL_L_X4Y114_SLICE_X5Y114_B3 = RIOB33_X105Y121_IOB_X1Y121_I;
  assign CLBLL_L_X4Y114_SLICE_X5Y114_B4 = CLBLM_R_X7Y114_SLICE_X8Y114_BQ;
  assign CLBLL_L_X4Y114_SLICE_X5Y114_B5 = 1'b1;
  assign CLBLL_L_X4Y114_SLICE_X5Y114_B6 = 1'b1;
  assign LIOI3_X0Y51_ILOGIC_X0Y52_D = LIOB33_X0Y51_IOB_X0Y52_I;
  assign CLBLM_R_X103Y172_SLICE_X162Y172_D6 = 1'b1;
  assign CLBLL_L_X4Y114_SLICE_X5Y114_C1 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLL_L_X4Y114_SLICE_X5Y114_C2 = CLBLM_R_X7Y119_SLICE_X9Y119_AQ;
  assign CLBLL_L_X4Y114_SLICE_X5Y114_C3 = CLBLM_L_X8Y120_SLICE_X10Y120_BQ;
  assign CLBLL_L_X4Y114_SLICE_X5Y114_C4 = CLBLM_R_X5Y121_SLICE_X6Y121_AQ;
  assign CLBLL_L_X4Y114_SLICE_X5Y114_C5 = CLBLL_L_X4Y114_SLICE_X5Y114_BO5;
  assign CLBLL_L_X4Y114_SLICE_X5Y114_C6 = CLBLL_L_X4Y112_SLICE_X5Y112_AQ;
  assign CLBLM_L_X8Y116_SLICE_X10Y116_C3 = CLBLL_L_X4Y119_SLICE_X4Y119_CQ;
  assign CLBLL_L_X4Y114_SLICE_X5Y114_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign LIOI3_X0Y51_ILOGIC_X0Y51_D = LIOB33_X0Y51_IOB_X0Y51_I;
  assign RIOB33_X105Y151_IOB_X1Y151_O = LIOB33_X0Y75_IOB_X0Y76_I;
  assign RIOB33_X105Y151_IOB_X1Y152_O = RIOB33_SING_X105Y100_IOB_X1Y100_I;
  assign RIOI3_SING_X105Y199_OLOGIC_X1Y199_D1 = CLBLM_R_X11Y128_SLICE_X15Y128_AQ;
  assign CLBLL_L_X4Y114_SLICE_X5Y114_D1 = CLBLL_L_X4Y116_SLICE_X5Y116_DQ;
  assign CLBLL_L_X4Y114_SLICE_X5Y114_D2 = CLBLL_L_X4Y113_SLICE_X5Y113_CQ;
  assign CLBLL_L_X4Y114_SLICE_X5Y114_D3 = CLBLM_R_X5Y116_SLICE_X6Y116_DQ;
  assign CLBLL_L_X4Y114_SLICE_X5Y114_D4 = 1'b1;
  assign CLBLL_L_X4Y114_SLICE_X5Y114_D5 = 1'b1;
  assign CLBLL_L_X4Y114_SLICE_X5Y114_D6 = CLBLL_L_X4Y112_SLICE_X4Y112_BQ;
  assign CLBLM_R_X7Y112_SLICE_X9Y112_B1 = CLBLM_R_X7Y128_SLICE_X8Y128_AQ;
  assign CLBLM_R_X7Y112_SLICE_X9Y112_B2 = CLBLM_L_X8Y112_SLICE_X11Y112_CO6;
  assign LIOI3_TBYTESRC_X0Y57_ILOGIC_X0Y58_D = LIOB33_X0Y57_IOB_X0Y58_I;
  assign LIOI3_TBYTESRC_X0Y57_ILOGIC_X0Y57_D = LIOB33_X0Y57_IOB_X0Y57_I;
  assign CLBLM_R_X7Y112_SLICE_X9Y112_B5 = RIOB33_X105Y141_IOB_X1Y142_I;
  assign LIOB33_X0Y183_IOB_X0Y184_O = RIOB33_X105Y135_IOB_X1Y136_I;
  assign LIOB33_X0Y183_IOB_X0Y183_O = RIOB33_X105Y135_IOB_X1Y135_I;
  assign CLBLM_L_X8Y116_SLICE_X10Y116_SR = CLBLM_R_X11Y123_SLICE_X14Y123_CO6;
  assign RIOI3_X105Y161_OLOGIC_X1Y162_D1 = CLBLM_R_X11Y117_SLICE_X14Y117_DO6;
  assign CLBLL_L_X4Y122_SLICE_X4Y122_B1 = LIOB33_X0Y65_IOB_X0Y65_I;
  assign CLBLL_L_X4Y122_SLICE_X4Y122_B2 = CLBLL_L_X2Y121_SLICE_X1Y121_BO6;
  assign CLBLL_L_X4Y122_SLICE_X4Y122_B3 = CLBLM_L_X8Y120_SLICE_X10Y120_D5Q;
  assign CLBLL_L_X4Y122_SLICE_X4Y122_B4 = RIOB33_X105Y129_IOB_X1Y129_I;
  assign CLBLL_L_X4Y122_SLICE_X4Y122_B5 = CLBLM_R_X3Y124_SLICE_X2Y124_AO5;
  assign CLBLM_L_X10Y119_SLICE_X13Y119_A1 = RIOB33_X105Y121_IOB_X1Y121_I;
  assign CLBLM_L_X10Y119_SLICE_X13Y119_A2 = CLBLM_R_X7Y120_SLICE_X9Y120_D5Q;
  assign CLBLM_L_X10Y119_SLICE_X13Y119_A3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y119_SLICE_X13Y119_A4 = CLBLM_L_X10Y119_SLICE_X13Y119_AQ;
  assign CLBLM_L_X10Y119_SLICE_X13Y119_A5 = CLBLM_L_X12Y120_SLICE_X16Y120_AO6;
  assign CLBLM_L_X10Y119_SLICE_X13Y119_A6 = CLBLM_R_X11Y118_SLICE_X14Y118_BQ;
  assign RIOI3_X105Y171_OLOGIC_X1Y172_T1 = 1'b1;
  assign CLBLL_L_X4Y122_SLICE_X4Y122_C1 = RIOB33_X105Y109_IOB_X1Y110_I;
  assign CLBLM_L_X10Y119_SLICE_X13Y119_B1 = 1'b1;
  assign CLBLM_L_X10Y119_SLICE_X13Y119_B2 = CLBLM_L_X8Y119_SLICE_X10Y119_BQ;
  assign CLBLM_L_X10Y119_SLICE_X13Y119_B3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y119_SLICE_X13Y119_B4 = CLBLM_L_X12Y120_SLICE_X17Y120_CO6;
  assign CLBLM_L_X10Y119_SLICE_X13Y119_B5 = CLBLM_R_X7Y113_SLICE_X9Y113_A5Q;
  assign CLBLM_L_X10Y119_SLICE_X13Y119_B6 = 1'b1;
  assign CLBLL_L_X4Y122_SLICE_X4Y122_C3 = CLBLL_L_X2Y122_SLICE_X0Y122_AO6;
  assign CLBLM_L_X10Y119_SLICE_X13Y119_C1 = CLBLM_R_X13Y119_SLICE_X18Y119_CQ;
  assign CLBLM_L_X10Y119_SLICE_X13Y119_C2 = CLBLM_L_X10Y119_SLICE_X13Y119_AQ;
  assign CLBLM_L_X10Y119_SLICE_X13Y119_C3 = CLBLM_L_X10Y119_SLICE_X13Y119_BQ;
  assign CLBLM_L_X10Y119_SLICE_X13Y119_C4 = CLBLM_R_X11Y118_SLICE_X14Y118_BQ;
  assign CLBLM_L_X10Y119_SLICE_X13Y119_C5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y119_SLICE_X13Y119_C6 = CLBLM_R_X11Y119_SLICE_X15Y119_CQ;
  assign CLBLL_L_X4Y122_SLICE_X4Y122_C4 = CLBLL_L_X4Y121_SLICE_X5Y121_DO6;
  assign CLBLM_L_X10Y119_SLICE_X13Y119_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLL_L_X4Y122_SLICE_X4Y122_C5 = CLBLM_R_X3Y123_SLICE_X3Y123_BO5;
  assign CLBLL_L_X4Y122_SLICE_X4Y122_C6 = CLBLL_L_X4Y122_SLICE_X4Y122_BO6;
  assign CLBLM_L_X10Y119_SLICE_X13Y119_D1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y119_SLICE_X13Y119_D2 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X10Y119_SLICE_X13Y119_D3 = CLBLM_L_X10Y114_SLICE_X13Y114_BO5;
  assign CLBLM_L_X10Y119_SLICE_X13Y119_D4 = CLBLM_L_X10Y119_SLICE_X13Y119_BQ;
  assign CLBLM_L_X10Y119_SLICE_X13Y119_D5 = CLBLL_L_X4Y117_SLICE_X5Y117_DQ;
  assign CLBLM_L_X10Y119_SLICE_X13Y119_D6 = 1'b1;
  assign CLBLL_L_X4Y115_SLICE_X4Y115_A1 = CLBLM_R_X5Y115_SLICE_X6Y115_CO5;
  assign CLBLL_L_X4Y115_SLICE_X4Y115_A2 = CLBLL_L_X4Y115_SLICE_X4Y115_DQ;
  assign CLBLL_L_X4Y115_SLICE_X4Y115_A3 = CLBLL_L_X4Y115_SLICE_X4Y115_AQ;
  assign CLBLL_L_X4Y115_SLICE_X4Y115_A4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLL_L_X4Y115_SLICE_X4Y115_A5 = CLBLL_L_X4Y111_SLICE_X4Y111_AQ;
  assign CLBLL_L_X4Y115_SLICE_X4Y115_A6 = 1'b1;
  assign CLBLM_L_X10Y119_SLICE_X12Y119_A1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y119_SLICE_X12Y119_A2 = CLBLM_L_X10Y119_SLICE_X12Y119_BQ;
  assign CLBLL_L_X4Y115_SLICE_X4Y115_B1 = 1'b1;
  assign CLBLL_L_X4Y115_SLICE_X4Y115_B2 = CLBLL_L_X4Y115_SLICE_X4Y115_DQ;
  assign CLBLM_L_X10Y119_SLICE_X12Y119_A6 = CLBLM_R_X5Y115_SLICE_X7Y115_DO6;
  assign CLBLL_L_X4Y115_SLICE_X4Y115_B3 = CLBLL_L_X2Y115_SLICE_X1Y115_AQ;
  assign CLBLL_L_X4Y115_SLICE_X4Y115_B4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLL_L_X4Y115_SLICE_X4Y115_B5 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLL_L_X4Y115_SLICE_X4Y115_B6 = 1'b1;
  assign CLBLM_L_X10Y119_SLICE_X12Y119_A3 = CLBLM_L_X10Y119_SLICE_X12Y119_AQ;
  assign CLBLM_L_X10Y119_SLICE_X12Y119_A4 = CLBLM_R_X3Y118_SLICE_X2Y118_AQ;
  assign CLBLL_L_X4Y115_SLICE_X4Y115_C1 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLL_L_X4Y115_SLICE_X4Y115_C2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLL_L_X4Y115_SLICE_X4Y115_C3 = CLBLM_R_X5Y117_SLICE_X6Y117_BQ;
  assign CLBLL_L_X4Y115_SLICE_X4Y115_C4 = CLBLM_L_X8Y115_SLICE_X10Y115_CQ;
  assign CLBLL_L_X4Y115_SLICE_X4Y115_C5 = CLBLM_R_X3Y115_SLICE_X2Y115_AQ;
  assign CLBLL_L_X4Y115_SLICE_X4Y115_C6 = 1'b1;
  assign CLBLM_L_X10Y119_SLICE_X12Y119_B1 = CLBLM_L_X8Y120_SLICE_X11Y120_BQ;
  assign CLBLM_L_X10Y119_SLICE_X12Y119_B2 = CLBLM_L_X10Y119_SLICE_X12Y119_BQ;
  assign CLBLM_L_X10Y119_SLICE_X12Y119_C1 = CLBLM_L_X8Y119_SLICE_X11Y119_BQ;
  assign CLBLM_L_X10Y119_SLICE_X12Y119_C2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y119_SLICE_X12Y119_C3 = CLBLM_R_X7Y114_SLICE_X8Y114_BQ;
  assign CLBLL_L_X4Y115_SLICE_X4Y115_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X10Y119_SLICE_X12Y119_C6 = CLBLM_L_X8Y119_SLICE_X10Y119_DO5;
  assign CLBLL_L_X4Y115_SLICE_X4Y115_D1 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLL_L_X4Y115_SLICE_X4Y115_D2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLL_L_X4Y115_SLICE_X4Y115_D3 = 1'b1;
  assign CLBLL_L_X4Y115_SLICE_X4Y115_D4 = CLBLM_R_X5Y115_SLICE_X6Y115_BQ;
  assign CLBLL_L_X4Y115_SLICE_X4Y115_D5 = 1'b1;
  assign CLBLL_L_X4Y115_SLICE_X4Y115_D6 = CLBLM_R_X3Y115_SLICE_X3Y115_AQ;
  assign CLBLM_L_X10Y119_SLICE_X12Y119_C5 = 1'b1;
  assign CLBLM_L_X10Y119_SLICE_X12Y119_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X10Y119_SLICE_X12Y119_D1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y119_SLICE_X12Y119_D2 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X10Y119_SLICE_X12Y119_D3 = RIOB33_X105Y121_IOB_X1Y121_I;
  assign CLBLM_L_X10Y119_SLICE_X12Y119_D4 = CLBLM_L_X8Y119_SLICE_X11Y119_CQ;
  assign CLBLM_L_X10Y119_SLICE_X12Y119_D5 = CLBLM_R_X7Y114_SLICE_X8Y114_BQ;
  assign CLBLM_L_X10Y119_SLICE_X12Y119_D6 = CLBLM_R_X13Y119_SLICE_X18Y119_BQ;
  assign CLBLL_L_X4Y122_SLICE_X4Y122_D1 = CLBLL_L_X4Y122_SLICE_X4Y122_AO6;
  assign CLBLL_L_X4Y122_SLICE_X4Y122_D2 = CLBLM_R_X5Y122_SLICE_X7Y122_CQ;
  assign CLBLL_L_X4Y122_SLICE_X4Y122_D3 = RIOB33_X105Y131_IOB_X1Y131_I;
  assign CLBLL_L_X4Y122_SLICE_X4Y122_D4 = 1'b1;
  assign CLBLL_L_X4Y122_SLICE_X4Y122_D5 = CLBLM_R_X3Y124_SLICE_X2Y124_AO5;
  assign CLBLL_L_X4Y122_SLICE_X4Y122_D6 = CLBLM_R_X5Y122_SLICE_X6Y122_BQ;
  assign RIOB33_X105Y153_IOB_X1Y154_O = RIOB33_X105Y101_IOB_X1Y102_I;
  assign CLBLL_L_X4Y115_SLICE_X5Y115_A1 = CLBLL_L_X4Y113_SLICE_X4Y113_DO6;
  assign CLBLL_L_X4Y115_SLICE_X5Y115_A2 = CLBLM_R_X11Y116_SLICE_X14Y116_CQ;
  assign CLBLL_L_X4Y115_SLICE_X5Y115_A3 = CLBLL_L_X4Y115_SLICE_X5Y115_AQ;
  assign CLBLL_L_X4Y115_SLICE_X5Y115_A4 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLL_L_X4Y115_SLICE_X5Y115_A5 = CLBLM_R_X3Y118_SLICE_X2Y118_AQ;
  assign CLBLL_L_X4Y115_SLICE_X5Y115_A6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign RIOB33_X105Y153_IOB_X1Y153_O = RIOB33_X105Y101_IOB_X1Y101_I;
  assign CLBLL_L_X4Y115_SLICE_X5Y115_B1 = CLBLL_L_X4Y113_SLICE_X5Y113_DO6;
  assign CLBLL_L_X4Y115_SLICE_X5Y115_B2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLL_L_X4Y115_SLICE_X5Y115_B3 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLL_L_X4Y115_SLICE_X5Y115_B4 = CLBLL_L_X4Y115_SLICE_X4Y115_DQ;
  assign CLBLL_L_X4Y115_SLICE_X5Y115_B5 = 1'b1;
  assign CLBLL_L_X4Y115_SLICE_X5Y115_B6 = CLBLM_R_X5Y116_SLICE_X6Y116_DQ;
  assign CLBLL_L_X4Y115_SLICE_X5Y115_C1 = CLBLM_R_X5Y115_SLICE_X7Y115_AQ;
  assign CLBLL_L_X4Y115_SLICE_X5Y115_C2 = CLBLM_R_X7Y118_SLICE_X9Y118_CQ;
  assign CLBLL_L_X4Y115_SLICE_X5Y115_C3 = 1'b1;
  assign CLBLL_L_X4Y115_SLICE_X5Y115_C4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLL_L_X4Y115_SLICE_X5Y115_C5 = 1'b1;
  assign CLBLL_L_X4Y115_SLICE_X5Y115_C6 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLL_L_X4Y115_SLICE_X5Y115_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLL_L_X4Y115_SLICE_X5Y115_D1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLL_L_X4Y115_SLICE_X5Y115_D2 = CLBLM_L_X10Y113_SLICE_X13Y113_BO6;
  assign CLBLL_L_X4Y115_SLICE_X5Y115_D3 = CLBLL_L_X4Y115_SLICE_X5Y115_DQ;
  assign CLBLL_L_X4Y115_SLICE_X5Y115_D4 = CLBLM_R_X3Y115_SLICE_X2Y115_BQ;
  assign CLBLL_L_X4Y115_SLICE_X5Y115_D5 = CLBLL_L_X4Y111_SLICE_X5Y111_AQ;
  assign CLBLL_L_X4Y115_SLICE_X5Y115_D6 = CLBLM_R_X7Y119_SLICE_X8Y119_D5Q;
  assign CLBLM_R_X11Y113_SLICE_X15Y113_A1 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X11Y113_SLICE_X15Y113_A2 = CLBLM_L_X10Y113_SLICE_X12Y113_DO6;
  assign CLBLM_R_X11Y113_SLICE_X15Y113_A3 = CLBLM_R_X11Y113_SLICE_X15Y113_AQ;
  assign CLBLM_R_X11Y113_SLICE_X15Y113_B1 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X11Y113_SLICE_X15Y113_B2 = CLBLM_R_X11Y113_SLICE_X15Y113_BQ;
  assign CLBLM_R_X11Y113_SLICE_X15Y113_B3 = CLBLM_L_X12Y115_SLICE_X16Y115_AQ;
  assign CLBLM_R_X11Y113_SLICE_X15Y113_B4 = CLBLM_L_X10Y113_SLICE_X12Y113_DO6;
  assign CLBLM_R_X11Y113_SLICE_X15Y113_B5 = CLBLM_L_X10Y113_SLICE_X13Y113_AO6;
  assign CLBLM_R_X11Y113_SLICE_X15Y113_B6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign LIOB33_X0Y185_IOB_X0Y185_O = RIOB33_X105Y137_IOB_X1Y137_I;
  assign LIOB33_X0Y185_IOB_X0Y186_O = RIOB33_X105Y143_IOB_X1Y143_I;
  assign CLBLM_R_X11Y113_SLICE_X15Y113_C1 = 1'b1;
  assign CLBLM_R_X11Y113_SLICE_X15Y113_C2 = CLBLM_L_X8Y113_SLICE_X11Y113_AQ;
  assign CLBLM_R_X11Y113_SLICE_X15Y113_C3 = 1'b1;
  assign CLBLM_R_X11Y113_SLICE_X15Y113_C4 = CLBLM_L_X8Y112_SLICE_X10Y112_BQ;
  assign CLBLM_R_X11Y113_SLICE_X15Y113_C5 = CLBLM_R_X11Y113_SLICE_X15Y113_AQ;
  assign CLBLM_R_X11Y113_SLICE_X15Y113_C6 = 1'b1;
  assign CLBLM_R_X11Y113_SLICE_X15Y113_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X11Y113_SLICE_X15Y113_D1 = CLBLM_L_X10Y112_SLICE_X12Y112_BQ;
  assign CLBLM_R_X11Y113_SLICE_X15Y113_D2 = 1'b1;
  assign CLBLM_R_X11Y113_SLICE_X15Y113_D3 = 1'b1;
  assign CLBLM_R_X11Y113_SLICE_X15Y113_D4 = CLBLM_R_X5Y109_SLICE_X7Y109_AQ;
  assign CLBLM_R_X11Y113_SLICE_X15Y113_D5 = 1'b1;
  assign CLBLM_R_X11Y113_SLICE_X15Y113_D6 = CLBLM_R_X3Y117_SLICE_X3Y117_BQ;
  assign RIOI3_TBYTESRC_X105Y119_ILOGIC_X1Y119_D = RIOB33_X105Y119_IOB_X1Y119_I;
  assign LIOI3_X0Y123_OLOGIC_X0Y124_D1 = CLBLL_L_X4Y116_SLICE_X4Y116_C5Q;
  assign CLBLM_R_X11Y113_SLICE_X14Y113_A1 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X11Y113_SLICE_X14Y113_A2 = CLBLM_L_X8Y112_SLICE_X10Y112_AQ;
  assign CLBLM_R_X11Y113_SLICE_X14Y113_A3 = CLBLM_R_X11Y113_SLICE_X14Y113_AQ;
  assign CLBLM_R_X11Y113_SLICE_X14Y113_A4 = CLBLM_L_X10Y113_SLICE_X12Y113_DO6;
  assign CLBLM_R_X11Y113_SLICE_X14Y113_A5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X11Y113_SLICE_X14Y113_A6 = CLBLM_L_X10Y121_SLICE_X13Y121_AQ;
  assign CLBLM_R_X11Y113_SLICE_X14Y113_B1 = CLBLM_R_X11Y114_SLICE_X14Y114_CQ;
  assign CLBLM_R_X11Y113_SLICE_X14Y113_B2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X11Y113_SLICE_X14Y113_B3 = 1'b1;
  assign CLBLM_R_X11Y113_SLICE_X14Y113_B4 = RIOB33_X105Y141_IOB_X1Y142_I;
  assign CLBLM_R_X11Y113_SLICE_X14Y113_B5 = CLBLM_R_X7Y128_SLICE_X8Y128_AQ;
  assign CLBLM_R_X11Y113_SLICE_X14Y113_B6 = CLBLM_R_X11Y113_SLICE_X14Y113_CO6;
  assign CLBLM_R_X11Y120_SLICE_X14Y120_C6 = CLBLM_L_X10Y120_SLICE_X12Y120_DQ;
  assign CLBLM_R_X11Y113_SLICE_X14Y113_C1 = CLBLM_R_X11Y113_SLICE_X14Y113_BQ;
  assign CLBLM_R_X11Y113_SLICE_X14Y113_C2 = CLBLM_R_X5Y111_SLICE_X7Y111_DO6;
  assign CLBLM_R_X11Y113_SLICE_X14Y113_C3 = CLBLM_L_X10Y122_SLICE_X13Y122_A5Q;
  assign CLBLM_R_X11Y113_SLICE_X14Y113_C4 = CLBLM_L_X10Y112_SLICE_X13Y112_CQ;
  assign CLBLM_R_X11Y113_SLICE_X14Y113_C5 = CLBLM_L_X10Y113_SLICE_X12Y113_AO5;
  assign CLBLM_R_X11Y113_SLICE_X14Y113_C6 = CLBLM_R_X11Y117_SLICE_X14Y117_BQ;
  assign CLBLM_R_X11Y113_SLICE_X14Y113_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X11Y113_SLICE_X14Y113_D1 = CLBLM_L_X8Y113_SLICE_X11Y113_BQ;
  assign CLBLM_R_X11Y113_SLICE_X14Y113_D2 = 1'b1;
  assign CLBLM_R_X11Y113_SLICE_X14Y113_D3 = CLBLM_L_X10Y112_SLICE_X13Y112_BQ;
  assign CLBLM_R_X11Y113_SLICE_X14Y113_D4 = CLBLM_L_X8Y111_SLICE_X10Y111_AQ;
  assign CLBLM_R_X11Y113_SLICE_X14Y113_D5 = CLBLM_R_X11Y114_SLICE_X14Y114_CQ;
  assign CLBLM_R_X11Y113_SLICE_X14Y113_D6 = 1'b1;
  assign LIOI3_X0Y123_OLOGIC_X0Y124_T1 = 1'b1;
  assign CLBLL_L_X4Y122_SLICE_X5Y122_A4 = CLBLL_L_X4Y123_SLICE_X5Y123_AO5;
  assign CLBLL_L_X4Y122_SLICE_X5Y122_A5 = CLBLM_R_X3Y124_SLICE_X2Y124_BO6;
  assign CLBLL_L_X4Y122_SLICE_X5Y122_A6 = CLBLM_R_X3Y122_SLICE_X3Y122_AO5;
  assign LIOI3_X0Y123_OLOGIC_X0Y123_D1 = CLBLM_R_X5Y117_SLICE_X6Y117_D5Q;
  assign CLBLM_L_X10Y120_SLICE_X13Y120_A1 = CLBLM_L_X10Y121_SLICE_X13Y121_DO6;
  assign CLBLM_L_X10Y120_SLICE_X13Y120_A2 = CLBLM_L_X10Y124_SLICE_X13Y124_BO5;
  assign CLBLM_L_X10Y120_SLICE_X13Y120_A3 = 1'b1;
  assign CLBLM_L_X10Y120_SLICE_X13Y120_A4 = CLBLL_L_X2Y113_SLICE_X1Y113_AQ;
  assign CLBLM_L_X10Y120_SLICE_X13Y120_A5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y120_SLICE_X13Y120_A6 = CLBLM_L_X10Y124_SLICE_X13Y124_AO5;
  assign RIOB33_X105Y187_IOB_X1Y187_O = CLBLM_L_X10Y114_SLICE_X12Y114_AQ;
  assign RIOB33_X105Y187_IOB_X1Y188_O = CLBLM_R_X11Y122_SLICE_X14Y122_AQ;
  assign CLBLM_L_X10Y120_SLICE_X13Y120_AX = CLBLM_L_X8Y118_SLICE_X11Y118_BO6;
  assign CLBLM_L_X10Y120_SLICE_X13Y120_B1 = CLBLM_L_X10Y120_SLICE_X13Y120_DO6;
  assign CLBLM_L_X10Y120_SLICE_X13Y120_B2 = CLBLM_L_X10Y124_SLICE_X13Y124_BO5;
  assign CLBLM_L_X10Y120_SLICE_X13Y120_B3 = 1'b1;
  assign CLBLM_L_X10Y120_SLICE_X13Y120_B4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y120_SLICE_X13Y120_B5 = CLBLM_R_X3Y112_SLICE_X3Y112_AQ;
  assign CLBLM_L_X10Y120_SLICE_X13Y120_B6 = CLBLM_L_X10Y124_SLICE_X13Y124_AO5;
  assign LIOI3_X0Y175_OLOGIC_X0Y176_D1 = RIOB33_X105Y127_IOB_X1Y128_I;
  assign CLBLM_L_X8Y110_SLICE_X11Y110_A1 = 1'b1;
  assign CLBLM_L_X8Y110_SLICE_X11Y110_A2 = 1'b1;
  assign CLBLM_L_X8Y110_SLICE_X11Y110_A3 = 1'b1;
  assign CLBLM_L_X8Y110_SLICE_X11Y110_A4 = 1'b1;
  assign CLBLM_L_X8Y110_SLICE_X11Y110_A5 = 1'b1;
  assign CLBLM_L_X8Y110_SLICE_X11Y110_A6 = 1'b1;
  assign CLBLM_L_X10Y120_SLICE_X13Y120_C1 = CLBLM_L_X10Y121_SLICE_X13Y121_AQ;
  assign CLBLM_L_X10Y120_SLICE_X13Y120_C2 = CLBLM_L_X10Y124_SLICE_X12Y124_AQ;
  assign CLBLM_L_X10Y120_SLICE_X13Y120_C3 = CLBLM_L_X10Y121_SLICE_X13Y121_CQ;
  assign CLBLM_L_X8Y110_SLICE_X11Y110_B1 = 1'b1;
  assign CLBLM_L_X8Y110_SLICE_X11Y110_B2 = 1'b1;
  assign CLBLM_L_X8Y110_SLICE_X11Y110_B3 = 1'b1;
  assign CLBLM_L_X8Y110_SLICE_X11Y110_B4 = 1'b1;
  assign CLBLM_L_X8Y110_SLICE_X11Y110_B5 = 1'b1;
  assign CLBLM_L_X8Y110_SLICE_X11Y110_B6 = 1'b1;
  assign CLBLL_L_X4Y116_SLICE_X4Y116_A1 = CLBLL_L_X4Y113_SLICE_X4Y113_AQ;
  assign CLBLL_L_X4Y116_SLICE_X4Y116_A2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLL_L_X4Y116_SLICE_X4Y116_A3 = CLBLL_L_X4Y116_SLICE_X4Y116_AQ;
  assign CLBLL_L_X4Y116_SLICE_X4Y116_A4 = CLBLL_L_X4Y116_SLICE_X5Y116_A5Q;
  assign CLBLL_L_X4Y116_SLICE_X4Y116_A5 = CLBLL_L_X2Y112_SLICE_X1Y112_BQ;
  assign CLBLL_L_X4Y116_SLICE_X4Y116_A6 = CLBLM_L_X8Y112_SLICE_X10Y112_CQ;
  assign CLBLM_L_X8Y110_SLICE_X11Y110_C3 = 1'b1;
  assign CLBLM_L_X8Y110_SLICE_X11Y110_C1 = 1'b1;
  assign CLBLM_L_X8Y110_SLICE_X11Y110_C6 = 1'b1;
  assign CLBLM_L_X8Y110_SLICE_X11Y110_C2 = 1'b1;
  assign CLBLL_L_X4Y116_SLICE_X4Y116_B1 = 1'b1;
  assign CLBLL_L_X4Y116_SLICE_X4Y116_B2 = CLBLL_L_X4Y116_SLICE_X4Y116_BQ;
  assign CLBLL_L_X4Y116_SLICE_X4Y116_B3 = CLBLL_L_X4Y119_SLICE_X5Y119_AQ;
  assign CLBLL_L_X4Y116_SLICE_X4Y116_B4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLL_L_X4Y116_SLICE_X4Y116_B5 = 1'b1;
  assign CLBLL_L_X4Y116_SLICE_X4Y116_B6 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLL_L_X4Y116_SLICE_X4Y116_C1 = RIOB33_X105Y101_IOB_X1Y102_I;
  assign CLBLL_L_X4Y116_SLICE_X4Y116_C2 = CLBLL_L_X4Y116_SLICE_X4Y116_AQ;
  assign CLBLL_L_X4Y116_SLICE_X4Y116_C3 = CLBLL_L_X4Y111_SLICE_X4Y111_CQ;
  assign CLBLM_L_X8Y110_SLICE_X11Y110_D1 = 1'b1;
  assign CLBLL_L_X4Y116_SLICE_X4Y116_C4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLL_L_X4Y116_SLICE_X4Y116_C6 = 1'b1;
  assign CLBLL_L_X4Y116_SLICE_X4Y116_C5 = 1'b1;
  assign CLBLM_L_X8Y110_SLICE_X11Y110_D2 = 1'b1;
  assign CLBLM_L_X8Y110_SLICE_X11Y110_D3 = 1'b1;
  assign CLBLL_L_X4Y116_SLICE_X4Y116_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X8Y110_SLICE_X11Y110_D4 = 1'b1;
  assign CLBLM_L_X8Y110_SLICE_X11Y110_D5 = 1'b1;
  assign CLBLM_L_X8Y110_SLICE_X11Y110_D6 = 1'b1;
  assign CLBLM_L_X8Y110_SLICE_X10Y110_A2 = CLBLL_L_X4Y110_SLICE_X5Y110_BQ;
  assign CLBLM_L_X8Y110_SLICE_X10Y110_A3 = CLBLM_L_X8Y110_SLICE_X10Y110_AQ;
  assign CLBLM_L_X10Y120_SLICE_X12Y120_C2 = CLBLM_L_X10Y120_SLICE_X12Y120_CQ;
  assign CLBLM_L_X10Y120_SLICE_X12Y120_C3 = CLBLM_L_X10Y120_SLICE_X12Y120_DQ;
  assign CLBLM_L_X10Y120_SLICE_X12Y120_C4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y120_SLICE_X12Y120_C5 = CLBLM_L_X8Y121_SLICE_X10Y121_BQ;
  assign CLBLM_L_X10Y120_SLICE_X12Y120_C6 = CLBLM_L_X12Y119_SLICE_X17Y119_AO5;
  assign CLBLM_L_X8Y110_SLICE_X10Y110_A4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y110_SLICE_X10Y110_A5 = 1'b1;
  assign CLBLM_L_X8Y110_SLICE_X10Y110_A6 = CLBLL_L_X4Y110_SLICE_X4Y110_A5Q;
  assign CLBLL_L_X4Y116_SLICE_X4Y116_D1 = CLBLM_R_X7Y119_SLICE_X8Y119_D5Q;
  assign CLBLL_L_X4Y116_SLICE_X4Y116_D2 = CLBLM_R_X7Y115_SLICE_X9Y115_C5Q;
  assign CLBLL_L_X4Y116_SLICE_X4Y116_D3 = CLBLL_L_X4Y116_SLICE_X4Y116_DQ;
  assign CLBLL_L_X4Y116_SLICE_X4Y116_D4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLL_L_X4Y116_SLICE_X4Y116_D5 = CLBLM_L_X10Y113_SLICE_X13Y113_BO6;
  assign CLBLL_L_X4Y116_SLICE_X4Y116_D6 = CLBLM_R_X3Y113_SLICE_X2Y113_BQ;
  assign CLBLM_L_X10Y120_SLICE_X12Y120_D2 = CLBLM_R_X11Y118_SLICE_X15Y118_CQ;
  assign CLBLM_L_X8Y110_SLICE_X10Y110_B1 = CLBLM_L_X10Y111_SLICE_X13Y111_BO6;
  assign CLBLM_L_X8Y110_SLICE_X10Y110_B2 = CLBLM_L_X8Y110_SLICE_X10Y110_BQ;
  assign CLBLM_L_X10Y120_SLICE_X12Y120_D5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y110_SLICE_X10Y110_B4 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X8Y110_SLICE_X10Y110_B5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y110_SLICE_X10Y110_B6 = CLBLM_L_X10Y115_SLICE_X12Y115_AQ;
  assign CLBLM_L_X10Y120_SLICE_X12Y120_D1 = CLBLM_R_X11Y119_SLICE_X14Y119_AO6;
  assign CLBLM_L_X8Y110_SLICE_X10Y110_C1 = CLBLM_R_X5Y111_SLICE_X6Y111_C5Q;
  assign CLBLM_L_X8Y110_SLICE_X10Y110_C2 = CLBLM_L_X10Y118_SLICE_X12Y118_BQ;
  assign CLBLM_L_X8Y110_SLICE_X10Y110_C3 = CLBLM_L_X10Y115_SLICE_X12Y115_DQ;
  assign CLBLM_L_X8Y110_SLICE_X10Y110_C4 = CLBLM_L_X10Y110_SLICE_X12Y110_BQ;
  assign CLBLM_L_X8Y110_SLICE_X10Y110_C5 = CLBLM_L_X8Y110_SLICE_X10Y110_DO6;
  assign CLBLM_L_X8Y110_SLICE_X10Y110_C6 = 1'b1;
  assign CLBLM_L_X8Y110_SLICE_X10Y110_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign LIOB33_X0Y193_IOB_X0Y193_O = LIOB33_X0Y55_IOB_X0Y56_I;
  assign CLBLM_L_X8Y110_SLICE_X10Y110_D1 = CLBLM_R_X7Y115_SLICE_X9Y115_BQ;
  assign CLBLM_L_X8Y110_SLICE_X10Y110_D2 = 1'b1;
  assign CLBLL_L_X4Y116_SLICE_X5Y116_A1 = CLBLM_R_X5Y115_SLICE_X6Y115_CO5;
  assign CLBLL_L_X4Y116_SLICE_X5Y116_A2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y110_SLICE_X10Y110_D3 = CLBLM_L_X8Y116_SLICE_X11Y116_BQ;
  assign CLBLM_L_X8Y110_SLICE_X10Y110_D4 = CLBLM_R_X7Y110_SLICE_X9Y110_BQ;
  assign CLBLM_L_X8Y110_SLICE_X10Y110_D5 = 1'b1;
  assign CLBLM_L_X8Y110_SLICE_X10Y110_D6 = CLBLM_L_X10Y116_SLICE_X13Y116_CQ;
  assign CLBLL_L_X4Y116_SLICE_X5Y116_A3 = CLBLL_L_X4Y116_SLICE_X5Y116_AQ;
  assign CLBLL_L_X4Y116_SLICE_X5Y116_A4 = CLBLM_R_X5Y115_SLICE_X6Y115_BQ;
  assign CLBLL_L_X4Y116_SLICE_X5Y116_A5 = CLBLM_R_X5Y115_SLICE_X7Y115_BQ;
  assign CLBLL_L_X4Y116_SLICE_X5Y116_A6 = 1'b1;
  assign CLBLL_L_X4Y116_SLICE_X5Y116_AX = CLBLL_L_X4Y116_SLICE_X5Y116_CO6;
  assign CLBLL_L_X4Y116_SLICE_X5Y116_B1 = CLBLL_L_X4Y110_SLICE_X5Y110_AQ;
  assign CLBLL_L_X4Y116_SLICE_X5Y116_B2 = CLBLL_L_X4Y116_SLICE_X5Y116_BQ;
  assign CLBLL_L_X4Y116_SLICE_X5Y116_B3 = CLBLM_R_X5Y115_SLICE_X6Y115_CO5;
  assign CLBLL_L_X4Y116_SLICE_X5Y116_B4 = CLBLL_L_X4Y116_SLICE_X5Y116_DQ;
  assign CLBLL_L_X4Y116_SLICE_X5Y116_B5 = 1'b1;
  assign CLBLL_L_X4Y116_SLICE_X5Y116_B6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLL_L_X4Y116_SLICE_X5Y116_C1 = RIOB33_X105Y121_IOB_X1Y121_I;
  assign CLBLL_L_X4Y116_SLICE_X5Y116_C2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLL_L_X4Y116_SLICE_X5Y116_C3 = CLBLM_R_X11Y116_SLICE_X15Y116_AQ;
  assign CLBLL_L_X4Y116_SLICE_X5Y116_C4 = CLBLM_R_X7Y118_SLICE_X9Y118_CQ;
  assign CLBLL_L_X4Y116_SLICE_X5Y116_C5 = CLBLM_R_X11Y113_SLICE_X14Y113_BQ;
  assign CLBLL_L_X4Y116_SLICE_X5Y116_C6 = 1'b1;
  assign CLBLL_L_X4Y122_SLICE_X5Y122_D3 = CLBLL_L_X4Y123_SLICE_X5Y123_AO5;
  assign LIOB33_X0Y187_IOB_X0Y187_O = RIOB33_X105Y143_IOB_X1Y144_I;
  assign CLBLL_L_X4Y116_SLICE_X5Y116_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign LIOB33_X0Y187_IOB_X0Y188_O = RIOB33_X105Y145_IOB_X1Y145_I;
  assign CLBLL_L_X4Y122_SLICE_X5Y122_D4 = RIOB33_X105Y131_IOB_X1Y131_I;
  assign CLBLL_L_X4Y116_SLICE_X5Y116_D1 = CLBLL_L_X4Y116_SLICE_X5Y116_AQ;
  assign CLBLL_L_X4Y116_SLICE_X5Y116_D2 = CLBLM_R_X5Y111_SLICE_X6Y111_CQ;
  assign CLBLL_L_X4Y116_SLICE_X5Y116_D3 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLL_L_X4Y116_SLICE_X5Y116_D4 = 1'b1;
  assign CLBLL_L_X4Y116_SLICE_X5Y116_D5 = 1'b1;
  assign CLBLL_L_X4Y116_SLICE_X5Y116_D6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X11Y114_SLICE_X15Y114_A1 = 1'b1;
  assign CLBLM_R_X11Y114_SLICE_X15Y114_A2 = 1'b1;
  assign CLBLM_R_X11Y114_SLICE_X15Y114_A3 = 1'b1;
  assign CLBLM_R_X11Y114_SLICE_X15Y114_A4 = 1'b1;
  assign CLBLM_R_X11Y114_SLICE_X15Y114_A5 = 1'b1;
  assign CLBLM_R_X11Y114_SLICE_X15Y114_A6 = 1'b1;
  assign CLBLM_R_X11Y114_SLICE_X15Y114_B1 = 1'b1;
  assign CLBLM_R_X11Y114_SLICE_X15Y114_B2 = 1'b1;
  assign CLBLM_R_X11Y114_SLICE_X15Y114_B3 = 1'b1;
  assign CLBLM_R_X11Y114_SLICE_X15Y114_B4 = 1'b1;
  assign CLBLM_R_X11Y114_SLICE_X15Y114_B5 = 1'b1;
  assign CLBLM_R_X11Y114_SLICE_X15Y114_B6 = 1'b1;
  assign CLBLM_R_X11Y114_SLICE_X15Y114_C1 = 1'b1;
  assign CLBLM_R_X11Y114_SLICE_X15Y114_C2 = 1'b1;
  assign CLBLM_R_X11Y114_SLICE_X15Y114_C3 = 1'b1;
  assign CLBLM_R_X11Y114_SLICE_X15Y114_C4 = 1'b1;
  assign CLBLM_R_X11Y114_SLICE_X15Y114_C5 = 1'b1;
  assign CLBLM_R_X11Y114_SLICE_X15Y114_C6 = 1'b1;
  assign CLBLM_R_X11Y114_SLICE_X15Y114_D1 = 1'b1;
  assign CLBLM_R_X11Y114_SLICE_X15Y114_D2 = 1'b1;
  assign CLBLM_R_X11Y114_SLICE_X15Y114_D3 = 1'b1;
  assign CLBLM_R_X11Y114_SLICE_X15Y114_D4 = 1'b1;
  assign CLBLM_R_X11Y114_SLICE_X15Y114_D5 = 1'b1;
  assign CLBLM_R_X11Y114_SLICE_X15Y114_D6 = 1'b1;
  assign CLBLM_R_X11Y114_SLICE_X14Y114_A1 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X11Y114_SLICE_X14Y114_A2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X11Y114_SLICE_X14Y114_A3 = CLBLM_R_X11Y114_SLICE_X14Y114_AQ;
  assign CLBLM_R_X11Y114_SLICE_X14Y114_A4 = CLBLM_R_X11Y117_SLICE_X14Y117_AQ;
  assign CLBLM_R_X11Y114_SLICE_X14Y114_A5 = CLBLM_R_X11Y114_SLICE_X14Y114_CQ;
  assign CLBLM_R_X11Y114_SLICE_X14Y114_A6 = CLBLM_L_X10Y113_SLICE_X12Y113_DO6;
  assign CLBLM_R_X13Y119_SLICE_X19Y119_A6 = 1'b1;
  assign CLBLM_R_X11Y114_SLICE_X14Y114_B1 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X11Y114_SLICE_X14Y114_B2 = CLBLM_R_X11Y114_SLICE_X14Y114_BQ;
  assign CLBLM_R_X11Y114_SLICE_X14Y114_B3 = CLBLM_L_X8Y113_SLICE_X11Y113_BQ;
  assign CLBLM_R_X11Y114_SLICE_X14Y114_B4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X11Y114_SLICE_X14Y114_B5 = CLBLM_L_X10Y120_SLICE_X13Y120_BQ;
  assign CLBLM_R_X11Y114_SLICE_X14Y114_B6 = CLBLM_L_X10Y113_SLICE_X12Y113_DO6;
  assign CLBLM_R_X11Y114_SLICE_X14Y114_C1 = CLBLM_L_X8Y113_SLICE_X11Y113_AQ;
  assign CLBLM_R_X11Y114_SLICE_X14Y114_C2 = CLBLM_R_X11Y114_SLICE_X14Y114_CQ;
  assign CLBLM_R_X11Y114_SLICE_X14Y114_C3 = CLBLM_L_X12Y115_SLICE_X16Y115_CQ;
  assign CLBLM_R_X11Y114_SLICE_X14Y114_C4 = CLBLM_L_X10Y113_SLICE_X12Y113_DO6;
  assign CLBLM_R_X11Y114_SLICE_X14Y114_C5 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X11Y114_SLICE_X14Y114_C6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X11Y114_SLICE_X14Y114_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLL_L_X52Y126_SLICE_X78Y126_B4 = 1'b1;
  assign RIOI3_X105Y101_ILOGIC_X1Y102_D = RIOB33_X105Y101_IOB_X1Y102_I;
  assign CLBLM_R_X11Y114_SLICE_X14Y114_D1 = CLBLM_L_X10Y114_SLICE_X13Y114_CQ;
  assign CLBLL_L_X52Y126_SLICE_X78Y126_B5 = 1'b1;
  assign CLBLM_R_X11Y114_SLICE_X14Y114_D2 = CLBLM_L_X8Y115_SLICE_X10Y115_C5Q;
  assign CLBLM_R_X11Y114_SLICE_X14Y114_D3 = CLBLM_R_X11Y114_SLICE_X14Y114_AQ;
  assign CLBLM_R_X11Y114_SLICE_X14Y114_D4 = RIOB33_X105Y103_IOB_X1Y104_I;
  assign CLBLM_R_X11Y114_SLICE_X14Y114_D5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLL_L_X52Y126_SLICE_X78Y126_B6 = 1'b1;
  assign CLBLM_R_X11Y114_SLICE_X14Y114_D6 = 1'b1;
  assign LIOI3_X0Y53_ILOGIC_X0Y54_D = LIOB33_X0Y53_IOB_X0Y54_I;
  assign LIOI3_X0Y53_ILOGIC_X0Y53_D = LIOB33_X0Y53_IOB_X0Y53_I;
  assign RIOI3_X105Y101_ILOGIC_X1Y101_D = RIOB33_X105Y101_IOB_X1Y101_I;
  assign CLBLM_R_X13Y119_SLICE_X19Y119_C1 = 1'b1;
  assign CLBLM_R_X13Y119_SLICE_X19Y119_C2 = 1'b1;
  assign CLBLL_L_X52Y126_SLICE_X78Y126_C4 = 1'b1;
  assign LIOI3_TBYTESRC_X0Y69_ILOGIC_X0Y70_D = LIOB33_X0Y69_IOB_X0Y70_I;
  assign LIOI3_TBYTESRC_X0Y69_ILOGIC_X0Y69_D = LIOB33_X0Y69_IOB_X0Y69_I;
  assign CLBLM_R_X13Y119_SLICE_X19Y119_C5 = 1'b1;
  assign LIOI3_X0Y183_OLOGIC_X0Y184_D1 = RIOB33_X105Y135_IOB_X1Y136_I;
  assign CLBLM_L_X10Y121_SLICE_X13Y121_A1 = CLBLM_L_X10Y124_SLICE_X13Y124_BO5;
  assign CLBLM_L_X10Y121_SLICE_X13Y121_A2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y121_SLICE_X13Y121_A3 = CLBLM_L_X10Y121_SLICE_X13Y121_AQ;
  assign CLBLM_L_X10Y121_SLICE_X13Y121_A4 = CLBLM_L_X10Y121_SLICE_X12Y121_CO6;
  assign CLBLM_L_X10Y121_SLICE_X13Y121_A5 = CLBLM_R_X7Y122_SLICE_X8Y122_DQ;
  assign CLBLM_L_X10Y121_SLICE_X13Y121_A6 = CLBLM_L_X10Y124_SLICE_X13Y124_AO5;
  assign CLBLM_L_X10Y121_SLICE_X13Y121_B1 = CLBLM_L_X10Y124_SLICE_X13Y124_BO5;
  assign CLBLM_L_X10Y121_SLICE_X13Y121_B2 = 1'b1;
  assign CLBLM_L_X10Y121_SLICE_X13Y121_B3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y121_SLICE_X13Y121_B4 = CLBLM_L_X10Y123_SLICE_X12Y123_DO6;
  assign CLBLM_L_X10Y121_SLICE_X13Y121_B5 = CLBLM_R_X11Y120_SLICE_X15Y120_BQ;
  assign CLBLM_L_X10Y121_SLICE_X13Y121_B6 = CLBLM_L_X10Y124_SLICE_X13Y124_AO5;
  assign CLBLM_R_X13Y120_SLICE_X19Y120_A2 = 1'b1;
  assign CLBLM_L_X8Y111_SLICE_X11Y111_A1 = CLBLM_L_X8Y111_SLICE_X11Y111_DO6;
  assign CLBLM_L_X8Y111_SLICE_X11Y111_A2 = CLBLM_L_X8Y111_SLICE_X10Y111_BO6;
  assign CLBLM_L_X8Y111_SLICE_X11Y111_A3 = CLBLM_L_X10Y111_SLICE_X12Y111_DO6;
  assign CLBLM_L_X8Y111_SLICE_X11Y111_A4 = CLBLM_L_X8Y111_SLICE_X11Y111_BO6;
  assign CLBLM_L_X8Y111_SLICE_X11Y111_A5 = CLBLM_L_X8Y113_SLICE_X11Y113_DO6;
  assign CLBLM_L_X8Y111_SLICE_X11Y111_A6 = CLBLM_L_X8Y111_SLICE_X11Y111_CO6;
  assign CLBLM_L_X10Y121_SLICE_X13Y121_C1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y121_SLICE_X13Y121_C2 = CLBLM_L_X10Y124_SLICE_X13Y124_AO5;
  assign CLBLM_L_X10Y121_SLICE_X13Y121_C3 = CLBLM_L_X10Y124_SLICE_X13Y124_BO5;
  assign CLBLM_L_X8Y111_SLICE_X11Y111_B1 = CLBLM_L_X8Y112_SLICE_X11Y112_BO5;
  assign CLBLL_L_X4Y117_SLICE_X4Y117_A1 = 1'b1;
  assign CLBLM_L_X8Y111_SLICE_X11Y111_B3 = CLBLM_R_X7Y111_SLICE_X9Y111_BO6;
  assign CLBLM_L_X8Y111_SLICE_X11Y111_B4 = CLBLM_R_X5Y119_SLICE_X7Y119_CO6;
  assign CLBLM_L_X8Y111_SLICE_X11Y111_B5 = CLBLM_L_X10Y118_SLICE_X12Y118_BQ;
  assign CLBLM_L_X8Y111_SLICE_X11Y111_B6 = CLBLL_L_X4Y119_SLICE_X4Y119_CQ;
  assign CLBLL_L_X4Y117_SLICE_X4Y117_A2 = CLBLM_R_X5Y114_SLICE_X6Y114_CQ;
  assign CLBLL_L_X4Y117_SLICE_X4Y117_A3 = CLBLL_L_X4Y117_SLICE_X4Y117_AQ;
  assign CLBLL_L_X4Y117_SLICE_X4Y117_A4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLL_L_X4Y117_SLICE_X4Y117_A5 = CLBLL_L_X4Y116_SLICE_X5Y116_BQ;
  assign CLBLL_L_X4Y117_SLICE_X4Y117_A6 = CLBLM_R_X5Y115_SLICE_X6Y115_CO5;
  assign CLBLM_L_X8Y111_SLICE_X11Y111_C2 = CLBLM_L_X10Y111_SLICE_X13Y111_CO5;
  assign CLBLM_L_X8Y111_SLICE_X11Y111_C3 = CLBLM_R_X5Y119_SLICE_X7Y119_CO6;
  assign CLBLM_L_X8Y111_SLICE_X11Y111_C4 = 1'b1;
  assign CLBLL_L_X4Y117_SLICE_X4Y117_B5 = 1'b1;
  assign CLBLL_L_X4Y117_SLICE_X4Y117_B6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y111_SLICE_X11Y111_C5 = CLBLM_R_X5Y111_SLICE_X7Y111_CO6;
  assign CLBLM_L_X8Y111_SLICE_X11Y111_C6 = CLBLM_R_X7Y115_SLICE_X9Y115_BQ;
  assign CLBLL_L_X4Y117_SLICE_X4Y117_B1 = 1'b1;
  assign CLBLL_L_X4Y117_SLICE_X4Y117_B2 = CLBLL_L_X4Y117_SLICE_X4Y117_BQ;
  assign CLBLL_L_X4Y117_SLICE_X4Y117_C2 = CLBLL_L_X2Y121_SLICE_X1Y121_BO5;
  assign CLBLL_L_X4Y117_SLICE_X4Y117_C1 = CLBLL_L_X4Y115_SLICE_X4Y115_AQ;
  assign CLBLL_L_X4Y117_SLICE_X4Y117_C4 = CLBLL_L_X2Y121_SLICE_X1Y121_BO6;
  assign CLBLM_L_X8Y111_SLICE_X11Y111_D1 = CLBLM_R_X7Y111_SLICE_X9Y111_AO5;
  assign CLBLM_L_X8Y111_SLICE_X11Y111_D2 = CLBLM_L_X10Y127_SLICE_X12Y127_AQ;
  assign CLBLM_L_X8Y111_SLICE_X11Y111_D3 = CLBLM_R_X5Y119_SLICE_X7Y119_CO6;
  assign CLBLL_L_X4Y117_SLICE_X4Y117_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X8Y111_SLICE_X11Y111_D4 = 1'b1;
  assign CLBLM_L_X8Y111_SLICE_X11Y111_D5 = CLBLM_R_X5Y111_SLICE_X7Y111_CO6;
  assign CLBLM_L_X8Y111_SLICE_X11Y111_D6 = CLBLM_L_X10Y111_SLICE_X12Y111_AO6;
  assign CLBLL_L_X4Y117_SLICE_X4Y117_C6 = CLBLL_L_X4Y111_SLICE_X4Y111_BQ;
  assign CLBLL_L_X4Y117_SLICE_X4Y117_D1 = CLBLL_L_X4Y116_SLICE_X5Y116_BQ;
  assign CLBLL_L_X4Y117_SLICE_X4Y117_D2 = 1'b1;
  assign CLBLM_L_X8Y111_SLICE_X10Y111_A1 = CLBLM_R_X5Y111_SLICE_X7Y111_BQ;
  assign CLBLM_L_X8Y111_SLICE_X10Y111_A2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y111_SLICE_X10Y111_A3 = CLBLM_L_X8Y111_SLICE_X10Y111_AQ;
  assign CLBLM_L_X8Y111_SLICE_X10Y111_A4 = CLBLM_L_X10Y113_SLICE_X12Y113_DO6;
  assign CLBLM_L_X8Y111_SLICE_X10Y111_A5 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X8Y111_SLICE_X10Y111_A6 = CLBLM_R_X11Y113_SLICE_X15Y113_BQ;
  assign CLBLL_L_X4Y117_SLICE_X4Y117_D3 = CLBLL_L_X4Y120_SLICE_X5Y120_BO6;
  assign CLBLL_L_X4Y117_SLICE_X4Y117_D4 = CLBLM_R_X3Y117_SLICE_X2Y117_DO6;
  assign CLBLL_L_X4Y117_SLICE_X4Y117_D5 = CLBLL_L_X4Y116_SLICE_X4Y116_DQ;
  assign CLBLL_L_X4Y117_SLICE_X4Y117_D6 = CLBLL_L_X2Y121_SLICE_X1Y121_AO6;
  assign CLBLM_L_X8Y111_SLICE_X10Y111_B1 = CLBLM_R_X5Y111_SLICE_X7Y111_CO6;
  assign CLBLM_L_X8Y111_SLICE_X10Y111_B2 = CLBLM_R_X7Y111_SLICE_X9Y111_AO5;
  assign CLBLM_L_X8Y111_SLICE_X10Y111_B3 = CLBLM_R_X5Y119_SLICE_X7Y119_CO6;
  assign CLBLM_L_X8Y111_SLICE_X10Y111_B4 = CLBLM_R_X7Y111_SLICE_X9Y111_BO5;
  assign CLBLM_L_X8Y111_SLICE_X10Y111_B5 = CLBLM_R_X5Y111_SLICE_X6Y111_C5Q;
  assign CLBLM_L_X8Y111_SLICE_X10Y111_B6 = CLBLM_R_X5Y114_SLICE_X6Y114_DQ;
  assign CLBLM_L_X10Y121_SLICE_X12Y121_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X10Y121_SLICE_X12Y121_D2 = CLBLM_L_X8Y121_SLICE_X10Y121_CQ;
  assign CLBLM_L_X10Y121_SLICE_X12Y121_D1 = CLBLM_L_X8Y115_SLICE_X10Y115_AQ;
  assign CLBLM_L_X8Y111_SLICE_X10Y111_C1 = CLBLM_R_X7Y110_SLICE_X8Y110_AQ;
  assign CLBLM_L_X8Y111_SLICE_X10Y111_C2 = CLBLM_L_X8Y118_SLICE_X10Y118_CQ;
  assign CLBLM_L_X8Y111_SLICE_X10Y111_C3 = 1'b1;
  assign CLBLM_L_X8Y111_SLICE_X10Y111_C4 = CLBLM_R_X5Y114_SLICE_X6Y114_AQ;
  assign CLBLM_L_X8Y111_SLICE_X10Y111_C5 = CLBLM_L_X8Y117_SLICE_X10Y117_BQ;
  assign CLBLM_L_X8Y111_SLICE_X10Y111_C6 = 1'b1;
  assign CLBLM_L_X10Y121_SLICE_X12Y121_D3 = CLBLM_L_X10Y119_SLICE_X13Y119_DQ;
  assign CLBLM_L_X10Y121_SLICE_X12Y121_D4 = CLBLM_L_X10Y126_SLICE_X12Y126_AQ;
  assign CLBLM_L_X8Y111_SLICE_X10Y111_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X10Y121_SLICE_X12Y121_D6 = CLBLL_L_X4Y117_SLICE_X5Y117_DQ;
  assign CLBLL_L_X4Y117_SLICE_X5Y117_A1 = CLBLM_L_X8Y112_SLICE_X10Y112_CQ;
  assign CLBLL_L_X4Y117_SLICE_X5Y117_A2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLL_L_X4Y117_SLICE_X5Y117_A3 = CLBLM_R_X3Y111_SLICE_X3Y111_BQ;
  assign CLBLL_L_X4Y117_SLICE_X5Y117_A4 = CLBLL_L_X4Y117_SLICE_X5Y117_AQ;
  assign CLBLL_L_X4Y117_SLICE_X5Y117_A5 = CLBLL_L_X2Y112_SLICE_X1Y112_BQ;
  assign CLBLL_L_X4Y117_SLICE_X5Y117_A6 = CLBLM_R_X5Y117_SLICE_X7Y117_BQ;
  assign CLBLM_L_X8Y111_SLICE_X10Y111_D2 = CLBLM_L_X8Y118_SLICE_X10Y118_CQ;
  assign CLBLM_L_X8Y111_SLICE_X10Y111_D3 = CLBLM_R_X11Y114_SLICE_X14Y114_BQ;
  assign CLBLM_L_X8Y111_SLICE_X10Y111_D4 = 1'b1;
  assign CLBLM_L_X8Y111_SLICE_X10Y111_D5 = 1'b1;
  assign CLBLM_L_X8Y111_SLICE_X10Y111_D6 = CLBLM_R_X11Y113_SLICE_X15Y113_BQ;
  assign CLBLM_L_X8Y111_SLICE_X10Y111_D1 = CLBLM_R_X7Y110_SLICE_X8Y110_AQ;
  assign CLBLL_L_X4Y117_SLICE_X5Y117_B1 = 1'b1;
  assign CLBLL_L_X4Y117_SLICE_X5Y117_B2 = CLBLL_L_X4Y117_SLICE_X5Y117_BQ;
  assign CLBLL_L_X4Y117_SLICE_X5Y117_B3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLL_L_X4Y117_SLICE_X5Y117_B4 = CLBLM_R_X11Y121_SLICE_X14Y121_CO6;
  assign CLBLL_L_X4Y117_SLICE_X5Y117_B5 = CLBLL_L_X4Y117_SLICE_X4Y117_AQ;
  assign CLBLL_L_X4Y117_SLICE_X5Y117_B6 = CLBLL_L_X4Y110_SLICE_X4Y110_CQ;
  assign CLBLL_L_X4Y117_SLICE_X5Y117_C1 = CLBLM_R_X3Y116_SLICE_X3Y116_BQ;
  assign CLBLL_L_X4Y117_SLICE_X5Y117_C2 = CLBLL_L_X4Y117_SLICE_X5Y117_CQ;
  assign CLBLL_L_X4Y117_SLICE_X5Y117_C3 = CLBLM_R_X7Y119_SLICE_X9Y119_BQ;
  assign CLBLL_L_X4Y117_SLICE_X5Y117_C4 = 1'b1;
  assign CLBLL_L_X4Y117_SLICE_X5Y117_C5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLL_L_X4Y117_SLICE_X5Y117_C6 = CLBLM_R_X11Y121_SLICE_X14Y121_CO6;
  assign CLBLL_L_X4Y117_SLICE_X5Y117_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X13Y119_SLICE_X18Y119_A6 = 1'b1;
  assign CLBLM_R_X11Y121_SLICE_X15Y121_C1 = 1'b1;
  assign CLBLM_R_X13Y120_SLICE_X19Y120_A3 = 1'b1;
  assign CLBLL_L_X4Y117_SLICE_X5Y117_D1 = CLBLL_L_X4Y116_SLICE_X5Y116_CO5;
  assign CLBLL_L_X4Y117_SLICE_X5Y117_D2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLL_L_X4Y117_SLICE_X5Y117_D3 = 1'b1;
  assign CLBLL_L_X4Y117_SLICE_X5Y117_D4 = CLBLL_L_X4Y115_SLICE_X5Y115_DQ;
  assign CLBLL_L_X4Y117_SLICE_X5Y117_D5 = CLBLM_L_X8Y115_SLICE_X10Y115_AQ;
  assign CLBLL_L_X4Y117_SLICE_X5Y117_D6 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X11Y121_SLICE_X15Y121_C2 = CLBLM_L_X10Y120_SLICE_X13Y120_A5Q;
  assign CLBLM_R_X11Y121_SLICE_X15Y121_C3 = 1'b1;
  assign RIOB33_X105Y175_IOB_X1Y175_O = CLBLM_L_X10Y128_SLICE_X13Y128_AO6;
  assign CLBLM_R_X11Y115_SLICE_X15Y115_A1 = CLBLM_R_X3Y118_SLICE_X2Y118_AQ;
  assign CLBLM_R_X11Y115_SLICE_X15Y115_A2 = CLBLM_R_X11Y115_SLICE_X15Y115_DQ;
  assign CLBLM_R_X11Y115_SLICE_X15Y115_A3 = CLBLM_R_X11Y115_SLICE_X15Y115_AQ;
  assign CLBLM_R_X11Y115_SLICE_X15Y115_A4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X11Y115_SLICE_X15Y115_A5 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_R_X11Y115_SLICE_X15Y115_A6 = CLBLM_R_X5Y112_SLICE_X7Y112_BO6;
  assign CLBLM_R_X11Y121_SLICE_X15Y121_C4 = CLBLM_R_X11Y120_SLICE_X15Y120_BQ;
  assign CLBLM_R_X11Y121_SLICE_X15Y121_C5 = 1'b1;
  assign CLBLM_R_X11Y115_SLICE_X15Y115_B1 = 1'b1;
  assign CLBLM_R_X11Y115_SLICE_X15Y115_B2 = CLBLM_R_X11Y115_SLICE_X15Y115_DQ;
  assign CLBLM_R_X11Y115_SLICE_X15Y115_B3 = CLBLM_L_X8Y113_SLICE_X11Y113_BQ;
  assign CLBLM_R_X11Y115_SLICE_X15Y115_B4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X11Y115_SLICE_X15Y115_B5 = CLBLM_R_X5Y111_SLICE_X7Y111_DO6;
  assign CLBLM_R_X11Y115_SLICE_X15Y115_B6 = CLBLM_R_X11Y115_SLICE_X15Y115_BQ;
  assign CLBLM_R_X11Y121_SLICE_X15Y121_C6 = 1'b1;
  assign CLBLM_R_X11Y115_SLICE_X15Y115_C1 = CLBLM_R_X5Y111_SLICE_X7Y111_DO6;
  assign CLBLM_R_X11Y115_SLICE_X15Y115_C2 = CLBLM_R_X11Y115_SLICE_X15Y115_CQ;
  assign CLBLM_R_X11Y115_SLICE_X15Y115_C3 = CLBLM_R_X11Y115_SLICE_X15Y115_BQ;
  assign CLBLM_R_X11Y115_SLICE_X15Y115_C4 = CLBLM_L_X10Y115_SLICE_X12Y115_DQ;
  assign CLBLM_R_X11Y115_SLICE_X15Y115_C5 = 1'b1;
  assign CLBLM_R_X11Y115_SLICE_X15Y115_C6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X11Y115_SLICE_X15Y115_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign LIOI3_X0Y183_OLOGIC_X0Y183_T1 = 1'b1;
  assign CLBLM_R_X13Y119_SLICE_X18Y119_B6 = CLBLM_R_X7Y114_SLICE_X8Y114_BQ;
  assign CLBLM_R_X11Y115_SLICE_X15Y115_D1 = CLBLM_R_X5Y111_SLICE_X7Y111_DO6;
  assign CLBLM_R_X11Y115_SLICE_X15Y115_D2 = CLBLM_R_X11Y115_SLICE_X15Y115_CQ;
  assign CLBLM_R_X11Y115_SLICE_X15Y115_D3 = CLBLM_R_X11Y115_SLICE_X15Y115_DQ;
  assign CLBLM_R_X11Y115_SLICE_X15Y115_D4 = 1'b1;
  assign CLBLM_R_X11Y115_SLICE_X15Y115_D5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X11Y115_SLICE_X15Y115_D6 = CLBLM_R_X11Y117_SLICE_X14Y117_BQ;
  assign CLBLM_R_X11Y115_SLICE_X14Y115_A1 = CLBLM_R_X11Y116_SLICE_X14Y116_BO5;
  assign CLBLM_R_X11Y115_SLICE_X14Y115_A2 = CLBLM_L_X10Y110_SLICE_X13Y110_CO5;
  assign CLBLM_R_X11Y115_SLICE_X14Y115_A3 = CLBLM_R_X11Y115_SLICE_X14Y115_AQ;
  assign CLBLM_R_X11Y115_SLICE_X14Y115_A4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X11Y115_SLICE_X14Y115_A5 = CLBLM_L_X10Y113_SLICE_X12Y113_DO6;
  assign CLBLM_R_X11Y115_SLICE_X14Y115_A6 = CLBLM_R_X11Y120_SLICE_X15Y120_CQ;
  assign LIOB33_SING_X0Y100_IOB_X0Y100_O = CLBLL_L_X2Y111_SLICE_X0Y111_BO6;
  assign CLBLL_L_X52Y126_SLICE_X79Y126_A2 = 1'b1;
  assign CLBLM_R_X11Y115_SLICE_X14Y115_B1 = 1'b1;
  assign CLBLM_R_X11Y115_SLICE_X14Y115_B2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X11Y115_SLICE_X14Y115_B3 = CLBLM_R_X7Y128_SLICE_X8Y128_AQ;
  assign CLBLM_R_X11Y115_SLICE_X14Y115_B4 = RIOB33_X105Y141_IOB_X1Y142_I;
  assign CLBLL_L_X52Y126_SLICE_X79Y126_A3 = 1'b1;
  assign CLBLM_R_X11Y115_SLICE_X14Y115_B5 = CLBLM_L_X10Y115_SLICE_X13Y115_BO6;
  assign CLBLM_R_X11Y115_SLICE_X14Y115_B6 = CLBLM_R_X11Y115_SLICE_X14Y115_DQ;
  assign CLBLM_R_X11Y121_SLICE_X15Y121_D1 = 1'b1;
  assign CLBLM_R_X11Y121_SLICE_X15Y121_D2 = 1'b1;
  assign CLBLL_L_X52Y126_SLICE_X79Y126_A4 = 1'b1;
  assign CLBLM_R_X11Y115_SLICE_X14Y115_C1 = CLBLM_R_X7Y128_SLICE_X8Y128_AQ;
  assign CLBLM_R_X11Y115_SLICE_X14Y115_C2 = 1'b1;
  assign CLBLM_R_X11Y115_SLICE_X14Y115_C3 = CLBLM_R_X7Y117_SLICE_X9Y117_CQ;
  assign CLBLM_R_X11Y115_SLICE_X14Y115_C4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLL_L_X52Y126_SLICE_X79Y126_A5 = 1'b1;
  assign CLBLM_R_X11Y115_SLICE_X14Y115_C5 = CLBLM_L_X10Y115_SLICE_X13Y115_AO6;
  assign CLBLM_R_X11Y115_SLICE_X14Y115_C6 = RIOB33_X105Y141_IOB_X1Y142_I;
  assign CLBLM_R_X11Y121_SLICE_X15Y121_D3 = 1'b1;
  assign CLBLM_R_X11Y121_SLICE_X15Y121_D4 = 1'b1;
  assign CLBLL_L_X52Y126_SLICE_X79Y126_A6 = 1'b1;
  assign CLBLM_R_X11Y115_SLICE_X14Y115_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X11Y121_SLICE_X15Y121_D5 = 1'b1;
  assign LIOB33_X0Y135_IOB_X0Y136_O = CLBLM_R_X7Y124_SLICE_X8Y124_CQ;
  assign CLBLM_R_X11Y115_SLICE_X14Y115_D1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X11Y115_SLICE_X14Y115_D2 = CLBLM_R_X7Y113_SLICE_X8Y113_DO6;
  assign CLBLM_R_X11Y115_SLICE_X14Y115_D3 = CLBLM_R_X3Y118_SLICE_X2Y118_AQ;
  assign CLBLM_R_X11Y115_SLICE_X14Y115_D4 = CLBLM_R_X11Y115_SLICE_X14Y115_DQ;
  assign CLBLM_R_X11Y115_SLICE_X14Y115_D5 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_R_X11Y115_SLICE_X14Y115_D6 = CLBLM_L_X8Y115_SLICE_X10Y115_C5Q;
  assign CLBLM_R_X11Y121_SLICE_X15Y121_D6 = 1'b1;
  assign CLBLM_R_X13Y119_SLICE_X18Y119_C6 = CLBLM_L_X12Y119_SLICE_X17Y119_AO6;
  assign LIOB33_X0Y135_IOB_X0Y135_O = CLBLL_L_X4Y123_SLICE_X4Y123_AQ;
  assign LIOI3_TBYTESRC_X0Y119_OLOGIC_X0Y120_D1 = CLBLM_R_X3Y116_SLICE_X3Y116_A5Q;
  assign RIOI3_X105Y185_OLOGIC_X1Y186_D1 = CLBLM_L_X12Y115_SLICE_X16Y115_BQ;
  assign RIOI3_X105Y153_OLOGIC_X1Y153_T1 = 1'b1;
  assign CLBLL_L_X52Y126_SLICE_X79Y126_B1 = 1'b1;
  assign CLBLM_R_X13Y119_SLICE_X18Y119_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLL_L_X52Y126_SLICE_X79Y126_B2 = 1'b1;
  assign CLBLL_L_X52Y126_SLICE_X79Y126_B3 = 1'b1;
  assign CLBLM_R_X13Y120_SLICE_X19Y120_A4 = 1'b1;
  assign CLBLL_L_X2Y110_SLICE_X0Y110_A6 = 1'b1;
  assign CLBLL_L_X52Y126_SLICE_X79Y126_B4 = 1'b1;
  assign CLBLL_L_X52Y126_SLICE_X79Y126_B5 = 1'b1;
  assign CLBLM_R_X11Y121_SLICE_X14Y121_A1 = CLBLM_L_X10Y119_SLICE_X13Y119_AQ;
  assign CLBLL_L_X52Y126_SLICE_X79Y126_B6 = 1'b1;
  assign CLBLM_R_X11Y121_SLICE_X14Y121_A2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X11Y121_SLICE_X14Y121_A3 = CLBLM_R_X11Y119_SLICE_X15Y119_CQ;
  assign CLBLM_R_X11Y121_SLICE_X14Y121_A4 = CLBLM_R_X7Y120_SLICE_X9Y120_AQ;
  assign CLBLL_L_X52Y126_SLICE_X79Y126_C1 = 1'b1;
  assign RIOI3_X105Y185_OLOGIC_X1Y186_T1 = 1'b1;
  assign CLBLM_R_X13Y119_SLICE_X18Y119_D4 = CLBLM_R_X11Y119_SLICE_X15Y119_CQ;
  assign CLBLL_L_X52Y126_SLICE_X79Y126_C2 = 1'b1;
  assign CLBLM_R_X13Y119_SLICE_X18Y119_D5 = CLBLM_R_X11Y120_SLICE_X15Y120_AQ;
  assign CLBLL_L_X2Y110_SLICE_X0Y110_B5 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLL_L_X52Y126_SLICE_X79Y126_C3 = 1'b1;
  assign CLBLM_R_X13Y119_SLICE_X18Y119_D6 = CLBLM_R_X11Y118_SLICE_X14Y118_BQ;
  assign CLBLM_L_X10Y122_SLICE_X13Y122_A1 = CLBLM_L_X10Y124_SLICE_X13Y124_BO5;
  assign CLBLM_L_X10Y122_SLICE_X13Y122_A2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y122_SLICE_X13Y122_A3 = CLBLM_L_X10Y112_SLICE_X13Y112_AQ;
  assign CLBLM_L_X10Y122_SLICE_X13Y122_A4 = CLBLM_L_X10Y122_SLICE_X12Y122_DO6;
  assign CLBLM_L_X10Y122_SLICE_X13Y122_A5 = 1'b1;
  assign CLBLM_L_X10Y122_SLICE_X13Y122_A6 = CLBLM_L_X10Y124_SLICE_X13Y124_AO5;
  assign CLBLL_L_X2Y110_SLICE_X0Y110_B6 = CLBLL_L_X4Y120_SLICE_X4Y120_AO6;
  assign CLBLL_L_X52Y126_SLICE_X79Y126_C4 = 1'b1;
  assign CLBLM_L_X10Y122_SLICE_X13Y122_AX = CLBLM_L_X10Y124_SLICE_X13Y124_AO6;
  assign CLBLL_L_X52Y126_SLICE_X79Y126_C5 = 1'b1;
  assign CLBLM_L_X10Y122_SLICE_X13Y122_B1 = CLBLM_L_X10Y124_SLICE_X13Y124_BO5;
  assign CLBLM_L_X10Y122_SLICE_X13Y122_B2 = CLBLM_L_X10Y122_SLICE_X13Y122_BQ;
  assign CLBLM_L_X10Y122_SLICE_X13Y122_B3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y122_SLICE_X13Y122_B4 = CLBLM_L_X10Y122_SLICE_X13Y122_DO6;
  assign CLBLM_L_X10Y122_SLICE_X13Y122_B5 = CLBLM_R_X7Y120_SLICE_X9Y120_DQ;
  assign CLBLM_L_X10Y122_SLICE_X13Y122_B6 = CLBLM_L_X10Y124_SLICE_X13Y124_AO5;
  assign CLBLL_L_X52Y126_SLICE_X79Y126_C6 = 1'b1;
  assign CLBLM_R_X7Y123_SLICE_X9Y123_C5 = CLBLM_R_X7Y124_SLICE_X9Y124_AQ;
  assign CLBLM_R_X7Y123_SLICE_X9Y123_C6 = CLBLM_R_X5Y120_SLICE_X6Y120_A5Q;
  assign CLBLM_L_X8Y112_SLICE_X11Y112_A1 = CLBLM_L_X8Y112_SLICE_X11Y112_DO6;
  assign CLBLM_L_X10Y122_SLICE_X13Y122_C2 = CLBLM_L_X10Y122_SLICE_X13Y122_CQ;
  assign CLBLM_L_X10Y122_SLICE_X13Y122_C3 = CLBLM_L_X10Y124_SLICE_X13Y124_BO5;
  assign CLBLM_L_X10Y122_SLICE_X13Y122_C4 = CLBLM_L_X10Y124_SLICE_X13Y124_AO5;
  assign CLBLM_L_X10Y122_SLICE_X13Y122_C5 = CLBLM_L_X10Y119_SLICE_X12Y119_AQ;
  assign CLBLM_L_X10Y122_SLICE_X13Y122_C6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y112_SLICE_X11Y112_A2 = CLBLM_R_X3Y118_SLICE_X2Y118_AQ;
  assign CLBLM_L_X8Y112_SLICE_X11Y112_A3 = CLBLM_R_X7Y111_SLICE_X9Y111_AO6;
  assign CLBLM_L_X10Y122_SLICE_X13Y122_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X8Y112_SLICE_X11Y112_A4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y112_SLICE_X11Y112_A5 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_L_X8Y112_SLICE_X11Y112_A6 = CLBLM_L_X8Y117_SLICE_X11Y117_CQ;
  assign CLBLL_L_X4Y118_SLICE_X4Y118_A1 = CLBLM_R_X5Y115_SLICE_X6Y115_CO6;
  assign CLBLL_L_X4Y118_SLICE_X4Y118_A2 = CLBLL_L_X4Y112_SLICE_X5Y112_AQ;
  assign CLBLM_L_X10Y122_SLICE_X13Y122_D1 = CLBLM_R_X11Y121_SLICE_X14Y121_BO6;
  assign CLBLM_L_X10Y122_SLICE_X13Y122_D2 = CLBLM_L_X10Y123_SLICE_X12Y123_CO6;
  assign CLBLM_L_X10Y122_SLICE_X13Y122_D3 = CLBLM_L_X8Y122_SLICE_X11Y122_DO6;
  assign CLBLM_L_X10Y122_SLICE_X13Y122_D4 = CLBLM_L_X10Y122_SLICE_X13Y122_AQ;
  assign CLBLM_L_X10Y122_SLICE_X13Y122_D5 = CLBLM_R_X11Y121_SLICE_X14Y121_BO5;
  assign CLBLM_L_X10Y122_SLICE_X13Y122_D6 = CLBLM_L_X8Y121_SLICE_X11Y121_AQ;
  assign CLBLL_L_X4Y118_SLICE_X4Y118_B1 = CLBLL_L_X2Y119_SLICE_X1Y119_AO5;
  assign CLBLL_L_X4Y118_SLICE_X4Y118_B2 = CLBLL_L_X4Y120_SLICE_X5Y120_BO6;
  assign CLBLL_L_X4Y118_SLICE_X4Y118_B3 = CLBLM_L_X10Y117_SLICE_X13Y117_CQ;
  assign CLBLL_L_X4Y118_SLICE_X4Y118_B4 = CLBLL_L_X2Y121_SLICE_X1Y121_AO6;
  assign CLBLL_L_X4Y118_SLICE_X4Y118_B5 = CLBLM_R_X3Y112_SLICE_X2Y112_AQ;
  assign CLBLM_L_X10Y122_SLICE_X12Y122_A1 = 1'b1;
  assign CLBLM_L_X10Y122_SLICE_X12Y122_A2 = CLBLM_R_X7Y122_SLICE_X8Y122_CQ;
  assign CLBLM_L_X10Y122_SLICE_X12Y122_A3 = 1'b1;
  assign CLBLM_L_X10Y122_SLICE_X12Y122_A4 = CLBLM_L_X10Y124_SLICE_X13Y124_BO6;
  assign CLBLM_L_X10Y122_SLICE_X12Y122_A5 = CLBLM_L_X10Y118_SLICE_X13Y118_AQ;
  assign CLBLM_L_X10Y122_SLICE_X12Y122_A6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLL_L_X4Y118_SLICE_X4Y118_C2 = CLBLM_R_X3Y118_SLICE_X3Y118_BO6;
  assign CLBLL_L_X4Y118_SLICE_X4Y118_C3 = CLBLL_L_X4Y121_SLICE_X4Y121_CO6;
  assign CLBLL_L_X4Y118_SLICE_X4Y118_C5 = CLBLL_L_X4Y120_SLICE_X5Y120_BO5;
  assign CLBLM_L_X10Y122_SLICE_X12Y122_B1 = CLBLM_R_X7Y119_SLICE_X9Y119_DO6;
  assign CLBLM_L_X10Y122_SLICE_X12Y122_B2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y122_SLICE_X12Y122_B3 = CLBLM_L_X10Y119_SLICE_X13Y119_AQ;
  assign CLBLM_L_X10Y122_SLICE_X12Y122_B4 = CLBLM_L_X10Y123_SLICE_X12Y123_AO6;
  assign CLBLM_L_X10Y122_SLICE_X12Y122_B5 = CLBLM_L_X10Y122_SLICE_X12Y122_CO5;
  assign CLBLM_L_X10Y122_SLICE_X12Y122_B6 = CLBLM_L_X8Y122_SLICE_X10Y122_CO6;
  assign CLBLM_L_X8Y112_SLICE_X11Y112_D2 = CLBLM_L_X12Y115_SLICE_X16Y115_CQ;
  assign CLBLL_L_X4Y118_SLICE_X4Y118_D1 = CLBLL_L_X4Y116_SLICE_X4Y116_AQ;
  assign CLBLL_L_X4Y118_SLICE_X4Y118_D2 = 1'b1;
  assign CLBLL_L_X4Y118_SLICE_X4Y118_D3 = CLBLL_L_X4Y118_SLICE_X5Y118_DO6;
  assign CLBLM_L_X10Y122_SLICE_X12Y122_C2 = 1'b1;
  assign CLBLM_L_X10Y122_SLICE_X12Y122_C3 = CLBLM_R_X7Y124_SLICE_X8Y124_AQ;
  assign CLBLM_L_X10Y122_SLICE_X12Y122_C4 = 1'b1;
  assign CLBLL_L_X4Y118_SLICE_X4Y118_D5 = CLBLM_R_X3Y121_SLICE_X2Y121_AO6;
  assign CLBLM_L_X8Y112_SLICE_X10Y112_A1 = CLBLM_R_X11Y114_SLICE_X14Y114_BQ;
  assign CLBLM_L_X8Y112_SLICE_X10Y112_A2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y112_SLICE_X10Y112_A3 = CLBLM_L_X8Y112_SLICE_X10Y112_AQ;
  assign CLBLM_L_X8Y112_SLICE_X10Y112_A4 = CLBLM_R_X7Y112_SLICE_X9Y112_BQ;
  assign CLBLM_L_X8Y112_SLICE_X10Y112_A5 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X8Y112_SLICE_X10Y112_A6 = CLBLM_L_X10Y113_SLICE_X12Y113_DO6;
  assign CLBLM_L_X8Y112_SLICE_X10Y112_B1 = CLBLM_R_X7Y112_SLICE_X8Y112_CQ;
  assign CLBLM_L_X8Y112_SLICE_X10Y112_B2 = CLBLM_L_X8Y112_SLICE_X10Y112_BQ;
  assign CLBLM_L_X8Y112_SLICE_X10Y112_B3 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X8Y112_SLICE_X10Y112_B4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y112_SLICE_X10Y112_B5 = CLBLM_L_X10Y113_SLICE_X12Y113_DO6;
  assign CLBLM_L_X8Y112_SLICE_X10Y112_B6 = CLBLM_R_X11Y113_SLICE_X15Y113_AQ;
  assign CLBLM_L_X10Y122_SLICE_X12Y122_D3 = CLBLM_L_X8Y122_SLICE_X11Y122_DO6;
  assign CLBLM_L_X10Y122_SLICE_X12Y122_D4 = CLBLM_L_X10Y123_SLICE_X12Y123_CO6;
  assign CLBLM_L_X10Y122_SLICE_X12Y122_D5 = CLBLM_R_X11Y121_SLICE_X14Y121_BO6;
  assign CLBLM_L_X10Y122_SLICE_X12Y122_D6 = CLBLM_L_X8Y120_SLICE_X11Y120_BQ;
  assign CLBLM_L_X10Y122_SLICE_X12Y122_D1 = CLBLM_L_X10Y122_SLICE_X13Y122_AQ;
  assign CLBLM_L_X10Y122_SLICE_X12Y122_D2 = CLBLM_R_X11Y121_SLICE_X14Y121_BO5;
  assign CLBLM_L_X8Y112_SLICE_X10Y112_C2 = CLBLM_L_X8Y112_SLICE_X10Y112_CQ;
  assign CLBLM_L_X8Y112_SLICE_X10Y112_C1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y112_SLICE_X10Y112_C3 = 1'b1;
  assign CLBLM_L_X8Y112_SLICE_X10Y112_C4 = CLBLM_L_X8Y112_SLICE_X10Y112_BQ;
  assign CLBLM_L_X8Y112_SLICE_X10Y112_C5 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLL_L_X4Y118_SLICE_X5Y118_A1 = CLBLM_R_X7Y119_SLICE_X9Y119_BQ;
  assign CLBLL_L_X4Y118_SLICE_X5Y118_A2 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLL_L_X4Y118_SLICE_X5Y118_A3 = CLBLL_L_X4Y118_SLICE_X5Y118_AQ;
  assign CLBLL_L_X4Y118_SLICE_X5Y118_A4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLL_L_X4Y118_SLICE_X5Y118_A5 = CLBLM_R_X3Y118_SLICE_X2Y118_AQ;
  assign CLBLL_L_X4Y118_SLICE_X5Y118_A6 = CLBLM_R_X5Y110_SLICE_X7Y110_BQ;
  assign CLBLM_L_X8Y112_SLICE_X10Y112_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLL_L_X4Y118_SLICE_X5Y118_B1 = CLBLM_L_X10Y113_SLICE_X13Y113_BO6;
  assign CLBLL_L_X4Y118_SLICE_X5Y118_B2 = CLBLL_L_X4Y118_SLICE_X5Y118_BQ;
  assign CLBLL_L_X4Y118_SLICE_X5Y118_B3 = CLBLM_R_X3Y111_SLICE_X3Y111_BQ;
  assign CLBLL_L_X4Y118_SLICE_X5Y118_B4 = CLBLM_R_X5Y122_SLICE_X6Y122_AQ;
  assign CLBLL_L_X4Y118_SLICE_X5Y118_B5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLL_L_X4Y118_SLICE_X5Y118_B6 = CLBLM_R_X7Y119_SLICE_X8Y119_D5Q;
  assign CLBLM_L_X8Y112_SLICE_X10Y112_D3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y112_SLICE_X10Y112_D4 = CLBLM_L_X10Y116_SLICE_X13Y116_CQ;
  assign CLBLM_L_X8Y112_SLICE_X10Y112_D5 = 1'b1;
  assign CLBLM_L_X8Y112_SLICE_X10Y112_D6 = CLBLM_R_X7Y109_SLICE_X8Y109_BQ;
  assign CLBLL_L_X4Y118_SLICE_X5Y118_C3 = CLBLM_R_X7Y119_SLICE_X8Y119_D5Q;
  assign CLBLL_L_X4Y118_SLICE_X5Y118_C1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLL_L_X4Y118_SLICE_X5Y118_C2 = CLBLL_L_X4Y118_SLICE_X5Y118_CQ;
  assign CLBLL_L_X4Y118_SLICE_X5Y118_C4 = CLBLL_L_X4Y117_SLICE_X5Y117_CQ;
  assign CLBLL_L_X4Y118_SLICE_X5Y118_C5 = CLBLM_L_X10Y113_SLICE_X13Y113_BO6;
  assign CLBLL_L_X4Y118_SLICE_X5Y118_C6 = CLBLL_L_X4Y118_SLICE_X5Y118_AQ;
  assign CLBLL_L_X4Y118_SLICE_X5Y118_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLL_L_X4Y118_SLICE_X5Y118_D1 = CLBLM_L_X8Y118_SLICE_X11Y118_AQ;
  assign CLBLL_L_X4Y118_SLICE_X5Y118_D2 = CLBLM_R_X11Y116_SLICE_X14Y116_AQ;
  assign CLBLL_L_X4Y118_SLICE_X5Y118_D3 = CLBLL_L_X2Y122_SLICE_X1Y122_DO6;
  assign CLBLL_L_X4Y118_SLICE_X5Y118_D4 = RIOB33_X105Y131_IOB_X1Y131_I;
  assign CLBLL_L_X4Y118_SLICE_X5Y118_D5 = RIOB33_X105Y131_IOB_X1Y132_I;
  assign CLBLL_L_X4Y118_SLICE_X5Y118_D6 = CLBLM_R_X3Y122_SLICE_X3Y122_AO6;
  assign LIOI3_X0Y177_OLOGIC_X0Y178_T1 = 1'b1;
  assign LIOI3_X0Y117_OLOGIC_X0Y118_D1 = CLBLL_L_X4Y116_SLICE_X4Y116_CQ;
  assign CLBLM_R_X11Y116_SLICE_X15Y116_A1 = CLBLM_R_X7Y113_SLICE_X8Y113_DO6;
  assign CLBLM_R_X11Y116_SLICE_X15Y116_A2 = CLBLM_R_X3Y118_SLICE_X2Y118_AQ;
  assign CLBLM_R_X11Y116_SLICE_X15Y116_A3 = CLBLM_R_X11Y116_SLICE_X15Y116_AQ;
  assign CLBLM_R_X11Y116_SLICE_X15Y116_A4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X11Y116_SLICE_X15Y116_A5 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_R_X11Y116_SLICE_X15Y116_A6 = CLBLM_R_X11Y119_SLICE_X14Y119_AQ;
  assign LIOI3_X0Y117_OLOGIC_X0Y118_T1 = 1'b1;
  assign LIOI3_X0Y177_OLOGIC_X0Y177_D1 = RIOB33_X105Y129_IOB_X1Y129_I;
  assign CLBLM_L_X8Y117_SLICE_X11Y117_B1 = 1'b1;
  assign CLBLM_R_X11Y116_SLICE_X15Y116_B1 = 1'b1;
  assign CLBLM_R_X11Y116_SLICE_X15Y116_B2 = 1'b1;
  assign CLBLM_R_X11Y116_SLICE_X15Y116_B3 = 1'b1;
  assign CLBLM_R_X11Y116_SLICE_X15Y116_B4 = 1'b1;
  assign CLBLM_L_X8Y117_SLICE_X11Y117_B2 = CLBLM_L_X8Y117_SLICE_X11Y117_BQ;
  assign CLBLM_R_X11Y116_SLICE_X15Y116_B5 = 1'b1;
  assign CLBLM_R_X11Y116_SLICE_X15Y116_B6 = 1'b1;
  assign LIOI3_X0Y117_OLOGIC_X0Y117_D1 = CLBLL_L_X4Y119_SLICE_X4Y119_BQ;
  assign CLBLM_L_X8Y117_SLICE_X11Y117_B3 = CLBLM_R_X5Y111_SLICE_X7Y111_DO6;
  assign CLBLM_R_X11Y116_SLICE_X15Y116_C1 = 1'b1;
  assign CLBLM_R_X11Y116_SLICE_X15Y116_C2 = 1'b1;
  assign CLBLM_R_X11Y116_SLICE_X15Y116_C3 = 1'b1;
  assign CLBLM_R_X11Y116_SLICE_X15Y116_C4 = 1'b1;
  assign CLBLM_R_X11Y116_SLICE_X15Y116_C5 = 1'b1;
  assign CLBLM_R_X11Y116_SLICE_X15Y116_C6 = 1'b1;
  assign RIOI3_X105Y161_OLOGIC_X1Y162_T1 = 1'b1;
  assign CLBLM_R_X11Y116_SLICE_X15Y116_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X8Y117_SLICE_X11Y117_B5 = CLBLM_L_X10Y116_SLICE_X13Y116_AO5;
  assign LIOI3_X0Y117_OLOGIC_X0Y117_T1 = 1'b1;
  assign RIOI3_X105Y161_OLOGIC_X1Y161_D1 = CLBLM_R_X11Y119_SLICE_X14Y119_CO5;
  assign CLBLM_R_X5Y125_SLICE_X7Y125_C4 = 1'b1;
  assign CLBLM_R_X11Y116_SLICE_X15Y116_D1 = 1'b1;
  assign CLBLM_R_X11Y116_SLICE_X15Y116_D2 = 1'b1;
  assign CLBLM_R_X11Y116_SLICE_X15Y116_D3 = 1'b1;
  assign CLBLM_R_X11Y116_SLICE_X15Y116_D4 = 1'b1;
  assign CLBLM_R_X5Y125_SLICE_X7Y125_C5 = 1'b1;
  assign CLBLM_R_X11Y116_SLICE_X15Y116_D5 = 1'b1;
  assign CLBLM_R_X11Y116_SLICE_X15Y116_D6 = 1'b1;
  assign CLBLM_R_X5Y125_SLICE_X7Y125_C6 = 1'b1;
  assign RIOI3_X105Y161_OLOGIC_X1Y161_T1 = 1'b1;
  assign CLBLM_R_X11Y116_SLICE_X14Y116_A1 = CLBLM_L_X10Y119_SLICE_X12Y119_CQ;
  assign CLBLM_R_X11Y116_SLICE_X14Y116_A2 = 1'b1;
  assign CLBLM_R_X11Y116_SLICE_X14Y116_A3 = CLBLM_R_X11Y116_SLICE_X14Y116_AQ;
  assign CLBLM_R_X11Y116_SLICE_X14Y116_A4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X11Y116_SLICE_X14Y116_A5 = CLBLM_L_X10Y116_SLICE_X12Y116_BQ;
  assign CLBLM_R_X11Y116_SLICE_X14Y116_A6 = CLBLM_R_X11Y121_SLICE_X14Y121_CO6;
  assign CLBLM_R_X11Y116_SLICE_X14Y116_B1 = CLBLM_R_X7Y119_SLICE_X9Y119_AQ;
  assign CLBLM_R_X11Y116_SLICE_X14Y116_B2 = CLBLM_R_X7Y120_SLICE_X9Y120_DQ;
  assign CLBLM_R_X11Y116_SLICE_X14Y116_B3 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X7Y123_SLICE_X8Y123_B5 = CLBLM_L_X10Y124_SLICE_X13Y124_BO6;
  assign CLBLM_R_X11Y116_SLICE_X14Y116_B4 = CLBLM_L_X8Y119_SLICE_X10Y119_CQ;
  assign CLBLM_R_X11Y116_SLICE_X14Y116_B5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X11Y116_SLICE_X14Y116_B6 = 1'b1;
  assign CLBLM_L_X8Y117_SLICE_X11Y117_C2 = CLBLM_L_X8Y117_SLICE_X11Y117_CQ;
  assign CLBLM_R_X7Y123_SLICE_X8Y123_B6 = CLBLM_R_X7Y122_SLICE_X8Y122_AQ;
  assign CLBLM_R_X11Y116_SLICE_X14Y116_C1 = CLBLM_L_X10Y116_SLICE_X12Y116_BQ;
  assign CLBLM_L_X8Y117_SLICE_X11Y117_C3 = CLBLM_R_X3Y118_SLICE_X2Y118_AQ;
  assign CLBLM_R_X11Y116_SLICE_X14Y116_C2 = CLBLM_R_X11Y116_SLICE_X14Y116_CQ;
  assign CLBLM_R_X11Y116_SLICE_X14Y116_C3 = CLBLM_L_X12Y115_SLICE_X16Y115_DQ;
  assign CLBLM_R_X11Y116_SLICE_X14Y116_C4 = CLBLM_R_X11Y119_SLICE_X14Y119_AO6;
  assign CLBLM_R_X11Y116_SLICE_X14Y116_C5 = CLBLM_L_X10Y116_SLICE_X13Y116_CO5;
  assign CLBLM_L_X8Y117_SLICE_X11Y117_C4 = CLBLM_R_X7Y120_SLICE_X9Y120_CQ;
  assign CLBLM_R_X11Y116_SLICE_X14Y116_C6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign RIOI3_TBYTETERM_X105Y187_OLOGIC_X1Y187_T1 = 1'b1;
  assign CLBLM_R_X11Y116_SLICE_X14Y116_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X11Y116_SLICE_X14Y116_D1 = CLBLM_R_X11Y118_SLICE_X15Y118_AQ;
  assign CLBLM_R_X11Y116_SLICE_X14Y116_D2 = 1'b1;
  assign CLBLM_R_X11Y116_SLICE_X14Y116_D3 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X11Y116_SLICE_X14Y116_D4 = CLBLL_L_X4Y114_SLICE_X5Y114_AQ;
  assign CLBLM_R_X11Y116_SLICE_X14Y116_D5 = 1'b1;
  assign CLBLM_R_X11Y116_SLICE_X14Y116_D6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y115_SLICE_X12Y115_B4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X5Y125_SLICE_X7Y125_D2 = 1'b1;
  assign CLBLM_L_X10Y115_SLICE_X12Y115_B5 = CLBLM_L_X10Y117_SLICE_X12Y117_AQ;
  assign CLBLM_L_X10Y115_SLICE_X12Y115_B6 = CLBLM_L_X8Y121_SLICE_X10Y121_CQ;
  assign CLBLM_R_X7Y123_SLICE_X8Y123_C4 = 1'b1;
  assign CLBLM_R_X5Y125_SLICE_X7Y125_D5 = 1'b1;
  assign CLBLM_R_X7Y123_SLICE_X8Y123_C5 = CLBLM_L_X10Y126_SLICE_X12Y126_AQ;
  assign CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_S0 = 1'b1;
  assign CLBLM_R_X5Y125_SLICE_X7Y125_D6 = 1'b1;
  assign CLBLM_R_X7Y123_SLICE_X8Y123_C6 = CLBLM_R_X11Y121_SLICE_X14Y121_CO6;
  assign CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_S1 = 1'b1;
  assign RIOB33_X105Y161_IOB_X1Y162_O = CLBLM_R_X11Y117_SLICE_X14Y117_DO6;
  assign RIOB33_X105Y161_IOB_X1Y161_O = CLBLM_R_X11Y119_SLICE_X14Y119_CO5;
  assign CLBLM_L_X10Y115_SLICE_X12Y115_C5 = CLBLM_L_X10Y117_SLICE_X13Y117_DQ;
  assign CLBLM_L_X10Y115_SLICE_X12Y115_C6 = CLBLM_R_X7Y114_SLICE_X8Y114_BQ;
  assign CLBLM_L_X10Y123_SLICE_X13Y123_A1 = CLBLM_L_X10Y124_SLICE_X13Y124_BO5;
  assign CLBLM_L_X10Y123_SLICE_X13Y123_A2 = CLBLM_L_X10Y124_SLICE_X13Y124_AO5;
  assign CLBLM_L_X10Y123_SLICE_X13Y123_A3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y123_SLICE_X13Y123_A4 = 1'b1;
  assign CLBLM_L_X10Y123_SLICE_X13Y123_A5 = CLBLM_L_X10Y120_SLICE_X13Y120_A5Q;
  assign CLBLM_L_X10Y123_SLICE_X13Y123_A6 = CLBLM_L_X10Y123_SLICE_X13Y123_CO6;
  assign CLBLM_L_X8Y128_SLICE_X11Y128_C3 = 1'b1;
  assign CLBLM_L_X10Y123_SLICE_X13Y123_B1 = CLBLM_L_X10Y123_SLICE_X12Y123_AO5;
  assign CLBLM_L_X10Y123_SLICE_X13Y123_B2 = CLBLM_R_X7Y123_SLICE_X9Y123_CO6;
  assign CLBLM_L_X10Y123_SLICE_X13Y123_B3 = RIOB33_X105Y121_IOB_X1Y121_I;
  assign CLBLM_L_X10Y123_SLICE_X13Y123_B4 = CLBLM_L_X10Y118_SLICE_X12Y118_B5Q;
  assign CLBLM_L_X10Y115_SLICE_X12Y115_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X10Y123_SLICE_X13Y123_B5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y123_SLICE_X13Y123_B6 = CLBLM_L_X8Y121_SLICE_X10Y121_AQ;
  assign CLBLM_R_X7Y123_SLICE_X8Y123_D2 = 1'b1;
  assign CLBLM_R_X7Y123_SLICE_X8Y123_D3 = 1'b1;
  assign CLBLM_L_X10Y123_SLICE_X13Y123_C1 = CLBLM_R_X11Y123_SLICE_X14Y123_BO6;
  assign CLBLM_L_X10Y123_SLICE_X13Y123_C2 = CLBLM_L_X10Y123_SLICE_X12Y123_CO6;
  assign CLBLM_L_X10Y123_SLICE_X13Y123_C3 = CLBLM_R_X11Y123_SLICE_X14Y123_AO6;
  assign CLBLM_L_X8Y113_SLICE_X11Y113_A4 = CLBLM_L_X10Y113_SLICE_X12Y113_DO6;
  assign CLBLM_L_X8Y113_SLICE_X11Y113_A5 = CLBLL_L_X4Y121_SLICE_X4Y121_AQ;
  assign CLBLM_L_X10Y123_SLICE_X13Y123_C4 = CLBLM_L_X10Y123_SLICE_X13Y123_AQ;
  assign CLBLM_L_X10Y123_SLICE_X13Y123_C5 = CLBLM_L_X8Y122_SLICE_X11Y122_DO6;
  assign CLBLM_L_X10Y123_SLICE_X13Y123_C6 = CLBLM_L_X8Y121_SLICE_X10Y121_AQ;
  assign CLBLM_L_X10Y123_SLICE_X13Y123_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X8Y113_SLICE_X11Y113_A1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLL_L_X4Y119_SLICE_X4Y119_A1 = 1'b1;
  assign CLBLL_L_X4Y119_SLICE_X4Y119_A2 = CLBLM_R_X5Y120_SLICE_X7Y120_AQ;
  assign CLBLL_L_X4Y119_SLICE_X4Y119_A3 = CLBLL_L_X4Y119_SLICE_X4Y119_AQ;
  assign CLBLM_L_X8Y113_SLICE_X11Y113_A6 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X10Y123_SLICE_X13Y123_D1 = CLBLM_R_X11Y123_SLICE_X14Y123_AO6;
  assign CLBLM_L_X10Y123_SLICE_X13Y123_D2 = CLBLM_L_X10Y122_SLICE_X13Y122_CQ;
  assign CLBLM_L_X10Y123_SLICE_X13Y123_D3 = CLBLM_L_X8Y122_SLICE_X11Y122_DO6;
  assign CLBLM_L_X10Y123_SLICE_X13Y123_D4 = CLBLM_R_X11Y123_SLICE_X14Y123_BO5;
  assign CLBLM_L_X10Y123_SLICE_X13Y123_D5 = CLBLM_L_X10Y123_SLICE_X13Y123_AQ;
  assign CLBLM_L_X10Y123_SLICE_X13Y123_D6 = CLBLM_L_X10Y121_SLICE_X13Y121_BQ;
  assign CLBLL_L_X4Y119_SLICE_X4Y119_B2 = CLBLL_L_X4Y119_SLICE_X4Y119_BQ;
  assign CLBLM_L_X8Y113_SLICE_X11Y113_B6 = CLBLL_L_X4Y115_SLICE_X4Y115_BQ;
  assign CLBLL_L_X4Y119_SLICE_X4Y119_B5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLL_L_X4Y119_SLICE_X4Y119_B6 = 1'b1;
  assign CLBLM_L_X8Y113_SLICE_X11Y113_C1 = CLBLM_R_X7Y111_SLICE_X9Y111_AO6;
  assign CLBLL_L_X4Y119_SLICE_X4Y119_C1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y123_SLICE_X12Y123_A1 = CLBLM_R_X7Y123_SLICE_X9Y123_BO5;
  assign CLBLM_L_X10Y123_SLICE_X12Y123_A2 = CLBLM_R_X7Y124_SLICE_X8Y124_AQ;
  assign CLBLM_L_X10Y123_SLICE_X12Y123_A3 = CLBLM_R_X5Y120_SLICE_X6Y120_A5Q;
  assign CLBLM_L_X10Y123_SLICE_X12Y123_A4 = CLBLM_L_X10Y124_SLICE_X12Y124_AQ;
  assign CLBLM_L_X10Y123_SLICE_X12Y123_A5 = CLBLM_R_X7Y120_SLICE_X9Y120_A5Q;
  assign CLBLM_L_X10Y123_SLICE_X12Y123_A6 = 1'b1;
  assign CLBLL_L_X4Y119_SLICE_X4Y119_C5 = CLBLL_L_X2Y117_SLICE_X0Y117_A5Q;
  assign CLBLL_L_X4Y119_SLICE_X4Y119_C6 = 1'b1;
  assign CLBLL_L_X4Y119_SLICE_X4Y119_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X10Y123_SLICE_X12Y123_B1 = CLBLM_L_X8Y122_SLICE_X11Y122_DO6;
  assign CLBLM_L_X10Y123_SLICE_X12Y123_B2 = CLBLM_L_X10Y122_SLICE_X13Y122_BQ;
  assign CLBLM_L_X10Y123_SLICE_X12Y123_B3 = CLBLM_L_X10Y122_SLICE_X13Y122_AQ;
  assign CLBLM_L_X10Y123_SLICE_X12Y123_B4 = CLBLM_L_X8Y121_SLICE_X11Y121_BQ;
  assign CLBLM_L_X10Y123_SLICE_X12Y123_B5 = CLBLM_R_X11Y121_SLICE_X14Y121_BO6;
  assign CLBLM_L_X10Y123_SLICE_X12Y123_B6 = CLBLM_R_X11Y121_SLICE_X14Y121_BO5;
  assign CLBLL_L_X4Y119_SLICE_X4Y119_D1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLL_L_X4Y119_SLICE_X4Y119_D2 = CLBLM_R_X3Y116_SLICE_X2Y116_DO6;
  assign CLBLL_L_X4Y119_SLICE_X4Y119_D3 = CLBLL_L_X4Y119_SLICE_X4Y119_DQ;
  assign CLBLL_L_X4Y119_SLICE_X4Y119_D4 = 1'b1;
  assign CLBLL_L_X4Y119_SLICE_X4Y119_D5 = CLBLL_L_X4Y119_SLICE_X4Y119_B5Q;
  assign CLBLL_L_X4Y119_SLICE_X4Y119_D6 = CLBLM_R_X11Y119_SLICE_X15Y119_AQ;
  assign CLBLM_L_X8Y113_SLICE_X10Y113_A1 = CLBLM_L_X8Y113_SLICE_X10Y113_DO6;
  assign CLBLM_L_X10Y123_SLICE_X12Y123_C4 = CLBLM_R_X7Y120_SLICE_X9Y120_A5Q;
  assign CLBLM_L_X8Y113_SLICE_X10Y113_A2 = CLBLL_L_X4Y112_SLICE_X4Y112_AQ;
  assign CLBLM_L_X10Y123_SLICE_X12Y123_C6 = CLBLM_R_X7Y124_SLICE_X8Y124_AQ;
  assign CLBLM_L_X8Y113_SLICE_X10Y113_A3 = 1'b1;
  assign CLBLM_L_X8Y113_SLICE_X10Y113_A4 = CLBLM_L_X8Y113_SLICE_X11Y113_BQ;
  assign CLBLM_L_X8Y113_SLICE_X10Y113_A5 = 1'b1;
  assign CLBLM_L_X8Y113_SLICE_X10Y113_A6 = CLBLM_L_X8Y113_SLICE_X10Y113_CO6;
  assign CLBLM_L_X10Y115_SLICE_X12Y115_D6 = CLBLM_R_X7Y119_SLICE_X8Y119_BQ;
  assign CLBLM_L_X8Y113_SLICE_X10Y113_B1 = 1'b1;
  assign CLBLM_L_X8Y113_SLICE_X10Y113_B2 = CLBLL_L_X4Y112_SLICE_X4Y112_AQ;
  assign CLBLM_L_X8Y113_SLICE_X10Y113_B3 = CLBLM_R_X7Y112_SLICE_X9Y112_AQ;
  assign CLBLM_L_X8Y113_SLICE_X10Y113_B4 = CLBLM_R_X5Y118_SLICE_X6Y118_BQ;
  assign CLBLM_L_X8Y113_SLICE_X10Y113_B5 = CLBLM_L_X8Y114_SLICE_X10Y114_AQ;
  assign CLBLM_L_X10Y123_SLICE_X12Y123_D2 = 1'b1;
  assign CLBLM_L_X10Y123_SLICE_X12Y123_D3 = CLBLM_L_X10Y121_SLICE_X13Y121_BQ;
  assign CLBLM_L_X10Y123_SLICE_X12Y123_D4 = CLBLM_L_X10Y123_SLICE_X12Y123_CO6;
  assign CLBLM_L_X10Y123_SLICE_X12Y123_D5 = 1'b1;
  assign CLBLM_L_X8Y113_SLICE_X10Y113_C2 = CLBLM_R_X7Y112_SLICE_X9Y112_AQ;
  assign CLBLM_L_X10Y123_SLICE_X12Y123_D6 = CLBLM_L_X10Y123_SLICE_X12Y123_BO6;
  assign CLBLM_L_X8Y113_SLICE_X10Y113_B6 = 1'b1;
  assign CLBLM_L_X8Y113_SLICE_X10Y113_C1 = CLBLM_L_X8Y114_SLICE_X10Y114_AQ;
  assign CLBLL_L_X4Y119_SLICE_X5Y119_A1 = CLBLM_R_X5Y120_SLICE_X6Y120_A5Q;
  assign CLBLM_L_X8Y113_SLICE_X10Y113_C3 = 1'b1;
  assign CLBLM_L_X8Y113_SLICE_X10Y113_C4 = CLBLM_L_X8Y112_SLICE_X10Y112_AQ;
  assign CLBLM_L_X8Y113_SLICE_X10Y113_C5 = 1'b1;
  assign CLBLM_L_X8Y113_SLICE_X10Y113_C6 = CLBLM_R_X11Y113_SLICE_X15Y113_AQ;
  assign CLBLL_L_X4Y119_SLICE_X5Y119_A3 = CLBLL_L_X4Y119_SLICE_X5Y119_AQ;
  assign CLBLL_L_X4Y119_SLICE_X5Y119_A4 = 1'b1;
  assign CLBLL_L_X4Y119_SLICE_X5Y119_A5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLL_L_X4Y119_SLICE_X5Y119_B5 = CLBLL_L_X4Y116_SLICE_X5Y116_AQ;
  assign CLBLL_L_X4Y119_SLICE_X5Y119_B6 = CLBLM_R_X7Y118_SLICE_X8Y118_CQ;
  assign CLBLL_L_X4Y119_SLICE_X5Y119_B1 = CLBLL_L_X4Y121_SLICE_X4Y121_DO5;
  assign CLBLL_L_X4Y119_SLICE_X5Y119_B2 = CLBLL_L_X4Y120_SLICE_X5Y120_BO6;
  assign CLBLL_L_X4Y119_SLICE_X5Y119_B3 = CLBLL_L_X4Y119_SLICE_X5Y119_AQ;
  assign CLBLM_L_X8Y113_SLICE_X10Y113_D1 = CLBLM_L_X8Y112_SLICE_X10Y112_BQ;
  assign CLBLM_L_X8Y113_SLICE_X10Y113_D2 = CLBLM_L_X8Y117_SLICE_X10Y117_BQ;
  assign CLBLM_L_X8Y113_SLICE_X10Y113_D3 = 1'b1;
  assign CLBLM_L_X8Y113_SLICE_X10Y113_D4 = CLBLM_R_X11Y113_SLICE_X14Y113_AQ;
  assign CLBLM_L_X8Y113_SLICE_X10Y113_D5 = 1'b1;
  assign CLBLM_L_X8Y113_SLICE_X10Y113_D6 = CLBLM_R_X5Y118_SLICE_X6Y118_BQ;
  assign CLBLL_L_X4Y119_SLICE_X5Y119_C1 = CLBLM_R_X3Y122_SLICE_X3Y122_AO6;
  assign CLBLL_L_X4Y119_SLICE_X5Y119_C4 = CLBLM_R_X7Y120_SLICE_X8Y120_AQ;
  assign CLBLL_L_X4Y119_SLICE_X5Y119_C5 = RIOB33_X105Y133_IOB_X1Y134_I;
  assign CLBLL_L_X4Y119_SLICE_X5Y119_C6 = RIOB33_X105Y131_IOB_X1Y131_I;
  assign CLBLL_L_X4Y119_SLICE_X5Y119_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X5Y125_SLICE_X6Y125_C4 = CLBLM_R_X7Y124_SLICE_X8Y124_CQ;
  assign CLBLL_L_X4Y119_SLICE_X5Y119_D1 = CLBLL_L_X2Y116_SLICE_X1Y116_AQ;
  assign CLBLL_L_X4Y119_SLICE_X5Y119_D2 = CLBLM_R_X5Y119_SLICE_X6Y119_DO6;
  assign CLBLL_L_X4Y119_SLICE_X5Y119_D3 = CLBLL_L_X4Y120_SLICE_X5Y120_BO5;
  assign CLBLL_L_X4Y119_SLICE_X5Y119_D4 = CLBLL_L_X4Y119_SLICE_X5Y119_CO6;
  assign CLBLL_L_X4Y119_SLICE_X5Y119_D5 = CLBLM_R_X3Y121_SLICE_X2Y121_AO5;
  assign CLBLL_L_X4Y119_SLICE_X5Y119_D6 = CLBLM_L_X8Y116_SLICE_X11Y116_AQ;
  assign CLBLM_R_X5Y125_SLICE_X6Y125_C5 = CLBLM_R_X7Y124_SLICE_X8Y124_BQ;
  assign CLBLM_R_X5Y125_SLICE_X6Y125_C6 = 1'b1;
  assign CLBLM_L_X8Y117_SLICE_X10Y117_C1 = CLBLM_L_X8Y117_SLICE_X10Y117_CQ;
  assign CLBLM_R_X11Y117_SLICE_X15Y117_A1 = CLBLM_R_X11Y118_SLICE_X15Y118_BQ;
  assign CLBLM_R_X11Y117_SLICE_X15Y117_A2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X11Y117_SLICE_X15Y117_A3 = CLBLM_R_X11Y117_SLICE_X15Y117_AQ;
  assign CLBLM_R_X11Y117_SLICE_X15Y117_A4 = CLBLM_R_X11Y119_SLICE_X14Y119_AO6;
  assign CLBLM_R_X11Y117_SLICE_X15Y117_A5 = CLBLM_L_X12Y119_SLICE_X17Y119_AO5;
  assign CLBLM_R_X11Y117_SLICE_X15Y117_A6 = CLBLM_L_X8Y117_SLICE_X11Y117_DQ;
  assign CLBLM_R_X11Y117_SLICE_X15Y117_B1 = 1'b1;
  assign CLBLM_R_X11Y117_SLICE_X15Y117_B2 = 1'b1;
  assign CLBLM_L_X8Y117_SLICE_X10Y117_C4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X11Y117_SLICE_X15Y117_B3 = 1'b1;
  assign CLBLM_R_X11Y117_SLICE_X15Y117_B4 = 1'b1;
  assign CLBLM_R_X11Y117_SLICE_X15Y117_B5 = 1'b1;
  assign CLBLM_R_X11Y117_SLICE_X15Y117_B6 = 1'b1;
  assign CLBLM_L_X8Y117_SLICE_X10Y117_C5 = CLBLM_L_X10Y117_SLICE_X12Y117_BQ;
  assign CLBLM_R_X11Y117_SLICE_X15Y117_C1 = 1'b1;
  assign CLBLM_R_X11Y117_SLICE_X15Y117_C2 = 1'b1;
  assign CLBLM_L_X8Y117_SLICE_X10Y117_C6 = CLBLM_R_X11Y115_SLICE_X14Y115_CQ;
  assign CLBLM_R_X11Y117_SLICE_X15Y117_C3 = 1'b1;
  assign CLBLM_R_X11Y117_SLICE_X15Y117_C4 = 1'b1;
  assign CLBLM_R_X11Y117_SLICE_X15Y117_C5 = 1'b1;
  assign CLBLM_R_X11Y117_SLICE_X15Y117_C6 = 1'b1;
  assign CLBLM_R_X11Y117_SLICE_X15Y117_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X11Y117_SLICE_X15Y117_D1 = 1'b1;
  assign CLBLM_R_X11Y117_SLICE_X15Y117_D2 = 1'b1;
  assign CLBLM_R_X11Y117_SLICE_X15Y117_D3 = 1'b1;
  assign CLBLM_L_X10Y126_SLICE_X12Y126_B3 = 1'b1;
  assign CLBLM_R_X11Y117_SLICE_X15Y117_D4 = 1'b1;
  assign CLBLM_R_X11Y117_SLICE_X15Y117_D5 = 1'b1;
  assign CLBLM_R_X11Y117_SLICE_X15Y117_D6 = 1'b1;
  assign CLBLM_L_X8Y117_SLICE_X10Y117_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X11Y117_SLICE_X14Y117_A1 = CLBLL_L_X4Y113_SLICE_X4Y113_AQ;
  assign CLBLM_R_X11Y117_SLICE_X14Y117_A2 = CLBLM_R_X11Y119_SLICE_X14Y119_AO6;
  assign CLBLM_R_X11Y117_SLICE_X14Y117_A3 = CLBLM_R_X11Y117_SLICE_X14Y117_AQ;
  assign CLBLM_R_X11Y117_SLICE_X14Y117_A4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X11Y117_SLICE_X14Y117_A5 = CLBLM_L_X10Y118_SLICE_X13Y118_AQ;
  assign CLBLM_R_X11Y117_SLICE_X14Y117_A6 = CLBLM_L_X12Y119_SLICE_X17Y119_AO5;
  assign CLBLM_R_X11Y117_SLICE_X14Y117_B1 = CLBLM_L_X8Y110_SLICE_X10Y110_AQ;
  assign CLBLM_R_X11Y117_SLICE_X14Y117_B2 = CLBLM_R_X11Y117_SLICE_X14Y117_BQ;
  assign CLBLM_R_X11Y117_SLICE_X14Y117_B3 = 1'b1;
  assign CLBLM_R_X11Y117_SLICE_X14Y117_B4 = CLBLM_R_X7Y117_SLICE_X8Y117_BQ;
  assign CLBLM_R_X11Y117_SLICE_X14Y117_B5 = CLBLM_R_X5Y111_SLICE_X7Y111_DO6;
  assign CLBLM_R_X11Y117_SLICE_X14Y117_B6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X11Y117_SLICE_X14Y117_C1 = CLBLM_R_X11Y118_SLICE_X14Y118_AQ;
  assign CLBLM_R_X11Y117_SLICE_X14Y117_C2 = CLBLM_R_X11Y117_SLICE_X14Y117_CQ;
  assign CLBLM_R_X11Y117_SLICE_X14Y117_C3 = CLBLM_R_X7Y113_SLICE_X9Y113_CO6;
  assign CLBLM_R_X11Y117_SLICE_X14Y117_C4 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_R_X11Y117_SLICE_X14Y117_C5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X11Y117_SLICE_X14Y117_C6 = CLBLM_R_X3Y118_SLICE_X2Y118_AQ;
  assign CLBLM_R_X11Y117_SLICE_X14Y117_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X11Y117_SLICE_X14Y117_D1 = CLBLM_R_X11Y115_SLICE_X15Y115_AQ;
  assign CLBLM_R_X11Y117_SLICE_X14Y117_D2 = CLBLM_R_X11Y117_SLICE_X14Y117_CQ;
  assign CLBLM_R_X11Y117_SLICE_X14Y117_D3 = CLBLM_R_X3Y117_SLICE_X3Y117_BQ;
  assign CLBLM_R_X11Y117_SLICE_X14Y117_D4 = CLBLM_L_X8Y117_SLICE_X11Y117_DQ;
  assign CLBLM_R_X11Y117_SLICE_X14Y117_D5 = CLBLL_L_X4Y111_SLICE_X4Y111_AQ;
  assign CLBLM_R_X11Y117_SLICE_X14Y117_D6 = 1'b1;
  assign CLBLL_L_X4Y123_SLICE_X4Y123_B3 = CLBLL_L_X2Y113_SLICE_X1Y113_C5Q;
  assign RIOB33_X105Y163_IOB_X1Y164_O = CLBLM_R_X7Y119_SLICE_X9Y119_DO5;
  assign RIOB33_X105Y163_IOB_X1Y163_O = CLBLM_R_X11Y117_SLICE_X14Y117_DO5;
  assign CLBLL_L_X4Y123_SLICE_X4Y123_B4 = CLBLL_L_X4Y119_SLICE_X4Y119_C5Q;
  assign CLBLL_L_X4Y123_SLICE_X4Y123_B5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLL_L_X4Y123_SLICE_X4Y123_B6 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLL_L_X4Y123_SLICE_X4Y123_C1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLL_L_X4Y123_SLICE_X4Y123_C2 = CLBLL_L_X4Y117_SLICE_X5Y117_DQ;
  assign CLBLM_L_X10Y124_SLICE_X13Y124_A1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y124_SLICE_X13Y124_A2 = CLBLM_L_X10Y123_SLICE_X13Y123_DO6;
  assign CLBLM_L_X10Y124_SLICE_X13Y124_A3 = CLBLM_L_X10Y120_SLICE_X13Y120_A5Q;
  assign CLBLM_L_X10Y124_SLICE_X13Y124_A4 = CLBLM_L_X10Y120_SLICE_X13Y120_AQ;
  assign CLBLM_L_X10Y124_SLICE_X13Y124_A5 = CLBLM_L_X10Y124_SLICE_X13Y124_CO5;
  assign CLBLM_L_X10Y124_SLICE_X13Y124_A6 = 1'b1;
  assign LIOB33_X0Y195_IOB_X0Y195_O = LIOB33_X0Y63_IOB_X0Y64_I;
  assign LIOB33_X0Y195_IOB_X0Y196_O = LIOB33_X0Y69_IOB_X0Y69_I;
  assign CLBLM_L_X10Y124_SLICE_X13Y124_AX = CLBLM_L_X10Y118_SLICE_X12Y118_B5Q;
  assign CLBLM_L_X10Y124_SLICE_X13Y124_B1 = CLBLM_R_X7Y124_SLICE_X8Y124_AQ;
  assign CLBLM_L_X10Y124_SLICE_X13Y124_B2 = CLBLM_L_X10Y123_SLICE_X13Y123_DO6;
  assign CLBLM_L_X10Y124_SLICE_X13Y124_B3 = CLBLM_R_X7Y120_SLICE_X9Y120_A5Q;
  assign CLBLM_L_X10Y124_SLICE_X13Y124_B4 = CLBLM_R_X5Y120_SLICE_X6Y120_A5Q;
  assign CLBLM_L_X10Y124_SLICE_X13Y124_B5 = CLBLM_L_X10Y124_SLICE_X12Y124_AQ;
  assign CLBLM_L_X10Y124_SLICE_X13Y124_B6 = 1'b1;
  assign CLBLL_L_X4Y120_SLICE_X4Y120_A1 = CLBLM_R_X5Y121_SLICE_X6Y121_DO6;
  assign CLBLL_L_X4Y120_SLICE_X4Y120_A2 = CLBLL_L_X4Y118_SLICE_X4Y118_BO6;
  assign CLBLL_L_X4Y120_SLICE_X4Y120_A3 = CLBLM_R_X3Y123_SLICE_X2Y123_BO6;
  assign CLBLM_L_X10Y124_SLICE_X13Y124_C1 = CLBLM_R_X5Y120_SLICE_X6Y120_A5Q;
  assign CLBLM_L_X10Y124_SLICE_X13Y124_C2 = CLBLM_R_X7Y124_SLICE_X8Y124_AQ;
  assign CLBLM_L_X10Y124_SLICE_X13Y124_C3 = CLBLM_L_X10Y118_SLICE_X12Y118_B5Q;
  assign CLBLM_L_X8Y114_SLICE_X11Y114_A4 = CLBLM_L_X10Y112_SLICE_X12Y112_CQ;
  assign CLBLM_L_X10Y124_SLICE_X13Y124_C4 = CLBLM_R_X7Y120_SLICE_X9Y120_A5Q;
  assign CLBLM_L_X10Y124_SLICE_X13Y124_C5 = CLBLM_L_X10Y124_SLICE_X12Y124_AQ;
  assign CLBLM_L_X10Y124_SLICE_X13Y124_C6 = 1'b1;
  assign CLBLM_L_X10Y124_SLICE_X13Y124_CE = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y124_SLICE_X13Y124_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLL_L_X4Y120_SLICE_X4Y120_A5 = CLBLM_R_X5Y120_SLICE_X6Y120_CO6;
  assign CLBLL_L_X4Y120_SLICE_X4Y120_A6 = CLBLL_L_X4Y120_SLICE_X4Y120_CO6;
  assign CLBLL_L_X4Y120_SLICE_X4Y120_B6 = CLBLL_L_X4Y121_SLICE_X5Y121_CO5;
  assign CLBLM_L_X8Y114_SLICE_X11Y114_B3 = CLBLM_L_X8Y114_SLICE_X11Y114_AQ;
  assign CLBLM_L_X8Y114_SLICE_X11Y114_B5 = 1'b1;
  assign CLBLL_L_X4Y120_SLICE_X4Y120_C1 = RIOB33_X105Y107_IOB_X1Y107_I;
  assign CLBLM_L_X10Y124_SLICE_X13Y124_D1 = 1'b1;
  assign CLBLM_L_X10Y124_SLICE_X13Y124_D2 = 1'b1;
  assign CLBLL_L_X4Y120_SLICE_X4Y120_C4 = CLBLM_R_X7Y118_SLICE_X8Y118_BQ;
  assign CLBLM_L_X10Y124_SLICE_X13Y124_D3 = 1'b1;
  assign CLBLL_L_X4Y120_SLICE_X4Y120_C6 = CLBLM_R_X3Y122_SLICE_X2Y122_BO5;
  assign CLBLM_L_X10Y124_SLICE_X13Y124_D4 = 1'b1;
  assign CLBLM_L_X10Y124_SLICE_X13Y124_D5 = 1'b1;
  assign CLBLM_L_X10Y124_SLICE_X13Y124_D6 = 1'b1;
  assign CLBLM_L_X10Y124_SLICE_X13Y124_SR = CLBLM_R_X11Y123_SLICE_X14Y123_CO6;
  assign CLBLM_L_X10Y124_SLICE_X12Y124_A1 = CLBLM_L_X8Y121_SLICE_X11Y121_DQ;
  assign CLBLM_L_X10Y124_SLICE_X12Y124_A2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y124_SLICE_X12Y124_A3 = CLBLM_L_X10Y124_SLICE_X12Y124_AQ;
  assign CLBLM_L_X10Y124_SLICE_X12Y124_A4 = CLBLM_L_X10Y124_SLICE_X13Y124_CO6;
  assign CLBLM_L_X10Y124_SLICE_X12Y124_A5 = RIOB33_X105Y121_IOB_X1Y121_I;
  assign CLBLM_L_X10Y124_SLICE_X12Y124_A6 = CLBLM_L_X10Y123_SLICE_X13Y123_DO6;
  assign CLBLM_L_X8Y114_SLICE_X11Y114_C6 = CLBLM_L_X8Y114_SLICE_X10Y114_BQ;
  assign CLBLM_L_X8Y114_SLICE_X11Y114_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLL_L_X4Y120_SLICE_X4Y120_D1 = RIOB33_X105Y107_IOB_X1Y108_I;
  assign CLBLL_L_X4Y120_SLICE_X4Y120_D2 = CLBLL_L_X2Y122_SLICE_X0Y122_AO6;
  assign CLBLM_L_X10Y124_SLICE_X12Y124_B2 = 1'b1;
  assign CLBLM_L_X10Y124_SLICE_X12Y124_B3 = 1'b1;
  assign CLBLM_L_X10Y124_SLICE_X12Y124_B4 = 1'b1;
  assign CLBLM_L_X10Y124_SLICE_X12Y124_B5 = 1'b1;
  assign CLBLM_L_X10Y124_SLICE_X12Y124_B6 = 1'b1;
  assign CLBLM_L_X8Y114_SLICE_X11Y114_D2 = CLBLM_L_X8Y114_SLICE_X11Y114_CQ;
  assign CLBLM_L_X8Y114_SLICE_X11Y114_D3 = CLBLM_L_X8Y115_SLICE_X11Y115_DQ;
  assign CLBLM_L_X8Y114_SLICE_X11Y114_D4 = CLBLM_L_X8Y120_SLICE_X11Y120_CQ;
  assign CLBLM_L_X8Y114_SLICE_X11Y114_D5 = 1'b1;
  assign CLBLM_L_X8Y114_SLICE_X11Y114_D6 = 1'b1;
  assign CLBLM_L_X8Y114_SLICE_X10Y114_A1 = CLBLM_L_X8Y117_SLICE_X10Y117_CQ;
  assign CLBLM_L_X10Y124_SLICE_X12Y124_C3 = 1'b1;
  assign CLBLM_L_X10Y124_SLICE_X12Y124_C4 = 1'b1;
  assign CLBLM_L_X10Y124_SLICE_X12Y124_C5 = 1'b1;
  assign CLBLM_L_X8Y114_SLICE_X10Y114_A2 = CLBLM_L_X8Y114_SLICE_X10Y114_DQ;
  assign CLBLM_L_X8Y114_SLICE_X10Y114_A3 = CLBLM_L_X8Y114_SLICE_X10Y114_AQ;
  assign CLBLM_L_X8Y114_SLICE_X10Y114_A4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y114_SLICE_X10Y114_A5 = CLBLM_R_X3Y118_SLICE_X2Y118_AQ;
  assign CLBLM_L_X8Y114_SLICE_X10Y114_A6 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_L_X8Y114_SLICE_X10Y114_B1 = CLBLM_R_X11Y115_SLICE_X14Y115_CQ;
  assign CLBLM_L_X8Y114_SLICE_X10Y114_B2 = CLBLM_L_X8Y112_SLICE_X10Y112_DQ;
  assign CLBLM_L_X8Y114_SLICE_X10Y114_B3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y114_SLICE_X10Y114_B4 = CLBLM_R_X3Y116_SLICE_X3Y116_BQ;
  assign CLBLM_L_X10Y124_SLICE_X12Y124_D1 = 1'b1;
  assign CLBLM_L_X10Y124_SLICE_X12Y124_D2 = 1'b1;
  assign CLBLM_L_X10Y124_SLICE_X12Y124_D3 = 1'b1;
  assign CLBLM_L_X10Y124_SLICE_X12Y124_D4 = 1'b1;
  assign CLBLM_L_X10Y124_SLICE_X12Y124_D5 = 1'b1;
  assign CLBLM_L_X10Y124_SLICE_X12Y124_D6 = 1'b1;
  assign CLBLM_L_X8Y114_SLICE_X10Y114_C3 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X8Y114_SLICE_X10Y114_C4 = CLBLM_L_X8Y114_SLICE_X11Y114_CQ;
  assign CLBLL_L_X4Y120_SLICE_X5Y120_A1 = CLBLL_L_X2Y120_SLICE_X0Y120_CO6;
  assign CLBLM_L_X8Y114_SLICE_X10Y114_C6 = 1'b1;
  assign CLBLL_L_X4Y120_SLICE_X5Y120_A3 = CLBLL_L_X4Y120_SLICE_X4Y120_AO6;
  assign CLBLL_L_X4Y120_SLICE_X5Y120_A4 = 1'b1;
  assign CLBLL_L_X4Y120_SLICE_X5Y120_A5 = CLBLL_L_X2Y119_SLICE_X0Y119_BO6;
  assign CLBLL_L_X4Y120_SLICE_X5Y120_A6 = 1'b1;
  assign CLBLL_L_X4Y120_SLICE_X5Y120_B1 = RIOB33_X105Y131_IOB_X1Y132_I;
  assign CLBLL_L_X4Y120_SLICE_X5Y120_B2 = CLBLM_R_X3Y122_SLICE_X3Y122_AO6;
  assign CLBLL_L_X4Y120_SLICE_X5Y120_B3 = RIOB33_X105Y133_IOB_X1Y134_I;
  assign CLBLM_L_X8Y114_SLICE_X10Y114_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLL_L_X4Y120_SLICE_X5Y120_B4 = RIOB33_X105Y131_IOB_X1Y131_I;
  assign CLBLL_L_X4Y120_SLICE_X5Y120_C2 = CLBLM_R_X3Y122_SLICE_X2Y122_BO5;
  assign CLBLL_L_X4Y120_SLICE_X5Y120_B5 = RIOB33_X105Y133_IOB_X1Y133_I;
  assign CLBLL_L_X4Y120_SLICE_X5Y120_B6 = 1'b1;
  assign CLBLM_L_X8Y114_SLICE_X10Y114_D1 = CLBLM_R_X3Y118_SLICE_X2Y118_AQ;
  assign CLBLM_L_X8Y114_SLICE_X10Y114_D2 = CLBLM_R_X5Y115_SLICE_X7Y115_CO6;
  assign CLBLM_L_X8Y114_SLICE_X10Y114_D3 = CLBLM_L_X8Y114_SLICE_X10Y114_DQ;
  assign CLBLM_L_X8Y114_SLICE_X10Y114_D4 = CLBLL_L_X4Y116_SLICE_X5Y116_DQ;
  assign CLBLM_L_X8Y114_SLICE_X10Y114_D5 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLL_L_X4Y120_SLICE_X5Y120_C6 = CLBLL_L_X4Y120_SLICE_X5Y120_BO6;
  assign CLBLM_L_X8Y114_SLICE_X10Y114_D6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLL_L_X4Y120_SLICE_X5Y120_D1 = CLBLL_L_X4Y122_SLICE_X5Y122_CO6;
  assign CLBLL_L_X4Y120_SLICE_X5Y120_D2 = CLBLM_R_X5Y120_SLICE_X6Y120_DO6;
  assign CLBLL_L_X4Y120_SLICE_X5Y120_D3 = CLBLL_L_X4Y119_SLICE_X5Y119_DO6;
  assign CLBLL_L_X4Y120_SLICE_X5Y120_D4 = CLBLL_L_X2Y121_SLICE_X1Y121_DO6;
  assign CLBLL_L_X4Y120_SLICE_X5Y120_D5 = CLBLL_L_X4Y122_SLICE_X4Y122_CO6;
  assign CLBLL_L_X4Y120_SLICE_X5Y120_D6 = CLBLL_L_X4Y117_SLICE_X4Y117_DO6;
  assign CLBLM_R_X11Y118_SLICE_X15Y118_A1 = CLBLM_R_X11Y118_SLICE_X15Y118_DO6;
  assign CLBLM_R_X11Y118_SLICE_X15Y118_A2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X11Y118_SLICE_X15Y118_A3 = 1'b1;
  assign CLBLM_R_X11Y118_SLICE_X15Y118_A4 = CLBLM_L_X12Y120_SLICE_X17Y120_CO5;
  assign CLBLM_R_X11Y118_SLICE_X15Y118_A5 = CLBLM_L_X8Y117_SLICE_X10Y117_AQ;
  assign CLBLM_R_X11Y118_SLICE_X15Y118_A6 = 1'b1;
  assign CLBLM_R_X11Y118_SLICE_X15Y118_B1 = CLBLM_R_X5Y116_SLICE_X7Y116_AQ;
  assign CLBLM_R_X11Y118_SLICE_X15Y118_B2 = CLBLM_R_X11Y118_SLICE_X15Y118_BQ;
  assign CLBLM_R_X11Y118_SLICE_X15Y118_B3 = CLBLM_R_X11Y117_SLICE_X14Y117_AQ;
  assign CLBLM_R_X11Y118_SLICE_X15Y118_B4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X11Y118_SLICE_X15Y118_B5 = CLBLM_R_X11Y119_SLICE_X14Y119_AO6;
  assign CLBLM_R_X11Y118_SLICE_X15Y118_B6 = CLBLM_L_X12Y119_SLICE_X17Y119_AO5;
  assign CLBLM_R_X11Y118_SLICE_X15Y118_C1 = CLBLL_L_X4Y114_SLICE_X4Y114_AQ;
  assign CLBLM_R_X11Y118_SLICE_X15Y118_C2 = CLBLM_R_X11Y119_SLICE_X14Y119_AO6;
  assign CLBLM_R_X11Y118_SLICE_X15Y118_C3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X11Y118_SLICE_X15Y118_C4 = CLBLM_L_X10Y118_SLICE_X13Y118_BQ;
  assign CLBLM_R_X11Y118_SLICE_X15Y118_C5 = CLBLM_L_X12Y119_SLICE_X17Y119_AO5;
  assign CLBLM_R_X11Y118_SLICE_X15Y118_C6 = CLBLM_R_X11Y118_SLICE_X15Y118_CQ;
  assign CLBLM_R_X11Y118_SLICE_X15Y118_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X11Y118_SLICE_X15Y118_D1 = 1'b1;
  assign CLBLM_R_X11Y118_SLICE_X15Y118_D2 = CLBLM_R_X11Y120_SLICE_X14Y120_AO5;
  assign CLBLM_R_X11Y118_SLICE_X15Y118_D3 = CLBLM_L_X12Y119_SLICE_X17Y119_DO6;
  assign CLBLM_R_X11Y118_SLICE_X15Y118_D4 = CLBLM_R_X11Y118_SLICE_X14Y118_DO5;
  assign CLBLM_R_X11Y118_SLICE_X15Y118_D5 = CLBLM_L_X10Y120_SLICE_X12Y120_CQ;
  assign CLBLM_R_X11Y118_SLICE_X15Y118_D6 = CLBLM_R_X11Y118_SLICE_X15Y118_AQ;
  assign CLBLM_R_X11Y118_SLICE_X14Y118_A1 = CLBLM_R_X11Y118_SLICE_X14Y118_DO6;
  assign CLBLM_R_X11Y118_SLICE_X14Y118_A2 = CLBLM_R_X3Y116_SLICE_X2Y116_AQ;
  assign CLBLM_R_X11Y118_SLICE_X14Y118_A3 = CLBLM_R_X11Y118_SLICE_X14Y118_AQ;
  assign CLBLM_R_X11Y118_SLICE_X14Y118_A4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X11Y118_SLICE_X14Y118_A5 = CLBLM_L_X10Y116_SLICE_X12Y116_DO5;
  assign CLBLM_R_X11Y118_SLICE_X14Y118_A6 = CLBLM_R_X11Y119_SLICE_X14Y119_AO6;
  assign CLBLM_R_X11Y118_SLICE_X14Y118_B1 = CLBLM_R_X11Y120_SLICE_X14Y120_DO6;
  assign CLBLM_R_X11Y118_SLICE_X14Y118_B2 = CLBLM_R_X11Y118_SLICE_X14Y118_BQ;
  assign CLBLM_R_X11Y118_SLICE_X14Y118_B3 = RIOB33_X105Y121_IOB_X1Y121_I;
  assign CLBLM_R_X11Y118_SLICE_X14Y118_B4 = CLBLM_R_X11Y119_SLICE_X14Y119_AO6;
  assign CLBLM_R_X11Y118_SLICE_X14Y118_B5 = CLBLM_R_X11Y115_SLICE_X14Y115_AQ;
  assign CLBLM_R_X11Y118_SLICE_X14Y118_B6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X11Y118_SLICE_X14Y118_C1 = CLBLM_L_X8Y114_SLICE_X10Y114_BQ;
  assign CLBLM_R_X11Y118_SLICE_X14Y118_C2 = CLBLM_R_X11Y118_SLICE_X14Y118_CQ;
  assign CLBLM_R_X11Y118_SLICE_X14Y118_C3 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_R_X11Y118_SLICE_X14Y118_C4 = CLBLM_R_X5Y115_SLICE_X7Y115_CO6;
  assign CLBLM_R_X11Y118_SLICE_X14Y118_C5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X11Y118_SLICE_X14Y118_C6 = CLBLM_R_X3Y118_SLICE_X2Y118_AQ;
  assign CLBLM_R_X11Y118_SLICE_X14Y118_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X11Y118_SLICE_X14Y118_D1 = CLBLM_L_X10Y116_SLICE_X12Y116_DO5;
  assign CLBLM_R_X11Y118_SLICE_X14Y118_D2 = CLBLM_R_X11Y118_SLICE_X14Y118_AQ;
  assign CLBLM_R_X11Y118_SLICE_X14Y118_D3 = CLBLM_L_X10Y119_SLICE_X13Y119_AQ;
  assign CLBLM_R_X11Y118_SLICE_X14Y118_D4 = CLBLM_R_X11Y118_SLICE_X14Y118_BQ;
  assign CLBLM_R_X11Y118_SLICE_X14Y118_D5 = CLBLM_R_X11Y120_SLICE_X14Y120_BO5;
  assign CLBLM_R_X11Y118_SLICE_X14Y118_D6 = 1'b1;
  assign LIOI3_X0Y179_OLOGIC_X0Y180_D1 = RIOB33_X105Y131_IOB_X1Y132_I;
  assign RIOB33_X105Y165_IOB_X1Y166_O = RIOB33_SING_X105Y149_IOB_X1Y149_I;
  assign RIOB33_X105Y165_IOB_X1Y165_O = RIOB33_X105Y125_IOB_X1Y125_I;
  assign CLBLL_L_X4Y123_SLICE_X5Y123_A1 = 1'b1;
  assign LIOI3_X0Y179_OLOGIC_X0Y180_T1 = 1'b1;
  assign LIOI3_X0Y121_OLOGIC_X0Y122_D1 = CLBLM_R_X5Y121_SLICE_X6Y121_A5Q;
  assign CLBLL_L_X4Y123_SLICE_X5Y123_A4 = RIOB33_X105Y133_IOB_X1Y133_I;
  assign LIOI3_X0Y179_OLOGIC_X0Y179_D1 = RIOB33_X105Y131_IOB_X1Y131_I;
  assign CLBLL_L_X4Y123_SLICE_X5Y123_A5 = RIOB33_X105Y133_IOB_X1Y134_I;
  assign LIOI3_X0Y121_OLOGIC_X0Y122_T1 = 1'b1;
  assign RIOI3_X105Y165_OLOGIC_X1Y166_D1 = RIOB33_SING_X105Y149_IOB_X1Y149_I;
  assign CLBLL_L_X4Y123_SLICE_X5Y123_A6 = 1'b1;
  assign LIOI3_X0Y179_OLOGIC_X0Y179_T1 = 1'b1;
  assign LIOI3_X0Y121_OLOGIC_X0Y121_D1 = CLBLM_L_X8Y123_SLICE_X11Y123_A5Q;
  assign RIOI3_X105Y165_OLOGIC_X1Y166_T1 = 1'b1;
  assign LIOB33_X0Y197_IOB_X0Y198_O = LIOB33_X0Y73_IOB_X0Y73_I;
  assign LIOB33_X0Y197_IOB_X0Y197_O = LIOB33_X0Y71_IOB_X0Y72_I;
  assign LIOI3_X0Y121_OLOGIC_X0Y121_T1 = 1'b1;
  assign RIOI3_X105Y165_OLOGIC_X1Y165_D1 = RIOB33_X105Y125_IOB_X1Y125_I;
  assign CLBLL_L_X4Y123_SLICE_X5Y123_B1 = 1'b1;
  assign CLBLL_L_X4Y123_SLICE_X5Y123_B2 = 1'b1;
  assign CLBLL_L_X4Y123_SLICE_X5Y123_B3 = 1'b1;
  assign RIOI3_X105Y165_OLOGIC_X1Y165_T1 = 1'b1;
  assign CLBLL_L_X4Y123_SLICE_X5Y123_B4 = 1'b1;
  assign CLBLL_L_X4Y123_SLICE_X5Y123_B5 = 1'b1;
  assign CLBLM_R_X13Y120_SLICE_X19Y120_B2 = 1'b1;
  assign CLBLL_L_X4Y123_SLICE_X5Y123_B6 = 1'b1;
  assign CLBLL_L_X4Y121_SLICE_X4Y121_A1 = 1'b1;
  assign CLBLL_L_X4Y121_SLICE_X4Y121_A2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLL_L_X4Y121_SLICE_X4Y121_A3 = CLBLL_L_X4Y121_SLICE_X4Y121_AQ;
  assign CLBLL_L_X4Y121_SLICE_X4Y121_A4 = CLBLM_R_X5Y124_SLICE_X6Y124_BQ;
  assign CLBLL_L_X4Y121_SLICE_X4Y121_A5 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLL_L_X4Y121_SLICE_X4Y121_A6 = CLBLL_L_X4Y115_SLICE_X4Y115_CQ;
  assign CLBLM_L_X8Y115_SLICE_X11Y115_A1 = CLBLM_L_X10Y111_SLICE_X13Y111_AQ;
  assign CLBLM_L_X8Y115_SLICE_X11Y115_A2 = CLBLM_R_X5Y119_SLICE_X7Y119_AO6;
  assign CLBLM_L_X8Y115_SLICE_X11Y115_A3 = CLBLM_L_X8Y115_SLICE_X11Y115_AQ;
  assign CLBLM_L_X8Y115_SLICE_X11Y115_A4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y115_SLICE_X11Y115_A5 = 1'b1;
  assign CLBLM_L_X8Y115_SLICE_X11Y115_A6 = CLBLM_R_X7Y116_SLICE_X9Y116_AQ;
  assign CLBLL_L_X4Y121_SLICE_X4Y121_B1 = CLBLM_R_X5Y122_SLICE_X6Y122_AQ;
  assign CLBLL_L_X4Y121_SLICE_X4Y121_B2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLL_L_X4Y121_SLICE_X4Y121_B3 = CLBLM_L_X8Y115_SLICE_X11Y115_BQ;
  assign CLBLL_L_X4Y121_SLICE_X4Y121_B4 = CLBLM_R_X7Y120_SLICE_X8Y120_CQ;
  assign CLBLL_L_X4Y121_SLICE_X4Y121_C1 = RIOB33_X105Y133_IOB_X1Y133_I;
  assign CLBLL_L_X4Y121_SLICE_X4Y121_C2 = CLBLM_R_X3Y122_SLICE_X3Y122_AO6;
  assign CLBLL_L_X4Y121_SLICE_X4Y121_B5 = CLBLM_R_X5Y121_SLICE_X6Y121_B5Q;
  assign CLBLL_L_X4Y121_SLICE_X4Y121_C4 = RIOB33_X105Y131_IOB_X1Y132_I;
  assign CLBLL_L_X4Y121_SLICE_X4Y121_B6 = CLBLL_L_X4Y117_SLICE_X4Y117_BQ;
  assign CLBLL_L_X4Y121_SLICE_X4Y121_C6 = 1'b1;
  assign CLBLL_L_X4Y121_SLICE_X4Y121_C3 = RIOB33_X105Y131_IOB_X1Y131_I;
  assign CLBLL_L_X4Y121_SLICE_X4Y121_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLL_L_X4Y121_SLICE_X4Y121_C5 = RIOB33_X105Y133_IOB_X1Y134_I;
  assign CLBLM_L_X8Y115_SLICE_X11Y115_C2 = CLBLM_R_X7Y119_SLICE_X9Y119_CQ;
  assign CLBLM_L_X8Y115_SLICE_X11Y115_C3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y115_SLICE_X11Y115_B5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y115_SLICE_X11Y115_B6 = CLBLM_L_X10Y115_SLICE_X12Y115_CQ;
  assign CLBLM_L_X8Y115_SLICE_X11Y115_C6 = 1'b1;
  assign CLBLM_L_X8Y115_SLICE_X11Y115_C1 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLL_L_X4Y121_SLICE_X4Y121_D1 = RIOB33_X105Y133_IOB_X1Y133_I;
  assign CLBLL_L_X4Y121_SLICE_X4Y121_D2 = CLBLM_R_X3Y122_SLICE_X3Y122_AO6;
  assign CLBLL_L_X4Y121_SLICE_X4Y121_D3 = RIOB33_X105Y131_IOB_X1Y131_I;
  assign CLBLL_L_X4Y121_SLICE_X4Y121_D4 = RIOB33_X105Y131_IOB_X1Y132_I;
  assign CLBLL_L_X4Y121_SLICE_X4Y121_D5 = RIOB33_X105Y133_IOB_X1Y134_I;
  assign CLBLL_L_X4Y121_SLICE_X4Y121_D6 = 1'b1;
  assign CLBLM_L_X8Y115_SLICE_X11Y115_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X8Y115_SLICE_X11Y115_D1 = CLBLM_L_X8Y115_SLICE_X11Y115_C5Q;
  assign CLBLM_L_X8Y115_SLICE_X11Y115_D4 = CLBLM_L_X10Y120_SLICE_X12Y120_BQ;
  assign CLBLM_L_X8Y115_SLICE_X11Y115_D2 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X8Y115_SLICE_X11Y115_D3 = 1'b1;
  assign CLBLM_L_X8Y115_SLICE_X11Y115_D5 = 1'b1;
  assign CLBLM_L_X8Y115_SLICE_X11Y115_D6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y126_SLICE_X13Y126_A6 = 1'b1;
  assign CLBLM_L_X8Y115_SLICE_X10Y115_A1 = CLBLM_L_X8Y115_SLICE_X10Y115_BO5;
  assign CLBLM_L_X8Y115_SLICE_X10Y115_A2 = 1'b1;
  assign CLBLM_L_X8Y115_SLICE_X10Y115_A3 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X8Y115_SLICE_X10Y115_A4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y115_SLICE_X10Y115_A5 = CLBLL_L_X4Y115_SLICE_X5Y115_CQ;
  assign CLBLM_L_X8Y115_SLICE_X10Y115_A6 = CLBLM_R_X7Y119_SLICE_X8Y119_BQ;
  assign CLBLM_L_X8Y115_SLICE_X10Y115_B1 = CLBLM_R_X7Y115_SLICE_X8Y115_CQ;
  assign CLBLM_L_X8Y115_SLICE_X10Y115_B2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y115_SLICE_X10Y115_B3 = RIOB33_X105Y121_IOB_X1Y121_I;
  assign CLBLM_L_X8Y115_SLICE_X10Y115_B4 = CLBLM_R_X7Y115_SLICE_X8Y115_AQ;
  assign CLBLL_L_X4Y121_SLICE_X5Y121_A1 = 1'b1;
  assign CLBLM_L_X8Y115_SLICE_X10Y115_B6 = 1'b1;
  assign CLBLL_L_X4Y121_SLICE_X5Y121_A2 = CLBLM_R_X7Y122_SLICE_X9Y122_BQ;
  assign CLBLM_L_X8Y115_SLICE_X10Y115_B5 = CLBLM_R_X11Y113_SLICE_X14Y113_AQ;
  assign CLBLL_L_X4Y121_SLICE_X5Y121_A3 = CLBLL_L_X4Y121_SLICE_X5Y121_AQ;
  assign CLBLL_L_X4Y121_SLICE_X5Y121_A4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLL_L_X4Y121_SLICE_X5Y121_A5 = CLBLL_L_X4Y119_SLICE_X4Y119_AQ;
  assign CLBLL_L_X4Y121_SLICE_X5Y121_A6 = CLBLM_R_X5Y115_SLICE_X6Y115_CO5;
  assign CLBLM_L_X8Y115_SLICE_X10Y115_C1 = CLBLM_R_X7Y122_SLICE_X9Y122_AQ;
  assign CLBLM_L_X8Y115_SLICE_X10Y115_C5 = CLBLM_L_X8Y114_SLICE_X10Y114_B5Q;
  assign CLBLM_L_X8Y115_SLICE_X10Y115_C6 = 1'b1;
  assign CLBLL_L_X4Y121_SLICE_X5Y121_B1 = RIOB33_X105Y129_IOB_X1Y129_I;
  assign CLBLL_L_X4Y121_SLICE_X5Y121_B2 = CLBLM_R_X7Y127_SLICE_X8Y127_AQ;
  assign CLBLL_L_X4Y121_SLICE_X5Y121_B3 = RIOB33_X105Y137_IOB_X1Y137_I;
  assign CLBLL_L_X4Y121_SLICE_X5Y121_B4 = CLBLL_L_X4Y120_SLICE_X5Y120_AO5;
  assign CLBLL_L_X4Y121_SLICE_X5Y121_C1 = CLBLM_L_X8Y121_SLICE_X10Y121_BQ;
  assign CLBLL_L_X4Y121_SLICE_X5Y121_B5 = CLBLM_R_X5Y120_SLICE_X7Y120_DO5;
  assign CLBLL_L_X4Y121_SLICE_X5Y121_B6 = 1'b1;
  assign CLBLL_L_X4Y121_SLICE_X5Y121_C2 = CLBLL_L_X4Y122_SLICE_X4Y122_AO5;
  assign CLBLL_L_X4Y121_SLICE_X5Y121_C3 = CLBLL_L_X4Y113_SLICE_X5Y113_AQ;
  assign CLBLL_L_X4Y121_SLICE_X5Y121_C4 = RIOB33_X105Y135_IOB_X1Y136_I;
  assign CLBLL_L_X4Y121_SLICE_X5Y121_C5 = RIOB33_X105Y131_IOB_X1Y131_I;
  assign CLBLL_L_X4Y121_SLICE_X5Y121_C6 = 1'b1;
  assign CLBLM_L_X8Y115_SLICE_X10Y115_D5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y115_SLICE_X10Y115_D6 = CLBLM_R_X7Y113_SLICE_X9Y113_CO6;
  assign CLBLL_L_X4Y121_SLICE_X5Y121_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X8Y115_SLICE_X10Y115_D1 = CLBLM_R_X3Y114_SLICE_X2Y114_AQ;
  assign CLBLM_L_X8Y115_SLICE_X10Y115_D2 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_L_X8Y115_SLICE_X10Y115_D3 = CLBLM_L_X8Y115_SLICE_X10Y115_DQ;
  assign CLBLM_L_X8Y115_SLICE_X10Y115_D4 = CLBLM_R_X3Y118_SLICE_X2Y118_AQ;
  assign CLBLL_L_X4Y121_SLICE_X5Y121_D1 = RIOB33_X105Y133_IOB_X1Y133_I;
  assign CLBLL_L_X4Y121_SLICE_X5Y121_D2 = RIOB33_X105Y131_IOB_X1Y132_I;
  assign CLBLL_L_X4Y121_SLICE_X5Y121_D3 = RIOB33_X105Y133_IOB_X1Y134_I;
  assign CLBLL_L_X4Y121_SLICE_X5Y121_D4 = CLBLM_R_X3Y122_SLICE_X3Y122_AO6;
  assign CLBLL_L_X4Y121_SLICE_X5Y121_D5 = RIOB33_X105Y131_IOB_X1Y131_I;
  assign CLBLL_L_X4Y121_SLICE_X5Y121_D6 = CLBLL_L_X4Y113_SLICE_X5Y113_BQ;
  assign CLBLM_R_X11Y119_SLICE_X15Y119_A1 = CLBLM_R_X11Y119_SLICE_X15Y119_DO6;
  assign CLBLM_R_X11Y119_SLICE_X15Y119_A2 = CLBLM_L_X12Y120_SLICE_X17Y120_CO5;
  assign CLBLM_R_X11Y119_SLICE_X15Y119_A3 = 1'b1;
  assign CLBLM_R_X11Y119_SLICE_X15Y119_A4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X11Y119_SLICE_X15Y119_A5 = 1'b1;
  assign CLBLM_R_X11Y119_SLICE_X15Y119_A6 = CLBLM_R_X7Y119_SLICE_X9Y119_AQ;
  assign CLBLM_R_X11Y119_SLICE_X15Y119_B1 = CLBLM_R_X5Y118_SLICE_X6Y118_CQ;
  assign CLBLM_R_X11Y119_SLICE_X15Y119_B2 = CLBLM_L_X12Y120_SLICE_X17Y120_CO5;
  assign CLBLM_R_X11Y119_SLICE_X15Y119_B3 = 1'b1;
  assign CLBLM_R_X11Y119_SLICE_X15Y119_B4 = CLBLM_L_X12Y119_SLICE_X16Y119_AO6;
  assign CLBLM_R_X11Y119_SLICE_X15Y119_B5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X11Y119_SLICE_X15Y119_B6 = CLBLM_R_X11Y120_SLICE_X14Y120_AO5;
  assign LIOI3_X0Y59_ILOGIC_X0Y60_D = LIOB33_X0Y59_IOB_X0Y60_I;
  assign LIOI3_X0Y59_ILOGIC_X0Y59_D = LIOB33_X0Y59_IOB_X0Y59_I;
  assign CLBLM_R_X7Y109_SLICE_X9Y109_A1 = 1'b1;
  assign CLBLM_R_X7Y109_SLICE_X9Y109_A2 = 1'b1;
  assign CLBLM_R_X7Y109_SLICE_X9Y109_A3 = 1'b1;
  assign CLBLM_R_X7Y109_SLICE_X9Y109_A4 = 1'b1;
  assign CLBLM_R_X7Y109_SLICE_X9Y109_A5 = 1'b1;
  assign CLBLM_R_X7Y109_SLICE_X9Y109_A6 = 1'b1;
  assign CLBLM_R_X11Y119_SLICE_X15Y119_C1 = CLBLM_L_X12Y120_SLICE_X16Y120_AO6;
  assign CLBLM_R_X11Y119_SLICE_X15Y119_C2 = CLBLM_R_X11Y119_SLICE_X15Y119_CQ;
  assign CLBLM_R_X11Y119_SLICE_X15Y119_C3 = RIOB33_X105Y121_IOB_X1Y121_I;
  assign CLBLM_R_X7Y109_SLICE_X9Y109_B1 = 1'b1;
  assign CLBLM_R_X7Y109_SLICE_X9Y109_B2 = 1'b1;
  assign CLBLM_R_X7Y109_SLICE_X9Y109_B3 = 1'b1;
  assign CLBLM_R_X7Y109_SLICE_X9Y109_B4 = 1'b1;
  assign CLBLM_R_X7Y109_SLICE_X9Y109_B5 = 1'b1;
  assign CLBLM_R_X7Y109_SLICE_X9Y109_B6 = 1'b1;
  assign CLBLM_R_X11Y119_SLICE_X15Y119_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X11Y119_SLICE_X15Y119_D5 = CLBLM_R_X11Y119_SLICE_X15Y119_AQ;
  assign CLBLM_R_X7Y109_SLICE_X9Y109_C1 = 1'b1;
  assign CLBLM_R_X7Y109_SLICE_X9Y109_C2 = 1'b1;
  assign CLBLM_R_X7Y109_SLICE_X9Y109_C3 = 1'b1;
  assign CLBLM_R_X7Y109_SLICE_X9Y109_C4 = 1'b1;
  assign CLBLM_R_X7Y109_SLICE_X9Y109_C5 = 1'b1;
  assign CLBLM_R_X7Y109_SLICE_X9Y109_C6 = 1'b1;
  assign CLBLM_R_X11Y119_SLICE_X15Y119_D6 = CLBLM_R_X11Y118_SLICE_X15Y118_BQ;
  assign CLBLM_R_X11Y119_SLICE_X14Y119_A1 = CLBLM_L_X10Y119_SLICE_X13Y119_AQ;
  assign CLBLM_R_X11Y119_SLICE_X14Y119_A2 = CLBLM_R_X11Y119_SLICE_X15Y119_CQ;
  assign CLBLM_R_X11Y119_SLICE_X14Y119_A3 = CLBLM_L_X10Y116_SLICE_X12Y116_DO5;
  assign CLBLM_R_X11Y119_SLICE_X14Y119_A4 = CLBLM_R_X13Y119_SLICE_X18Y119_CQ;
  assign CLBLM_R_X11Y119_SLICE_X14Y119_A5 = CLBLM_R_X11Y118_SLICE_X14Y118_BQ;
  assign CLBLM_R_X11Y119_SLICE_X14Y119_A6 = 1'b1;
  assign CLBLM_R_X7Y109_SLICE_X9Y109_D1 = 1'b1;
  assign CLBLM_R_X7Y109_SLICE_X9Y109_D2 = 1'b1;
  assign CLBLM_R_X7Y109_SLICE_X9Y109_D3 = 1'b1;
  assign CLBLM_R_X7Y109_SLICE_X9Y109_D4 = 1'b1;
  assign CLBLM_R_X7Y109_SLICE_X9Y109_D5 = 1'b1;
  assign CLBLM_R_X7Y109_SLICE_X9Y109_D6 = 1'b1;
  assign CLBLM_R_X11Y119_SLICE_X14Y119_AX = CLBLM_L_X10Y118_SLICE_X13Y118_BQ;
  assign CLBLM_R_X11Y119_SLICE_X14Y119_B1 = CLBLM_L_X10Y119_SLICE_X13Y119_AQ;
  assign CLBLM_R_X11Y119_SLICE_X14Y119_B2 = CLBLM_R_X11Y119_SLICE_X15Y119_CQ;
  assign CLBLM_R_X11Y119_SLICE_X14Y119_B3 = CLBLM_R_X7Y120_SLICE_X9Y120_AQ;
  assign CLBLM_R_X11Y119_SLICE_X14Y119_B4 = CLBLM_R_X13Y119_SLICE_X18Y119_CQ;
  assign CLBLM_R_X11Y119_SLICE_X14Y119_B5 = CLBLM_R_X11Y118_SLICE_X14Y118_BQ;
  assign CLBLM_R_X7Y109_SLICE_X8Y109_A1 = CLBLM_R_X7Y109_SLICE_X8Y109_CQ;
  assign CLBLM_R_X7Y109_SLICE_X8Y109_A2 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_R_X7Y109_SLICE_X8Y109_A3 = CLBLM_R_X7Y109_SLICE_X8Y109_AQ;
  assign CLBLM_R_X7Y109_SLICE_X8Y109_A4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y109_SLICE_X8Y109_A5 = 1'b1;
  assign CLBLM_R_X7Y109_SLICE_X8Y109_A6 = CLBLM_R_X3Y118_SLICE_X2Y118_AQ;
  assign CLBLM_R_X11Y119_SLICE_X14Y119_C1 = CLBLM_R_X5Y119_SLICE_X6Y119_AQ;
  assign CLBLM_R_X11Y119_SLICE_X14Y119_C2 = CLBLM_L_X10Y120_SLICE_X12Y120_AQ;
  assign CLBLM_R_X11Y119_SLICE_X14Y119_C3 = CLBLM_R_X11Y115_SLICE_X14Y115_DQ;
  assign CLBLM_R_X7Y109_SLICE_X8Y109_B1 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X7Y109_SLICE_X8Y109_B2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y109_SLICE_X8Y109_B3 = CLBLM_R_X5Y109_SLICE_X7Y109_AQ;
  assign CLBLL_L_X2Y109_SLICE_X0Y109_C4 = 1'b1;
  assign CLBLM_R_X7Y109_SLICE_X8Y109_B4 = CLBLM_R_X5Y110_SLICE_X7Y110_CQ;
  assign CLBLM_R_X7Y109_SLICE_X8Y109_B5 = 1'b1;
  assign CLBLM_R_X7Y109_SLICE_X8Y109_B6 = 1'b1;
  assign CLBLM_R_X11Y119_SLICE_X14Y119_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X11Y119_SLICE_X14Y119_D1 = CLBLM_R_X11Y118_SLICE_X15Y118_AQ;
  assign CLBLM_R_X7Y109_SLICE_X8Y109_C1 = CLBLM_R_X5Y111_SLICE_X6Y111_C5Q;
  assign CLBLM_R_X7Y109_SLICE_X8Y109_C2 = CLBLM_R_X7Y109_SLICE_X8Y109_CQ;
  assign CLBLM_R_X7Y109_SLICE_X8Y109_C3 = 1'b1;
  assign CLBLM_R_X7Y109_SLICE_X8Y109_C4 = 1'b1;
  assign CLBLM_R_X7Y109_SLICE_X8Y109_C5 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X7Y109_SLICE_X8Y109_C6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X11Y119_SLICE_X14Y119_D2 = CLBLM_L_X10Y119_SLICE_X13Y119_AQ;
  assign CLBLM_R_X11Y119_SLICE_X14Y119_D3 = CLBLM_R_X11Y120_SLICE_X15Y120_AQ;
  assign CLBLM_R_X11Y119_SLICE_X14Y119_D4 = CLBLM_R_X11Y119_SLICE_X15Y119_CQ;
  assign CLBLM_R_X7Y109_SLICE_X8Y109_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X11Y119_SLICE_X14Y119_D6 = CLBLM_R_X11Y118_SLICE_X14Y118_BQ;
  assign CLBLM_R_X11Y119_SLICE_X14Y119_SR = CLBLM_R_X11Y123_SLICE_X14Y123_CO6;
  assign CLBLM_R_X13Y120_SLICE_X19Y120_B3 = 1'b1;
  assign CLBLM_R_X13Y120_SLICE_X19Y120_B4 = 1'b1;
  assign CLBLM_R_X7Y109_SLICE_X8Y109_D1 = 1'b1;
  assign CLBLM_R_X7Y109_SLICE_X8Y109_D2 = 1'b1;
  assign CLBLM_R_X7Y109_SLICE_X8Y109_D3 = 1'b1;
  assign CLBLM_R_X7Y109_SLICE_X8Y109_D4 = 1'b1;
  assign CLBLM_R_X7Y109_SLICE_X8Y109_D5 = 1'b1;
  assign CLBLM_R_X7Y109_SLICE_X8Y109_D6 = 1'b1;
  assign CLBLM_R_X13Y120_SLICE_X19Y120_B5 = 1'b1;
  assign CLBLM_R_X13Y120_SLICE_X19Y120_B6 = 1'b1;
  assign CLBLM_L_X8Y128_SLICE_X11Y128_B3 = 1'b1;
  assign CLBLM_R_X103Y172_SLICE_X162Y172_D4 = 1'b1;
  assign CLBLM_L_X8Y128_SLICE_X11Y128_B6 = 1'b1;
  assign CLBLM_L_X10Y126_SLICE_X12Y126_A6 = 1'b1;
  assign CLBLM_R_X13Y120_SLICE_X19Y120_C5 = 1'b1;
  assign CLBLM_L_X8Y128_SLICE_X11Y128_C1 = 1'b1;
  assign CLBLM_L_X10Y126_SLICE_X13Y126_A1 = 1'b1;
  assign CLBLM_L_X8Y128_SLICE_X11Y128_C2 = 1'b1;
  assign CLBLM_L_X10Y126_SLICE_X13Y126_A2 = 1'b1;
  assign CLBLM_L_X10Y126_SLICE_X13Y126_A3 = 1'b1;
  assign CLBLM_L_X10Y126_SLICE_X13Y126_A4 = 1'b1;
  assign CLBLM_L_X10Y126_SLICE_X13Y126_A5 = 1'b1;
  assign CLBLL_L_X4Y122_SLICE_X4Y122_A1 = 1'b1;
  assign CLBLL_L_X4Y122_SLICE_X4Y122_A2 = RIOB33_X105Y131_IOB_X1Y132_I;
  assign CLBLL_L_X4Y122_SLICE_X4Y122_A3 = RIOB33_X105Y133_IOB_X1Y133_I;
  assign CLBLM_L_X10Y126_SLICE_X13Y126_B1 = 1'b1;
  assign CLBLM_L_X10Y126_SLICE_X13Y126_B2 = 1'b1;
  assign CLBLM_L_X10Y126_SLICE_X13Y126_B3 = 1'b1;
  assign CLBLM_L_X10Y126_SLICE_X13Y126_B4 = 1'b1;
  assign CLBLM_L_X10Y126_SLICE_X13Y126_B5 = 1'b1;
  assign CLBLM_L_X10Y126_SLICE_X13Y126_B6 = 1'b1;
  assign CLBLL_L_X4Y122_SLICE_X4Y122_A4 = CLBLM_R_X3Y122_SLICE_X3Y122_AO6;
  assign CLBLL_L_X4Y122_SLICE_X4Y122_A5 = RIOB33_X105Y133_IOB_X1Y134_I;
  assign CLBLL_L_X4Y122_SLICE_X4Y122_A6 = 1'b1;
  assign CLBLM_L_X10Y126_SLICE_X13Y126_C1 = 1'b1;
  assign CLBLL_L_X4Y122_SLICE_X4Y122_B6 = RIOB33_X105Y137_IOB_X1Y137_I;
  assign CLBLM_L_X10Y126_SLICE_X13Y126_C2 = 1'b1;
  assign CLBLM_L_X10Y126_SLICE_X13Y126_C3 = 1'b1;
  assign CLBLM_L_X10Y126_SLICE_X13Y126_C4 = 1'b1;
  assign CLBLM_L_X10Y126_SLICE_X13Y126_C5 = 1'b1;
  assign CLBLL_L_X4Y122_SLICE_X4Y122_C2 = CLBLL_L_X4Y123_SLICE_X4Y123_CQ;
  assign CLBLM_L_X10Y124_SLICE_X12Y124_C2 = 1'b1;
  assign CLBLM_L_X10Y126_SLICE_X13Y126_C6 = 1'b1;
  assign CLBLM_L_X8Y116_SLICE_X11Y116_A2 = CLBLM_R_X11Y121_SLICE_X14Y121_CO6;
  assign CLBLM_L_X8Y116_SLICE_X11Y116_A3 = CLBLM_L_X8Y116_SLICE_X11Y116_AQ;
  assign CLBLM_L_X8Y116_SLICE_X11Y116_A4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y116_SLICE_X11Y116_A6 = CLBLM_L_X8Y111_SLICE_X10Y111_AQ;
  assign CLBLM_L_X10Y126_SLICE_X13Y126_D1 = 1'b1;
  assign CLBLM_L_X10Y126_SLICE_X13Y126_D2 = 1'b1;
  assign CLBLM_L_X10Y126_SLICE_X13Y126_D3 = 1'b1;
  assign CLBLM_L_X10Y126_SLICE_X13Y126_D4 = 1'b1;
  assign CLBLM_L_X10Y126_SLICE_X13Y126_D5 = 1'b1;
  assign CLBLM_L_X10Y126_SLICE_X13Y126_D6 = 1'b1;
  assign CLBLM_L_X8Y116_SLICE_X11Y116_B3 = CLBLM_R_X7Y110_SLICE_X9Y110_BQ;
  assign CLBLM_L_X8Y116_SLICE_X11Y116_B5 = CLBLM_L_X8Y118_SLICE_X11Y118_AQ;
  assign CLBLM_L_X8Y116_SLICE_X11Y116_B6 = CLBLM_R_X5Y111_SLICE_X7Y111_DO6;
  assign CLBLM_L_X8Y116_SLICE_X11Y116_C1 = CLBLM_R_X11Y119_SLICE_X14Y119_AO6;
  assign CLBLM_L_X8Y116_SLICE_X11Y116_C2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y126_SLICE_X12Y126_A1 = 1'b1;
  assign CLBLM_L_X10Y126_SLICE_X12Y126_A2 = 1'b1;
  assign CLBLM_L_X10Y126_SLICE_X12Y126_A3 = 1'b1;
  assign CLBLM_L_X10Y126_SLICE_X12Y126_A4 = 1'b1;
  assign CLBLM_L_X10Y126_SLICE_X12Y126_A5 = 1'b1;
  assign CLBLM_L_X8Y116_SLICE_X11Y116_C5 = CLBLM_L_X8Y119_SLICE_X10Y119_BQ;
  assign CLBLM_L_X8Y116_SLICE_X11Y116_C6 = 1'b1;
  assign CLBLM_L_X8Y116_SLICE_X11Y116_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X8Y116_SLICE_X11Y116_D1 = CLBLM_R_X7Y116_SLICE_X8Y116_AQ;
  assign CLBLM_L_X8Y116_SLICE_X11Y116_D2 = 1'b1;
  assign CLBLM_L_X8Y116_SLICE_X11Y116_D3 = CLBLM_L_X8Y116_SLICE_X11Y116_DQ;
  assign CLBLM_L_X8Y116_SLICE_X11Y116_D5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y126_SLICE_X12Y126_B4 = 1'b1;
  assign CLBLM_L_X10Y126_SLICE_X12Y126_B5 = 1'b1;
  assign CLBLM_L_X10Y126_SLICE_X12Y126_B6 = 1'b1;
  assign CLBLM_L_X8Y116_SLICE_X11Y116_D6 = CLBLM_L_X10Y115_SLICE_X12Y115_DQ;
  assign CLBLM_L_X8Y116_SLICE_X11Y116_D4 = CLBLM_R_X5Y111_SLICE_X7Y111_DO6;
  assign CLBLM_L_X10Y126_SLICE_X12Y126_B1 = 1'b1;
  assign CLBLM_L_X10Y126_SLICE_X12Y126_B2 = 1'b1;
  assign CLBLL_L_X4Y113_SLICE_X4Y113_A5 = 1'b1;
  assign CLBLM_L_X10Y126_SLICE_X12Y126_C2 = 1'b1;
  assign CLBLM_L_X10Y126_SLICE_X12Y126_C3 = 1'b1;
  assign CLBLM_L_X10Y126_SLICE_X12Y126_C4 = 1'b1;
  assign CLBLM_L_X10Y126_SLICE_X12Y126_C5 = 1'b1;
  assign CLBLM_L_X10Y126_SLICE_X12Y126_C6 = 1'b1;
  assign CLBLM_L_X8Y116_SLICE_X10Y116_A1 = CLBLM_R_X7Y116_SLICE_X9Y116_CO6;
  assign CLBLM_L_X8Y116_SLICE_X10Y116_AX = CLBLM_R_X7Y116_SLICE_X8Y116_AQ;
  assign CLBLM_L_X8Y116_SLICE_X10Y116_A2 = CLBLM_R_X7Y115_SLICE_X9Y115_B5Q;
  assign CLBLM_L_X8Y116_SLICE_X10Y116_A3 = CLBLM_L_X8Y117_SLICE_X10Y117_AQ;
  assign CLBLM_L_X8Y116_SLICE_X10Y116_A4 = CLBLM_L_X8Y110_SLICE_X10Y110_CO6;
  assign CLBLM_L_X8Y128_SLICE_X11Y128_D3 = 1'b1;
  assign CLBLM_L_X8Y116_SLICE_X10Y116_A6 = CLBLM_L_X8Y116_SLICE_X10Y116_CO6;
  assign CLBLL_L_X4Y122_SLICE_X5Y122_A1 = RIOB33_X105Y135_IOB_X1Y135_I;
  assign CLBLL_L_X4Y122_SLICE_X5Y122_A2 = RIOB33_X105Y135_IOB_X1Y136_I;
  assign CLBLL_L_X4Y122_SLICE_X5Y122_A3 = RIOB33_X105Y131_IOB_X1Y131_I;
  assign CLBLL_L_X4Y122_SLICE_X5Y122_B1 = RIOB33_X105Y135_IOB_X1Y135_I;
  assign CLBLL_L_X4Y122_SLICE_X5Y122_B2 = CLBLL_L_X4Y121_SLICE_X5Y121_BO6;
  assign CLBLL_L_X4Y122_SLICE_X5Y122_B3 = CLBLM_R_X7Y113_SLICE_X9Y113_AQ;
  assign CLBLL_L_X4Y122_SLICE_X5Y122_B4 = CLBLL_L_X4Y123_SLICE_X5Y123_AO5;
  assign CLBLL_L_X4Y122_SLICE_X5Y122_B5 = RIOB33_X105Y129_IOB_X1Y130_I;
  assign CLBLM_L_X8Y116_SLICE_X10Y116_B4 = CLBLM_R_X7Y110_SLICE_X9Y110_BQ;
  assign CLBLM_L_X8Y116_SLICE_X10Y116_B5 = CLBLM_L_X8Y115_SLICE_X11Y115_AQ;
  assign CLBLM_L_X8Y116_SLICE_X10Y116_B6 = CLBLM_L_X10Y115_SLICE_X12Y115_DQ;
  assign CLBLM_L_X8Y116_SLICE_X10Y116_C1 = CLBLM_L_X8Y115_SLICE_X11Y115_AQ;
  assign CLBLM_L_X8Y116_SLICE_X10Y116_C2 = 1'b1;
  assign CLBLL_L_X4Y122_SLICE_X5Y122_B6 = CLBLL_L_X4Y121_SLICE_X5Y121_CO6;
  assign CLBLM_L_X8Y116_SLICE_X10Y116_C4 = CLBLM_R_X7Y116_SLICE_X9Y116_AQ;
  assign CLBLM_L_X8Y116_SLICE_X10Y116_C5 = CLBLM_L_X8Y116_SLICE_X10Y116_DO6;
  assign CLBLL_L_X4Y122_SLICE_X5Y122_C6 = RIOB33_X105Y135_IOB_X1Y136_I;
  assign CLBLM_L_X8Y116_SLICE_X10Y116_C6 = CLBLM_L_X10Y127_SLICE_X12Y127_AQ;
  assign CLBLM_L_X8Y116_SLICE_X10Y116_CE = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y116_SLICE_X10Y116_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLL_L_X4Y122_SLICE_X5Y122_C3 = CLBLL_L_X4Y123_SLICE_X5Y123_AO5;
  assign CLBLL_L_X4Y122_SLICE_X5Y122_C2 = RIOB33_X105Y135_IOB_X1Y135_I;
  assign CLBLL_L_X4Y122_SLICE_X5Y122_C4 = RIOB33_X105Y131_IOB_X1Y131_I;
  assign CLBLL_L_X4Y122_SLICE_X5Y122_C5 = CLBLM_R_X3Y122_SLICE_X3Y122_AO5;
  assign CLBLL_L_X4Y113_SLICE_X4Y113_B3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y116_SLICE_X10Y116_D1 = CLBLM_R_X11Y115_SLICE_X15Y115_CQ;
  assign CLBLM_L_X8Y116_SLICE_X10Y116_D2 = CLBLM_L_X8Y115_SLICE_X11Y115_CQ;
  assign CLBLM_L_X8Y116_SLICE_X10Y116_D3 = CLBLM_L_X10Y122_SLICE_X13Y122_A5Q;
  assign CLBLL_L_X4Y113_SLICE_X4Y113_B4 = CLBLL_L_X4Y111_SLICE_X5Y111_BQ;
  assign CLBLM_L_X8Y116_SLICE_X10Y116_D4 = 1'b1;
  assign CLBLM_L_X8Y116_SLICE_X10Y116_D5 = CLBLM_R_X7Y116_SLICE_X8Y116_CQ;
  assign CLBLM_L_X8Y116_SLICE_X10Y116_D6 = 1'b1;
  assign CLBLL_L_X4Y122_SLICE_X5Y122_D1 = RIOB33_X105Y129_IOB_X1Y130_I;
  assign CLBLL_L_X4Y113_SLICE_X4Y113_B5 = 1'b1;
  assign CLBLL_L_X4Y122_SLICE_X5Y122_D2 = RIOB33_X105Y135_IOB_X1Y135_I;
  assign CLBLL_L_X4Y122_SLICE_X5Y122_D5 = CLBLL_L_X4Y121_SLICE_X5Y121_BO6;
  assign CLBLL_L_X4Y122_SLICE_X5Y122_D6 = RIOB33_X105Y135_IOB_X1Y136_I;
  assign CLBLL_L_X4Y113_SLICE_X4Y113_B6 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X10Y126_SLICE_X12Y126_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X10Y124_SLICE_X12Y124_C6 = 1'b1;
  assign CLBLM_R_X11Y122_SLICE_X15Y122_C1 = 1'b1;
  assign CLBLM_R_X11Y120_SLICE_X15Y120_A1 = CLBLM_R_X11Y120_SLICE_X14Y120_AO5;
  assign CLBLM_R_X11Y120_SLICE_X15Y120_A2 = CLBLM_L_X12Y120_SLICE_X17Y120_CO5;
  assign CLBLM_R_X11Y120_SLICE_X15Y120_A3 = CLBLM_R_X11Y120_SLICE_X15Y120_AQ;
  assign CLBLM_R_X11Y120_SLICE_X15Y120_A4 = CLBLM_L_X10Y121_SLICE_X13Y121_CQ;
  assign CLBLM_R_X11Y120_SLICE_X15Y120_A5 = CLBLM_L_X12Y120_SLICE_X16Y120_BO6;
  assign CLBLM_R_X11Y120_SLICE_X15Y120_A6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X11Y122_SLICE_X15Y122_C2 = 1'b1;
  assign CLBLM_L_X10Y126_SLICE_X12Y126_D1 = 1'b1;
  assign CLBLM_R_X11Y122_SLICE_X15Y122_C3 = 1'b1;
  assign CLBLM_R_X11Y120_SLICE_X15Y120_B1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X11Y120_SLICE_X15Y120_B2 = CLBLM_R_X11Y120_SLICE_X15Y120_BQ;
  assign CLBLM_L_X10Y126_SLICE_X12Y126_D2 = 1'b1;
  assign CLBLM_R_X11Y120_SLICE_X15Y120_B3 = CLBLM_R_X11Y120_SLICE_X14Y120_AO6;
  assign CLBLM_R_X11Y120_SLICE_X15Y120_B4 = CLBLM_R_X5Y120_SLICE_X7Y120_BQ;
  assign CLBLM_R_X11Y120_SLICE_X15Y120_B5 = CLBLM_L_X12Y120_SLICE_X17Y120_CO5;
  assign CLBLM_R_X11Y120_SLICE_X15Y120_B6 = CLBLM_R_X11Y120_SLICE_X14Y120_BO6;
  assign CLBLM_L_X10Y126_SLICE_X12Y126_D3 = 1'b1;
  assign CLBLM_R_X11Y122_SLICE_X15Y122_C4 = 1'b1;
  assign CLBLM_R_X7Y110_SLICE_X9Y110_A1 = CLBLM_L_X10Y112_SLICE_X12Y112_DQ;
  assign CLBLM_R_X7Y110_SLICE_X9Y110_A2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y126_SLICE_X12Y126_D4 = 1'b1;
  assign CLBLM_R_X7Y110_SLICE_X9Y110_A3 = CLBLM_R_X7Y110_SLICE_X9Y110_AQ;
  assign CLBLM_R_X7Y110_SLICE_X9Y110_A4 = CLBLM_R_X3Y118_SLICE_X2Y118_AQ;
  assign CLBLM_R_X7Y110_SLICE_X9Y110_A5 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_R_X7Y110_SLICE_X9Y110_A6 = CLBLM_R_X5Y113_SLICE_X7Y113_A5Q;
  assign CLBLM_L_X10Y126_SLICE_X12Y126_D5 = 1'b1;
  assign CLBLM_R_X11Y120_SLICE_X15Y120_C1 = CLBLM_L_X12Y121_SLICE_X16Y121_AQ;
  assign CLBLM_R_X7Y110_SLICE_X9Y110_B1 = CLBLM_R_X5Y111_SLICE_X7Y111_DO6;
  assign CLBLM_R_X7Y110_SLICE_X9Y110_B2 = CLBLM_R_X7Y110_SLICE_X9Y110_BQ;
  assign CLBLM_L_X10Y126_SLICE_X12Y126_D6 = 1'b1;
  assign CLBLM_R_X7Y110_SLICE_X9Y110_B3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y110_SLICE_X9Y110_B4 = 1'b1;
  assign CLBLM_R_X7Y110_SLICE_X9Y110_B5 = CLBLM_L_X8Y117_SLICE_X10Y117_AQ;
  assign CLBLM_R_X7Y110_SLICE_X9Y110_B6 = CLBLM_R_X5Y116_SLICE_X7Y116_CQ;
  assign CLBLM_R_X11Y120_SLICE_X15Y120_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X7Y110_SLICE_X9Y110_C1 = 1'b1;
  assign CLBLM_R_X7Y110_SLICE_X9Y110_C2 = CLBLM_R_X7Y110_SLICE_X9Y110_CQ;
  assign CLBLM_R_X7Y110_SLICE_X9Y110_C3 = 1'b1;
  assign CLBLM_R_X7Y110_SLICE_X9Y110_C4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y110_SLICE_X9Y110_C5 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X7Y110_SLICE_X9Y110_C6 = CLBLM_R_X7Y115_SLICE_X9Y115_BQ;
  assign CLBLM_R_X11Y120_SLICE_X15Y120_D3 = CLBLM_R_X11Y121_SLICE_X15Y121_AO6;
  assign CLBLM_R_X11Y120_SLICE_X15Y120_D4 = CLBLM_L_X12Y120_SLICE_X17Y120_DO5;
  assign CLBLM_R_X7Y110_SLICE_X9Y110_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X11Y120_SLICE_X14Y120_A1 = CLBLM_R_X11Y118_SLICE_X14Y118_BQ;
  assign CLBLM_R_X11Y120_SLICE_X14Y120_A2 = CLBLM_R_X13Y119_SLICE_X18Y119_CQ;
  assign CLBLM_R_X11Y120_SLICE_X14Y120_A3 = CLBLM_R_X7Y120_SLICE_X9Y120_AQ;
  assign CLBLM_R_X11Y120_SLICE_X14Y120_A4 = CLBLM_L_X10Y119_SLICE_X13Y119_AQ;
  assign CLBLM_R_X7Y110_SLICE_X9Y110_D1 = 1'b1;
  assign CLBLM_R_X7Y110_SLICE_X9Y110_D2 = 1'b1;
  assign CLBLM_R_X7Y110_SLICE_X9Y110_D3 = 1'b1;
  assign CLBLM_R_X7Y110_SLICE_X9Y110_D4 = 1'b1;
  assign CLBLM_R_X7Y110_SLICE_X9Y110_D5 = 1'b1;
  assign CLBLM_R_X7Y110_SLICE_X9Y110_D6 = 1'b1;
  assign CLBLM_R_X11Y120_SLICE_X14Y120_A5 = CLBLM_R_X11Y119_SLICE_X15Y119_CQ;
  assign CLBLM_R_X11Y120_SLICE_X14Y120_A6 = 1'b1;
  assign CLBLM_R_X11Y120_SLICE_X14Y120_AX = CLBLM_R_X11Y118_SLICE_X14Y118_BQ;
  assign CLBLM_R_X11Y120_SLICE_X14Y120_B1 = CLBLM_L_X12Y120_SLICE_X16Y120_AO6;
  assign CLBLM_R_X11Y120_SLICE_X14Y120_B2 = CLBLM_R_X13Y119_SLICE_X18Y119_CQ;
  assign CLBLM_R_X11Y120_SLICE_X14Y120_B3 = CLBLM_R_X7Y120_SLICE_X9Y120_AQ;
  assign CLBLM_R_X7Y110_SLICE_X8Y110_A1 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_R_X7Y110_SLICE_X8Y110_A2 = CLBLM_R_X7Y110_SLICE_X8Y110_BQ;
  assign CLBLM_R_X7Y110_SLICE_X8Y110_A3 = CLBLM_R_X7Y110_SLICE_X8Y110_AQ;
  assign CLBLM_R_X7Y110_SLICE_X8Y110_A4 = CLBLM_R_X3Y118_SLICE_X2Y118_AQ;
  assign CLBLM_R_X7Y110_SLICE_X8Y110_A5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y110_SLICE_X8Y110_A6 = CLBLM_R_X7Y118_SLICE_X8Y118_CQ;
  assign CLBLM_R_X11Y120_SLICE_X14Y120_C1 = CLBLM_R_X7Y120_SLICE_X9Y120_AQ;
  assign CLBLM_R_X11Y120_SLICE_X14Y120_C2 = CLBLM_R_X11Y119_SLICE_X14Y119_AO5;
  assign CLBLM_R_X11Y120_SLICE_X14Y120_C3 = RIOB33_X105Y121_IOB_X1Y121_I;
  assign CLBLM_R_X7Y110_SLICE_X8Y110_B1 = CLBLM_R_X7Y111_SLICE_X8Y111_CQ;
  assign CLBLM_R_X7Y110_SLICE_X8Y110_B2 = CLBLM_R_X7Y110_SLICE_X8Y110_BQ;
  assign CLBLM_R_X7Y110_SLICE_X8Y110_B3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y110_SLICE_X8Y110_B4 = CLBLM_R_X7Y115_SLICE_X8Y115_BQ;
  assign CLBLM_R_X7Y110_SLICE_X8Y110_B5 = CLBLM_R_X3Y118_SLICE_X2Y118_AQ;
  assign CLBLM_R_X7Y110_SLICE_X8Y110_B6 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_R_X11Y120_SLICE_X14Y120_CE = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X11Y120_SLICE_X14Y120_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X11Y120_SLICE_X14Y120_D1 = CLBLM_R_X11Y119_SLICE_X15Y119_CQ;
  assign CLBLM_R_X7Y110_SLICE_X8Y110_C1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y110_SLICE_X8Y110_C2 = CLBLM_R_X7Y110_SLICE_X8Y110_CQ;
  assign CLBLM_R_X7Y110_SLICE_X8Y110_C3 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X7Y110_SLICE_X8Y110_C4 = CLBLM_L_X8Y113_SLICE_X11Y113_CQ;
  assign CLBLM_R_X7Y110_SLICE_X8Y110_C5 = CLBLM_R_X7Y110_SLICE_X8Y110_DO6;
  assign CLBLM_R_X7Y110_SLICE_X8Y110_C6 = CLBLM_L_X8Y118_SLICE_X10Y118_DQ;
  assign CLBLM_R_X11Y120_SLICE_X14Y120_D2 = CLBLM_L_X12Y120_SLICE_X16Y120_AO6;
  assign CLBLM_R_X11Y120_SLICE_X14Y120_D3 = CLBLM_R_X11Y118_SLICE_X14Y118_BQ;
  assign CLBLL_L_X2Y111_SLICE_X0Y111_A5 = RIOB33_X105Y137_IOB_X1Y137_I;
  assign CLBLM_R_X7Y110_SLICE_X8Y110_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X11Y120_SLICE_X14Y120_D6 = CLBLM_R_X11Y120_SLICE_X15Y120_BQ;
  assign CLBLM_R_X11Y120_SLICE_X14Y120_SR = CLBLM_R_X11Y123_SLICE_X14Y123_CO6;
  assign CLBLL_L_X2Y111_SLICE_X0Y111_A6 = 1'b1;
  assign CLBLM_R_X11Y122_SLICE_X15Y122_D6 = 1'b1;
  assign CLBLM_R_X7Y110_SLICE_X8Y110_D1 = CLBLM_L_X10Y112_SLICE_X13Y112_CQ;
  assign CLBLM_R_X7Y110_SLICE_X8Y110_D2 = CLBLM_R_X7Y110_SLICE_X8Y110_CQ;
  assign CLBLM_R_X7Y110_SLICE_X8Y110_D3 = CLBLL_L_X4Y110_SLICE_X5Y110_AQ;
  assign CLBLM_R_X7Y110_SLICE_X8Y110_D4 = CLBLM_L_X8Y110_SLICE_X10Y110_BQ;
  assign CLBLM_R_X7Y110_SLICE_X8Y110_D5 = CLBLM_R_X5Y111_SLICE_X7Y111_DO6;
  assign CLBLM_R_X7Y110_SLICE_X8Y110_D6 = 1'b1;
  assign CLBLM_R_X11Y122_SLICE_X14Y122_A1 = 1'b1;
  assign LIOB33_X0Y189_IOB_X0Y190_O = RIOB33_X105Y147_IOB_X1Y147_I;
  assign CLBLM_R_X11Y122_SLICE_X14Y122_A2 = CLBLM_L_X10Y122_SLICE_X13Y122_CQ;
  assign CLBLM_R_X11Y122_SLICE_X14Y122_A3 = CLBLM_R_X11Y122_SLICE_X14Y122_AQ;
  assign CLBLM_R_X11Y122_SLICE_X14Y122_A4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign LIOB33_X0Y189_IOB_X0Y189_O = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_L_X10Y127_SLICE_X13Y127_A1 = 1'b1;
  assign CLBLL_L_X4Y123_SLICE_X4Y123_A1 = CLBLL_L_X4Y123_SLICE_X4Y123_CQ;
  assign CLBLL_L_X4Y123_SLICE_X4Y123_A2 = CLBLM_R_X7Y124_SLICE_X8Y124_BQ;
  assign CLBLM_L_X10Y127_SLICE_X13Y127_A4 = 1'b1;
  assign CLBLM_L_X10Y127_SLICE_X13Y127_A5 = 1'b1;
  assign CLBLM_L_X10Y127_SLICE_X13Y127_A6 = 1'b1;
  assign CLBLL_L_X4Y123_SLICE_X4Y123_A3 = CLBLL_L_X4Y123_SLICE_X4Y123_AQ;
  assign CLBLL_L_X4Y123_SLICE_X4Y123_A4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLL_L_X4Y123_SLICE_X4Y123_A5 = CLBLM_R_X7Y124_SLICE_X8Y124_DO5;
  assign CLBLL_L_X4Y123_SLICE_X4Y123_A6 = CLBLM_R_X7Y124_SLICE_X8Y124_A5Q;
  assign CLBLM_L_X10Y127_SLICE_X13Y127_B2 = 1'b1;
  assign CLBLM_L_X10Y127_SLICE_X13Y127_B3 = 1'b1;
  assign CLBLM_L_X10Y127_SLICE_X13Y127_B4 = 1'b1;
  assign CLBLM_L_X10Y127_SLICE_X13Y127_B5 = 1'b1;
  assign CLBLM_L_X10Y127_SLICE_X13Y127_B6 = 1'b1;
  assign CLBLL_L_X4Y123_SLICE_X4Y123_B1 = CLBLM_R_X5Y125_SLICE_X6Y125_BO5;
  assign CLBLL_L_X4Y123_SLICE_X4Y123_B2 = CLBLL_L_X4Y123_SLICE_X4Y123_BQ;
  assign CLBLM_L_X10Y127_SLICE_X13Y127_C1 = 1'b1;
  assign CLBLM_L_X10Y127_SLICE_X13Y127_C2 = 1'b1;
  assign CLBLM_L_X10Y127_SLICE_X13Y127_C3 = 1'b1;
  assign CLBLM_L_X10Y127_SLICE_X13Y127_C4 = 1'b1;
  assign CLBLM_L_X10Y127_SLICE_X13Y127_C5 = 1'b1;
  assign CLBLM_L_X10Y127_SLICE_X13Y127_C6 = 1'b1;
  assign CLBLL_L_X4Y123_SLICE_X4Y123_C3 = CLBLM_R_X3Y116_SLICE_X2Y116_DO6;
  assign CLBLL_L_X4Y123_SLICE_X4Y123_C4 = CLBLM_R_X5Y116_SLICE_X6Y116_A5Q;
  assign CLBLL_L_X4Y123_SLICE_X4Y123_C5 = CLBLL_L_X4Y123_SLICE_X4Y123_CQ;
  assign CLBLL_L_X4Y123_SLICE_X4Y123_C6 = 1'b1;
  assign CLBLM_L_X8Y117_SLICE_X11Y117_A2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y117_SLICE_X11Y117_A3 = RIOB33_X105Y135_IOB_X1Y135_I;
  assign CLBLM_L_X8Y117_SLICE_X11Y117_A4 = RIOB33_X105Y131_IOB_X1Y131_I;
  assign CLBLM_L_X8Y117_SLICE_X11Y117_A6 = CLBLM_L_X10Y114_SLICE_X13Y114_A5Q;
  assign CLBLM_L_X10Y127_SLICE_X13Y127_D1 = 1'b1;
  assign CLBLM_L_X10Y127_SLICE_X13Y127_D2 = 1'b1;
  assign CLBLM_L_X10Y127_SLICE_X13Y127_D3 = 1'b1;
  assign CLBLM_L_X10Y127_SLICE_X13Y127_D4 = 1'b1;
  assign CLBLM_L_X10Y127_SLICE_X13Y127_D5 = 1'b1;
  assign CLBLM_L_X10Y127_SLICE_X13Y127_D6 = 1'b1;
  assign CLBLM_L_X8Y128_SLICE_X10Y128_D6 = 1'b1;
  assign CLBLM_L_X8Y117_SLICE_X11Y117_B4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y117_SLICE_X11Y117_B6 = CLBLM_R_X7Y121_SLICE_X9Y121_A5Q;
  assign CLBLL_L_X4Y123_SLICE_X4Y123_D1 = RIOB33_X105Y131_IOB_X1Y132_I;
  assign CLBLM_L_X8Y117_SLICE_X11Y117_C1 = CLBLM_R_X7Y116_SLICE_X8Y116_DO6;
  assign CLBLM_L_X10Y127_SLICE_X12Y127_A1 = 1'b1;
  assign CLBLM_L_X10Y127_SLICE_X12Y127_A2 = 1'b1;
  assign CLBLM_L_X10Y127_SLICE_X12Y127_A3 = 1'b1;
  assign CLBLM_L_X10Y127_SLICE_X12Y127_A4 = 1'b1;
  assign CLBLM_L_X10Y127_SLICE_X12Y127_A5 = 1'b1;
  assign CLBLM_L_X8Y117_SLICE_X11Y117_C5 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_L_X8Y117_SLICE_X11Y117_C6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y117_SLICE_X11Y117_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X8Y117_SLICE_X11Y117_D1 = CLBLM_R_X7Y116_SLICE_X8Y116_DO6;
  assign CLBLM_L_X8Y117_SLICE_X11Y117_D2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y117_SLICE_X11Y117_D3 = CLBLM_L_X8Y117_SLICE_X11Y117_DQ;
  assign CLBLM_L_X8Y117_SLICE_X11Y117_D4 = CLBLM_R_X3Y118_SLICE_X2Y118_AQ;
  assign CLBLM_L_X10Y127_SLICE_X12Y127_B3 = 1'b1;
  assign CLBLM_L_X10Y127_SLICE_X12Y127_B4 = 1'b1;
  assign CLBLM_L_X10Y127_SLICE_X12Y127_B5 = 1'b1;
  assign CLBLM_L_X10Y127_SLICE_X12Y127_B6 = 1'b1;
  assign CLBLM_L_X8Y117_SLICE_X11Y117_D5 = CLBLM_R_X7Y118_SLICE_X8Y118_AQ;
  assign CLBLM_L_X8Y117_SLICE_X11Y117_D6 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_L_X10Y127_SLICE_X12Y127_B2 = 1'b1;
  assign CLBLM_L_X10Y127_SLICE_X12Y127_C1 = 1'b1;
  assign CLBLM_L_X10Y127_SLICE_X12Y127_C2 = 1'b1;
  assign CLBLM_L_X10Y127_SLICE_X12Y127_C3 = 1'b1;
  assign CLBLM_L_X10Y127_SLICE_X12Y127_C4 = 1'b1;
  assign CLBLM_L_X10Y127_SLICE_X12Y127_C5 = 1'b1;
  assign CLBLM_L_X10Y127_SLICE_X12Y127_C6 = 1'b1;
  assign CLBLL_L_X4Y123_SLICE_X5Y123_A2 = 1'b1;
  assign CLBLL_L_X4Y123_SLICE_X5Y123_A3 = RIOB33_X105Y131_IOB_X1Y132_I;
  assign CLBLM_L_X8Y117_SLICE_X10Y117_A2 = CLBLM_R_X7Y121_SLICE_X8Y121_AQ;
  assign CLBLM_L_X10Y127_SLICE_X12Y127_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X8Y117_SLICE_X10Y117_A4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLL_L_X2Y109_SLICE_X0Y109_A1 = 1'b1;
  assign CLBLL_L_X2Y109_SLICE_X0Y109_A2 = 1'b1;
  assign CLBLL_L_X2Y109_SLICE_X0Y109_A3 = 1'b1;
  assign CLBLL_L_X2Y109_SLICE_X0Y109_A5 = 1'b1;
  assign CLBLM_L_X10Y127_SLICE_X12Y127_D1 = 1'b1;
  assign CLBLM_L_X10Y127_SLICE_X12Y127_D2 = 1'b1;
  assign CLBLM_L_X10Y127_SLICE_X12Y127_D3 = 1'b1;
  assign CLBLM_L_X10Y127_SLICE_X12Y127_D4 = 1'b1;
  assign CLBLM_L_X10Y127_SLICE_X12Y127_D5 = 1'b1;
  assign CLBLM_L_X10Y127_SLICE_X12Y127_D6 = 1'b1;
  assign CLBLL_L_X4Y123_SLICE_X5Y123_C1 = 1'b1;
  assign CLBLL_L_X4Y123_SLICE_X5Y123_C2 = 1'b1;
  assign CLBLL_L_X4Y123_SLICE_X5Y123_C3 = 1'b1;
  assign CLBLL_L_X4Y123_SLICE_X5Y123_C5 = 1'b1;
  assign CLBLL_L_X2Y109_SLICE_X0Y109_B1 = 1'b1;
  assign CLBLL_L_X2Y109_SLICE_X0Y109_B2 = 1'b1;
  assign CLBLM_L_X8Y117_SLICE_X10Y117_C2 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_L_X8Y117_SLICE_X10Y117_C3 = CLBLM_R_X3Y118_SLICE_X2Y118_AQ;
  assign CLBLL_L_X2Y109_SLICE_X0Y109_B3 = 1'b1;
  assign CLBLL_L_X2Y109_SLICE_X0Y109_C3 = 1'b1;
  assign CLBLL_L_X2Y109_SLICE_X0Y109_C5 = 1'b1;
  assign CLBLL_L_X4Y123_SLICE_X5Y123_D1 = 1'b1;
  assign CLBLL_L_X4Y123_SLICE_X5Y123_D2 = 1'b1;
  assign CLBLL_L_X2Y109_SLICE_X0Y109_C6 = 1'b1;
  assign CLBLL_L_X4Y123_SLICE_X5Y123_D3 = 1'b1;
  assign CLBLL_L_X4Y123_SLICE_X5Y123_D4 = 1'b1;
  assign CLBLL_L_X4Y123_SLICE_X5Y123_D5 = 1'b1;
  assign CLBLM_L_X8Y117_SLICE_X10Y117_D1 = CLBLM_L_X8Y117_SLICE_X10Y117_BQ;
  assign CLBLM_L_X8Y117_SLICE_X10Y117_D2 = CLBLM_R_X3Y116_SLICE_X3Y116_BQ;
  assign CLBLM_L_X8Y117_SLICE_X10Y117_D3 = CLBLM_L_X8Y115_SLICE_X10Y115_DQ;
  assign CLBLM_L_X8Y117_SLICE_X10Y117_D4 = RIOB33_X105Y121_IOB_X1Y121_I;
  assign CLBLM_L_X8Y117_SLICE_X10Y117_D5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y117_SLICE_X10Y117_D6 = 1'b1;
  assign CLBLL_L_X4Y123_SLICE_X5Y123_D6 = 1'b1;
  assign CLBLL_L_X2Y109_SLICE_X0Y109_D1 = 1'b1;
  assign CLBLL_L_X2Y109_SLICE_X0Y109_D2 = 1'b1;
  assign CLBLL_L_X2Y109_SLICE_X0Y109_D3 = 1'b1;
  assign CLBLL_L_X2Y109_SLICE_X0Y109_D4 = 1'b1;
  assign CLBLL_L_X2Y109_SLICE_X0Y109_D5 = 1'b1;
  assign CLBLL_L_X2Y109_SLICE_X0Y109_D6 = 1'b1;
  assign CLBLM_L_X8Y118_SLICE_X11Y118_A3 = CLBLM_L_X8Y118_SLICE_X11Y118_AQ;
  assign CLBLM_L_X8Y118_SLICE_X11Y118_A4 = CLBLM_R_X11Y121_SLICE_X14Y121_CO6;
  assign LIOI3_TBYTESRC_X0Y107_OLOGIC_X0Y107_D1 = CLBLL_L_X2Y109_SLICE_X0Y109_AO6;
  assign CLBLM_L_X8Y118_SLICE_X11Y118_A5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign LIOI3_TBYTESRC_X0Y107_OLOGIC_X0Y107_T1 = 1'b1;
  assign CLBLM_L_X8Y118_SLICE_X11Y118_A6 = 1'b1;
  assign CLBLM_R_X11Y121_SLICE_X15Y121_A1 = CLBLM_L_X10Y119_SLICE_X13Y119_AQ;
  assign CLBLM_R_X11Y121_SLICE_X15Y121_A2 = CLBLM_R_X7Y120_SLICE_X9Y120_AQ;
  assign CLBLM_R_X11Y121_SLICE_X15Y121_A3 = CLBLM_R_X11Y118_SLICE_X14Y118_AQ;
  assign CLBLM_R_X11Y121_SLICE_X15Y121_A4 = CLBLM_R_X11Y121_SLICE_X15Y121_BO6;
  assign CLBLM_R_X11Y121_SLICE_X15Y121_A5 = CLBLM_R_X11Y119_SLICE_X15Y119_CQ;
  assign CLBLL_L_X2Y109_SLICE_X1Y109_A1 = 1'b1;
  assign CLBLL_L_X2Y109_SLICE_X1Y109_A2 = 1'b1;
  assign CLBLL_L_X2Y109_SLICE_X1Y109_A3 = 1'b1;
  assign CLBLL_L_X2Y109_SLICE_X1Y109_A4 = 1'b1;
  assign CLBLL_L_X2Y109_SLICE_X1Y109_A5 = 1'b1;
  assign CLBLL_L_X2Y109_SLICE_X1Y109_A6 = 1'b1;
  assign CLBLM_R_X11Y121_SLICE_X15Y121_A6 = CLBLM_R_X11Y121_SLICE_X15Y121_CO6;
  assign CLBLM_R_X11Y121_SLICE_X15Y121_B1 = CLBLM_R_X11Y119_SLICE_X15Y119_CQ;
  assign CLBLL_L_X2Y109_SLICE_X1Y109_B1 = 1'b1;
  assign CLBLL_L_X2Y109_SLICE_X1Y109_B2 = 1'b1;
  assign CLBLL_L_X2Y109_SLICE_X1Y109_B3 = 1'b1;
  assign CLBLL_L_X2Y109_SLICE_X1Y109_B4 = 1'b1;
  assign CLBLL_L_X2Y109_SLICE_X1Y109_B5 = 1'b1;
  assign CLBLL_L_X2Y109_SLICE_X1Y109_B6 = 1'b1;
  assign CLBLM_L_X8Y118_SLICE_X11Y118_B1 = CLBLM_R_X5Y124_SLICE_X6Y124_CQ;
  assign CLBLM_R_X7Y111_SLICE_X9Y111_A1 = CLBLM_R_X3Y119_SLICE_X2Y119_AO6;
  assign CLBLM_R_X7Y111_SLICE_X9Y111_A2 = CLBLL_L_X4Y120_SLICE_X4Y120_BO6;
  assign CLBLL_L_X2Y109_SLICE_X1Y109_C1 = 1'b1;
  assign CLBLL_L_X2Y109_SLICE_X1Y109_C2 = 1'b1;
  assign CLBLL_L_X2Y109_SLICE_X1Y109_C3 = 1'b1;
  assign CLBLL_L_X2Y109_SLICE_X1Y109_C4 = 1'b1;
  assign CLBLL_L_X2Y109_SLICE_X1Y109_C5 = 1'b1;
  assign CLBLL_L_X2Y109_SLICE_X1Y109_C6 = 1'b1;
  assign CLBLM_L_X8Y118_SLICE_X11Y118_B2 = CLBLM_L_X8Y114_SLICE_X10Y114_BQ;
  assign CLBLM_L_X8Y118_SLICE_X11Y118_B3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y111_SLICE_X9Y111_A5 = CLBLL_L_X4Y120_SLICE_X4Y120_AO6;
  assign CLBLM_R_X7Y111_SLICE_X9Y111_A6 = 1'b1;
  assign CLBLM_L_X8Y118_SLICE_X11Y118_B4 = RIOB33_X105Y121_IOB_X1Y121_I;
  assign CLBLM_R_X7Y111_SLICE_X9Y111_B1 = CLBLL_L_X4Y110_SLICE_X5Y110_AQ;
  assign CLBLM_R_X7Y111_SLICE_X9Y111_B2 = CLBLM_L_X8Y117_SLICE_X11Y117_BQ;
  assign CLBLL_L_X2Y109_SLICE_X1Y109_D1 = 1'b1;
  assign CLBLL_L_X2Y109_SLICE_X1Y109_D2 = 1'b1;
  assign CLBLL_L_X2Y109_SLICE_X1Y109_D3 = 1'b1;
  assign CLBLL_L_X2Y109_SLICE_X1Y109_D4 = 1'b1;
  assign CLBLL_L_X2Y109_SLICE_X1Y109_D5 = 1'b1;
  assign CLBLL_L_X2Y109_SLICE_X1Y109_D6 = 1'b1;
  assign CLBLM_L_X8Y118_SLICE_X11Y118_B5 = CLBLM_L_X8Y117_SLICE_X11Y117_CQ;
  assign CLBLM_L_X8Y118_SLICE_X11Y118_B6 = 1'b1;
  assign CLBLM_R_X7Y111_SLICE_X9Y111_C1 = 1'b1;
  assign CLBLM_R_X7Y111_SLICE_X9Y111_C2 = CLBLL_L_X4Y119_SLICE_X4Y119_CQ;
  assign CLBLM_R_X7Y111_SLICE_X9Y111_C3 = 1'b1;
  assign CLBLM_R_X7Y111_SLICE_X9Y111_C4 = CLBLM_R_X7Y111_SLICE_X8Y111_CQ;
  assign CLBLM_R_X7Y111_SLICE_X9Y111_C6 = CLBLM_R_X7Y111_SLICE_X9Y111_BO6;
  assign CLBLM_R_X7Y111_SLICE_X9Y111_D1 = CLBLM_R_X7Y110_SLICE_X9Y110_AQ;
  assign CLBLM_R_X7Y111_SLICE_X9Y111_D2 = CLBLM_R_X5Y117_SLICE_X7Y117_DO6;
  assign CLBLM_R_X7Y111_SLICE_X9Y111_D3 = CLBLM_R_X5Y114_SLICE_X6Y114_AQ;
  assign CLBLM_R_X7Y111_SLICE_X9Y111_D4 = CLBLM_R_X3Y119_SLICE_X2Y119_AO6;
  assign CLBLM_R_X7Y111_SLICE_X9Y111_D5 = 1'b1;
  assign CLBLM_R_X7Y111_SLICE_X9Y111_D6 = 1'b1;
  assign CLBLM_R_X11Y121_SLICE_X14Y121_A5 = CLBLM_R_X11Y118_SLICE_X14Y118_BQ;
  assign CLBLM_R_X11Y121_SLICE_X14Y121_A6 = CLBLM_R_X13Y119_SLICE_X18Y119_CQ;
  assign CLBLM_R_X11Y121_SLICE_X14Y121_B1 = CLBLM_L_X10Y122_SLICE_X12Y122_CO6;
  assign CLBLM_R_X11Y121_SLICE_X14Y121_B2 = CLBLM_L_X10Y121_SLICE_X13Y121_CQ;
  assign CLBLM_R_X11Y121_SLICE_X14Y121_B3 = CLBLM_L_X10Y120_SLICE_X13Y120_BQ;
  assign CLBLM_R_X7Y111_SLICE_X8Y111_A1 = 1'b1;
  assign CLBLM_R_X7Y111_SLICE_X8Y111_A2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y111_SLICE_X8Y111_A3 = CLBLM_R_X7Y111_SLICE_X8Y111_AQ;
  assign CLBLM_R_X7Y111_SLICE_X8Y111_A4 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X7Y111_SLICE_X8Y111_A5 = CLBLM_R_X5Y111_SLICE_X7Y111_AQ;
  assign CLBLM_R_X7Y111_SLICE_X8Y111_A6 = 1'b1;
  assign CLBLM_R_X7Y124_SLICE_X8Y124_B5 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X11Y121_SLICE_X14Y121_C1 = 1'b1;
  assign CLBLM_R_X7Y124_SLICE_X8Y124_B6 = CLBLM_R_X7Y124_SLICE_X8Y124_A5Q;
  assign CLBLM_R_X7Y111_SLICE_X8Y111_B1 = CLBLM_R_X3Y115_SLICE_X3Y115_DQ;
  assign CLBLM_R_X7Y111_SLICE_X8Y111_B2 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X7Y111_SLICE_X8Y111_B3 = 1'b1;
  assign CLBLM_R_X7Y111_SLICE_X8Y111_B4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y111_SLICE_X8Y111_B5 = 1'b1;
  assign CLBLM_R_X7Y111_SLICE_X8Y111_B6 = CLBLM_R_X7Y111_SLICE_X8Y111_BQ;
  assign CLBLM_R_X11Y121_SLICE_X14Y121_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X11Y121_SLICE_X14Y121_D1 = 1'b1;
  assign CLBLM_R_X11Y121_SLICE_X14Y121_D2 = CLBLM_L_X8Y122_SLICE_X11Y122_DO6;
  assign CLBLM_R_X7Y111_SLICE_X8Y111_C1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y111_SLICE_X8Y111_C2 = CLBLM_R_X7Y111_SLICE_X9Y111_CO6;
  assign CLBLM_R_X7Y111_SLICE_X8Y111_C3 = CLBLM_R_X7Y111_SLICE_X8Y111_BQ;
  assign CLBLM_R_X7Y111_SLICE_X8Y111_C4 = CLBLM_R_X7Y128_SLICE_X8Y128_AQ;
  assign CLBLM_R_X7Y111_SLICE_X8Y111_C5 = 1'b1;
  assign CLBLM_R_X7Y111_SLICE_X8Y111_C6 = RIOB33_X105Y141_IOB_X1Y142_I;
  assign CLBLM_R_X11Y121_SLICE_X14Y121_D3 = CLBLM_L_X10Y123_SLICE_X12Y123_CO6;
  assign CLBLM_R_X11Y121_SLICE_X14Y121_D4 = CLBLM_L_X10Y121_SLICE_X13Y121_CQ;
  assign CLBLM_R_X11Y121_SLICE_X14Y121_D5 = CLBLM_L_X8Y121_SLICE_X11Y121_CQ;
  assign CLBLM_R_X7Y111_SLICE_X8Y111_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X11Y121_SLICE_X14Y121_D6 = 1'b1;
  assign CLBLM_L_X10Y116_SLICE_X12Y116_B3 = CLBLL_L_X4Y116_SLICE_X4Y116_DQ;
  assign CLBLM_R_X7Y111_SLICE_X8Y111_D1 = 1'b1;
  assign CLBLM_L_X10Y116_SLICE_X12Y116_B4 = 1'b1;
  assign CLBLM_R_X7Y111_SLICE_X8Y111_D2 = CLBLM_R_X7Y110_SLICE_X9Y110_CQ;
  assign CLBLM_R_X7Y111_SLICE_X8Y111_D3 = CLBLM_R_X7Y111_SLICE_X8Y111_BQ;
  assign CLBLM_R_X7Y111_SLICE_X8Y111_D4 = CLBLM_R_X5Y115_SLICE_X7Y115_A5Q;
  assign CLBLM_R_X7Y111_SLICE_X8Y111_D5 = 1'b1;
  assign CLBLM_R_X7Y111_SLICE_X8Y111_D6 = CLBLM_R_X7Y111_SLICE_X8Y111_AQ;
  assign CLBLM_R_X13Y120_SLICE_X19Y120_A6 = 1'b1;
  assign LIOI3_SING_X0Y50_ILOGIC_X0Y50_D = LIOB33_SING_X0Y50_IOB_X0Y50_I;
  assign CLBLM_R_X7Y124_SLICE_X8Y124_C4 = CLBLM_R_X7Y122_SLICE_X8Y122_CQ;
  assign CLBLM_R_X7Y124_SLICE_X8Y124_C5 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign LIOI3_X0Y61_ILOGIC_X0Y62_D = LIOB33_X0Y61_IOB_X0Y62_I;
  assign LIOI3_X0Y61_ILOGIC_X0Y61_D = LIOB33_X0Y61_IOB_X0Y61_I;
  assign CLBLM_R_X7Y124_SLICE_X8Y124_C6 = CLBLM_R_X7Y125_SLICE_X8Y125_AO6;
  assign RIOI3_X105Y105_ILOGIC_X1Y106_D = RIOB33_X105Y105_IOB_X1Y106_I;
  assign CLBLM_L_X8Y118_SLICE_X11Y118_D1 = 1'b1;
  assign CLBLM_L_X10Y116_SLICE_X12Y116_C1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign RIOI3_X105Y105_ILOGIC_X1Y105_D = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X10Y116_SLICE_X12Y116_C2 = CLBLM_L_X10Y116_SLICE_X13Y116_BQ;
  assign CLBLM_L_X8Y118_SLICE_X11Y118_D3 = 1'b1;
  assign CLBLM_L_X10Y116_SLICE_X12Y116_C3 = CLBLM_L_X10Y114_SLICE_X12Y114_BO5;
  assign CLBLM_R_X11Y128_SLICE_X15Y128_D5 = 1'b1;
  assign CLBLM_L_X10Y116_SLICE_X12Y116_C4 = 1'b1;
  assign CLBLM_L_X8Y118_SLICE_X11Y118_D5 = 1'b1;
  assign CLBLL_L_X52Y126_SLICE_X78Y126_A1 = 1'b1;
  assign CLBLL_L_X52Y126_SLICE_X78Y126_A2 = 1'b1;
  assign CLBLL_L_X52Y126_SLICE_X78Y126_A3 = 1'b1;
  assign CLBLL_L_X52Y126_SLICE_X78Y126_A4 = RIOB33_X105Y123_IOB_X1Y124_I;
  assign CLBLM_L_X10Y128_SLICE_X13Y128_A3 = CLBLM_L_X10Y124_SLICE_X13Y124_AQ;
  assign CLBLM_L_X10Y128_SLICE_X13Y128_A4 = RIOB33_X105Y143_IOB_X1Y143_I;
  assign CLBLM_L_X10Y128_SLICE_X13Y128_A5 = CLBLM_L_X8Y122_SLICE_X11Y122_A5Q;
  assign CLBLM_L_X10Y128_SLICE_X13Y128_A6 = 1'b1;
  assign CLBLL_L_X52Y126_SLICE_X78Y126_A5 = 1'b1;
  assign CLBLL_L_X52Y126_SLICE_X78Y126_A6 = 1'b1;
  assign CLBLM_L_X10Y116_SLICE_X12Y116_C6 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X10Y128_SLICE_X13Y128_A1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y128_SLICE_X13Y128_B1 = 1'b1;
  assign CLBLM_L_X10Y128_SLICE_X13Y128_B2 = 1'b1;
  assign CLBLM_L_X10Y128_SLICE_X13Y128_B3 = 1'b1;
  assign CLBLM_L_X10Y128_SLICE_X13Y128_B4 = 1'b1;
  assign CLBLM_L_X10Y128_SLICE_X13Y128_B5 = 1'b1;
  assign CLBLM_L_X10Y128_SLICE_X13Y128_B6 = 1'b1;
  assign CLBLL_L_X52Y126_SLICE_X78Y126_B1 = 1'b1;
  assign CLBLL_L_X52Y126_SLICE_X78Y126_B2 = 1'b1;
  assign CLBLL_L_X52Y126_SLICE_X78Y126_B3 = 1'b1;
  assign CLBLM_L_X10Y128_SLICE_X13Y128_C1 = 1'b1;
  assign CLBLM_L_X10Y128_SLICE_X13Y128_C2 = 1'b1;
  assign CLBLM_L_X10Y128_SLICE_X13Y128_C3 = 1'b1;
  assign CLBLM_L_X10Y128_SLICE_X13Y128_C4 = 1'b1;
  assign CLBLM_L_X10Y128_SLICE_X13Y128_C5 = 1'b1;
  assign CLBLM_L_X10Y128_SLICE_X13Y128_C6 = 1'b1;
  assign CLBLL_L_X52Y126_SLICE_X78Y126_C3 = 1'b1;
  assign CLBLL_L_X52Y126_SLICE_X78Y126_C1 = 1'b1;
  assign CLBLL_L_X52Y126_SLICE_X78Y126_C2 = 1'b1;
  assign CLBLM_L_X8Y118_SLICE_X11Y118_A1 = CLBLM_L_X10Y119_SLICE_X13Y119_DQ;
  assign CLBLM_L_X8Y118_SLICE_X11Y118_A2 = CLBLM_L_X10Y118_SLICE_X12Y118_BQ;
  assign CLBLL_L_X52Y126_SLICE_X78Y126_C5 = 1'b1;
  assign CLBLL_L_X52Y126_SLICE_X78Y126_C6 = 1'b1;
  assign CLBLM_L_X10Y128_SLICE_X13Y128_D1 = 1'b1;
  assign CLBLM_L_X10Y128_SLICE_X13Y128_D2 = 1'b1;
  assign CLBLM_L_X10Y128_SLICE_X13Y128_D3 = 1'b1;
  assign CLBLM_L_X10Y128_SLICE_X13Y128_D4 = 1'b1;
  assign CLBLM_L_X10Y128_SLICE_X13Y128_D5 = 1'b1;
  assign CLBLM_L_X10Y128_SLICE_X13Y128_D6 = 1'b1;
  assign CLBLL_L_X52Y126_SLICE_X78Y126_D5 = 1'b1;
  assign CLBLL_L_X52Y126_SLICE_X78Y126_D3 = 1'b1;
  assign CLBLL_L_X52Y126_SLICE_X78Y126_D4 = 1'b1;
  assign CLBLM_L_X8Y118_SLICE_X11Y118_C1 = 1'b1;
  assign CLBLM_L_X8Y118_SLICE_X11Y118_C2 = 1'b1;
  assign CLBLM_L_X8Y118_SLICE_X11Y118_C3 = 1'b1;
  assign CLBLM_L_X8Y118_SLICE_X11Y118_C4 = 1'b1;
  assign CLBLM_L_X8Y118_SLICE_X11Y118_C5 = 1'b1;
  assign CLBLM_L_X10Y128_SLICE_X12Y128_A5 = 1'b1;
  assign CLBLM_L_X8Y118_SLICE_X11Y118_C6 = 1'b1;
  assign CLBLM_L_X8Y118_SLICE_X11Y118_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X10Y128_SLICE_X12Y128_A1 = 1'b1;
  assign CLBLM_L_X10Y128_SLICE_X12Y128_A2 = 1'b1;
  assign CLBLM_L_X10Y128_SLICE_X12Y128_A3 = 1'b1;
  assign CLBLM_L_X8Y118_SLICE_X10Y118_A3 = CLBLM_L_X8Y118_SLICE_X10Y118_AQ;
  assign CLBLM_L_X10Y128_SLICE_X12Y128_A4 = 1'b1;
  assign CLBLM_L_X10Y128_SLICE_X12Y128_B3 = 1'b1;
  assign CLBLM_L_X10Y128_SLICE_X12Y128_B4 = 1'b1;
  assign CLBLM_L_X10Y128_SLICE_X12Y128_B5 = 1'b1;
  assign CLBLM_L_X10Y128_SLICE_X12Y128_B6 = 1'b1;
  assign CLBLM_L_X8Y118_SLICE_X11Y118_D2 = 1'b1;
  assign CLBLM_L_X8Y118_SLICE_X10Y118_A4 = CLBLM_R_X11Y121_SLICE_X14Y121_CO6;
  assign CLBLM_L_X8Y118_SLICE_X11Y118_D4 = 1'b1;
  assign CLBLL_L_X52Y126_SLICE_X79Y126_A1 = 1'b1;
  assign CLBLM_L_X10Y128_SLICE_X12Y128_C1 = 1'b1;
  assign CLBLM_L_X10Y128_SLICE_X12Y128_C2 = 1'b1;
  assign CLBLM_L_X10Y128_SLICE_X12Y128_C3 = 1'b1;
  assign CLBLM_L_X10Y128_SLICE_X12Y128_C4 = 1'b1;
  assign CLBLM_L_X10Y128_SLICE_X12Y128_C5 = 1'b1;
  assign CLBLM_L_X10Y128_SLICE_X12Y128_C6 = 1'b1;
  assign CLBLL_L_X2Y110_SLICE_X0Y110_A1 = 1'b1;
  assign CLBLL_L_X2Y110_SLICE_X0Y110_A2 = 1'b1;
  assign CLBLL_L_X2Y110_SLICE_X0Y110_A3 = CLBLM_R_X3Y111_SLICE_X3Y111_CO6;
  assign CLBLL_L_X2Y110_SLICE_X0Y110_A4 = CLBLL_L_X2Y110_SLICE_X0Y110_BO6;
  assign CLBLL_L_X2Y110_SLICE_X0Y110_A5 = CLBLL_L_X4Y121_SLICE_X5Y121_BO5;
  assign CLBLM_L_X8Y118_SLICE_X10Y118_A6 = CLBLM_L_X8Y119_SLICE_X11Y119_CQ;
  assign CLBLM_L_X10Y128_SLICE_X12Y128_D1 = 1'b1;
  assign CLBLM_L_X10Y128_SLICE_X12Y128_D2 = 1'b1;
  assign CLBLM_L_X10Y128_SLICE_X12Y128_D3 = 1'b1;
  assign CLBLM_L_X10Y128_SLICE_X12Y128_D4 = 1'b1;
  assign CLBLM_L_X10Y128_SLICE_X12Y128_D5 = 1'b1;
  assign CLBLM_L_X10Y128_SLICE_X12Y128_D6 = 1'b1;
  assign CLBLL_L_X2Y110_SLICE_X0Y110_B1 = LIOB33_X0Y51_IOB_X0Y51_I;
  assign CLBLL_L_X2Y110_SLICE_X0Y110_B2 = CLBLM_R_X3Y111_SLICE_X2Y111_CO6;
  assign CLBLL_L_X2Y110_SLICE_X0Y110_B3 = CLBLL_L_X2Y120_SLICE_X0Y120_CO6;
  assign CLBLL_L_X2Y110_SLICE_X0Y110_B4 = LIOB33_X0Y53_IOB_X0Y53_I;
  assign CLBLL_L_X2Y110_SLICE_X0Y110_C2 = 1'b1;
  assign CLBLL_L_X2Y110_SLICE_X0Y110_C1 = 1'b1;
  assign CLBLL_L_X2Y110_SLICE_X0Y110_C3 = 1'b1;
  assign CLBLL_L_X2Y110_SLICE_X0Y110_C5 = 1'b1;
  assign CLBLL_L_X2Y110_SLICE_X0Y110_C6 = 1'b1;
  assign CLBLM_L_X8Y118_SLICE_X10Y118_B1 = 1'b1;
  assign CLBLM_L_X8Y118_SLICE_X10Y118_B2 = CLBLM_L_X8Y118_SLICE_X10Y118_BQ;
  assign CLBLL_L_X2Y110_SLICE_X0Y110_C4 = 1'b1;
  assign CLBLL_L_X52Y126_SLICE_X79Y126_D4 = 1'b1;
  assign CLBLM_L_X8Y118_SLICE_X10Y118_B3 = CLBLM_R_X11Y121_SLICE_X14Y121_CO6;
  assign CLBLL_L_X52Y126_SLICE_X79Y126_D5 = 1'b1;
  assign CLBLL_L_X52Y126_SLICE_X79Y126_D6 = 1'b1;
  assign CLBLL_L_X52Y126_SLICE_X79Y126_D1 = 1'b1;
  assign CLBLL_L_X52Y126_SLICE_X79Y126_D2 = 1'b1;
  assign CLBLM_L_X8Y118_SLICE_X10Y118_B4 = CLBLM_L_X10Y112_SLICE_X12Y112_CQ;
  assign CLBLL_L_X2Y110_SLICE_X0Y110_D1 = 1'b1;
  assign CLBLL_L_X2Y110_SLICE_X0Y110_D2 = 1'b1;
  assign CLBLM_L_X8Y118_SLICE_X10Y118_B5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLL_L_X2Y110_SLICE_X0Y110_D3 = 1'b1;
  assign CLBLL_L_X2Y110_SLICE_X0Y110_D4 = 1'b1;
  assign CLBLL_L_X2Y110_SLICE_X0Y110_D5 = 1'b1;
  assign CLBLL_L_X2Y110_SLICE_X0Y110_D6 = 1'b1;
  assign CLBLM_L_X8Y118_SLICE_X10Y118_B6 = CLBLM_L_X10Y116_SLICE_X12Y116_CQ;
  assign RIOB33_X105Y173_IOB_X1Y173_O = CLBLM_R_X103Y172_SLICE_X163Y172_AO5;
  assign CLBLM_L_X8Y128_SLICE_X10Y128_D5 = 1'b1;
  assign CLBLL_L_X2Y110_SLICE_X1Y110_A1 = 1'b1;
  assign CLBLL_L_X2Y110_SLICE_X1Y110_A2 = 1'b1;
  assign CLBLL_L_X2Y110_SLICE_X1Y110_A3 = 1'b1;
  assign CLBLL_L_X2Y110_SLICE_X1Y110_A4 = 1'b1;
  assign CLBLL_L_X2Y110_SLICE_X1Y110_A5 = 1'b1;
  assign CLBLL_L_X2Y110_SLICE_X1Y110_A6 = 1'b1;
  assign CLBLM_R_X11Y122_SLICE_X15Y122_A1 = 1'b1;
  assign CLBLM_L_X8Y118_SLICE_X10Y118_C1 = CLBLM_L_X8Y115_SLICE_X11Y115_BQ;
  assign CLBLM_R_X11Y122_SLICE_X15Y122_A2 = 1'b1;
  assign CLBLL_L_X2Y110_SLICE_X1Y110_B1 = 1'b1;
  assign CLBLL_L_X2Y110_SLICE_X1Y110_B2 = 1'b1;
  assign CLBLL_L_X2Y110_SLICE_X1Y110_B3 = 1'b1;
  assign CLBLL_L_X2Y110_SLICE_X1Y110_B4 = 1'b1;
  assign CLBLL_L_X2Y110_SLICE_X1Y110_B5 = 1'b1;
  assign CLBLL_L_X2Y110_SLICE_X1Y110_B6 = 1'b1;
  assign CLBLM_L_X8Y118_SLICE_X10Y118_C2 = CLBLM_L_X8Y118_SLICE_X10Y118_CQ;
  assign CLBLM_L_X8Y118_SLICE_X10Y118_C3 = CLBLM_R_X11Y118_SLICE_X15Y118_CQ;
  assign CLBLM_R_X11Y122_SLICE_X15Y122_B1 = 1'b1;
  assign CLBLL_L_X2Y110_SLICE_X1Y110_C1 = 1'b1;
  assign CLBLL_L_X2Y110_SLICE_X1Y110_C2 = 1'b1;
  assign CLBLM_L_X8Y118_SLICE_X10Y118_C4 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLL_L_X2Y110_SLICE_X1Y110_C3 = 1'b1;
  assign CLBLL_L_X2Y110_SLICE_X1Y110_C4 = 1'b1;
  assign CLBLL_L_X2Y110_SLICE_X1Y110_C5 = 1'b1;
  assign CLBLL_L_X2Y110_SLICE_X1Y110_C6 = 1'b1;
  assign CLBLM_L_X8Y118_SLICE_X10Y118_C5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y112_SLICE_X9Y112_A1 = CLBLM_R_X3Y118_SLICE_X2Y118_AQ;
  assign CLBLM_R_X7Y112_SLICE_X9Y112_A2 = CLBLM_R_X7Y110_SLICE_X9Y110_BQ;
  assign CLBLM_R_X7Y112_SLICE_X9Y112_A3 = CLBLM_R_X7Y112_SLICE_X9Y112_AQ;
  assign CLBLM_R_X7Y112_SLICE_X9Y112_A4 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_L_X8Y118_SLICE_X10Y118_C6 = CLBLM_R_X3Y118_SLICE_X2Y118_AQ;
  assign CLBLM_R_X7Y112_SLICE_X9Y112_A6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLL_L_X2Y110_SLICE_X1Y110_D1 = 1'b1;
  assign CLBLL_L_X2Y110_SLICE_X1Y110_D2 = 1'b1;
  assign CLBLL_L_X2Y110_SLICE_X1Y110_D3 = 1'b1;
  assign CLBLL_L_X2Y110_SLICE_X1Y110_D4 = 1'b1;
  assign CLBLL_L_X2Y110_SLICE_X1Y110_D5 = 1'b1;
  assign CLBLL_L_X2Y110_SLICE_X1Y110_D6 = 1'b1;
  assign CLBLM_R_X7Y112_SLICE_X9Y112_B3 = 1'b1;
  assign CLBLM_R_X7Y112_SLICE_X9Y112_B4 = CLBLM_R_X5Y122_SLICE_X7Y122_BQ;
  assign CLBLM_R_X7Y112_SLICE_X9Y112_B6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y112_SLICE_X9Y112_C1 = 1'b1;
  assign CLBLM_R_X7Y112_SLICE_X9Y112_C2 = CLBLM_R_X7Y112_SLICE_X9Y112_CQ;
  assign CLBLM_R_X7Y112_SLICE_X9Y112_C3 = CLBLM_R_X5Y111_SLICE_X7Y111_DO6;
  assign CLBLM_R_X7Y112_SLICE_X9Y112_C4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y112_SLICE_X9Y112_C5 = CLBLM_L_X10Y115_SLICE_X12Y115_AQ;
  assign CLBLM_R_X7Y112_SLICE_X9Y112_C6 = CLBLM_R_X3Y115_SLICE_X3Y115_CQ;
  assign CLBLM_L_X8Y118_SLICE_X10Y118_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X7Y112_SLICE_X9Y112_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X7Y112_SLICE_X9Y112_D1 = CLBLM_R_X7Y109_SLICE_X8Y109_AQ;
  assign CLBLM_R_X7Y112_SLICE_X9Y112_D2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y112_SLICE_X9Y112_D3 = 1'b1;
  assign CLBLM_R_X7Y112_SLICE_X9Y112_D4 = CLBLM_R_X5Y116_SLICE_X7Y116_CQ;
  assign CLBLM_R_X7Y112_SLICE_X9Y112_D5 = CLBLM_R_X3Y118_SLICE_X2Y118_AQ;
  assign CLBLM_R_X7Y112_SLICE_X9Y112_D6 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_R_X11Y122_SLICE_X14Y122_A5 = CLBLM_R_X7Y128_SLICE_X8Y128_AQ;
  assign CLBLM_R_X11Y122_SLICE_X14Y122_A6 = RIOB33_X105Y141_IOB_X1Y142_I;
  assign CLBLM_R_X11Y122_SLICE_X14Y122_B1 = CLBLM_R_X11Y123_SLICE_X14Y123_BO5;
  assign CLBLM_R_X11Y122_SLICE_X14Y122_B2 = CLBLM_L_X10Y121_SLICE_X13Y121_BQ;
  assign CLBLM_R_X11Y122_SLICE_X14Y122_B3 = CLBLM_R_X11Y123_SLICE_X14Y123_AO5;
  assign CLBLM_R_X7Y112_SLICE_X8Y112_A1 = CLBLM_R_X3Y118_SLICE_X2Y118_AQ;
  assign CLBLM_R_X7Y112_SLICE_X8Y112_A2 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_R_X7Y112_SLICE_X8Y112_A3 = CLBLM_R_X7Y112_SLICE_X8Y112_AQ;
  assign CLBLM_R_X7Y112_SLICE_X8Y112_A4 = CLBLM_R_X7Y112_SLICE_X9Y112_BQ;
  assign CLBLM_R_X7Y112_SLICE_X8Y112_A5 = CLBLM_R_X3Y112_SLICE_X3Y112_BQ;
  assign CLBLM_R_X7Y112_SLICE_X8Y112_A6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X11Y122_SLICE_X14Y122_C1 = 1'b1;
  assign CLBLM_R_X11Y122_SLICE_X14Y122_C2 = 1'b1;
  assign CLBLM_R_X7Y112_SLICE_X8Y112_B1 = CLBLM_R_X7Y113_SLICE_X9Y113_DO6;
  assign CLBLM_R_X7Y112_SLICE_X8Y112_B2 = CLBLM_R_X7Y112_SLICE_X8Y112_BQ;
  assign CLBLM_R_X7Y112_SLICE_X8Y112_B3 = CLBLM_R_X7Y109_SLICE_X8Y109_BQ;
  assign CLBLM_R_X7Y112_SLICE_X8Y112_B4 = CLBLM_R_X5Y115_SLICE_X7Y115_A5Q;
  assign CLBLM_R_X7Y112_SLICE_X8Y112_B5 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X7Y112_SLICE_X8Y112_B6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X11Y122_SLICE_X14Y122_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X11Y122_SLICE_X14Y122_D1 = 1'b1;
  assign CLBLM_L_X8Y118_SLICE_X10Y118_D1 = CLBLM_L_X8Y120_SLICE_X11Y120_AQ;
  assign CLBLM_R_X7Y112_SLICE_X8Y112_C1 = CLBLM_R_X5Y111_SLICE_X7Y111_CO5;
  assign CLBLM_R_X7Y112_SLICE_X8Y112_C2 = CLBLM_R_X7Y112_SLICE_X8Y112_CQ;
  assign CLBLM_R_X7Y112_SLICE_X8Y112_C3 = CLBLM_R_X3Y118_SLICE_X2Y118_AQ;
  assign CLBLM_L_X8Y118_SLICE_X10Y118_D2 = CLBLM_L_X10Y122_SLICE_X12Y122_BQ;
  assign CLBLM_R_X7Y112_SLICE_X8Y112_C4 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_R_X7Y112_SLICE_X8Y112_C5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y112_SLICE_X8Y112_C6 = CLBLL_L_X2Y112_SLICE_X1Y112_BQ;
  assign CLBLM_R_X11Y122_SLICE_X14Y122_D3 = 1'b1;
  assign CLBLM_L_X8Y118_SLICE_X10Y118_D3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y112_SLICE_X8Y112_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X11Y122_SLICE_X14Y122_D6 = 1'b1;
  assign CLBLM_L_X8Y118_SLICE_X10Y118_D4 = CLBLM_R_X7Y111_SLICE_X8Y111_CQ;
  assign CLBLM_R_X7Y112_SLICE_X8Y112_D1 = CLBLM_R_X7Y109_SLICE_X8Y109_AQ;
  assign CLBLM_R_X7Y112_SLICE_X8Y112_D2 = CLBLM_R_X5Y116_SLICE_X7Y116_CQ;
  assign CLBLM_L_X8Y118_SLICE_X10Y118_D5 = CLBLM_L_X10Y116_SLICE_X12Y116_CQ;
  assign CLBLM_R_X7Y112_SLICE_X8Y112_D3 = CLBLM_R_X7Y115_SLICE_X8Y115_DO6;
  assign CLBLM_R_X7Y112_SLICE_X8Y112_D4 = CLBLM_R_X5Y110_SLICE_X7Y110_AO5;
  assign CLBLM_R_X7Y112_SLICE_X8Y112_D5 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X7Y112_SLICE_X8Y112_D6 = CLBLL_L_X2Y120_SLICE_X0Y120_CO6;
  assign CLBLM_L_X8Y118_SLICE_X10Y118_D6 = 1'b1;
  assign LIOI3_X0Y75_ILOGIC_X0Y76_D = LIOB33_X0Y75_IOB_X0Y76_I;
  assign LIOI3_X0Y75_ILOGIC_X0Y75_D = LIOB33_X0Y75_IOB_X0Y75_I;
  assign CLBLM_L_X8Y119_SLICE_X11Y119_A1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y119_SLICE_X11Y119_A2 = CLBLM_R_X11Y121_SLICE_X14Y121_CO6;
  assign CLBLM_L_X8Y119_SLICE_X11Y119_A3 = CLBLM_L_X8Y119_SLICE_X11Y119_AQ;
  assign CLBLM_L_X8Y119_SLICE_X11Y119_A4 = CLBLM_L_X10Y120_SLICE_X12Y120_AQ;
  assign CLBLM_L_X8Y119_SLICE_X11Y119_A5 = CLBLM_R_X7Y119_SLICE_X8Y119_BQ;
  assign CLBLM_L_X8Y119_SLICE_X11Y119_A6 = 1'b1;
  assign CLBLM_L_X8Y119_SLICE_X11Y119_B1 = CLBLM_L_X8Y118_SLICE_X11Y118_BO5;
  assign CLBLM_L_X8Y119_SLICE_X11Y119_B2 = 1'b1;
  assign CLBLM_L_X8Y119_SLICE_X11Y119_B3 = CLBLM_L_X12Y120_SLICE_X17Y120_AQ;
  assign CLBLM_L_X8Y119_SLICE_X11Y119_B4 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X8Y119_SLICE_X11Y119_B5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y119_SLICE_X11Y119_B6 = CLBLM_L_X8Y121_SLICE_X10Y121_CQ;
  assign CLBLM_L_X8Y119_SLICE_X11Y119_C1 = CLBLM_R_X7Y116_SLICE_X8Y116_BQ;
  assign CLBLM_L_X8Y119_SLICE_X11Y119_C2 = CLBLM_L_X10Y119_SLICE_X13Y119_DQ;
  assign CLBLM_L_X8Y119_SLICE_X11Y119_C3 = CLBLM_R_X7Y121_SLICE_X9Y121_A5Q;
  assign CLBLM_L_X8Y119_SLICE_X11Y119_C4 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X8Y119_SLICE_X11Y119_C5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y119_SLICE_X11Y119_C6 = 1'b1;
  assign CLBLM_L_X8Y119_SLICE_X11Y119_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X8Y119_SLICE_X11Y119_D1 = CLBLM_L_X8Y116_SLICE_X11Y116_BQ;
  assign CLBLM_L_X8Y119_SLICE_X11Y119_D2 = CLBLM_L_X10Y123_SLICE_X12Y123_AO6;
  assign CLBLM_L_X8Y119_SLICE_X11Y119_D3 = CLBLM_L_X8Y122_SLICE_X11Y122_CO6;
  assign CLBLM_L_X8Y119_SLICE_X11Y119_D4 = CLBLM_R_X5Y118_SLICE_X7Y118_CO6;
  assign CLBLM_L_X8Y119_SLICE_X11Y119_D5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y119_SLICE_X11Y119_D6 = CLBLM_R_X3Y117_SLICE_X3Y117_BQ;
  assign CLBLM_L_X8Y119_SLICE_X10Y119_A1 = RIOB33_X105Y131_IOB_X1Y131_I;
  assign CLBLM_L_X8Y119_SLICE_X10Y119_A2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y119_SLICE_X10Y119_A3 = RIOB33_X105Y135_IOB_X1Y135_I;
  assign CLBLL_L_X2Y111_SLICE_X0Y111_A1 = RIOB33_X105Y129_IOB_X1Y129_I;
  assign CLBLL_L_X2Y111_SLICE_X0Y111_A2 = RIOB33_X105Y127_IOB_X1Y128_I;
  assign CLBLL_L_X2Y111_SLICE_X0Y111_A3 = CLBLL_L_X4Y120_SLICE_X4Y120_AO6;
  assign CLBLM_L_X8Y119_SLICE_X10Y119_A4 = RIOB33_X105Y135_IOB_X1Y136_I;
  assign CLBLM_L_X8Y119_SLICE_X10Y119_A5 = CLBLM_L_X8Y121_SLICE_X10Y121_DO6;
  assign CLBLM_L_X8Y119_SLICE_X10Y119_A6 = CLBLM_L_X10Y119_SLICE_X13Y119_CQ;
  assign CLBLM_L_X8Y119_SLICE_X10Y119_AX = CLBLM_L_X8Y119_SLICE_X10Y119_DO6;
  assign CLBLL_L_X2Y111_SLICE_X0Y111_A4 = CLBLM_R_X3Y119_SLICE_X2Y119_AO6;
  assign CLBLM_L_X8Y119_SLICE_X10Y119_B1 = CLBLM_L_X12Y120_SLICE_X17Y120_CO6;
  assign CLBLL_L_X2Y111_SLICE_X0Y111_B1 = CLBLL_L_X2Y119_SLICE_X0Y119_BO6;
  assign CLBLL_L_X2Y111_SLICE_X0Y111_B2 = RIOB33_X105Y127_IOB_X1Y128_I;
  assign CLBLL_L_X2Y111_SLICE_X0Y111_B3 = CLBLL_L_X4Y121_SLICE_X5Y121_BO5;
  assign CLBLL_L_X2Y111_SLICE_X0Y111_B4 = RIOB33_X105Y129_IOB_X1Y129_I;
  assign CLBLL_L_X2Y111_SLICE_X0Y111_B5 = RIOB33_X105Y137_IOB_X1Y137_I;
  assign CLBLL_L_X2Y111_SLICE_X0Y111_B6 = 1'b1;
  assign CLBLM_L_X8Y119_SLICE_X10Y119_B2 = 1'b1;
  assign CLBLM_L_X8Y119_SLICE_X10Y119_B3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y119_SLICE_X10Y119_C1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLL_L_X2Y111_SLICE_X0Y111_C1 = CLBLL_L_X2Y120_SLICE_X0Y120_CO6;
  assign CLBLL_L_X2Y111_SLICE_X0Y111_C2 = CLBLM_R_X3Y120_SLICE_X3Y120_BO6;
  assign CLBLL_L_X2Y111_SLICE_X0Y111_C3 = RIOB33_X105Y127_IOB_X1Y128_I;
  assign CLBLL_L_X2Y111_SLICE_X0Y111_C4 = RIOB33_X105Y137_IOB_X1Y137_I;
  assign CLBLL_L_X2Y111_SLICE_X0Y111_C5 = RIOB33_X105Y129_IOB_X1Y129_I;
  assign CLBLL_L_X2Y111_SLICE_X0Y111_C6 = 1'b1;
  assign CLBLM_L_X8Y119_SLICE_X10Y119_C2 = CLBLM_L_X10Y119_SLICE_X13Y119_CQ;
  assign CLBLM_L_X8Y119_SLICE_X10Y119_C3 = CLBLM_L_X8Y120_SLICE_X10Y120_DQ;
  assign CLBLM_L_X8Y119_SLICE_X10Y119_C4 = 1'b1;
  assign CLBLM_L_X8Y119_SLICE_X10Y119_C5 = CLBLM_L_X12Y120_SLICE_X17Y120_CO6;
  assign CLBLM_L_X8Y119_SLICE_X10Y119_C6 = 1'b1;
  assign CLBLM_L_X8Y119_SLICE_X10Y119_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLL_L_X2Y111_SLICE_X0Y111_D1 = RIOB33_X105Y137_IOB_X1Y137_I;
  assign CLBLL_L_X2Y111_SLICE_X0Y111_D2 = CLBLL_L_X2Y120_SLICE_X1Y120_DO6;
  assign CLBLL_L_X2Y111_SLICE_X0Y111_D3 = RIOB33_X105Y127_IOB_X1Y128_I;
  assign CLBLL_L_X2Y111_SLICE_X0Y111_D4 = CLBLL_L_X4Y120_SLICE_X5Y120_DO6;
  assign CLBLL_L_X2Y111_SLICE_X0Y111_D5 = RIOB33_X105Y129_IOB_X1Y129_I;
  assign CLBLL_L_X2Y111_SLICE_X0Y111_D6 = 1'b1;
  assign CLBLM_L_X8Y119_SLICE_X10Y119_D1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y119_SLICE_X10Y119_D4 = CLBLM_L_X8Y110_SLICE_X10Y110_AQ;
  assign CLBLM_L_X8Y119_SLICE_X10Y119_D5 = CLBLM_L_X10Y119_SLICE_X12Y119_AQ;
  assign CLBLM_L_X8Y119_SLICE_X10Y119_D6 = 1'b1;
  assign CLBLL_L_X2Y111_SLICE_X1Y111_A1 = 1'b1;
  assign CLBLL_L_X2Y111_SLICE_X1Y111_A2 = 1'b1;
  assign CLBLL_L_X2Y111_SLICE_X1Y111_A3 = 1'b1;
  assign CLBLL_L_X2Y111_SLICE_X1Y111_A4 = 1'b1;
  assign CLBLL_L_X2Y111_SLICE_X1Y111_A5 = 1'b1;
  assign CLBLL_L_X2Y111_SLICE_X1Y111_A6 = 1'b1;
  assign CLBLM_R_X11Y123_SLICE_X15Y123_A1 = 1'b1;
  assign CLBLM_R_X11Y123_SLICE_X15Y123_A2 = 1'b1;
  assign CLBLM_R_X11Y123_SLICE_X15Y123_A3 = 1'b1;
  assign CLBLL_L_X2Y111_SLICE_X1Y111_B1 = 1'b1;
  assign CLBLL_L_X2Y111_SLICE_X1Y111_B2 = 1'b1;
  assign CLBLL_L_X2Y111_SLICE_X1Y111_B3 = 1'b1;
  assign CLBLL_L_X2Y111_SLICE_X1Y111_B4 = 1'b1;
  assign CLBLL_L_X2Y111_SLICE_X1Y111_B5 = 1'b1;
  assign CLBLL_L_X2Y111_SLICE_X1Y111_B6 = 1'b1;
  assign CLBLM_R_X11Y123_SLICE_X15Y123_A4 = 1'b1;
  assign CLBLM_R_X11Y123_SLICE_X15Y123_A5 = 1'b1;
  assign CLBLM_R_X11Y123_SLICE_X15Y123_A6 = 1'b1;
  assign CLBLL_L_X2Y111_SLICE_X1Y111_C1 = 1'b1;
  assign CLBLL_L_X2Y111_SLICE_X1Y111_C2 = 1'b1;
  assign CLBLL_L_X2Y111_SLICE_X1Y111_C3 = 1'b1;
  assign CLBLL_L_X2Y111_SLICE_X1Y111_C4 = 1'b1;
  assign CLBLL_L_X2Y111_SLICE_X1Y111_C5 = 1'b1;
  assign CLBLL_L_X2Y111_SLICE_X1Y111_C6 = 1'b1;
  assign CLBLM_R_X7Y113_SLICE_X9Y113_A1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y113_SLICE_X9Y113_A2 = CLBLL_L_X2Y120_SLICE_X0Y120_CO6;
  assign CLBLM_R_X7Y113_SLICE_X9Y113_A3 = CLBLM_R_X11Y114_SLICE_X14Y114_BQ;
  assign CLBLM_R_X7Y113_SLICE_X9Y113_A4 = CLBLM_L_X8Y114_SLICE_X10Y114_AQ;
  assign CLBLM_R_X7Y113_SLICE_X9Y113_A5 = CLBLM_L_X10Y113_SLICE_X13Y113_BO6;
  assign CLBLM_R_X7Y113_SLICE_X9Y113_A6 = 1'b1;
  assign CLBLL_L_X2Y111_SLICE_X1Y111_D1 = 1'b1;
  assign CLBLL_L_X2Y111_SLICE_X1Y111_D2 = 1'b1;
  assign CLBLL_L_X2Y111_SLICE_X1Y111_D3 = 1'b1;
  assign CLBLL_L_X2Y111_SLICE_X1Y111_D4 = 1'b1;
  assign CLBLL_L_X2Y111_SLICE_X1Y111_D5 = 1'b1;
  assign CLBLL_L_X2Y111_SLICE_X1Y111_D6 = 1'b1;
  assign CLBLM_R_X7Y113_SLICE_X9Y113_B1 = CLBLM_R_X5Y113_SLICE_X6Y113_DO6;
  assign CLBLM_R_X7Y113_SLICE_X9Y113_B2 = CLBLM_R_X7Y113_SLICE_X9Y113_BQ;
  assign CLBLM_R_X7Y113_SLICE_X9Y113_B3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y113_SLICE_X9Y113_B4 = CLBLM_R_X3Y118_SLICE_X2Y118_AQ;
  assign CLBLM_R_X7Y113_SLICE_X9Y113_B5 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_R_X7Y113_SLICE_X9Y113_B6 = CLBLM_R_X11Y117_SLICE_X14Y117_CQ;
  assign CLBLM_R_X7Y113_SLICE_X9Y113_C1 = CLBLM_R_X5Y113_SLICE_X6Y113_AQ;
  assign CLBLM_R_X7Y113_SLICE_X9Y113_C2 = CLBLM_R_X5Y116_SLICE_X7Y116_CQ;
  assign CLBLM_R_X7Y113_SLICE_X9Y113_C3 = RIOB33_X105Y121_IOB_X1Y121_I;
  assign CLBLM_R_X7Y113_SLICE_X9Y113_C4 = CLBLM_R_X3Y116_SLICE_X3Y116_BQ;
  assign CLBLM_R_X7Y113_SLICE_X9Y113_C5 = CLBLM_R_X7Y112_SLICE_X9Y112_DO6;
  assign CLBLM_R_X7Y113_SLICE_X9Y113_C6 = CLBLM_R_X5Y111_SLICE_X7Y111_CO5;
  assign CLBLM_R_X7Y113_SLICE_X9Y113_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X11Y123_SLICE_X14Y123_A1 = CLBLM_L_X10Y122_SLICE_X13Y122_AQ;
  assign CLBLM_R_X11Y123_SLICE_X14Y123_A2 = CLBLM_L_X10Y122_SLICE_X13Y122_BQ;
  assign CLBLM_R_X11Y123_SLICE_X14Y123_A3 = CLBLM_R_X11Y121_SLICE_X14Y121_BO5;
  assign CLBLM_R_X7Y113_SLICE_X9Y113_D1 = 1'b1;
  assign CLBLM_R_X7Y113_SLICE_X9Y113_D2 = 1'b1;
  assign CLBLM_R_X7Y113_SLICE_X9Y113_D3 = CLBLM_R_X7Y114_SLICE_X8Y114_CO6;
  assign CLBLM_R_X7Y113_SLICE_X9Y113_D4 = CLBLM_R_X11Y116_SLICE_X14Y116_DQ;
  assign CLBLM_R_X7Y113_SLICE_X9Y113_D5 = CLBLM_L_X8Y112_SLICE_X10Y112_DQ;
  assign CLBLM_R_X7Y113_SLICE_X9Y113_D6 = CLBLM_R_X7Y112_SLICE_X8Y112_BQ;
  assign CLBLM_R_X11Y123_SLICE_X14Y123_B1 = CLBLM_L_X10Y122_SLICE_X13Y122_AQ;
  assign CLBLM_R_X11Y123_SLICE_X14Y123_B2 = CLBLM_R_X11Y121_SLICE_X14Y121_BO6;
  assign CLBLM_R_X11Y123_SLICE_X14Y123_B3 = CLBLM_L_X10Y122_SLICE_X13Y122_BQ;
  assign CLBLM_R_X11Y123_SLICE_X14Y123_B4 = CLBLM_L_X10Y122_SLICE_X13Y122_CQ;
  assign CLBLM_R_X11Y123_SLICE_X14Y123_B5 = CLBLM_L_X10Y121_SLICE_X13Y121_BQ;
  assign CLBLM_R_X11Y123_SLICE_X14Y123_B6 = 1'b1;
  assign CLBLM_R_X7Y113_SLICE_X8Y113_A1 = CLBLM_R_X7Y113_SLICE_X8Y113_BO5;
  assign CLBLM_R_X7Y113_SLICE_X8Y113_A2 = CLBLM_R_X3Y115_SLICE_X3Y115_DQ;
  assign CLBLM_R_X7Y113_SLICE_X8Y113_A3 = 1'b1;
  assign CLBLM_R_X7Y113_SLICE_X8Y113_A4 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X7Y113_SLICE_X8Y113_A5 = CLBLM_L_X8Y116_SLICE_X11Y116_A5Q;
  assign CLBLM_R_X7Y113_SLICE_X8Y113_A6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X11Y123_SLICE_X14Y123_C1 = CLBLM_R_X7Y128_SLICE_X8Y128_AQ;
  assign CLBLM_R_X11Y123_SLICE_X14Y123_C2 = 1'b1;
  assign CLBLM_R_X11Y123_SLICE_X14Y123_C3 = 1'b1;
  assign CLBLM_R_X7Y113_SLICE_X8Y113_B1 = RIOB33_X105Y121_IOB_X1Y121_I;
  assign CLBLM_R_X7Y113_SLICE_X8Y113_B2 = CLBLM_R_X7Y118_SLICE_X9Y118_CQ;
  assign CLBLM_R_X7Y113_SLICE_X8Y113_B3 = CLBLM_L_X8Y120_SLICE_X11Y120_CQ;
  assign CLBLM_R_X7Y113_SLICE_X8Y113_B4 = CLBLM_R_X7Y113_SLICE_X9Y113_BQ;
  assign CLBLM_R_X7Y113_SLICE_X8Y113_B5 = CLBLM_R_X7Y114_SLICE_X8Y114_AQ;
  assign CLBLM_R_X7Y113_SLICE_X8Y113_B6 = 1'b1;
  assign CLBLM_R_X11Y123_SLICE_X14Y123_D1 = 1'b1;
  assign CLBLM_R_X11Y123_SLICE_X14Y123_D2 = 1'b1;
  assign CLBLM_R_X11Y123_SLICE_X14Y123_D3 = 1'b1;
  assign CLBLM_R_X7Y113_SLICE_X8Y113_C1 = CLBLM_R_X7Y109_SLICE_X8Y109_AQ;
  assign CLBLM_R_X7Y113_SLICE_X8Y113_C2 = CLBLM_R_X5Y116_SLICE_X7Y116_CQ;
  assign CLBLM_R_X7Y113_SLICE_X8Y113_C3 = CLBLL_L_X2Y120_SLICE_X1Y120_DO6;
  assign CLBLM_R_X7Y113_SLICE_X8Y113_C4 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X7Y113_SLICE_X8Y113_C5 = CLBLM_R_X5Y112_SLICE_X6Y112_BO5;
  assign CLBLM_R_X7Y113_SLICE_X8Y113_C6 = CLBLM_R_X5Y110_SLICE_X7Y110_AO5;
  assign CLBLM_R_X11Y123_SLICE_X14Y123_D4 = 1'b1;
  assign CLBLM_R_X11Y123_SLICE_X14Y123_D5 = 1'b1;
  assign CLBLM_R_X11Y123_SLICE_X14Y123_D6 = 1'b1;
  assign CLBLM_R_X7Y113_SLICE_X8Y113_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign LIOI3_TBYTESRC_X0Y119_OLOGIC_X0Y119_D1 = CLBLM_L_X8Y114_SLICE_X10Y114_CQ;
  assign LIOI3_TBYTESRC_X0Y119_OLOGIC_X0Y119_T1 = 1'b1;
  assign CLBLM_R_X7Y113_SLICE_X8Y113_D1 = CLBLM_R_X7Y109_SLICE_X8Y109_AQ;
  assign CLBLM_R_X7Y113_SLICE_X8Y113_D2 = CLBLM_R_X5Y116_SLICE_X7Y116_CQ;
  assign CLBLM_R_X7Y113_SLICE_X8Y113_D3 = CLBLL_L_X4Y120_SLICE_X4Y120_AO6;
  assign CLBLM_R_X7Y113_SLICE_X8Y113_D4 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X7Y113_SLICE_X8Y113_D5 = CLBLM_R_X7Y113_SLICE_X8Y113_BO5;
  assign CLBLM_R_X7Y113_SLICE_X8Y113_D6 = CLBLM_R_X5Y110_SLICE_X7Y110_AO5;
  assign CLBLM_R_X7Y124_SLICE_X8Y124_D5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X103Y169_SLICE_X163Y169_C5 = 1'b1;
  assign CLBLM_L_X8Y120_SLICE_X11Y120_A1 = CLBLM_L_X8Y121_SLICE_X10Y121_DO6;
  assign CLBLM_L_X8Y120_SLICE_X11Y120_A2 = RIOB33_X105Y135_IOB_X1Y135_I;
  assign CLBLM_L_X8Y120_SLICE_X11Y120_A3 = RIOB33_X105Y131_IOB_X1Y131_I;
  assign CLBLM_L_X8Y120_SLICE_X11Y120_A4 = RIOB33_X105Y135_IOB_X1Y136_I;
  assign CLBLM_L_X8Y120_SLICE_X11Y120_A5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y120_SLICE_X11Y120_A6 = CLBLM_L_X8Y122_SLICE_X11Y122_A5Q;
  assign CLBLM_L_X8Y120_SLICE_X11Y120_B1 = CLBLM_L_X8Y115_SLICE_X10Y115_DQ;
  assign CLBLM_L_X8Y120_SLICE_X11Y120_B2 = CLBLM_L_X8Y120_SLICE_X11Y120_BQ;
  assign CLBLM_L_X8Y120_SLICE_X11Y120_B3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y120_SLICE_X11Y120_B4 = CLBLM_L_X10Y123_SLICE_X12Y123_AO6;
  assign CLBLM_L_X8Y120_SLICE_X11Y120_B5 = CLBLM_R_X7Y123_SLICE_X9Y123_CO6;
  assign CLBLM_L_X8Y120_SLICE_X11Y120_B6 = CLBLM_L_X10Y121_SLICE_X12Y121_BQ;
  assign CLBLM_R_X11Y122_SLICE_X15Y122_A3 = 1'b1;
  assign CLBLM_L_X8Y120_SLICE_X11Y120_C1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y120_SLICE_X11Y120_C2 = CLBLM_L_X8Y120_SLICE_X10Y120_A5Q;
  assign CLBLM_L_X8Y120_SLICE_X11Y120_C3 = CLBLM_L_X8Y115_SLICE_X11Y115_DQ;
  assign CLBLM_L_X8Y120_SLICE_X11Y120_C4 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X8Y120_SLICE_X11Y120_C5 = CLBLM_R_X7Y124_SLICE_X8Y124_AQ;
  assign CLBLM_L_X8Y120_SLICE_X11Y120_C6 = 1'b1;
  assign CLBLM_L_X8Y120_SLICE_X11Y120_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X10Y127_SLICE_X13Y127_A2 = 1'b1;
  assign RIOB33_X105Y177_IOB_X1Y177_O = CLBLM_R_X103Y177_SLICE_X163Y177_AO6;
  assign CLBLM_L_X8Y120_SLICE_X11Y120_D1 = CLBLM_L_X10Y126_SLICE_X12Y126_AQ;
  assign CLBLM_L_X8Y120_SLICE_X11Y120_D2 = 1'b1;
  assign CLBLM_L_X8Y120_SLICE_X11Y120_D3 = CLBLL_L_X4Y117_SLICE_X5Y117_DQ;
  assign CLBLM_L_X8Y120_SLICE_X11Y120_D4 = 1'b1;
  assign CLBLM_L_X8Y120_SLICE_X11Y120_D5 = 1'b1;
  assign CLBLM_L_X8Y120_SLICE_X11Y120_D6 = 1'b1;
  assign CLBLM_L_X10Y127_SLICE_X13Y127_A3 = 1'b1;
  assign CLBLM_R_X11Y122_SLICE_X15Y122_A4 = 1'b1;
  assign CLBLL_L_X2Y112_SLICE_X0Y112_A1 = 1'b1;
  assign CLBLL_L_X2Y112_SLICE_X0Y112_A2 = 1'b1;
  assign CLBLL_L_X2Y112_SLICE_X0Y112_A3 = 1'b1;
  assign CLBLL_L_X2Y112_SLICE_X0Y112_A4 = 1'b1;
  assign CLBLL_L_X2Y112_SLICE_X0Y112_A5 = 1'b1;
  assign CLBLL_L_X2Y112_SLICE_X0Y112_A6 = 1'b1;
  assign CLBLM_L_X8Y120_SLICE_X10Y120_A1 = CLBLM_L_X12Y120_SLICE_X17Y120_CO6;
  assign CLBLM_L_X8Y120_SLICE_X10Y120_A6 = 1'b1;
  assign CLBLM_L_X8Y120_SLICE_X10Y120_A2 = CLBLM_L_X8Y120_SLICE_X11Y120_CQ;
  assign CLBLL_L_X2Y112_SLICE_X0Y112_B1 = 1'b1;
  assign CLBLL_L_X2Y112_SLICE_X0Y112_B2 = 1'b1;
  assign CLBLL_L_X2Y112_SLICE_X0Y112_B3 = 1'b1;
  assign CLBLL_L_X2Y112_SLICE_X0Y112_B4 = 1'b1;
  assign CLBLL_L_X2Y112_SLICE_X0Y112_B5 = 1'b1;
  assign CLBLL_L_X2Y112_SLICE_X0Y112_B6 = 1'b1;
  assign CLBLM_L_X8Y120_SLICE_X10Y120_B1 = CLBLM_L_X10Y121_SLICE_X12Y121_BQ;
  assign CLBLM_L_X8Y120_SLICE_X10Y120_B2 = 1'b1;
  assign CLBLL_L_X2Y112_SLICE_X0Y112_C1 = 1'b1;
  assign CLBLL_L_X2Y112_SLICE_X0Y112_C2 = 1'b1;
  assign CLBLL_L_X2Y112_SLICE_X0Y112_C3 = 1'b1;
  assign CLBLL_L_X2Y112_SLICE_X0Y112_C4 = 1'b1;
  assign CLBLL_L_X2Y112_SLICE_X0Y112_C5 = 1'b1;
  assign CLBLL_L_X2Y112_SLICE_X0Y112_C6 = 1'b1;
  assign CLBLM_L_X8Y120_SLICE_X10Y120_B5 = 1'b1;
  assign CLBLM_L_X8Y120_SLICE_X10Y120_B6 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X8Y120_SLICE_X10Y120_C1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y120_SLICE_X10Y120_C2 = CLBLM_L_X8Y120_SLICE_X10Y120_CQ;
  assign CLBLM_L_X8Y120_SLICE_X10Y120_C3 = CLBLM_R_X7Y118_SLICE_X9Y118_AQ;
  assign CLBLM_L_X8Y120_SLICE_X10Y120_C4 = CLBLM_L_X8Y120_SLICE_X10Y120_A5Q;
  assign CLBLM_L_X8Y120_SLICE_X10Y120_C5 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLL_L_X2Y112_SLICE_X0Y112_D1 = 1'b1;
  assign CLBLL_L_X2Y112_SLICE_X0Y112_D2 = 1'b1;
  assign CLBLL_L_X2Y112_SLICE_X0Y112_D3 = 1'b1;
  assign CLBLL_L_X2Y112_SLICE_X0Y112_D4 = 1'b1;
  assign CLBLL_L_X2Y112_SLICE_X0Y112_D5 = 1'b1;
  assign CLBLL_L_X2Y112_SLICE_X0Y112_D6 = 1'b1;
  assign CLBLM_L_X8Y120_SLICE_X10Y120_D1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y120_SLICE_X10Y120_D2 = CLBLL_L_X2Y120_SLICE_X1Y120_DO6;
  assign CLBLM_L_X8Y120_SLICE_X10Y120_D3 = CLBLM_L_X8Y122_SLICE_X11Y122_BQ;
  assign CLBLM_L_X8Y120_SLICE_X10Y120_D4 = CLBLM_R_X7Y112_SLICE_X9Y112_AQ;
  assign CLBLM_L_X8Y120_SLICE_X10Y120_D6 = 1'b1;
  assign CLBLM_L_X8Y120_SLICE_X10Y120_D5 = CLBLL_L_X4Y120_SLICE_X5Y120_DO6;
  assign CLBLM_R_X11Y122_SLICE_X15Y122_A6 = 1'b1;
  assign RIOI3_TBYTETERM_X105Y137_ILOGIC_X1Y138_D = RIOB33_X105Y137_IOB_X1Y138_I;
  assign RIOI3_TBYTETERM_X105Y137_ILOGIC_X1Y137_D = RIOB33_X105Y137_IOB_X1Y137_I;
  assign CLBLL_L_X2Y112_SLICE_X1Y112_A1 = CLBLM_L_X8Y112_SLICE_X10Y112_CQ;
  assign CLBLL_L_X2Y112_SLICE_X1Y112_A2 = CLBLL_L_X2Y112_SLICE_X1Y112_BQ;
  assign CLBLL_L_X2Y112_SLICE_X1Y112_A3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLL_L_X2Y112_SLICE_X1Y112_A4 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLL_L_X2Y112_SLICE_X1Y112_A5 = 1'b1;
  assign CLBLL_L_X2Y112_SLICE_X1Y112_A6 = CLBLM_R_X3Y114_SLICE_X2Y114_BQ;
  assign CLBLL_L_X2Y112_SLICE_X1Y112_AX = CLBLL_L_X2Y112_SLICE_X1Y112_CO6;
  assign CLBLL_L_X2Y112_SLICE_X1Y112_B1 = CLBLM_R_X3Y112_SLICE_X3Y112_B5Q;
  assign CLBLL_L_X2Y112_SLICE_X1Y112_B2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLL_L_X2Y112_SLICE_X1Y112_B3 = 1'b1;
  assign CLBLL_L_X2Y112_SLICE_X1Y112_B4 = 1'b1;
  assign CLBLL_L_X2Y112_SLICE_X1Y112_B5 = CLBLL_L_X2Y113_SLICE_X1Y113_CQ;
  assign CLBLL_L_X2Y112_SLICE_X1Y112_B6 = CLBLM_L_X8Y112_SLICE_X10Y112_CQ;
  assign CLBLL_L_X2Y112_SLICE_X1Y112_C1 = CLBLM_L_X10Y113_SLICE_X13Y113_BO6;
  assign CLBLL_L_X2Y112_SLICE_X1Y112_C2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLL_L_X2Y112_SLICE_X1Y112_C3 = CLBLM_R_X3Y112_SLICE_X2Y112_CO6;
  assign CLBLL_L_X2Y112_SLICE_X1Y112_C4 = CLBLL_L_X2Y112_SLICE_X1Y112_A5Q;
  assign CLBLL_L_X2Y112_SLICE_X1Y112_C5 = CLBLM_R_X5Y119_SLICE_X6Y119_B5Q;
  assign CLBLL_L_X2Y112_SLICE_X1Y112_C6 = 1'b1;
  assign CLBLL_L_X2Y112_SLICE_X1Y112_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X7Y114_SLICE_X9Y114_A1 = CLBLM_R_X7Y114_SLICE_X9Y114_DO6;
  assign CLBLM_R_X7Y114_SLICE_X9Y114_A2 = CLBLL_L_X4Y115_SLICE_X5Y115_CQ;
  assign CLBLM_R_X7Y114_SLICE_X9Y114_A3 = CLBLM_R_X5Y115_SLICE_X7Y115_BQ;
  assign CLBLM_R_X7Y114_SLICE_X9Y114_A4 = CLBLM_R_X7Y114_SLICE_X9Y114_BO6;
  assign CLBLL_L_X2Y112_SLICE_X1Y112_D1 = 1'b1;
  assign CLBLL_L_X2Y112_SLICE_X1Y112_D2 = 1'b1;
  assign CLBLL_L_X2Y112_SLICE_X1Y112_D3 = 1'b1;
  assign CLBLL_L_X2Y112_SLICE_X1Y112_D4 = 1'b1;
  assign CLBLL_L_X2Y112_SLICE_X1Y112_D5 = 1'b1;
  assign CLBLL_L_X2Y112_SLICE_X1Y112_D6 = 1'b1;
  assign CLBLM_R_X7Y114_SLICE_X9Y114_A5 = CLBLM_R_X5Y119_SLICE_X6Y119_BQ;
  assign CLBLM_R_X7Y114_SLICE_X9Y114_A6 = CLBLM_R_X7Y114_SLICE_X9Y114_CO6;
  assign CLBLM_R_X7Y114_SLICE_X9Y114_B1 = CLBLM_R_X7Y115_SLICE_X8Y115_CQ;
  assign CLBLM_R_X7Y114_SLICE_X9Y114_B2 = CLBLL_L_X4Y114_SLICE_X5Y114_AQ;
  assign CLBLM_R_X7Y114_SLICE_X9Y114_B3 = CLBLM_R_X7Y109_SLICE_X8Y109_BQ;
  assign CLBLM_R_X7Y114_SLICE_X9Y114_B4 = 1'b1;
  assign CLBLM_R_X7Y114_SLICE_X9Y114_B5 = 1'b1;
  assign CLBLM_R_X7Y114_SLICE_X9Y114_B6 = CLBLM_L_X8Y114_SLICE_X11Y114_BQ;
  assign CLBLM_R_X7Y114_SLICE_X9Y114_C1 = CLBLM_L_X8Y114_SLICE_X10Y114_C5Q;
  assign CLBLM_R_X7Y114_SLICE_X9Y114_C2 = CLBLM_L_X8Y112_SLICE_X10Y112_DQ;
  assign CLBLM_R_X7Y114_SLICE_X9Y114_C3 = CLBLM_L_X8Y114_SLICE_X10Y114_BQ;
  assign CLBLM_R_X7Y114_SLICE_X9Y114_C4 = 1'b1;
  assign CLBLM_R_X7Y114_SLICE_X9Y114_C5 = 1'b1;
  assign CLBLM_R_X7Y114_SLICE_X9Y114_C6 = CLBLM_R_X7Y119_SLICE_X9Y119_CQ;
  assign CLBLM_R_X13Y120_SLICE_X19Y120_D6 = 1'b1;
  assign CLBLM_R_X7Y114_SLICE_X9Y114_D1 = CLBLM_R_X7Y120_SLICE_X8Y120_DQ;
  assign CLBLM_R_X7Y114_SLICE_X9Y114_D2 = CLBLM_R_X11Y116_SLICE_X14Y116_DQ;
  assign CLBLM_R_X7Y114_SLICE_X9Y114_D3 = CLBLM_L_X8Y114_SLICE_X10Y114_B5Q;
  assign CLBLM_R_X7Y114_SLICE_X9Y114_D4 = 1'b1;
  assign CLBLM_R_X7Y114_SLICE_X9Y114_D5 = 1'b1;
  assign CLBLM_R_X7Y114_SLICE_X9Y114_D6 = CLBLM_R_X5Y110_SLICE_X7Y110_CQ;
  assign CLBLM_R_X7Y114_SLICE_X8Y114_A1 = CLBLM_R_X7Y114_SLICE_X8Y114_DO6;
  assign CLBLM_R_X7Y114_SLICE_X8Y114_A2 = CLBLM_R_X3Y118_SLICE_X2Y118_AQ;
  assign CLBLM_R_X7Y114_SLICE_X8Y114_A3 = CLBLM_R_X7Y114_SLICE_X8Y114_AQ;
  assign CLBLM_R_X7Y114_SLICE_X8Y114_A4 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_R_X7Y114_SLICE_X8Y114_A5 = CLBLM_L_X8Y120_SLICE_X10Y120_BQ;
  assign CLBLM_R_X7Y114_SLICE_X8Y114_A6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y114_SLICE_X8Y114_B1 = CLBLM_L_X10Y115_SLICE_X12Y115_CQ;
  assign CLBLM_R_X7Y114_SLICE_X8Y114_B2 = CLBLM_R_X7Y112_SLICE_X8Y112_BQ;
  assign CLBLM_R_X7Y114_SLICE_X8Y114_B3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y114_SLICE_X8Y114_B4 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X7Y114_SLICE_X8Y114_B5 = CLBLM_R_X5Y109_SLICE_X6Y109_BQ;
  assign CLBLM_R_X7Y114_SLICE_X8Y114_B6 = CLBLM_R_X7Y114_SLICE_X8Y114_CO6;
  assign CLBLM_R_X7Y114_SLICE_X8Y114_C1 = CLBLM_R_X3Y116_SLICE_X3Y116_BQ;
  assign CLBLM_R_X7Y114_SLICE_X8Y114_C2 = CLBLM_R_X7Y114_SLICE_X9Y114_AO6;
  assign CLBLM_R_X7Y114_SLICE_X8Y114_C3 = CLBLM_R_X7Y118_SLICE_X9Y118_CQ;
  assign CLBLM_R_X7Y114_SLICE_X8Y114_C4 = CLBLM_L_X8Y114_SLICE_X11Y114_DO6;
  assign CLBLM_R_X7Y114_SLICE_X8Y114_C5 = CLBLM_L_X8Y115_SLICE_X10Y115_CQ;
  assign CLBLM_R_X7Y114_SLICE_X8Y114_C6 = CLBLL_L_X4Y115_SLICE_X4Y115_C5Q;
  assign CLBLM_R_X7Y114_SLICE_X8Y114_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign LIOB33_X0Y139_IOB_X0Y140_O = CLBLL_L_X4Y123_SLICE_X4Y123_BQ;
  assign CLBLM_R_X7Y114_SLICE_X8Y114_D1 = CLBLM_R_X3Y116_SLICE_X3Y116_BQ;
  assign CLBLM_R_X7Y114_SLICE_X8Y114_D2 = CLBLM_R_X7Y120_SLICE_X9Y120_CQ;
  assign CLBLM_R_X7Y114_SLICE_X8Y114_D3 = CLBLM_R_X7Y122_SLICE_X8Y122_DQ;
  assign CLBLM_R_X7Y114_SLICE_X8Y114_D4 = CLBLM_R_X5Y114_SLICE_X7Y114_BO5;
  assign CLBLM_R_X7Y114_SLICE_X8Y114_D5 = CLBLM_R_X5Y114_SLICE_X7Y114_AQ;
  assign CLBLM_R_X7Y114_SLICE_X8Y114_D6 = RIOB33_X105Y121_IOB_X1Y121_I;
  assign LIOB33_X0Y139_IOB_X0Y139_O = CLBLM_R_X5Y124_SLICE_X6Y124_AQ;
  assign CLBLM_R_X11Y122_SLICE_X15Y122_B2 = 1'b1;
  assign CLBLM_R_X11Y122_SLICE_X15Y122_B3 = 1'b1;
  assign CLBLM_R_X11Y122_SLICE_X15Y122_B4 = 1'b1;
  assign CLBLM_L_X10Y127_SLICE_X12Y127_A6 = 1'b1;
  assign CLBLM_L_X10Y127_SLICE_X12Y127_AX = CLBLM_L_X10Y128_SLICE_X13Y128_AO5;
  assign CLBLM_L_X8Y121_SLICE_X11Y121_A1 = CLBLM_L_X8Y120_SLICE_X11Y120_BQ;
  assign CLBLM_L_X8Y121_SLICE_X11Y121_A2 = CLBLM_L_X10Y123_SLICE_X12Y123_AO6;
  assign CLBLM_L_X8Y121_SLICE_X11Y121_A3 = CLBLM_L_X8Y121_SLICE_X11Y121_AQ;
  assign CLBLM_L_X8Y121_SLICE_X11Y121_A4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y121_SLICE_X11Y121_A5 = CLBLM_L_X8Y119_SLICE_X11Y119_C5Q;
  assign CLBLM_L_X8Y121_SLICE_X11Y121_A6 = CLBLM_R_X7Y123_SLICE_X9Y123_CO6;
  assign CLBLM_R_X11Y122_SLICE_X15Y122_B5 = 1'b1;
  assign CLBLM_L_X10Y127_SLICE_X12Y127_B1 = 1'b1;
  assign RIOB33_X105Y179_IOB_X1Y179_O = CLBLM_R_X11Y128_SLICE_X14Y128_AO5;
  assign CLBLM_L_X8Y121_SLICE_X11Y121_B1 = CLBLM_L_X10Y123_SLICE_X12Y123_AO6;
  assign CLBLM_L_X8Y121_SLICE_X11Y121_B2 = CLBLM_L_X8Y121_SLICE_X11Y121_BQ;
  assign CLBLM_L_X8Y121_SLICE_X11Y121_B3 = CLBLM_L_X8Y121_SLICE_X11Y121_AQ;
  assign CLBLM_L_X8Y121_SLICE_X11Y121_B4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y121_SLICE_X11Y121_B5 = CLBLM_R_X3Y118_SLICE_X2Y118_AQ;
  assign CLBLM_L_X8Y121_SLICE_X11Y121_B6 = CLBLM_R_X7Y123_SLICE_X9Y123_CO6;
  assign CLBLM_L_X8Y121_SLICE_X11Y121_C1 = CLBLM_L_X8Y121_SLICE_X10Y121_AQ;
  assign CLBLM_L_X8Y121_SLICE_X11Y121_C2 = CLBLM_L_X8Y121_SLICE_X11Y121_CQ;
  assign CLBLM_L_X8Y121_SLICE_X11Y121_C3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y121_SLICE_X11Y121_C4 = CLBLM_R_X7Y123_SLICE_X9Y123_CO6;
  assign CLBLM_L_X8Y121_SLICE_X11Y121_C5 = CLBLM_L_X10Y123_SLICE_X12Y123_AO6;
  assign CLBLM_L_X8Y121_SLICE_X11Y121_C6 = CLBLM_R_X5Y121_SLICE_X6Y121_AQ;
  assign CLBLM_R_X11Y122_SLICE_X15Y122_B6 = 1'b1;
  assign CLBLM_L_X8Y121_SLICE_X11Y121_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X8Y121_SLICE_X11Y121_D1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y121_SLICE_X11Y121_D2 = CLBLM_L_X10Y119_SLICE_X13Y119_DQ;
  assign CLBLM_L_X8Y121_SLICE_X11Y121_D3 = CLBLM_L_X8Y121_SLICE_X11Y121_DQ;
  assign CLBLM_L_X8Y121_SLICE_X11Y121_D4 = CLBLM_R_X7Y122_SLICE_X9Y122_AQ;
  assign CLBLM_L_X8Y121_SLICE_X11Y121_D5 = CLBLM_L_X8Y120_SLICE_X11Y120_DO6;
  assign CLBLM_L_X8Y121_SLICE_X11Y121_D6 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLL_L_X2Y113_SLICE_X0Y113_A1 = RIOB33_X105Y129_IOB_X1Y129_I;
  assign CLBLL_L_X2Y113_SLICE_X0Y113_A2 = CLBLL_L_X2Y113_SLICE_X1Y113_CQ;
  assign CLBLL_L_X2Y113_SLICE_X0Y113_A3 = RIOB33_X105Y137_IOB_X1Y137_I;
  assign CLBLL_L_X2Y113_SLICE_X0Y113_A4 = CLBLL_L_X4Y120_SLICE_X4Y120_BO6;
  assign CLBLL_L_X2Y113_SLICE_X0Y113_A5 = RIOB33_X105Y127_IOB_X1Y128_I;
  assign CLBLL_L_X2Y113_SLICE_X0Y113_A6 = 1'b1;
  assign CLBLM_L_X8Y121_SLICE_X10Y121_A1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y121_SLICE_X10Y121_A2 = CLBLM_L_X8Y114_SLICE_X10Y114_CQ;
  assign CLBLL_L_X2Y113_SLICE_X0Y113_B1 = 1'b1;
  assign CLBLL_L_X2Y113_SLICE_X0Y113_B2 = 1'b1;
  assign CLBLL_L_X2Y113_SLICE_X0Y113_B3 = 1'b1;
  assign CLBLL_L_X2Y113_SLICE_X0Y113_B4 = 1'b1;
  assign CLBLL_L_X2Y113_SLICE_X0Y113_B5 = 1'b1;
  assign CLBLL_L_X2Y113_SLICE_X0Y113_B6 = 1'b1;
  assign CLBLM_L_X8Y121_SLICE_X10Y121_A3 = CLBLM_L_X8Y121_SLICE_X10Y121_AQ;
  assign CLBLM_L_X8Y121_SLICE_X10Y121_B1 = CLBLM_L_X8Y119_SLICE_X11Y119_DQ;
  assign CLBLL_L_X2Y113_SLICE_X0Y113_C1 = 1'b1;
  assign CLBLL_L_X2Y113_SLICE_X0Y113_C2 = 1'b1;
  assign CLBLL_L_X2Y113_SLICE_X0Y113_C3 = 1'b1;
  assign CLBLL_L_X2Y113_SLICE_X0Y113_C4 = 1'b1;
  assign CLBLL_L_X2Y113_SLICE_X0Y113_C5 = 1'b1;
  assign CLBLL_L_X2Y113_SLICE_X0Y113_C6 = 1'b1;
  assign CLBLM_L_X8Y121_SLICE_X10Y121_B5 = RIOB33_X105Y121_IOB_X1Y121_I;
  assign CLBLM_L_X8Y121_SLICE_X10Y121_B2 = CLBLM_L_X8Y121_SLICE_X10Y121_BQ;
  assign CLBLM_L_X8Y121_SLICE_X10Y121_C1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y121_SLICE_X10Y121_C2 = CLBLM_L_X8Y121_SLICE_X11Y121_DQ;
  assign CLBLM_L_X8Y121_SLICE_X10Y121_C3 = 1'b1;
  assign CLBLM_L_X8Y121_SLICE_X10Y121_C4 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X8Y121_SLICE_X10Y121_C5 = CLBLM_R_X7Y117_SLICE_X9Y117_DQ;
  assign CLBLM_L_X8Y121_SLICE_X10Y121_C6 = 1'b1;
  assign CLBLL_L_X2Y113_SLICE_X0Y113_D1 = 1'b1;
  assign CLBLL_L_X2Y113_SLICE_X0Y113_D2 = 1'b1;
  assign CLBLL_L_X2Y113_SLICE_X0Y113_D3 = 1'b1;
  assign CLBLL_L_X2Y113_SLICE_X0Y113_D4 = 1'b1;
  assign CLBLL_L_X2Y113_SLICE_X0Y113_D5 = 1'b1;
  assign CLBLL_L_X2Y113_SLICE_X0Y113_D6 = 1'b1;
  assign CLBLM_L_X8Y121_SLICE_X10Y121_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X8Y121_SLICE_X10Y121_D1 = RIOB33_X105Y137_IOB_X1Y137_I;
  assign CLBLM_L_X8Y121_SLICE_X10Y121_D2 = RIOB33_X105Y131_IOB_X1Y132_I;
  assign CLBLM_L_X8Y121_SLICE_X10Y121_D3 = RIOB33_X105Y133_IOB_X1Y133_I;
  assign CLBLM_L_X8Y121_SLICE_X10Y121_D4 = RIOB33_X105Y127_IOB_X1Y128_I;
  assign CLBLM_L_X8Y121_SLICE_X10Y121_D5 = RIOB33_X105Y133_IOB_X1Y134_I;
  assign CLBLM_L_X8Y121_SLICE_X10Y121_D6 = RIOB33_X105Y129_IOB_X1Y130_I;
  assign CLBLM_R_X11Y123_SLICE_X15Y123_B2 = 1'b1;
  assign CLBLM_R_X11Y123_SLICE_X15Y123_B3 = 1'b1;
  assign CLBLM_R_X11Y123_SLICE_X15Y123_B4 = 1'b1;
  assign CLBLM_R_X11Y123_SLICE_X15Y123_B5 = 1'b1;
  assign CLBLM_R_X11Y123_SLICE_X15Y123_B6 = 1'b1;
  assign CLBLL_L_X2Y113_SLICE_X1Y113_A1 = CLBLM_R_X7Y120_SLICE_X9Y120_DQ;
  assign CLBLL_L_X2Y113_SLICE_X1Y113_A2 = 1'b1;
  assign CLBLL_L_X2Y113_SLICE_X1Y113_A3 = LIOB33_X0Y79_IOB_X0Y79_I;
  assign CLBLL_L_X2Y113_SLICE_X1Y113_A4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLL_L_X2Y113_SLICE_X1Y113_A5 = 1'b1;
  assign CLBLL_L_X2Y113_SLICE_X1Y113_A6 = CLBLL_L_X2Y113_SLICE_X1Y113_AQ;
  assign CLBLL_L_X2Y113_SLICE_X1Y113_B1 = 1'b1;
  assign CLBLL_L_X2Y113_SLICE_X1Y113_B2 = CLBLL_L_X4Y113_SLICE_X4Y113_BQ;
  assign CLBLL_L_X2Y113_SLICE_X1Y113_B3 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLL_L_X2Y113_SLICE_X1Y113_B4 = CLBLL_L_X4Y116_SLICE_X4Y116_C5Q;
  assign CLBLL_L_X2Y113_SLICE_X1Y113_B5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLL_L_X2Y113_SLICE_X1Y113_B6 = CLBLM_R_X5Y112_SLICE_X6Y112_DO6;
  assign CLBLL_L_X2Y113_SLICE_X1Y113_C1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLL_L_X2Y113_SLICE_X1Y113_C2 = CLBLL_L_X4Y113_SLICE_X4Y113_BQ;
  assign CLBLL_L_X2Y113_SLICE_X1Y113_C3 = CLBLL_L_X2Y119_SLICE_X0Y119_BO6;
  assign CLBLL_L_X2Y113_SLICE_X1Y113_C4 = CLBLM_R_X3Y114_SLICE_X3Y114_BQ;
  assign CLBLL_L_X2Y113_SLICE_X1Y113_C5 = CLBLL_L_X2Y114_SLICE_X1Y114_DO6;
  assign CLBLL_L_X2Y113_SLICE_X1Y113_C6 = 1'b1;
  assign CLBLM_R_X11Y123_SLICE_X15Y123_C1 = 1'b1;
  assign CLBLM_R_X11Y123_SLICE_X15Y123_C2 = 1'b1;
  assign CLBLL_L_X2Y113_SLICE_X1Y113_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign LIOI3_X0Y125_OLOGIC_X0Y126_D1 = CLBLM_R_X5Y124_SLICE_X6Y124_CQ;
  assign CLBLM_R_X11Y123_SLICE_X15Y123_C3 = 1'b1;
  assign CLBLL_L_X2Y113_SLICE_X1Y113_D1 = 1'b1;
  assign CLBLL_L_X2Y113_SLICE_X1Y113_D2 = 1'b1;
  assign CLBLL_L_X2Y113_SLICE_X1Y113_D3 = 1'b1;
  assign CLBLL_L_X2Y113_SLICE_X1Y113_D4 = 1'b1;
  assign CLBLL_L_X2Y113_SLICE_X1Y113_D5 = 1'b1;
  assign CLBLL_L_X2Y113_SLICE_X1Y113_D6 = 1'b1;
  assign CLBLM_R_X7Y115_SLICE_X9Y115_A1 = CLBLM_R_X7Y112_SLICE_X8Y112_AQ;
  assign CLBLM_R_X7Y115_SLICE_X9Y115_A2 = CLBLM_R_X7Y117_SLICE_X9Y117_BQ;
  assign CLBLM_R_X7Y115_SLICE_X9Y115_A3 = CLBLM_R_X7Y115_SLICE_X9Y115_AQ;
  assign CLBLM_R_X7Y115_SLICE_X9Y115_A4 = CLBLM_R_X5Y117_SLICE_X7Y117_CO6;
  assign CLBLM_R_X7Y115_SLICE_X9Y115_A5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y115_SLICE_X9Y115_A6 = 1'b1;
  assign CLBLM_R_X7Y115_SLICE_X9Y115_B1 = CLBLM_R_X7Y117_SLICE_X8Y117_A5Q;
  assign CLBLM_R_X7Y115_SLICE_X9Y115_B2 = CLBLM_R_X3Y115_SLICE_X3Y115_BQ;
  assign CLBLM_R_X7Y115_SLICE_X9Y115_B3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y115_SLICE_X9Y115_B4 = CLBLM_R_X7Y115_SLICE_X8Y115_A5Q;
  assign CLBLM_R_X7Y115_SLICE_X9Y115_B5 = CLBLM_R_X5Y118_SLICE_X7Y118_AQ;
  assign CLBLM_R_X7Y115_SLICE_X9Y115_B6 = 1'b1;
  assign CLBLM_R_X7Y115_SLICE_X9Y115_C1 = CLBLM_R_X7Y115_SLICE_X8Y115_AQ;
  assign CLBLM_R_X7Y115_SLICE_X9Y115_C2 = CLBLM_R_X7Y115_SLICE_X8Y115_A5Q;
  assign CLBLM_R_X7Y115_SLICE_X9Y115_C3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y115_SLICE_X9Y115_C4 = CLBLM_R_X3Y115_SLICE_X3Y115_CQ;
  assign CLBLM_R_X7Y115_SLICE_X9Y115_C5 = RIOB33_X105Y103_IOB_X1Y103_I;
  assign CLBLM_R_X7Y115_SLICE_X9Y115_C6 = 1'b1;
  assign CLBLM_R_X7Y115_SLICE_X9Y115_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X7Y115_SLICE_X9Y115_D1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y115_SLICE_X9Y115_D2 = CLBLM_L_X8Y123_SLICE_X11Y123_A5Q;
  assign CLBLM_R_X7Y115_SLICE_X9Y115_D3 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X7Y115_SLICE_X9Y115_D4 = CLBLM_R_X7Y114_SLICE_X8Y114_CO6;
  assign CLBLM_R_X7Y115_SLICE_X9Y115_D5 = 1'b1;
  assign CLBLM_R_X7Y115_SLICE_X9Y115_D6 = CLBLM_R_X7Y112_SLICE_X8Y112_BQ;
  assign CLBLM_R_X7Y115_SLICE_X8Y115_A1 = CLBLM_R_X3Y118_SLICE_X2Y118_AQ;
  assign CLBLM_R_X7Y115_SLICE_X8Y115_A2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y115_SLICE_X8Y115_A3 = CLBLM_R_X7Y115_SLICE_X8Y115_AQ;
  assign CLBLM_R_X7Y115_SLICE_X8Y115_A4 = CLBLM_R_X5Y114_SLICE_X7Y114_CO6;
  assign CLBLM_R_X7Y115_SLICE_X8Y115_A5 = CLBLM_R_X5Y119_SLICE_X6Y119_BQ;
  assign CLBLM_R_X7Y115_SLICE_X8Y115_A6 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign LIOI3_X0Y125_OLOGIC_X0Y126_T1 = 1'b1;
  assign CLBLM_R_X7Y115_SLICE_X8Y115_AX = CLBLM_L_X8Y117_SLICE_X10Y117_DO6;
  assign CLBLM_R_X7Y115_SLICE_X8Y115_B1 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X7Y115_SLICE_X8Y115_B2 = CLBLM_R_X7Y113_SLICE_X8Y113_BO6;
  assign CLBLM_R_X7Y115_SLICE_X8Y115_B3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y115_SLICE_X8Y115_B4 = 1'b1;
  assign CLBLM_R_X7Y115_SLICE_X8Y115_B5 = CLBLM_R_X7Y115_SLICE_X9Y115_AQ;
  assign CLBLM_R_X7Y115_SLICE_X8Y115_B6 = CLBLL_L_X4Y115_SLICE_X5Y115_BQ;
  assign CLBLM_R_X11Y123_SLICE_X15Y123_D1 = 1'b1;
  assign CLBLM_R_X11Y123_SLICE_X15Y123_D2 = 1'b1;
  assign CLBLM_R_X7Y115_SLICE_X8Y115_C1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y115_SLICE_X8Y115_C2 = 1'b1;
  assign CLBLM_R_X7Y115_SLICE_X8Y115_C3 = CLBLM_R_X7Y122_SLICE_X8Y122_BQ;
  assign CLBLM_R_X7Y115_SLICE_X8Y115_C4 = 1'b1;
  assign CLBLM_R_X7Y115_SLICE_X8Y115_C5 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X7Y115_SLICE_X8Y115_C6 = CLBLL_L_X4Y115_SLICE_X4Y115_C5Q;
  assign CLBLM_R_X11Y123_SLICE_X15Y123_D3 = 1'b1;
  assign CLBLM_R_X11Y123_SLICE_X15Y123_D4 = 1'b1;
  assign CLBLM_R_X7Y115_SLICE_X8Y115_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X11Y123_SLICE_X15Y123_D5 = 1'b1;
  assign CLBLM_R_X7Y115_SLICE_X8Y115_D1 = CLBLM_L_X8Y114_SLICE_X10Y114_BQ;
  assign CLBLM_R_X7Y115_SLICE_X8Y115_D2 = RIOB33_X105Y121_IOB_X1Y121_I;
  assign CLBLM_R_X7Y115_SLICE_X8Y115_D3 = CLBLM_R_X5Y111_SLICE_X7Y111_BQ;
  assign CLBLM_R_X7Y115_SLICE_X8Y115_D4 = CLBLL_L_X4Y114_SLICE_X5Y114_AQ;
  assign CLBLM_R_X7Y115_SLICE_X8Y115_D5 = CLBLM_R_X5Y116_SLICE_X7Y116_A5Q;
  assign CLBLM_R_X7Y115_SLICE_X8Y115_D6 = 1'b1;
  assign CLBLM_R_X11Y123_SLICE_X15Y123_D6 = 1'b1;
  assign LIOI3_X0Y189_OLOGIC_X0Y190_D1 = RIOB33_X105Y147_IOB_X1Y147_I;
  assign CLBLM_R_X11Y122_SLICE_X15Y122_C5 = 1'b1;
  assign LIOI3_X0Y125_OLOGIC_X0Y125_D1 = CLBLM_R_X7Y115_SLICE_X9Y115_CQ;
  assign LIOI3_X0Y189_OLOGIC_X0Y190_T1 = 1'b1;
  assign LIOI3_X0Y127_OLOGIC_X0Y128_D1 = CLBLL_L_X2Y117_SLICE_X0Y117_A5Q;
  assign LIOI3_X0Y189_OLOGIC_X0Y189_D1 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign LIOI3_X0Y127_OLOGIC_X0Y128_T1 = 1'b1;
  assign RIOI3_X105Y173_OLOGIC_X1Y174_D1 = CLBLM_R_X103Y174_SLICE_X163Y174_AO6;
  assign CLBLM_R_X11Y122_SLICE_X15Y122_C6 = 1'b1;
  assign LIOI3_X0Y189_OLOGIC_X0Y189_T1 = 1'b1;
  assign LIOI3_X0Y127_OLOGIC_X0Y127_D1 = CLBLL_L_X4Y121_SLICE_X4Y121_BQ;
  assign RIOB33_X105Y181_IOB_X1Y182_O = CLBLM_R_X11Y119_SLICE_X14Y119_CO5;
  assign CLBLM_R_X11Y123_SLICE_X14Y123_A4 = CLBLM_L_X10Y122_SLICE_X13Y122_CQ;
  assign RIOB33_X105Y181_IOB_X1Y181_O = CLBLM_R_X11Y119_SLICE_X14Y119_CO6;
  assign RIOI3_X105Y173_OLOGIC_X1Y174_T1 = 1'b1;
  assign CLBLM_R_X11Y123_SLICE_X14Y123_A5 = CLBLM_L_X10Y121_SLICE_X13Y121_BQ;
  assign CLBLM_R_X11Y123_SLICE_X14Y123_A6 = 1'b1;
  assign LIOI3_X0Y127_OLOGIC_X0Y127_T1 = 1'b1;
  assign LIOB33_X0Y137_IOB_X0Y138_O = CLBLM_R_X5Y125_SLICE_X6Y125_AQ;
  assign RIOI3_X105Y173_OLOGIC_X1Y173_D1 = CLBLM_R_X103Y172_SLICE_X163Y172_AO5;
  assign LIOI3_TBYTESRC_X0Y131_OLOGIC_X0Y132_D1 = CLBLM_R_X7Y128_SLICE_X8Y128_AQ;
  assign RIOI3_X105Y173_OLOGIC_X1Y173_T1 = 1'b1;
  assign CLBLM_L_X8Y122_SLICE_X11Y122_A1 = CLBLM_R_X5Y122_SLICE_X7Y122_CQ;
  assign CLBLM_L_X8Y122_SLICE_X11Y122_A2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y122_SLICE_X11Y122_A3 = CLBLM_L_X8Y122_SLICE_X11Y122_AQ;
  assign CLBLM_L_X8Y122_SLICE_X11Y122_A4 = CLBLM_L_X8Y121_SLICE_X11Y121_BQ;
  assign CLBLM_L_X8Y122_SLICE_X11Y122_A5 = CLBLM_L_X10Y123_SLICE_X12Y123_AO6;
  assign CLBLM_L_X8Y122_SLICE_X11Y122_A6 = CLBLM_R_X7Y123_SLICE_X9Y123_CO6;
  assign CLBLM_R_X7Y125_SLICE_X9Y125_C4 = 1'b1;
  assign CLBLM_L_X8Y122_SLICE_X11Y122_AX = CLBLM_L_X8Y115_SLICE_X10Y115_BO6;
  assign LIOB33_X0Y137_IOB_X0Y137_O = CLBLM_R_X5Y124_SLICE_X6Y124_BQ;
  assign CLBLM_L_X8Y122_SLICE_X11Y122_B1 = CLBLM_R_X7Y123_SLICE_X9Y123_CO6;
  assign CLBLM_L_X8Y122_SLICE_X11Y122_B2 = CLBLM_L_X8Y122_SLICE_X11Y122_BQ;
  assign CLBLM_L_X8Y122_SLICE_X11Y122_B3 = CLBLM_R_X5Y123_SLICE_X6Y123_CQ;
  assign CLBLM_L_X8Y122_SLICE_X11Y122_B4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y122_SLICE_X11Y122_B5 = CLBLM_L_X10Y123_SLICE_X12Y123_AO6;
  assign CLBLM_L_X8Y122_SLICE_X11Y122_B6 = CLBLM_L_X8Y121_SLICE_X11Y121_CQ;
  assign CLBLM_R_X7Y125_SLICE_X9Y125_C5 = 1'b1;
  assign CLBLM_R_X7Y125_SLICE_X9Y125_C6 = 1'b1;
  assign LIOI3_TBYTESRC_X0Y131_OLOGIC_X0Y131_D1 = CLBLM_R_X7Y128_SLICE_X8Y128_AO5;
  assign CLBLM_L_X8Y122_SLICE_X11Y122_C1 = CLBLM_R_X5Y120_SLICE_X6Y120_A5Q;
  assign CLBLM_L_X8Y122_SLICE_X11Y122_C2 = CLBLM_R_X7Y124_SLICE_X8Y124_AQ;
  assign CLBLM_L_X8Y122_SLICE_X11Y122_C3 = CLBLM_L_X10Y124_SLICE_X12Y124_AQ;
  assign CLBLM_L_X8Y122_SLICE_X11Y122_C4 = CLBLM_R_X7Y123_SLICE_X9Y123_BO5;
  assign CLBLM_L_X8Y122_SLICE_X11Y122_C5 = CLBLM_L_X8Y119_SLICE_X11Y119_DQ;
  assign CLBLM_L_X8Y122_SLICE_X11Y122_C6 = CLBLM_R_X7Y120_SLICE_X9Y120_A5Q;
  assign RIOI3_TBYTETERM_X105Y163_OLOGIC_X1Y164_T1 = 1'b1;
  assign CLBLM_L_X8Y122_SLICE_X11Y122_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign LIOI3_TBYTESRC_X0Y131_OLOGIC_X0Y131_T1 = 1'b1;
  assign RIOI3_TBYTETERM_X105Y163_OLOGIC_X1Y163_D1 = CLBLM_R_X11Y117_SLICE_X14Y117_DO5;
  assign CLBLM_L_X8Y122_SLICE_X11Y122_D1 = CLBLM_R_X7Y120_SLICE_X9Y120_A5Q;
  assign CLBLL_L_X2Y114_SLICE_X0Y114_A1 = 1'b1;
  assign CLBLL_L_X2Y114_SLICE_X0Y114_A2 = 1'b1;
  assign CLBLL_L_X2Y114_SLICE_X0Y114_A3 = 1'b1;
  assign CLBLM_L_X8Y122_SLICE_X11Y122_D5 = CLBLM_L_X8Y119_SLICE_X11Y119_DQ;
  assign CLBLM_L_X8Y122_SLICE_X11Y122_D6 = CLBLM_R_X7Y124_SLICE_X8Y124_AQ;
  assign CLBLL_L_X2Y114_SLICE_X0Y114_A4 = 1'b1;
  assign CLBLL_L_X2Y114_SLICE_X0Y114_A5 = 1'b1;
  assign CLBLL_L_X2Y114_SLICE_X0Y114_A6 = 1'b1;
  assign CLBLM_L_X8Y122_SLICE_X11Y122_D2 = CLBLM_L_X8Y122_SLICE_X10Y122_AO5;
  assign CLBLM_L_X8Y122_SLICE_X11Y122_D3 = 1'b1;
  assign CLBLL_L_X2Y114_SLICE_X0Y114_B1 = 1'b1;
  assign CLBLL_L_X2Y114_SLICE_X0Y114_B2 = 1'b1;
  assign CLBLM_L_X8Y122_SLICE_X10Y122_A1 = CLBLM_L_X10Y118_SLICE_X12Y118_B5Q;
  assign CLBLM_L_X8Y122_SLICE_X10Y122_A4 = CLBLM_R_X7Y124_SLICE_X8Y124_AQ;
  assign CLBLL_L_X2Y114_SLICE_X0Y114_B3 = 1'b1;
  assign CLBLL_L_X2Y114_SLICE_X0Y114_B4 = 1'b1;
  assign CLBLL_L_X2Y114_SLICE_X0Y114_B5 = 1'b1;
  assign CLBLL_L_X2Y114_SLICE_X0Y114_B6 = 1'b1;
  assign CLBLM_L_X8Y122_SLICE_X10Y122_A6 = 1'b1;
  assign CLBLM_L_X8Y122_SLICE_X10Y122_A2 = CLBLM_R_X7Y120_SLICE_X9Y120_A5Q;
  assign CLBLL_L_X2Y114_SLICE_X0Y114_C1 = 1'b1;
  assign CLBLM_L_X8Y122_SLICE_X10Y122_AX = CLBLM_R_X7Y122_SLICE_X9Y122_BQ;
  assign CLBLL_L_X2Y114_SLICE_X0Y114_C2 = 1'b1;
  assign CLBLM_L_X8Y122_SLICE_X10Y122_B1 = CLBLM_L_X8Y120_SLICE_X10Y120_DQ;
  assign CLBLM_L_X8Y122_SLICE_X10Y122_B2 = RIOB33_X105Y127_IOB_X1Y128_I;
  assign CLBLL_L_X2Y114_SLICE_X0Y114_C3 = 1'b1;
  assign CLBLL_L_X2Y114_SLICE_X0Y114_C4 = 1'b1;
  assign CLBLL_L_X2Y114_SLICE_X0Y114_C5 = 1'b1;
  assign CLBLL_L_X2Y114_SLICE_X0Y114_C6 = 1'b1;
  assign CLBLM_L_X8Y122_SLICE_X10Y122_B4 = RIOB33_X105Y129_IOB_X1Y129_I;
  assign CLBLM_L_X8Y122_SLICE_X10Y122_B5 = RIOB33_X105Y137_IOB_X1Y137_I;
  assign CLBLM_L_X8Y122_SLICE_X10Y122_B6 = 1'b1;
  assign CLBLM_L_X8Y122_SLICE_X10Y122_C1 = CLBLM_L_X8Y122_SLICE_X10Y122_AO6;
  assign CLBLL_L_X2Y114_SLICE_X0Y114_D1 = 1'b1;
  assign CLBLL_L_X2Y114_SLICE_X0Y114_D2 = 1'b1;
  assign CLBLL_L_X2Y114_SLICE_X0Y114_D3 = 1'b1;
  assign CLBLL_L_X2Y114_SLICE_X0Y114_D4 = 1'b1;
  assign CLBLL_L_X2Y114_SLICE_X0Y114_D5 = 1'b1;
  assign CLBLL_L_X2Y114_SLICE_X0Y114_D6 = 1'b1;
  assign CLBLM_L_X8Y122_SLICE_X10Y122_C2 = CLBLM_R_X7Y122_SLICE_X8Y122_CQ;
  assign CLBLM_L_X8Y122_SLICE_X10Y122_C3 = CLBLM_L_X10Y118_SLICE_X12Y118_B5Q;
  assign CLBLM_L_X8Y122_SLICE_X10Y122_C6 = CLBLM_L_X10Y122_SLICE_X12Y122_BQ;
  assign CLBLM_L_X8Y122_SLICE_X10Y122_CE = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y122_SLICE_X10Y122_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X8Y122_SLICE_X10Y122_D1 = CLBLM_R_X5Y120_SLICE_X6Y120_A5Q;
  assign CLBLM_L_X8Y122_SLICE_X10Y122_D2 = CLBLM_R_X5Y111_SLICE_X7Y111_CO5;
  assign CLBLM_L_X8Y122_SLICE_X10Y122_D3 = CLBLM_L_X8Y119_SLICE_X11Y119_DQ;
  assign CLBLM_L_X8Y122_SLICE_X10Y122_D4 = CLBLM_R_X7Y120_SLICE_X9Y120_A5Q;
  assign CLBLM_L_X8Y122_SLICE_X10Y122_D5 = CLBLM_L_X10Y124_SLICE_X12Y124_AQ;
  assign CLBLM_L_X8Y122_SLICE_X10Y122_D6 = CLBLM_R_X7Y124_SLICE_X8Y124_AQ;
  assign CLBLM_R_X7Y125_SLICE_X9Y125_D5 = 1'b1;
  assign CLBLM_R_X7Y125_SLICE_X9Y125_D6 = 1'b1;
  assign CLBLM_L_X8Y122_SLICE_X10Y122_SR = CLBLM_R_X11Y123_SLICE_X14Y123_CO6;
  assign CLBLM_R_X11Y123_SLICE_X14Y123_C5 = 1'b1;
  assign CLBLM_R_X11Y123_SLICE_X14Y123_C6 = RIOB33_X105Y141_IOB_X1Y142_I;
  assign CLBLL_L_X2Y114_SLICE_X1Y114_A1 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLL_L_X2Y114_SLICE_X1Y114_A2 = CLBLM_R_X5Y115_SLICE_X7Y115_AQ;
  assign CLBLL_L_X2Y114_SLICE_X1Y114_A3 = CLBLL_L_X2Y114_SLICE_X1Y114_AQ;
  assign CLBLL_L_X2Y114_SLICE_X1Y114_A4 = CLBLM_R_X3Y114_SLICE_X3Y114_AQ;
  assign CLBLL_L_X2Y114_SLICE_X1Y114_A5 = CLBLL_L_X2Y114_SLICE_X1Y114_CO5;
  assign CLBLL_L_X2Y114_SLICE_X1Y114_A6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLL_L_X2Y114_SLICE_X1Y114_B1 = CLBLL_L_X2Y115_SLICE_X1Y115_BQ;
  assign CLBLL_L_X2Y114_SLICE_X1Y114_B2 = CLBLM_R_X3Y114_SLICE_X2Y114_CQ;
  assign CLBLL_L_X2Y114_SLICE_X1Y114_B3 = CLBLL_L_X2Y114_SLICE_X1Y114_AQ;
  assign CLBLL_L_X2Y114_SLICE_X1Y114_B4 = CLBLM_R_X3Y114_SLICE_X2Y114_AQ;
  assign CLBLL_L_X2Y114_SLICE_X1Y114_B5 = CLBLM_R_X5Y119_SLICE_X7Y119_AO6;
  assign CLBLL_L_X2Y114_SLICE_X1Y114_B6 = 1'b1;
  assign CLBLL_L_X2Y114_SLICE_X1Y114_C1 = CLBLM_R_X3Y114_SLICE_X2Y114_CQ;
  assign CLBLL_L_X2Y114_SLICE_X1Y114_C2 = CLBLM_R_X3Y114_SLICE_X2Y114_AQ;
  assign CLBLL_L_X2Y114_SLICE_X1Y114_C3 = CLBLM_R_X5Y111_SLICE_X7Y111_DO6;
  assign CLBLL_L_X2Y114_SLICE_X1Y114_C4 = CLBLL_L_X2Y115_SLICE_X1Y115_BQ;
  assign CLBLL_L_X2Y114_SLICE_X1Y114_C5 = CLBLL_L_X2Y114_SLICE_X1Y114_AQ;
  assign CLBLL_L_X2Y114_SLICE_X1Y114_C6 = 1'b1;
  assign CLBLL_L_X2Y114_SLICE_X1Y114_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLL_L_X2Y114_SLICE_X1Y114_D1 = CLBLM_R_X3Y114_SLICE_X2Y114_CQ;
  assign CLBLL_L_X2Y114_SLICE_X1Y114_D2 = CLBLM_L_X8Y116_SLICE_X10Y116_AO6;
  assign CLBLL_L_X2Y114_SLICE_X1Y114_D3 = CLBLM_R_X5Y111_SLICE_X7Y111_DO6;
  assign CLBLL_L_X2Y114_SLICE_X1Y114_D4 = CLBLL_L_X2Y115_SLICE_X1Y115_BQ;
  assign CLBLL_L_X2Y114_SLICE_X1Y114_D5 = CLBLL_L_X2Y114_SLICE_X1Y114_AQ;
  assign CLBLL_L_X2Y114_SLICE_X1Y114_D6 = CLBLM_R_X3Y114_SLICE_X2Y114_AQ;
  assign CLBLM_R_X7Y116_SLICE_X9Y116_A1 = CLBLM_R_X7Y116_SLICE_X9Y116_AQ;
  assign CLBLM_R_X7Y116_SLICE_X9Y116_A2 = CLBLM_R_X5Y119_SLICE_X7Y119_AO6;
  assign CLBLM_R_X7Y116_SLICE_X9Y116_A3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y116_SLICE_X9Y116_A4 = CLBLM_R_X7Y119_SLICE_X8Y119_AQ;
  assign CLBLM_R_X7Y116_SLICE_X9Y116_A5 = 1'b1;
  assign CLBLM_R_X7Y116_SLICE_X9Y116_A6 = CLBLM_R_X7Y116_SLICE_X9Y116_CO6;
  assign CLBLM_R_X7Y116_SLICE_X9Y116_B1 = CLBLM_R_X7Y116_SLICE_X9Y116_DO6;
  assign CLBLM_R_X7Y116_SLICE_X9Y116_B2 = CLBLM_R_X7Y117_SLICE_X9Y117_BQ;
  assign CLBLM_R_X7Y116_SLICE_X9Y116_B3 = CLBLM_L_X8Y116_SLICE_X10Y116_BO6;
  assign CLBLM_R_X7Y116_SLICE_X9Y116_B4 = CLBLM_L_X8Y116_SLICE_X11Y116_BQ;
  assign CLBLM_R_X7Y116_SLICE_X9Y116_B5 = CLBLM_R_X7Y116_SLICE_X8Y116_AQ;
  assign CLBLM_R_X7Y116_SLICE_X9Y116_B6 = CLBLM_R_X7Y117_SLICE_X8Y117_BQ;
  assign CLBLM_R_X7Y116_SLICE_X9Y116_C1 = CLBLM_R_X7Y116_SLICE_X8Y116_AQ;
  assign CLBLM_R_X7Y116_SLICE_X9Y116_C2 = CLBLM_L_X10Y114_SLICE_X13Y114_DQ;
  assign CLBLM_R_X7Y116_SLICE_X9Y116_C3 = CLBLL_L_X2Y114_SLICE_X1Y114_BO5;
  assign CLBLM_R_X7Y116_SLICE_X9Y116_C4 = CLBLM_L_X8Y116_SLICE_X11Y116_DQ;
  assign CLBLM_R_X7Y116_SLICE_X9Y116_C5 = 1'b1;
  assign CLBLM_R_X7Y116_SLICE_X9Y116_C6 = CLBLM_R_X7Y116_SLICE_X9Y116_BO6;
  assign LIOI3_X0Y67_ILOGIC_X0Y68_D = LIOB33_X0Y67_IOB_X0Y68_I;
  assign LIOI3_X0Y67_ILOGIC_X0Y67_D = LIOB33_X0Y67_IOB_X0Y67_I;
  assign CLBLM_R_X7Y116_SLICE_X9Y116_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign RIOI3_X105Y103_ILOGIC_X1Y104_D = RIOB33_X105Y103_IOB_X1Y104_I;
  assign CLBLM_R_X7Y116_SLICE_X9Y116_D1 = CLBLM_R_X7Y115_SLICE_X9Y115_AQ;
  assign CLBLM_R_X7Y116_SLICE_X9Y116_D2 = CLBLM_R_X7Y117_SLICE_X9Y117_AQ;
  assign CLBLM_R_X7Y116_SLICE_X9Y116_D3 = 1'b1;
  assign CLBLM_R_X7Y116_SLICE_X9Y116_D4 = CLBLM_R_X7Y116_SLICE_X8Y116_CQ;
  assign CLBLM_R_X7Y116_SLICE_X9Y116_D5 = CLBLM_R_X7Y116_SLICE_X9Y116_AQ;
  assign CLBLM_R_X7Y116_SLICE_X9Y116_D6 = 1'b1;
  assign RIOI3_X105Y111_ILOGIC_X1Y112_D = RIOB33_X105Y111_IOB_X1Y112_I;
  assign RIOI3_X105Y111_ILOGIC_X1Y111_D = RIOB33_X105Y111_IOB_X1Y111_I;
  assign RIOI3_X105Y103_ILOGIC_X1Y103_D = RIOB33_X105Y103_IOB_X1Y103_I;
  assign CLBLM_R_X7Y116_SLICE_X8Y116_A1 = CLBLM_R_X7Y117_SLICE_X8Y117_BQ;
  assign CLBLM_R_X7Y116_SLICE_X8Y116_A2 = CLBLM_L_X8Y116_SLICE_X11Y116_AQ;
  assign CLBLM_R_X7Y116_SLICE_X8Y116_A3 = CLBLM_R_X7Y116_SLICE_X8Y116_AQ;
  assign CLBLM_R_X7Y116_SLICE_X8Y116_A4 = CLBLM_R_X5Y117_SLICE_X7Y117_CO6;
  assign CLBLM_R_X7Y116_SLICE_X8Y116_A5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y116_SLICE_X8Y116_A6 = 1'b1;
  assign CLBLM_R_X7Y116_SLICE_X8Y116_B1 = CLBLM_L_X8Y120_SLICE_X10Y120_A5Q;
  assign CLBLM_R_X7Y116_SLICE_X8Y116_B2 = CLBLL_L_X4Y116_SLICE_X5Y116_DQ;
  assign CLBLM_R_X7Y116_SLICE_X8Y116_B3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y116_SLICE_X8Y116_B4 = CLBLM_R_X7Y115_SLICE_X8Y115_DO5;
  assign CLBLM_R_X7Y116_SLICE_X8Y116_B5 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X7Y116_SLICE_X8Y116_B6 = 1'b1;
  assign CLBLM_R_X7Y125_SLICE_X8Y125_B5 = 1'b1;
  assign CLBLM_R_X7Y125_SLICE_X8Y125_B6 = 1'b1;
  assign CLBLM_R_X11Y122_SLICE_X15Y122_D1 = 1'b1;
  assign CLBLM_R_X7Y116_SLICE_X8Y116_C1 = CLBLM_R_X11Y115_SLICE_X15Y115_CQ;
  assign CLBLM_R_X7Y116_SLICE_X8Y116_C2 = CLBLM_R_X7Y116_SLICE_X8Y116_CQ;
  assign CLBLM_R_X7Y116_SLICE_X8Y116_C3 = 1'b1;
  assign CLBLM_R_X7Y116_SLICE_X8Y116_C4 = CLBLM_R_X5Y116_SLICE_X6Y116_A5Q;
  assign CLBLM_R_X7Y116_SLICE_X8Y116_C5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y116_SLICE_X8Y116_C6 = CLBLM_R_X5Y111_SLICE_X7Y111_DO6;
  assign CLBLM_R_X7Y116_SLICE_X8Y116_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X7Y116_SLICE_X8Y116_D1 = CLBLM_R_X7Y109_SLICE_X8Y109_AQ;
  assign CLBLM_R_X7Y116_SLICE_X8Y116_D2 = CLBLL_L_X4Y120_SLICE_X4Y120_AO6;
  assign CLBLM_R_X7Y116_SLICE_X8Y116_D3 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X7Y116_SLICE_X8Y116_D4 = CLBLM_R_X5Y116_SLICE_X7Y116_CQ;
  assign CLBLM_R_X7Y116_SLICE_X8Y116_D5 = 1'b1;
  assign CLBLM_R_X7Y116_SLICE_X8Y116_D6 = CLBLM_R_X7Y115_SLICE_X8Y115_DO5;
  assign CLBLM_R_X11Y122_SLICE_X15Y122_D2 = 1'b1;
  assign LIOI3_X0Y185_OLOGIC_X0Y186_D1 = RIOB33_X105Y143_IOB_X1Y143_I;
  assign RIOB33_X105Y183_IOB_X1Y184_O = CLBLM_R_X11Y117_SLICE_X14Y117_DO5;
  assign RIOB33_X105Y183_IOB_X1Y183_O = CLBLM_R_X11Y117_SLICE_X14Y117_DO6;
  assign CLBLM_R_X7Y125_SLICE_X8Y125_C4 = 1'b1;
  assign CLBLM_R_X7Y125_SLICE_X8Y125_C5 = 1'b1;
  assign CLBLM_R_X11Y122_SLICE_X15Y122_D3 = 1'b1;
  assign CLBLM_R_X11Y113_SLICE_X15Y113_A4 = CLBLM_L_X10Y112_SLICE_X13Y112_BQ;
  assign CLBLM_R_X7Y125_SLICE_X8Y125_C6 = 1'b1;
  assign LIOB33_X0Y117_IOB_X0Y118_O = CLBLL_L_X4Y116_SLICE_X4Y116_CQ;
  assign CLBLM_R_X11Y113_SLICE_X15Y113_A5 = CLBLM_R_X11Y119_SLICE_X15Y119_BQ;
  assign LIOB33_X0Y117_IOB_X0Y117_O = CLBLL_L_X4Y119_SLICE_X4Y119_BQ;
  assign CLBLM_L_X8Y118_SLICE_X11Y118_D6 = 1'b1;
  assign CLBLM_R_X11Y113_SLICE_X15Y113_A6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X11Y122_SLICE_X15Y122_D4 = 1'b1;
  assign LIOI3_X0Y185_OLOGIC_X0Y186_T1 = 1'b1;
  assign CLBLM_L_X8Y123_SLICE_X11Y123_A1 = CLBLM_R_X11Y120_SLICE_X15Y120_AQ;
  assign CLBLM_L_X8Y123_SLICE_X11Y123_A2 = 1'b1;
  assign CLBLM_L_X8Y123_SLICE_X11Y123_A3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y123_SLICE_X11Y123_A4 = CLBLL_L_X4Y123_SLICE_X4Y123_AQ;
  assign CLBLM_L_X8Y123_SLICE_X11Y123_A5 = RIOB33_X105Y125_IOB_X1Y126_I;
  assign CLBLM_L_X8Y123_SLICE_X11Y123_A6 = 1'b1;
  assign CLBLM_R_X11Y122_SLICE_X15Y122_D5 = 1'b1;
  assign CLBLM_L_X8Y123_SLICE_X11Y123_B1 = 1'b1;
  assign CLBLM_L_X8Y123_SLICE_X11Y123_B2 = 1'b1;
  assign CLBLM_L_X8Y123_SLICE_X11Y123_B3 = 1'b1;
  assign CLBLM_L_X8Y123_SLICE_X11Y123_B4 = 1'b1;
  assign CLBLM_L_X8Y123_SLICE_X11Y123_B5 = 1'b1;
  assign CLBLM_L_X8Y123_SLICE_X11Y123_B6 = 1'b1;
  assign CLBLM_L_X8Y123_SLICE_X11Y123_C1 = 1'b1;
  assign CLBLM_L_X8Y123_SLICE_X11Y123_C2 = 1'b1;
  assign CLBLM_L_X8Y123_SLICE_X11Y123_C3 = 1'b1;
  assign CLBLM_L_X8Y123_SLICE_X11Y123_C4 = 1'b1;
  assign CLBLM_L_X8Y123_SLICE_X11Y123_C5 = 1'b1;
  assign CLBLM_L_X8Y123_SLICE_X11Y123_C6 = 1'b1;
  assign CLBLM_L_X8Y123_SLICE_X11Y123_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLL_L_X2Y115_SLICE_X0Y115_A1 = 1'b1;
  assign CLBLL_L_X2Y115_SLICE_X0Y115_A2 = 1'b1;
  assign CLBLL_L_X2Y115_SLICE_X0Y115_A3 = 1'b1;
  assign CLBLL_L_X2Y115_SLICE_X0Y115_A4 = 1'b1;
  assign CLBLL_L_X2Y115_SLICE_X0Y115_A5 = 1'b1;
  assign CLBLL_L_X2Y115_SLICE_X0Y115_A6 = 1'b1;
  assign CLBLM_L_X8Y123_SLICE_X11Y123_D1 = 1'b1;
  assign CLBLM_L_X8Y123_SLICE_X11Y123_D2 = 1'b1;
  assign CLBLL_L_X2Y115_SLICE_X0Y115_B1 = 1'b1;
  assign CLBLL_L_X2Y115_SLICE_X0Y115_B2 = 1'b1;
  assign CLBLL_L_X2Y115_SLICE_X0Y115_B3 = 1'b1;
  assign CLBLL_L_X2Y115_SLICE_X0Y115_B4 = 1'b1;
  assign CLBLL_L_X2Y115_SLICE_X0Y115_B5 = 1'b1;
  assign CLBLL_L_X2Y115_SLICE_X0Y115_B6 = 1'b1;
  assign CLBLM_L_X8Y123_SLICE_X11Y123_D4 = 1'b1;
  assign CLBLM_L_X8Y123_SLICE_X10Y123_A1 = CLBLM_L_X8Y123_SLICE_X10Y123_B5Q;
  assign CLBLM_L_X8Y123_SLICE_X10Y123_A2 = CLBLM_L_X8Y123_SLICE_X10Y123_BQ;
  assign CLBLL_L_X2Y115_SLICE_X0Y115_C1 = 1'b1;
  assign CLBLL_L_X2Y115_SLICE_X0Y115_C2 = 1'b1;
  assign CLBLL_L_X2Y115_SLICE_X0Y115_C3 = 1'b1;
  assign CLBLL_L_X2Y115_SLICE_X0Y115_C4 = 1'b1;
  assign CLBLL_L_X2Y115_SLICE_X0Y115_C5 = 1'b1;
  assign CLBLL_L_X2Y115_SLICE_X0Y115_C6 = 1'b1;
  assign CLBLM_L_X8Y123_SLICE_X10Y123_A3 = CLBLM_R_X7Y118_SLICE_X9Y118_DO6;
  assign CLBLM_L_X8Y123_SLICE_X10Y123_A4 = 1'b1;
  assign CLBLM_L_X8Y123_SLICE_X10Y123_A5 = CLBLM_L_X8Y123_SLICE_X10Y123_A5Q;
  assign CLBLM_L_X8Y123_SLICE_X10Y123_A6 = 1'b1;
  assign CLBLM_L_X8Y123_SLICE_X10Y123_B1 = CLBLM_L_X8Y123_SLICE_X10Y123_B5Q;
  assign CLBLM_L_X8Y123_SLICE_X10Y123_B2 = CLBLM_L_X8Y123_SLICE_X10Y123_BQ;
  assign CLBLM_L_X8Y123_SLICE_X10Y123_B3 = CLBLM_R_X7Y118_SLICE_X9Y118_DO6;
  assign CLBLL_L_X2Y115_SLICE_X0Y115_D1 = 1'b1;
  assign CLBLL_L_X2Y115_SLICE_X0Y115_D2 = 1'b1;
  assign CLBLL_L_X2Y115_SLICE_X0Y115_D3 = 1'b1;
  assign CLBLL_L_X2Y115_SLICE_X0Y115_D4 = 1'b1;
  assign CLBLL_L_X2Y115_SLICE_X0Y115_D5 = 1'b1;
  assign CLBLL_L_X2Y115_SLICE_X0Y115_D6 = 1'b1;
  assign CLBLM_L_X8Y123_SLICE_X10Y123_B5 = CLBLM_L_X8Y123_SLICE_X10Y123_A5Q;
  assign CLBLM_L_X8Y123_SLICE_X10Y123_B6 = 1'b1;
  assign CLBLM_L_X8Y123_SLICE_X10Y123_C1 = 1'b1;
  assign CLBLM_L_X8Y123_SLICE_X10Y123_C2 = 1'b1;
  assign CLBLM_L_X8Y123_SLICE_X10Y123_C3 = 1'b1;
  assign CLBLM_L_X8Y123_SLICE_X10Y123_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X8Y123_SLICE_X10Y123_C4 = 1'b1;
  assign CLBLM_L_X8Y123_SLICE_X10Y123_C5 = 1'b1;
  assign CLBLM_L_X8Y123_SLICE_X10Y123_C6 = 1'b1;
  assign CLBLM_L_X8Y123_SLICE_X10Y123_D1 = 1'b1;
  assign CLBLM_L_X8Y123_SLICE_X10Y123_D2 = 1'b1;
  assign CLBLM_L_X8Y123_SLICE_X10Y123_D3 = 1'b1;
  assign CLBLM_L_X8Y123_SLICE_X10Y123_D4 = 1'b1;
  assign CLBLM_L_X8Y123_SLICE_X10Y123_D5 = 1'b1;
  assign CLBLM_L_X8Y123_SLICE_X10Y123_D6 = 1'b1;
  assign CLBLL_L_X2Y115_SLICE_X1Y115_A1 = CLBLM_R_X5Y113_SLICE_X6Y113_BQ;
  assign CLBLL_L_X2Y115_SLICE_X1Y115_A2 = CLBLM_L_X8Y112_SLICE_X10Y112_CQ;
  assign CLBLL_L_X2Y115_SLICE_X1Y115_A3 = CLBLL_L_X2Y115_SLICE_X1Y115_AQ;
  assign CLBLL_L_X2Y115_SLICE_X1Y115_A4 = CLBLM_R_X3Y113_SLICE_X2Y113_AQ;
  assign CLBLL_L_X2Y115_SLICE_X1Y115_A5 = CLBLL_L_X2Y112_SLICE_X1Y112_BQ;
  assign CLBLL_L_X2Y115_SLICE_X1Y115_A6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y119_SLICE_X10Y119_B4 = CLBLM_L_X8Y115_SLICE_X10Y115_AQ;
  assign CLBLM_L_X8Y119_SLICE_X10Y119_B5 = CLBLM_L_X8Y120_SLICE_X10Y120_AQ;
  assign LIOI3_X0Y65_ILOGIC_X0Y66_D = LIOB33_X0Y65_IOB_X0Y66_I;
  assign CLBLL_L_X2Y115_SLICE_X1Y115_B1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLL_L_X2Y115_SLICE_X1Y115_B2 = CLBLL_L_X2Y115_SLICE_X1Y115_BQ;
  assign CLBLL_L_X2Y115_SLICE_X1Y115_B3 = CLBLM_R_X3Y123_SLICE_X3Y123_AQ;
  assign CLBLL_L_X2Y115_SLICE_X1Y115_B4 = CLBLM_R_X5Y115_SLICE_X7Y115_AQ;
  assign CLBLL_L_X2Y115_SLICE_X1Y115_B5 = CLBLL_L_X2Y114_SLICE_X1Y114_CO6;
  assign CLBLL_L_X2Y115_SLICE_X1Y115_B6 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X8Y119_SLICE_X10Y119_B6 = 1'b1;
  assign LIOI3_TBYTETERM_X0Y187_OLOGIC_X0Y188_T1 = 1'b1;
  assign LIOI3_X0Y185_OLOGIC_X0Y185_T1 = 1'b1;
  assign CLBLL_L_X2Y115_SLICE_X1Y115_C1 = 1'b1;
  assign CLBLL_L_X2Y115_SLICE_X1Y115_C2 = 1'b1;
  assign CLBLL_L_X2Y115_SLICE_X1Y115_C3 = 1'b1;
  assign CLBLL_L_X2Y115_SLICE_X1Y115_C4 = 1'b1;
  assign CLBLL_L_X2Y115_SLICE_X1Y115_C5 = 1'b1;
  assign CLBLL_L_X2Y115_SLICE_X1Y115_C6 = 1'b1;
  assign LIOI3_X0Y65_ILOGIC_X0Y65_D = LIOB33_X0Y65_IOB_X0Y65_I;
  assign CLBLL_L_X2Y115_SLICE_X1Y115_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLL_L_X2Y115_SLICE_X1Y115_D1 = 1'b1;
  assign CLBLL_L_X2Y115_SLICE_X1Y115_D2 = 1'b1;
  assign CLBLL_L_X2Y115_SLICE_X1Y115_D3 = 1'b1;
  assign CLBLL_L_X2Y115_SLICE_X1Y115_D4 = 1'b1;
  assign CLBLL_L_X2Y115_SLICE_X1Y115_D5 = 1'b1;
  assign CLBLL_L_X2Y115_SLICE_X1Y115_D6 = 1'b1;
  assign CLBLM_R_X7Y117_SLICE_X9Y117_A1 = CLBLM_R_X5Y117_SLICE_X7Y117_CO6;
  assign CLBLM_R_X7Y117_SLICE_X9Y117_A2 = 1'b1;
  assign CLBLM_R_X7Y117_SLICE_X9Y117_A3 = CLBLM_R_X7Y117_SLICE_X9Y117_AQ;
  assign CLBLM_R_X7Y117_SLICE_X9Y117_A4 = CLBLM_R_X7Y116_SLICE_X8Y116_CQ;
  assign CLBLM_R_X7Y117_SLICE_X9Y117_A5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y117_SLICE_X9Y117_A6 = CLBLM_L_X10Y122_SLICE_X13Y122_A5Q;
  assign CLBLM_R_X7Y117_SLICE_X9Y117_B1 = CLBLM_R_X5Y121_SLICE_X7Y121_A5Q;
  assign CLBLM_R_X7Y117_SLICE_X9Y117_B2 = CLBLM_R_X7Y117_SLICE_X9Y117_BQ;
  assign CLBLM_R_X7Y117_SLICE_X9Y117_B3 = CLBLM_R_X7Y117_SLICE_X9Y117_AQ;
  assign CLBLM_L_X8Y118_SLICE_X10Y118_A1 = 1'b1;
  assign CLBLM_R_X7Y117_SLICE_X9Y117_B4 = 1'b1;
  assign CLBLM_R_X7Y117_SLICE_X9Y117_B5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y117_SLICE_X9Y117_B6 = CLBLM_R_X5Y117_SLICE_X7Y117_CO6;
  assign CLBLM_R_X7Y117_SLICE_X9Y117_C1 = CLBLM_R_X3Y115_SLICE_X2Y115_BQ;
  assign CLBLM_R_X7Y117_SLICE_X9Y117_C2 = CLBLM_R_X7Y117_SLICE_X9Y117_CQ;
  assign CLBLM_R_X7Y117_SLICE_X9Y117_C3 = CLBLM_L_X8Y112_SLICE_X10Y112_CQ;
  assign CLBLM_R_X7Y117_SLICE_X9Y117_C4 = CLBLM_R_X11Y117_SLICE_X15Y117_AQ;
  assign CLBLM_R_X7Y117_SLICE_X9Y117_C5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y117_SLICE_X9Y117_C6 = CLBLL_L_X2Y112_SLICE_X1Y112_BQ;
  assign CLBLM_R_X7Y117_SLICE_X9Y117_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign LIOI3_TBYTETERM_X0Y187_OLOGIC_X0Y187_D1 = RIOB33_X105Y143_IOB_X1Y144_I;
  assign CLBLM_R_X7Y117_SLICE_X9Y117_D1 = CLBLM_R_X5Y115_SLICE_X6Y115_CO5;
  assign CLBLM_R_X7Y117_SLICE_X9Y117_D2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y117_SLICE_X9Y117_D3 = CLBLM_R_X7Y117_SLICE_X9Y117_DQ;
  assign CLBLM_L_X8Y118_SLICE_X10Y118_A2 = CLBLM_R_X5Y110_SLICE_X7Y110_CQ;
  assign CLBLM_R_X7Y117_SLICE_X9Y117_D4 = 1'b1;
  assign CLBLM_R_X7Y117_SLICE_X9Y117_D5 = CLBLL_L_X2Y113_SLICE_X1Y113_BQ;
  assign CLBLM_R_X7Y117_SLICE_X9Y117_D6 = CLBLM_L_X8Y115_SLICE_X11Y115_AQ;
  assign CLBLM_R_X7Y117_SLICE_X8Y117_A1 = CLBLM_R_X3Y118_SLICE_X2Y118_AQ;
  assign CLBLM_R_X7Y117_SLICE_X8Y117_A2 = CLBLM_R_X5Y112_SLICE_X7Y112_BO6;
  assign CLBLM_R_X7Y117_SLICE_X8Y117_A3 = CLBLM_R_X7Y117_SLICE_X8Y117_AQ;
  assign CLBLM_R_X7Y117_SLICE_X8Y117_A4 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_R_X7Y117_SLICE_X8Y117_A5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y117_SLICE_X8Y117_A6 = CLBLL_L_X4Y117_SLICE_X5Y117_BQ;
  assign CLBLM_R_X7Y117_SLICE_X8Y117_AX = CLBLM_R_X7Y117_SLICE_X8Y117_DO6;
  assign CLBLM_R_X7Y117_SLICE_X8Y117_B1 = CLBLM_R_X5Y117_SLICE_X6Y117_DQ;
  assign CLBLM_R_X7Y117_SLICE_X8Y117_B2 = CLBLM_R_X7Y117_SLICE_X8Y117_BQ;
  assign CLBLM_R_X7Y117_SLICE_X8Y117_B3 = CLBLM_R_X5Y117_SLICE_X7Y117_CO6;
  assign CLBLM_R_X7Y117_SLICE_X8Y117_B4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y117_SLICE_X8Y117_B5 = CLBLM_R_X7Y115_SLICE_X9Y115_AQ;
  assign CLBLM_R_X7Y117_SLICE_X8Y117_B6 = 1'b1;
  assign CLBLM_R_X7Y117_SLICE_X8Y117_C1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y117_SLICE_X8Y117_C2 = 1'b1;
  assign CLBLM_R_X7Y117_SLICE_X8Y117_C3 = CLBLL_L_X2Y113_SLICE_X1Y113_BQ;
  assign CLBLM_R_X7Y117_SLICE_X8Y117_C4 = CLBLM_R_X7Y114_SLICE_X8Y114_DO6;
  assign CLBLM_R_X7Y117_SLICE_X8Y117_C5 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X7Y117_SLICE_X8Y117_C6 = CLBLM_L_X8Y119_SLICE_X11Y119_AQ;
  assign RIOB33_X105Y185_IOB_X1Y186_O = CLBLM_L_X12Y115_SLICE_X16Y115_BQ;
  assign CLBLM_R_X7Y117_SLICE_X8Y117_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign RIOB33_X105Y185_IOB_X1Y185_O = CLBLM_R_X7Y119_SLICE_X9Y119_DO5;
  assign CLBLM_L_X8Y119_SLICE_X10Y119_D2 = CLBLM_L_X8Y114_SLICE_X10Y114_C5Q;
  assign CLBLM_R_X7Y117_SLICE_X8Y117_D1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y119_SLICE_X10Y119_D3 = RIOB33_X105Y121_IOB_X1Y121_I;
  assign CLBLM_R_X7Y117_SLICE_X8Y117_D2 = CLBLM_L_X8Y115_SLICE_X10Y115_CQ;
  assign CLBLM_R_X7Y117_SLICE_X8Y117_D3 = CLBLM_R_X7Y117_SLICE_X8Y117_AQ;
  assign CLBLM_R_X7Y117_SLICE_X8Y117_D4 = CLBLM_L_X8Y118_SLICE_X10Y118_D5Q;
  assign CLBLM_R_X7Y117_SLICE_X8Y117_D5 = RIOB33_X105Y121_IOB_X1Y121_I;
  assign CLBLM_R_X7Y117_SLICE_X8Y117_D6 = 1'b1;
  assign LIOI3_TBYTETERM_X0Y187_OLOGIC_X0Y187_T1 = 1'b1;
  assign CLBLM_L_X8Y118_SLICE_X10Y118_A5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign RIOI3_SING_X105Y149_ILOGIC_X1Y149_D = RIOB33_SING_X105Y149_IOB_X1Y149_I;
  assign CLBLL_L_X2Y116_SLICE_X0Y116_A1 = 1'b1;
  assign CLBLL_L_X2Y116_SLICE_X0Y116_A2 = 1'b1;
  assign CLBLL_L_X2Y116_SLICE_X0Y116_A3 = 1'b1;
  assign CLBLL_L_X2Y116_SLICE_X0Y116_A4 = 1'b1;
  assign CLBLL_L_X2Y116_SLICE_X0Y116_A5 = 1'b1;
  assign CLBLL_L_X2Y116_SLICE_X0Y116_A6 = 1'b1;
  assign CLBLL_L_X2Y116_SLICE_X0Y116_B1 = 1'b1;
  assign CLBLL_L_X2Y116_SLICE_X0Y116_B2 = 1'b1;
  assign CLBLL_L_X2Y116_SLICE_X0Y116_B3 = 1'b1;
  assign CLBLL_L_X2Y116_SLICE_X0Y116_B4 = 1'b1;
  assign CLBLL_L_X2Y116_SLICE_X0Y116_B5 = 1'b1;
  assign CLBLL_L_X2Y116_SLICE_X0Y116_B6 = 1'b1;
  assign CLBLM_R_X7Y128_SLICE_X8Y128_B6 = 1'b1;
  assign LIOI3_X0Y191_OLOGIC_X0Y192_D1 = LIOB33_X0Y51_IOB_X0Y52_I;
  assign CLBLL_L_X2Y116_SLICE_X0Y116_C1 = 1'b1;
  assign CLBLL_L_X2Y116_SLICE_X0Y116_C2 = 1'b1;
  assign CLBLL_L_X2Y116_SLICE_X0Y116_C3 = 1'b1;
  assign CLBLL_L_X2Y116_SLICE_X0Y116_C4 = 1'b1;
  assign CLBLL_L_X2Y116_SLICE_X0Y116_C5 = 1'b1;
  assign CLBLL_L_X2Y116_SLICE_X0Y116_C6 = 1'b1;
  assign LIOI3_X0Y191_OLOGIC_X0Y192_T1 = 1'b1;
  assign LIOI3_X0Y129_OLOGIC_X0Y130_D1 = CLBLL_L_X52Y126_SLICE_X78Y126_AO6;
  assign CLBLL_L_X2Y116_SLICE_X0Y116_D1 = 1'b1;
  assign CLBLL_L_X2Y116_SLICE_X0Y116_D2 = 1'b1;
  assign CLBLL_L_X2Y116_SLICE_X0Y116_D3 = 1'b1;
  assign CLBLL_L_X2Y116_SLICE_X0Y116_D4 = 1'b1;
  assign CLBLL_L_X2Y116_SLICE_X0Y116_D5 = 1'b1;
  assign CLBLL_L_X2Y116_SLICE_X0Y116_D6 = 1'b1;
  assign LIOI3_X0Y191_OLOGIC_X0Y191_D1 = RIOB33_X105Y147_IOB_X1Y148_I;
  assign LIOI3_X0Y129_OLOGIC_X0Y130_T1 = 1'b1;
  assign RIOI3_X105Y175_OLOGIC_X1Y176_D1 = CLBLM_R_X103Y174_SLICE_X163Y174_AO5;
  assign CLBLM_R_X7Y124_SLICE_X9Y124_C4 = 1'b1;
  assign LIOI3_X0Y191_OLOGIC_X0Y191_T1 = 1'b1;
  assign LIOI3_X0Y129_OLOGIC_X0Y129_D1 = CLBLM_R_X3Y115_SLICE_X3Y115_CQ;
  assign RIOI3_X105Y175_OLOGIC_X1Y176_T1 = 1'b1;
  assign CLBLL_L_X2Y116_SLICE_X1Y116_A1 = CLBLL_L_X2Y115_SLICE_X1Y115_BQ;
  assign CLBLL_L_X2Y116_SLICE_X1Y116_A2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLL_L_X2Y116_SLICE_X1Y116_A3 = CLBLL_L_X2Y116_SLICE_X1Y116_AQ;
  assign CLBLL_L_X2Y116_SLICE_X1Y116_A4 = CLBLM_R_X3Y113_SLICE_X2Y113_BQ;
  assign CLBLL_L_X2Y116_SLICE_X1Y116_A5 = CLBLL_L_X2Y112_SLICE_X1Y112_BQ;
  assign CLBLL_L_X2Y116_SLICE_X1Y116_A6 = CLBLM_L_X8Y112_SLICE_X10Y112_CQ;
  assign LIOI3_X0Y129_OLOGIC_X0Y129_T1 = 1'b1;
  assign RIOI3_X105Y175_OLOGIC_X1Y175_D1 = CLBLM_L_X10Y128_SLICE_X13Y128_AO6;
  assign CLBLM_R_X7Y124_SLICE_X9Y124_C5 = 1'b1;
  assign CLBLL_L_X2Y116_SLICE_X1Y116_B1 = 1'b1;
  assign CLBLL_L_X2Y116_SLICE_X1Y116_B2 = 1'b1;
  assign CLBLL_L_X2Y116_SLICE_X1Y116_B3 = 1'b1;
  assign CLBLL_L_X2Y116_SLICE_X1Y116_B4 = 1'b1;
  assign CLBLL_L_X2Y116_SLICE_X1Y116_B5 = 1'b1;
  assign CLBLL_L_X2Y116_SLICE_X1Y116_B6 = 1'b1;
  assign LIOI3_TBYTESRC_X0Y143_OLOGIC_X0Y144_D1 = LIOB33_X0Y57_IOB_X0Y57_I;
  assign LIOI3_X0Y151_OLOGIC_X0Y152_D1 = LIOB33_X0Y65_IOB_X0Y66_I;
  assign RIOI3_X105Y175_OLOGIC_X1Y175_T1 = 1'b1;
  assign CLBLL_L_X2Y116_SLICE_X1Y116_C1 = 1'b1;
  assign CLBLL_L_X2Y116_SLICE_X1Y116_C2 = 1'b1;
  assign CLBLL_L_X2Y116_SLICE_X1Y116_C3 = 1'b1;
  assign CLBLL_L_X2Y116_SLICE_X1Y116_C4 = 1'b1;
  assign CLBLL_L_X2Y116_SLICE_X1Y116_C5 = 1'b1;
  assign CLBLL_L_X2Y116_SLICE_X1Y116_C6 = 1'b1;
  assign LIOI3_TBYTESRC_X0Y143_OLOGIC_X0Y144_T1 = 1'b1;
  assign RIOI3_TBYTETERM_X105Y187_OLOGIC_X1Y188_D1 = CLBLM_R_X11Y122_SLICE_X14Y122_AQ;
  assign CLBLL_L_X2Y116_SLICE_X1Y116_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X11Y128_SLICE_X15Y128_A1 = CLBLM_L_X8Y121_SLICE_X11Y121_CQ;
  assign CLBLM_R_X11Y128_SLICE_X15Y128_A2 = RIOB33_X105Y141_IOB_X1Y142_I;
  assign CLBLM_R_X11Y128_SLICE_X15Y128_A3 = CLBLM_R_X11Y128_SLICE_X15Y128_AQ;
  assign CLBLM_R_X7Y124_SLICE_X9Y124_C6 = 1'b1;
  assign CLBLL_L_X2Y116_SLICE_X1Y116_D1 = 1'b1;
  assign CLBLL_L_X2Y116_SLICE_X1Y116_D2 = 1'b1;
  assign CLBLL_L_X2Y116_SLICE_X1Y116_D3 = 1'b1;
  assign CLBLL_L_X2Y116_SLICE_X1Y116_D4 = 1'b1;
  assign CLBLL_L_X2Y116_SLICE_X1Y116_D5 = 1'b1;
  assign CLBLL_L_X2Y116_SLICE_X1Y116_D6 = 1'b1;
  assign CLBLM_R_X11Y128_SLICE_X15Y128_A4 = 1'b1;
  assign CLBLM_R_X11Y128_SLICE_X15Y128_A5 = CLBLM_R_X7Y128_SLICE_X8Y128_AQ;
  assign CLBLM_R_X11Y128_SLICE_X15Y128_A6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X11Y128_SLICE_X15Y128_B1 = 1'b1;
  assign CLBLM_R_X11Y128_SLICE_X15Y128_B2 = 1'b1;
  assign CLBLM_R_X11Y128_SLICE_X15Y128_B3 = 1'b1;
  assign CLBLM_R_X11Y128_SLICE_X15Y128_B4 = 1'b1;
  assign CLBLM_R_X7Y118_SLICE_X9Y118_A1 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X7Y118_SLICE_X9Y118_A2 = CLBLM_R_X7Y113_SLICE_X9Y113_A5Q;
  assign CLBLM_R_X7Y118_SLICE_X9Y118_A3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y118_SLICE_X9Y118_A4 = CLBLM_L_X10Y127_SLICE_X12Y127_AQ;
  assign CLBLM_R_X7Y118_SLICE_X9Y118_A5 = CLBLM_R_X7Y115_SLICE_X9Y115_C5Q;
  assign CLBLM_R_X7Y118_SLICE_X9Y118_A6 = CLBLM_R_X3Y115_SLICE_X3Y115_CQ;
  assign CLBLM_R_X11Y128_SLICE_X15Y128_C1 = 1'b1;
  assign CLBLM_R_X11Y128_SLICE_X15Y128_C2 = 1'b1;
  assign CLBLM_R_X11Y128_SLICE_X15Y128_C3 = 1'b1;
  assign CLBLM_R_X7Y118_SLICE_X9Y118_B1 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X7Y118_SLICE_X9Y118_B2 = CLBLM_L_X10Y118_SLICE_X12Y118_CO6;
  assign CLBLM_R_X7Y118_SLICE_X9Y118_B3 = 1'b1;
  assign CLBLM_R_X7Y118_SLICE_X9Y118_B4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y118_SLICE_X9Y118_B5 = CLBLM_R_X7Y117_SLICE_X9Y117_AQ;
  assign CLBLM_R_X7Y118_SLICE_X9Y118_B6 = CLBLM_R_X7Y118_SLICE_X9Y118_BQ;
  assign CLBLM_R_X11Y128_SLICE_X15Y128_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X11Y128_SLICE_X15Y128_D1 = 1'b1;
  assign CLBLM_R_X7Y118_SLICE_X9Y118_C1 = 1'b1;
  assign CLBLM_R_X7Y118_SLICE_X9Y118_C2 = CLBLM_L_X8Y114_SLICE_X11Y114_BQ;
  assign CLBLM_R_X7Y118_SLICE_X9Y118_C3 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X7Y118_SLICE_X9Y118_C4 = CLBLM_R_X7Y118_SLICE_X9Y118_BQ;
  assign CLBLM_R_X7Y118_SLICE_X9Y118_C5 = 1'b1;
  assign CLBLM_R_X7Y118_SLICE_X9Y118_C6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X11Y128_SLICE_X15Y128_D3 = 1'b1;
  assign CLBLM_R_X11Y128_SLICE_X15Y128_D4 = 1'b1;
  assign CLBLM_R_X7Y118_SLICE_X9Y118_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X11Y128_SLICE_X14Y128_A1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X11Y128_SLICE_X14Y128_A2 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X11Y128_SLICE_X14Y128_A3 = RIOB33_X105Y143_IOB_X1Y143_I;
  assign CLBLM_R_X11Y128_SLICE_X14Y128_A4 = CLBLM_L_X8Y119_SLICE_X11Y119_CQ;
  assign CLBLM_R_X11Y128_SLICE_X14Y128_A5 = CLBLM_R_X11Y120_SLICE_X14Y120_AQ;
  assign CLBLM_R_X7Y118_SLICE_X9Y118_D1 = CLBLM_R_X7Y116_SLICE_X9Y116_BO6;
  assign CLBLM_R_X7Y118_SLICE_X9Y118_D2 = CLBLL_L_X4Y120_SLICE_X4Y120_BO6;
  assign CLBLM_R_X7Y118_SLICE_X9Y118_D3 = CLBLL_L_X4Y121_SLICE_X4Y121_CO6;
  assign CLBLM_R_X7Y118_SLICE_X9Y118_D4 = CLBLM_L_X10Y118_SLICE_X13Y118_DO6;
  assign CLBLM_R_X7Y118_SLICE_X9Y118_D5 = CLBLM_L_X8Y116_SLICE_X11Y116_DQ;
  assign CLBLM_R_X7Y118_SLICE_X9Y118_D6 = CLBLM_R_X5Y110_SLICE_X7Y110_DO5;
  assign CLBLM_R_X11Y128_SLICE_X14Y128_A6 = 1'b1;
  assign CLBLM_R_X11Y128_SLICE_X14Y128_B1 = 1'b1;
  assign CLBLM_R_X11Y128_SLICE_X14Y128_B2 = 1'b1;
  assign CLBLM_R_X11Y128_SLICE_X14Y128_B3 = 1'b1;
  assign CLBLM_R_X11Y128_SLICE_X14Y128_B4 = 1'b1;
  assign CLBLM_R_X7Y118_SLICE_X8Y118_A1 = 1'b1;
  assign CLBLM_R_X7Y118_SLICE_X8Y118_A2 = CLBLL_L_X4Y114_SLICE_X4Y114_BQ;
  assign CLBLM_R_X7Y118_SLICE_X8Y118_A3 = CLBLM_R_X7Y118_SLICE_X8Y118_AQ;
  assign CLBLM_R_X7Y118_SLICE_X8Y118_A4 = CLBLM_L_X8Y119_SLICE_X11Y119_BQ;
  assign CLBLM_R_X7Y118_SLICE_X8Y118_A5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y118_SLICE_X8Y118_A6 = CLBLM_R_X11Y121_SLICE_X14Y121_CO6;
  assign CLBLM_R_X11Y128_SLICE_X14Y128_C1 = 1'b1;
  assign CLBLM_R_X11Y128_SLICE_X14Y128_C2 = 1'b1;
  assign CLBLM_R_X7Y124_SLICE_X9Y124_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X7Y118_SLICE_X8Y118_B1 = CLBLM_R_X5Y116_SLICE_X6Y116_DQ;
  assign CLBLM_R_X7Y118_SLICE_X8Y118_B2 = CLBLM_R_X7Y118_SLICE_X8Y118_BQ;
  assign CLBLM_R_X7Y118_SLICE_X8Y118_B3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y118_SLICE_X8Y118_B4 = 1'b1;
  assign CLBLM_R_X7Y118_SLICE_X8Y118_B5 = CLBLM_R_X5Y115_SLICE_X6Y115_CO5;
  assign CLBLM_R_X7Y118_SLICE_X8Y118_B6 = CLBLM_R_X7Y119_SLICE_X9Y119_AQ;
  assign CLBLM_R_X11Y128_SLICE_X14Y128_D1 = 1'b1;
  assign CLBLM_R_X11Y128_SLICE_X14Y128_D2 = 1'b1;
  assign CLBLM_R_X11Y128_SLICE_X14Y128_D3 = 1'b1;
  assign CLBLM_R_X7Y118_SLICE_X8Y118_C1 = CLBLM_R_X5Y115_SLICE_X6Y115_CO5;
  assign CLBLM_R_X7Y118_SLICE_X8Y118_C2 = CLBLM_R_X7Y118_SLICE_X8Y118_CQ;
  assign CLBLM_R_X7Y118_SLICE_X8Y118_C3 = CLBLM_R_X5Y116_SLICE_X6Y116_DQ;
  assign CLBLM_R_X7Y118_SLICE_X8Y118_C4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y118_SLICE_X8Y118_C5 = CLBLM_L_X8Y116_SLICE_X10Y116_AQ;
  assign CLBLM_R_X7Y118_SLICE_X8Y118_C6 = 1'b1;
  assign CLBLM_R_X11Y128_SLICE_X14Y128_D4 = 1'b1;
  assign CLBLM_R_X11Y128_SLICE_X14Y128_D5 = 1'b1;
  assign CLBLM_R_X11Y128_SLICE_X14Y128_D6 = 1'b1;
  assign CLBLM_R_X7Y118_SLICE_X8Y118_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X7Y118_SLICE_X8Y118_D1 = CLBLM_R_X7Y113_SLICE_X8Y113_CO6;
  assign CLBLM_R_X7Y118_SLICE_X8Y118_D2 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_R_X7Y118_SLICE_X8Y118_D3 = CLBLM_R_X7Y118_SLICE_X8Y118_DQ;
  assign CLBLM_R_X7Y118_SLICE_X8Y118_D4 = CLBLM_R_X5Y117_SLICE_X6Y117_D5Q;
  assign CLBLM_R_X7Y118_SLICE_X8Y118_D5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y118_SLICE_X8Y118_D6 = CLBLM_R_X3Y118_SLICE_X2Y118_AQ;
  assign LIOI3_X0Y151_OLOGIC_X0Y151_D1 = LIOB33_X0Y65_IOB_X0Y65_I;
  assign CLBLM_R_X11Y122_SLICE_X15Y122_A5 = 1'b1;
  assign CLBLM_R_X11Y122_SLICE_X14Y122_B4 = CLBLM_L_X8Y122_SLICE_X11Y122_AQ;
  assign LIOI3_X0Y71_ILOGIC_X0Y72_D = LIOB33_X0Y71_IOB_X0Y72_I;
  assign LIOI3_X0Y71_ILOGIC_X0Y71_D = LIOB33_X0Y71_IOB_X0Y71_I;
  assign CLBLM_R_X11Y122_SLICE_X14Y122_B5 = CLBLM_L_X10Y123_SLICE_X12Y123_CO6;
  assign RIOI3_X105Y115_ILOGIC_X1Y116_D = RIOB33_X105Y115_IOB_X1Y116_I;
  assign RIOI3_X105Y115_ILOGIC_X1Y115_D = RIOB33_X105Y115_IOB_X1Y115_I;
  assign RIOI3_SING_X105Y150_OLOGIC_X1Y150_D1 = LIOB33_X0Y75_IOB_X0Y75_I;
  assign CLBLM_R_X11Y122_SLICE_X14Y122_B6 = CLBLM_L_X8Y122_SLICE_X11Y122_DO6;
  assign CLBLL_L_X2Y117_SLICE_X0Y117_A1 = CLBLL_L_X2Y117_SLICE_X0Y117_CQ;
  assign CLBLL_L_X2Y117_SLICE_X0Y117_A2 = CLBLM_R_X3Y117_SLICE_X2Y117_BO6;
  assign CLBLL_L_X2Y117_SLICE_X0Y117_A3 = CLBLL_L_X2Y117_SLICE_X0Y117_AQ;
  assign CLBLL_L_X2Y117_SLICE_X0Y117_A4 = CLBLL_L_X4Y117_SLICE_X4Y117_BQ;
  assign CLBLL_L_X2Y117_SLICE_X0Y117_A5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLL_L_X2Y117_SLICE_X0Y117_A6 = CLBLL_L_X2Y114_SLICE_X1Y114_DO6;
  assign CLBLL_L_X2Y117_SLICE_X0Y117_AX = CLBLL_L_X2Y117_SLICE_X0Y117_DO5;
  assign CLBLL_L_X2Y117_SLICE_X0Y117_B1 = CLBLL_L_X2Y117_SLICE_X0Y117_DO6;
  assign CLBLL_L_X2Y117_SLICE_X0Y117_B2 = CLBLM_R_X3Y117_SLICE_X2Y117_BO6;
  assign CLBLL_L_X2Y117_SLICE_X0Y117_B3 = CLBLL_L_X2Y117_SLICE_X1Y117_CO6;
  assign CLBLL_L_X2Y117_SLICE_X0Y117_B4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLL_L_X2Y117_SLICE_X0Y117_B5 = CLBLM_R_X3Y116_SLICE_X3Y116_AQ;
  assign CLBLL_L_X2Y117_SLICE_X0Y117_B6 = CLBLL_L_X2Y117_SLICE_X0Y117_BQ;
  assign CLBLM_L_X10Y128_SLICE_X13Y128_A2 = 1'b1;
  assign CLBLL_L_X2Y117_SLICE_X0Y117_C1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLL_L_X2Y117_SLICE_X0Y117_C2 = CLBLL_L_X2Y117_SLICE_X0Y117_CQ;
  assign CLBLL_L_X2Y117_SLICE_X0Y117_C3 = CLBLL_L_X2Y117_SLICE_X0Y117_BQ;
  assign CLBLL_L_X2Y117_SLICE_X0Y117_C4 = CLBLL_L_X2Y114_SLICE_X1Y114_DO6;
  assign CLBLL_L_X2Y117_SLICE_X0Y117_C5 = 1'b1;
  assign CLBLL_L_X2Y117_SLICE_X0Y117_C6 = CLBLM_R_X3Y117_SLICE_X2Y117_BO6;
  assign RIOI3_X105Y153_OLOGIC_X1Y154_D1 = RIOB33_X105Y101_IOB_X1Y102_I;
  assign CLBLL_L_X2Y117_SLICE_X0Y117_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLL_L_X2Y117_SLICE_X0Y117_D1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLL_L_X2Y117_SLICE_X0Y117_D2 = CLBLL_L_X2Y117_SLICE_X0Y117_CQ;
  assign CLBLL_L_X2Y117_SLICE_X0Y117_D3 = CLBLL_L_X2Y117_SLICE_X0Y117_AQ;
  assign CLBLL_L_X2Y117_SLICE_X0Y117_D4 = CLBLL_L_X2Y117_SLICE_X0Y117_BQ;
  assign CLBLL_L_X2Y117_SLICE_X0Y117_D5 = CLBLL_L_X2Y117_SLICE_X1Y117_BQ;
  assign CLBLL_L_X2Y117_SLICE_X0Y117_D6 = 1'b1;
  assign CLBLL_L_X2Y117_SLICE_X1Y117_A1 = CLBLM_R_X3Y116_SLICE_X2Y116_BQ;
  assign CLBLL_L_X2Y117_SLICE_X1Y117_A2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLL_L_X2Y117_SLICE_X1Y117_A3 = CLBLL_L_X2Y117_SLICE_X1Y117_AQ;
  assign CLBLL_L_X2Y117_SLICE_X1Y117_A4 = CLBLM_R_X5Y116_SLICE_X6Y116_BQ;
  assign CLBLL_L_X2Y117_SLICE_X1Y117_A5 = CLBLL_L_X2Y112_SLICE_X1Y112_BQ;
  assign CLBLL_L_X2Y117_SLICE_X1Y117_A6 = CLBLM_L_X8Y112_SLICE_X10Y112_CQ;
  assign CLBLM_R_X7Y124_SLICE_X9Y124_D2 = 1'b1;
  assign LIOI3_X0Y141_OLOGIC_X0Y142_D1 = LIOB33_X0Y53_IOB_X0Y54_I;
  assign LIOI3_TBYTESRC_X0Y181_OLOGIC_X0Y181_T1 = 1'b1;
  assign CLBLL_L_X2Y117_SLICE_X1Y117_B1 = CLBLL_L_X2Y117_SLICE_X1Y117_DO6;
  assign CLBLL_L_X2Y117_SLICE_X1Y117_B2 = CLBLL_L_X2Y117_SLICE_X1Y117_BQ;
  assign CLBLL_L_X2Y117_SLICE_X1Y117_B3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLL_L_X2Y117_SLICE_X1Y117_B4 = CLBLM_L_X10Y117_SLICE_X12Y117_AQ;
  assign CLBLL_L_X2Y117_SLICE_X1Y117_B5 = CLBLM_R_X3Y117_SLICE_X2Y117_BO6;
  assign CLBLL_L_X2Y117_SLICE_X1Y117_B6 = CLBLL_L_X2Y117_SLICE_X0Y117_AQ;
  assign RIOI3_X105Y153_OLOGIC_X1Y154_T1 = 1'b1;
  assign CLBLL_L_X2Y117_SLICE_X1Y117_C1 = CLBLL_L_X2Y117_SLICE_X0Y117_AQ;
  assign CLBLL_L_X2Y117_SLICE_X1Y117_C2 = CLBLM_R_X5Y111_SLICE_X7Y111_DO6;
  assign CLBLL_L_X2Y117_SLICE_X1Y117_C3 = CLBLL_L_X2Y117_SLICE_X0Y117_CQ;
  assign CLBLL_L_X2Y117_SLICE_X1Y117_C4 = CLBLL_L_X2Y117_SLICE_X1Y117_BQ;
  assign CLBLL_L_X2Y117_SLICE_X1Y117_C5 = CLBLL_L_X2Y114_SLICE_X1Y114_BO5;
  assign CLBLL_L_X2Y117_SLICE_X1Y117_C6 = CLBLM_L_X8Y116_SLICE_X10Y116_AO6;
  assign CLBLL_L_X2Y117_SLICE_X1Y117_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign LIOB33_X0Y103_IOB_X0Y104_O = CLBLL_L_X2Y111_SLICE_X0Y111_CO5;
  assign LIOB33_X0Y103_IOB_X0Y103_O = CLBLL_L_X2Y113_SLICE_X0Y113_AO6;
  assign CLBLL_L_X2Y117_SLICE_X1Y117_D1 = CLBLM_R_X5Y111_SLICE_X7Y111_DO6;
  assign CLBLL_L_X2Y117_SLICE_X1Y117_D2 = 1'b1;
  assign CLBLL_L_X2Y117_SLICE_X1Y117_D3 = CLBLM_L_X8Y116_SLICE_X10Y116_AO6;
  assign CLBLL_L_X2Y117_SLICE_X1Y117_D4 = CLBLL_L_X2Y117_SLICE_X0Y117_CQ;
  assign CLBLL_L_X2Y117_SLICE_X1Y117_D5 = CLBLL_L_X2Y114_SLICE_X1Y114_BO5;
  assign CLBLL_L_X2Y117_SLICE_X1Y117_D6 = 1'b1;
  assign CLBLM_R_X7Y119_SLICE_X9Y119_A1 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X7Y119_SLICE_X9Y119_A2 = CLBLM_L_X10Y118_SLICE_X13Y118_CQ;
  assign CLBLM_R_X7Y119_SLICE_X9Y119_A3 = 1'b1;
  assign CLBLM_R_X7Y119_SLICE_X9Y119_A4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y119_SLICE_X9Y119_A5 = 1'b1;
  assign CLBLM_R_X7Y119_SLICE_X9Y119_A6 = CLBLM_L_X8Y120_SLICE_X10Y120_BQ;
  assign RIOI3_X105Y127_ILOGIC_X1Y128_D = RIOB33_X105Y127_IOB_X1Y128_I;
  assign CLBLM_R_X7Y119_SLICE_X9Y119_B1 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X7Y119_SLICE_X9Y119_B2 = CLBLM_L_X10Y118_SLICE_X13Y118_CQ;
  assign CLBLM_R_X7Y119_SLICE_X9Y119_B3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y119_SLICE_X9Y119_B4 = CLBLM_L_X8Y117_SLICE_X10Y117_DO5;
  assign CLBLM_R_X7Y119_SLICE_X9Y119_B5 = CLBLM_R_X5Y119_SLICE_X6Y119_AQ;
  assign CLBLM_R_X7Y119_SLICE_X9Y119_B6 = 1'b1;
  assign RIOB33_X105Y189_IOB_X1Y190_O = CLBLM_R_X13Y119_SLICE_X18Y119_AQ;
  assign RIOB33_X105Y189_IOB_X1Y189_O = CLBLM_L_X8Y122_SLICE_X10Y122_AQ;
  assign RIOI3_X105Y153_OLOGIC_X1Y153_D1 = RIOB33_X105Y101_IOB_X1Y101_I;
  assign CLBLM_R_X5Y109_SLICE_X7Y109_A1 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_R_X5Y109_SLICE_X7Y109_A2 = CLBLM_R_X5Y112_SLICE_X7Y112_AO6;
  assign CLBLM_R_X5Y109_SLICE_X7Y109_A3 = CLBLM_R_X5Y109_SLICE_X7Y109_AQ;
  assign CLBLM_R_X5Y109_SLICE_X7Y109_A4 = CLBLM_R_X3Y118_SLICE_X2Y118_AQ;
  assign CLBLM_R_X5Y109_SLICE_X7Y109_A5 = CLBLM_R_X5Y109_SLICE_X6Y109_AQ;
  assign CLBLM_R_X5Y109_SLICE_X7Y109_A6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y119_SLICE_X9Y119_C1 = CLBLM_L_X8Y114_SLICE_X10Y114_C5Q;
  assign CLBLM_R_X7Y119_SLICE_X9Y119_C2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y119_SLICE_X9Y119_C3 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X5Y109_SLICE_X7Y109_B1 = 1'b1;
  assign CLBLM_R_X5Y109_SLICE_X7Y109_B2 = 1'b1;
  assign CLBLM_R_X5Y109_SLICE_X7Y109_B3 = 1'b1;
  assign CLBLM_R_X5Y109_SLICE_X7Y109_B4 = 1'b1;
  assign CLBLM_R_X5Y109_SLICE_X7Y109_B5 = 1'b1;
  assign CLBLM_R_X5Y109_SLICE_X7Y109_B6 = 1'b1;
  assign CLBLM_R_X7Y119_SLICE_X9Y119_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X7Y119_SLICE_X9Y119_D1 = CLBLM_R_X3Y115_SLICE_X2Y115_BQ;
  assign CLBLM_R_X5Y109_SLICE_X7Y109_C1 = 1'b1;
  assign CLBLM_R_X5Y109_SLICE_X7Y109_C2 = 1'b1;
  assign CLBLM_R_X5Y109_SLICE_X7Y109_C3 = 1'b1;
  assign CLBLM_R_X5Y109_SLICE_X7Y109_C4 = 1'b1;
  assign CLBLM_R_X5Y109_SLICE_X7Y109_C5 = 1'b1;
  assign CLBLM_R_X5Y109_SLICE_X7Y109_C6 = 1'b1;
  assign CLBLM_R_X7Y119_SLICE_X9Y119_D3 = CLBLM_R_X5Y110_SLICE_X7Y110_AQ;
  assign CLBLM_R_X7Y119_SLICE_X9Y119_D4 = CLBLL_L_X2Y120_SLICE_X0Y120_CO6;
  assign CLBLM_R_X5Y109_SLICE_X7Y109_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X7Y119_SLICE_X8Y119_A1 = 1'b1;
  assign CLBLM_R_X7Y119_SLICE_X8Y119_A2 = CLBLM_R_X11Y121_SLICE_X14Y121_CO6;
  assign CLBLM_R_X7Y119_SLICE_X8Y119_A3 = CLBLM_R_X7Y119_SLICE_X8Y119_AQ;
  assign CLBLM_R_X7Y119_SLICE_X8Y119_A4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y119_SLICE_X8Y119_A5 = CLBLM_R_X7Y120_SLICE_X8Y120_AQ;
  assign CLBLM_R_X5Y109_SLICE_X7Y109_D1 = 1'b1;
  assign CLBLM_R_X5Y109_SLICE_X7Y109_D2 = 1'b1;
  assign CLBLM_R_X5Y109_SLICE_X7Y109_D3 = 1'b1;
  assign CLBLM_R_X5Y109_SLICE_X7Y109_D4 = 1'b1;
  assign CLBLM_R_X5Y109_SLICE_X7Y109_D5 = 1'b1;
  assign CLBLM_R_X5Y109_SLICE_X7Y109_D6 = 1'b1;
  assign CLBLM_R_X7Y119_SLICE_X8Y119_A6 = CLBLM_L_X10Y118_SLICE_X13Y118_CQ;
  assign CLBLM_R_X7Y119_SLICE_X8Y119_B1 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X7Y119_SLICE_X8Y119_B2 = CLBLM_R_X7Y117_SLICE_X8Y117_DO5;
  assign CLBLM_R_X7Y119_SLICE_X8Y119_B3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y119_SLICE_X8Y119_B4 = CLBLM_R_X7Y119_SLICE_X9Y119_BQ;
  assign CLBLM_R_X5Y109_SLICE_X6Y109_A1 = CLBLM_R_X5Y109_SLICE_X6Y109_CQ;
  assign CLBLM_R_X5Y109_SLICE_X6Y109_A2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X5Y109_SLICE_X6Y109_A3 = CLBLM_R_X5Y109_SLICE_X6Y109_AQ;
  assign CLBLM_R_X5Y109_SLICE_X6Y109_A4 = CLBLM_R_X3Y118_SLICE_X2Y118_AQ;
  assign CLBLM_R_X5Y109_SLICE_X6Y109_A5 = 1'b1;
  assign CLBLM_R_X5Y109_SLICE_X6Y109_A6 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_R_X7Y119_SLICE_X8Y119_C1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y119_SLICE_X8Y119_C2 = CLBLM_R_X7Y119_SLICE_X8Y119_CQ;
  assign CLBLM_R_X7Y119_SLICE_X8Y119_C3 = CLBLL_L_X4Y120_SLICE_X4Y120_AO6;
  assign CLBLM_R_X7Y119_SLICE_X8Y119_C4 = CLBLM_L_X8Y119_SLICE_X11Y119_BQ;
  assign CLBLM_R_X5Y109_SLICE_X6Y109_B1 = CLBLM_R_X3Y117_SLICE_X3Y117_B5Q;
  assign CLBLM_R_X5Y109_SLICE_X6Y109_B2 = CLBLM_R_X5Y109_SLICE_X6Y109_BQ;
  assign CLBLM_R_X5Y109_SLICE_X6Y109_B3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X5Y109_SLICE_X6Y109_B4 = CLBLM_R_X3Y118_SLICE_X2Y118_AQ;
  assign CLBLM_R_X5Y109_SLICE_X6Y109_B5 = 1'b1;
  assign CLBLM_R_X5Y109_SLICE_X6Y109_B6 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_R_X7Y119_SLICE_X8Y119_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X7Y119_SLICE_X8Y119_D1 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X7Y119_SLICE_X8Y119_D2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X5Y109_SLICE_X6Y109_C1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X5Y109_SLICE_X6Y109_C2 = CLBLM_R_X3Y118_SLICE_X2Y118_AQ;
  assign CLBLM_R_X5Y109_SLICE_X6Y109_C3 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_R_X5Y109_SLICE_X6Y109_C4 = CLBLM_R_X5Y110_SLICE_X6Y110_CO6;
  assign CLBLM_R_X5Y109_SLICE_X6Y109_C5 = CLBLM_R_X5Y109_SLICE_X6Y109_CQ;
  assign CLBLM_R_X5Y109_SLICE_X6Y109_C6 = CLBLM_L_X10Y110_SLICE_X12Y110_BQ;
  assign CLBLM_R_X7Y119_SLICE_X8Y119_D3 = CLBLM_R_X7Y119_SLICE_X8Y119_DQ;
  assign CLBLM_R_X7Y119_SLICE_X8Y119_D4 = CLBLM_R_X11Y122_SLICE_X14Y122_AQ;
  assign CLBLM_R_X7Y119_SLICE_X8Y119_D5 = CLBLM_R_X7Y118_SLICE_X9Y118_AQ;
  assign CLBLM_R_X5Y109_SLICE_X6Y109_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X7Y119_SLICE_X8Y119_D6 = 1'b1;
  assign CLBLM_R_X11Y122_SLICE_X14Y122_C5 = 1'b1;
  assign CLBLM_R_X5Y109_SLICE_X6Y109_D1 = 1'b1;
  assign CLBLM_R_X5Y109_SLICE_X6Y109_D2 = 1'b1;
  assign CLBLM_R_X5Y109_SLICE_X6Y109_D3 = 1'b1;
  assign CLBLM_R_X5Y109_SLICE_X6Y109_D4 = 1'b1;
  assign CLBLM_R_X5Y109_SLICE_X6Y109_D5 = 1'b1;
  assign CLBLM_R_X5Y109_SLICE_X6Y109_D6 = 1'b1;
  assign CLBLM_R_X11Y122_SLICE_X14Y122_C6 = 1'b1;
  assign LIOI3_X0Y115_OLOGIC_X0Y116_D1 = CLBLM_L_X8Y123_SLICE_X11Y123_AQ;
  assign CLBLM_L_X10Y128_SLICE_X12Y128_A6 = 1'b1;
  assign CLBLL_L_X2Y118_SLICE_X0Y118_A1 = RIOB33_X105Y135_IOB_X1Y136_I;
  assign CLBLL_L_X2Y118_SLICE_X0Y118_A2 = CLBLM_R_X3Y122_SLICE_X3Y122_AO5;
  assign CLBLL_L_X2Y118_SLICE_X0Y118_A3 = CLBLL_L_X4Y117_SLICE_X4Y117_AQ;
  assign CLBLL_L_X2Y118_SLICE_X0Y118_A4 = CLBLL_L_X2Y121_SLICE_X1Y121_BO6;
  assign CLBLL_L_X2Y118_SLICE_X0Y118_A5 = RIOB33_X105Y113_IOB_X1Y113_I;
  assign CLBLL_L_X2Y118_SLICE_X0Y118_A6 = RIOB33_X105Y135_IOB_X1Y135_I;
  assign CLBLM_L_X10Y128_SLICE_X12Y128_B1 = 1'b1;
  assign CLBLM_L_X10Y128_SLICE_X12Y128_B2 = 1'b1;
  assign CLBLL_L_X2Y118_SLICE_X0Y118_B1 = CLBLM_R_X3Y124_SLICE_X2Y124_AO5;
  assign CLBLL_L_X2Y118_SLICE_X0Y118_B2 = LIOB33_X0Y67_IOB_X0Y68_I;
  assign CLBLL_L_X2Y118_SLICE_X0Y118_B3 = CLBLL_L_X2Y120_SLICE_X1Y120_AO6;
  assign CLBLL_L_X2Y118_SLICE_X0Y118_B4 = CLBLL_L_X2Y121_SLICE_X1Y121_BO6;
  assign CLBLL_L_X2Y118_SLICE_X0Y118_B5 = CLBLM_R_X5Y119_SLICE_X6Y119_CQ;
  assign CLBLL_L_X2Y118_SLICE_X0Y118_B6 = CLBLL_L_X2Y113_SLICE_X0Y113_AO5;
  assign CLBLM_L_X8Y116_SLICE_X10Y116_B1 = CLBLM_R_X11Y115_SLICE_X15Y115_CQ;
  assign LIOI3_X0Y115_OLOGIC_X0Y116_T1 = 1'b1;
  assign CLBLL_L_X2Y118_SLICE_X0Y118_C1 = CLBLM_R_X3Y122_SLICE_X3Y122_AO6;
  assign CLBLL_L_X2Y118_SLICE_X0Y118_C2 = RIOB33_X105Y133_IOB_X1Y133_I;
  assign CLBLL_L_X2Y118_SLICE_X0Y118_C3 = RIOB33_X105Y131_IOB_X1Y131_I;
  assign CLBLL_L_X2Y118_SLICE_X0Y118_C4 = RIOB33_X105Y133_IOB_X1Y134_I;
  assign CLBLL_L_X2Y118_SLICE_X0Y118_C5 = RIOB33_X105Y131_IOB_X1Y132_I;
  assign CLBLL_L_X2Y118_SLICE_X0Y118_C6 = CLBLM_R_X7Y119_SLICE_X8Y119_AQ;
  assign CLBLL_L_X2Y118_SLICE_X0Y118_D1 = CLBLL_L_X2Y118_SLICE_X0Y118_AO6;
  assign CLBLL_L_X2Y118_SLICE_X0Y118_D2 = CLBLL_L_X2Y117_SLICE_X1Y117_AQ;
  assign CLBLL_L_X2Y118_SLICE_X0Y118_D3 = CLBLL_L_X2Y118_SLICE_X0Y118_CO6;
  assign CLBLL_L_X2Y118_SLICE_X0Y118_D4 = CLBLM_R_X3Y117_SLICE_X2Y117_CO6;
  assign CLBLL_L_X2Y118_SLICE_X0Y118_D5 = CLBLM_R_X3Y121_SLICE_X2Y121_AO6;
  assign CLBLL_L_X2Y118_SLICE_X0Y118_D6 = CLBLL_L_X2Y118_SLICE_X0Y118_BO6;
  assign CLBLM_L_X8Y116_SLICE_X10Y116_B2 = CLBLM_L_X10Y110_SLICE_X12Y110_BQ;
  assign CLBLM_L_X8Y116_SLICE_X10Y116_B3 = CLBLM_L_X8Y117_SLICE_X10Y117_AQ;
  assign CLBLL_L_X2Y118_SLICE_X1Y118_A1 = CLBLL_L_X2Y112_SLICE_X1Y112_A5Q;
  assign CLBLL_L_X2Y118_SLICE_X1Y118_A2 = CLBLL_L_X2Y121_SLICE_X0Y121_BO6;
  assign CLBLL_L_X2Y118_SLICE_X1Y118_A3 = CLBLM_R_X5Y115_SLICE_X6Y115_AQ;
  assign CLBLL_L_X2Y118_SLICE_X1Y118_A4 = CLBLM_R_X3Y122_SLICE_X3Y122_AO6;
  assign CLBLL_L_X2Y118_SLICE_X1Y118_A5 = CLBLM_R_X3Y124_SLICE_X2Y124_AO6;
  assign CLBLL_L_X2Y118_SLICE_X1Y118_A6 = CLBLL_L_X2Y120_SLICE_X1Y120_AO6;
  assign LIOB33_X0Y105_IOB_X0Y106_O = CLBLL_L_X2Y111_SLICE_X0Y111_DO5;
  assign LIOB33_X0Y105_IOB_X0Y105_O = CLBLL_L_X2Y111_SLICE_X0Y111_DO6;
  assign LIOI3_X0Y115_OLOGIC_X0Y115_D1 = CLBLM_R_X11Y114_SLICE_X14Y114_DQ;
  assign CLBLL_L_X2Y118_SLICE_X1Y118_B1 = CLBLM_R_X3Y122_SLICE_X2Y122_BO5;
  assign CLBLL_L_X2Y118_SLICE_X1Y118_B2 = CLBLM_R_X3Y118_SLICE_X2Y118_CO6;
  assign CLBLL_L_X2Y118_SLICE_X1Y118_B3 = 1'b1;
  assign CLBLL_L_X2Y118_SLICE_X1Y118_B4 = CLBLM_R_X5Y116_SLICE_X7Y116_AQ;
  assign CLBLL_L_X2Y118_SLICE_X1Y118_B5 = CLBLL_L_X2Y118_SLICE_X1Y118_AO6;
  assign CLBLL_L_X2Y118_SLICE_X1Y118_B6 = CLBLL_L_X2Y118_SLICE_X1Y118_CO6;
  assign CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_CE = 1'b1;
  assign CLBLL_L_X2Y118_SLICE_X1Y118_C1 = CLBLM_R_X3Y124_SLICE_X2Y124_AO6;
  assign CLBLL_L_X2Y118_SLICE_X1Y118_C2 = CLBLL_L_X4Y118_SLICE_X5Y118_BQ;
  assign CLBLL_L_X2Y118_SLICE_X1Y118_C3 = CLBLL_L_X2Y121_SLICE_X1Y121_BO5;
  assign CLBLL_L_X2Y118_SLICE_X1Y118_C4 = 1'b1;
  assign CLBLL_L_X2Y118_SLICE_X1Y118_C5 = RIOB33_X105Y105_IOB_X1Y106_I;
  assign CLBLL_L_X2Y118_SLICE_X1Y118_C6 = CLBLL_L_X2Y121_SLICE_X1Y121_BO6;
  assign CLBLL_L_X2Y118_SLICE_X1Y118_D1 = 1'b1;
  assign CLBLL_L_X2Y118_SLICE_X1Y118_D2 = 1'b1;
  assign CLBLL_L_X2Y118_SLICE_X1Y118_D3 = 1'b1;
  assign CLBLL_L_X2Y118_SLICE_X1Y118_D4 = 1'b1;
  assign CLBLL_L_X2Y118_SLICE_X1Y118_D5 = 1'b1;
  assign CLBLL_L_X2Y118_SLICE_X1Y118_D6 = 1'b1;
  assign RIOB33_X105Y191_IOB_X1Y192_O = CLBLM_L_X12Y115_SLICE_X16Y115_AQ;
  assign RIOB33_X105Y191_IOB_X1Y191_O = CLBLM_L_X8Y116_SLICE_X10Y116_AQ;
  assign CLBLM_R_X7Y120_SLICE_X9Y120_A1 = CLBLM_R_X11Y120_SLICE_X14Y120_CO6;
  assign CLBLM_R_X7Y120_SLICE_X9Y120_A2 = CLBLM_R_X7Y117_SLICE_X8Y117_AQ;
  assign CLBLM_R_X7Y120_SLICE_X9Y120_A3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y120_SLICE_X9Y120_A4 = CLBLM_R_X7Y117_SLICE_X9Y117_BQ;
  assign CLBLM_R_X7Y120_SLICE_X9Y120_A5 = CLBLM_R_X7Y122_SLICE_X9Y122_DO6;
  assign CLBLM_R_X7Y120_SLICE_X9Y120_A6 = 1'b1;
  assign LIOI3_X0Y115_OLOGIC_X0Y115_T1 = 1'b1;
  assign CLBLM_R_X7Y120_SLICE_X9Y120_B1 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_R_X7Y120_SLICE_X9Y120_B2 = CLBLM_R_X7Y120_SLICE_X9Y120_BQ;
  assign CLBLM_R_X7Y120_SLICE_X9Y120_B3 = CLBLL_L_X4Y113_SLICE_X5Y113_BQ;
  assign CLBLM_R_X7Y120_SLICE_X9Y120_B4 = CLBLM_L_X10Y118_SLICE_X12Y118_AQ;
  assign CLBLM_R_X7Y120_SLICE_X9Y120_B5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y120_SLICE_X9Y120_B6 = CLBLM_R_X3Y118_SLICE_X2Y118_AQ;
  assign LIOI3_X0Y195_OLOGIC_X0Y196_D1 = LIOB33_X0Y69_IOB_X0Y69_I;
  assign CLBLM_R_X5Y110_SLICE_X7Y110_A1 = CLBLM_R_X5Y110_SLICE_X7Y110_DO6;
  assign CLBLM_R_X5Y110_SLICE_X7Y110_A2 = CLBLM_R_X3Y118_SLICE_X2Y118_AQ;
  assign CLBLM_R_X5Y110_SLICE_X7Y110_A3 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_R_X5Y110_SLICE_X7Y110_A4 = CLBLM_L_X8Y112_SLICE_X11Y112_AQ;
  assign CLBLM_R_X5Y110_SLICE_X7Y110_A5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X5Y110_SLICE_X7Y110_A6 = 1'b1;
  assign CLBLM_R_X7Y120_SLICE_X9Y120_C1 = 1'b1;
  assign CLBLM_R_X7Y120_SLICE_X9Y120_C2 = CLBLM_R_X7Y120_SLICE_X9Y120_CQ;
  assign CLBLM_R_X7Y120_SLICE_X9Y120_C3 = CLBLM_L_X8Y120_SLICE_X10Y120_AQ;
  assign CLBLM_R_X5Y110_SLICE_X7Y110_B1 = CLBLM_R_X7Y110_SLICE_X8Y110_BQ;
  assign CLBLM_R_X5Y110_SLICE_X7Y110_B2 = CLBLM_R_X5Y110_SLICE_X7Y110_BQ;
  assign CLBLM_R_X5Y110_SLICE_X7Y110_B3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X5Y110_SLICE_X7Y110_B4 = CLBLM_R_X3Y118_SLICE_X2Y118_AQ;
  assign CLBLM_R_X5Y110_SLICE_X7Y110_B5 = CLBLM_R_X3Y117_SLICE_X3Y117_B5Q;
  assign CLBLM_R_X5Y110_SLICE_X7Y110_B6 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_R_X7Y120_SLICE_X9Y120_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X7Y120_SLICE_X9Y120_D1 = CLBLM_L_X10Y118_SLICE_X12Y118_AQ;
  assign CLBLM_R_X5Y110_SLICE_X7Y110_C1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X5Y110_SLICE_X7Y110_C2 = CLBLM_R_X7Y112_SLICE_X8Y112_BQ;
  assign CLBLM_R_X5Y110_SLICE_X7Y110_C3 = 1'b1;
  assign CLBLM_R_X5Y110_SLICE_X7Y110_C4 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X5Y110_SLICE_X7Y110_C5 = 1'b1;
  assign CLBLM_R_X5Y110_SLICE_X7Y110_C6 = CLBLL_L_X2Y114_SLICE_X1Y114_AQ;
  assign CLBLM_R_X7Y120_SLICE_X9Y120_D3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y120_SLICE_X9Y120_D4 = CLBLM_R_X7Y121_SLICE_X8Y121_BQ;
  assign CLBLM_R_X5Y110_SLICE_X7Y110_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X7Y120_SLICE_X8Y120_A1 = CLBLM_R_X5Y120_SLICE_X6Y120_A5Q;
  assign CLBLM_R_X7Y120_SLICE_X8Y120_A2 = CLBLM_R_X7Y124_SLICE_X8Y124_AQ;
  assign CLBLM_R_X7Y120_SLICE_X8Y120_A3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y120_SLICE_X8Y120_A4 = CLBLM_R_X7Y120_SLICE_X9Y120_A5Q;
  assign CLBLM_R_X7Y120_SLICE_X8Y120_A5 = CLBLM_R_X3Y110_SLICE_X2Y110_AQ;
  assign CLBLM_R_X5Y110_SLICE_X7Y110_D1 = CLBLM_R_X3Y120_SLICE_X3Y120_BO6;
  assign CLBLM_R_X5Y110_SLICE_X7Y110_D2 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X5Y110_SLICE_X7Y110_D3 = CLBLM_R_X7Y109_SLICE_X8Y109_AQ;
  assign CLBLM_R_X5Y110_SLICE_X7Y110_D4 = CLBLM_R_X5Y116_SLICE_X7Y116_CQ;
  assign CLBLM_R_X5Y110_SLICE_X7Y110_D5 = CLBLM_R_X5Y110_SLICE_X7Y110_AQ;
  assign CLBLM_R_X5Y110_SLICE_X7Y110_D6 = 1'b1;
  assign CLBLM_R_X7Y120_SLICE_X8Y120_A6 = CLBLM_L_X10Y124_SLICE_X12Y124_AQ;
  assign CLBLM_R_X7Y120_SLICE_X8Y120_B1 = 1'b1;
  assign CLBLM_R_X7Y120_SLICE_X8Y120_B2 = CLBLM_R_X7Y120_SLICE_X8Y120_BQ;
  assign CLBLM_R_X7Y120_SLICE_X8Y120_B3 = CLBLM_R_X5Y115_SLICE_X6Y115_CO5;
  assign CLBLM_R_X7Y120_SLICE_X8Y120_B4 = CLBLM_L_X8Y120_SLICE_X10Y120_BQ;
  assign CLBLM_R_X5Y110_SLICE_X6Y110_A1 = CLBLM_R_X5Y110_SLICE_X6Y110_DO6;
  assign CLBLM_R_X5Y110_SLICE_X6Y110_A2 = 1'b1;
  assign CLBLM_R_X5Y110_SLICE_X6Y110_A3 = RIOB33_X105Y141_IOB_X1Y142_I;
  assign CLBLM_R_X5Y110_SLICE_X6Y110_A4 = CLBLM_R_X7Y128_SLICE_X8Y128_AQ;
  assign CLBLM_R_X5Y110_SLICE_X6Y110_A5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X5Y110_SLICE_X6Y110_A6 = CLBLM_R_X5Y111_SLICE_X6Y111_CQ;
  assign CLBLM_R_X7Y120_SLICE_X8Y120_C1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y120_SLICE_X8Y120_C2 = CLBLM_R_X7Y120_SLICE_X8Y120_CQ;
  assign CLBLM_R_X7Y120_SLICE_X8Y120_C3 = 1'b1;
  assign CLBLM_R_X5Y110_SLICE_X6Y110_B1 = CLBLL_L_X2Y120_SLICE_X1Y120_DO6;
  assign CLBLM_R_X5Y110_SLICE_X6Y110_B2 = CLBLM_R_X5Y117_SLICE_X7Y117_DO6;
  assign CLBLM_R_X5Y110_SLICE_X6Y110_B3 = CLBLM_R_X5Y109_SLICE_X6Y109_CQ;
  assign CLBLM_R_X5Y110_SLICE_X6Y110_B4 = CLBLM_R_X7Y112_SLICE_X8Y112_BQ;
  assign CLBLM_R_X5Y110_SLICE_X6Y110_B5 = RIOB33_X105Y121_IOB_X1Y121_I;
  assign CLBLM_R_X5Y110_SLICE_X6Y110_B6 = CLBLL_L_X4Y110_SLICE_X5Y110_DO6;
  assign CLBLM_R_X7Y120_SLICE_X8Y120_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X7Y120_SLICE_X8Y120_D1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y120_SLICE_X8Y120_D2 = 1'b1;
  assign CLBLM_R_X5Y110_SLICE_X6Y110_C1 = 1'b1;
  assign CLBLM_R_X5Y110_SLICE_X6Y110_C2 = CLBLM_R_X5Y111_SLICE_X7Y111_CO5;
  assign CLBLM_R_X5Y110_SLICE_X6Y110_C3 = CLBLL_L_X2Y120_SLICE_X0Y120_CO6;
  assign CLBLM_R_X5Y110_SLICE_X6Y110_C4 = CLBLM_R_X3Y120_SLICE_X3Y120_BO6;
  assign CLBLM_R_X5Y110_SLICE_X6Y110_C5 = CLBLM_R_X5Y117_SLICE_X7Y117_DO6;
  assign CLBLM_R_X5Y110_SLICE_X6Y110_C6 = CLBLL_L_X4Y120_SLICE_X5Y120_AO6;
  assign CLBLM_R_X7Y120_SLICE_X8Y120_D3 = CLBLM_L_X8Y120_SLICE_X11Y120_CQ;
  assign CLBLM_R_X7Y120_SLICE_X8Y120_D4 = 1'b1;
  assign CLBLM_R_X7Y120_SLICE_X8Y120_D5 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X5Y110_SLICE_X6Y110_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X7Y120_SLICE_X8Y120_D6 = CLBLM_R_X7Y123_SLICE_X9Y123_AQ;
  assign LIOI3_TBYTESRC_X0Y157_OLOGIC_X0Y157_D1 = RIOB33_X105Y115_IOB_X1Y115_I;
  assign CLBLM_R_X5Y110_SLICE_X6Y110_D1 = CLBLM_R_X5Y111_SLICE_X6Y111_C5Q;
  assign CLBLM_R_X5Y110_SLICE_X6Y110_D2 = CLBLM_R_X5Y110_SLICE_X6Y110_AQ;
  assign CLBLM_R_X5Y110_SLICE_X6Y110_D3 = CLBLM_R_X5Y111_SLICE_X7Y111_DO6;
  assign CLBLM_R_X5Y110_SLICE_X6Y110_D4 = CLBLM_R_X7Y111_SLICE_X9Y111_BO5;
  assign CLBLM_R_X5Y110_SLICE_X6Y110_D5 = 1'b1;
  assign CLBLM_R_X5Y110_SLICE_X6Y110_D6 = CLBLM_R_X5Y114_SLICE_X6Y114_DQ;
  assign LIOI3_TBYTESRC_X0Y157_OLOGIC_X0Y157_T1 = 1'b1;
  assign CLBLM_R_X11Y122_SLICE_X14Y122_D2 = 1'b1;
  assign CLBLM_R_X7Y122_SLICE_X9Y122_D1 = CLBLM_R_X7Y124_SLICE_X8Y124_AQ;
  assign CLBLM_R_X7Y122_SLICE_X9Y122_D2 = CLBLM_L_X10Y124_SLICE_X12Y124_AQ;
  assign CLBLM_R_X11Y122_SLICE_X14Y122_D4 = 1'b1;
  assign CLBLL_L_X2Y119_SLICE_X0Y119_A1 = CLBLM_R_X3Y124_SLICE_X2Y124_AO5;
  assign CLBLL_L_X2Y119_SLICE_X0Y119_A2 = CLBLL_L_X2Y113_SLICE_X1Y113_CQ;
  assign CLBLL_L_X2Y119_SLICE_X0Y119_A3 = CLBLL_L_X2Y120_SLICE_X1Y120_AO6;
  assign CLBLL_L_X2Y119_SLICE_X0Y119_A4 = RIOB33_X105Y137_IOB_X1Y137_I;
  assign CLBLL_L_X2Y119_SLICE_X0Y119_A5 = RIOB33_X105Y129_IOB_X1Y129_I;
  assign CLBLL_L_X2Y119_SLICE_X0Y119_A6 = CLBLM_R_X5Y119_SLICE_X6Y119_CQ;
  assign CLBLL_L_X2Y119_SLICE_X0Y119_B1 = CLBLL_L_X2Y119_SLICE_X0Y119_DO6;
  assign CLBLL_L_X2Y119_SLICE_X0Y119_B2 = CLBLM_R_X7Y119_SLICE_X8Y119_AQ;
  assign CLBLL_L_X2Y119_SLICE_X0Y119_B3 = CLBLM_R_X3Y121_SLICE_X2Y121_DO6;
  assign CLBLL_L_X2Y119_SLICE_X0Y119_B4 = CLBLL_L_X2Y120_SLICE_X0Y120_BO6;
  assign CLBLL_L_X2Y119_SLICE_X0Y119_B5 = CLBLL_L_X2Y120_SLICE_X0Y120_AO5;
  assign CLBLL_L_X2Y119_SLICE_X0Y119_B6 = CLBLL_L_X2Y119_SLICE_X0Y119_CO6;
  assign CLBLM_R_X11Y122_SLICE_X14Y122_C3 = 1'b1;
  assign CLBLM_R_X11Y122_SLICE_X14Y122_D5 = 1'b1;
  assign CLBLL_L_X2Y119_SLICE_X0Y119_C1 = CLBLL_L_X2Y119_SLICE_X0Y119_AO6;
  assign CLBLL_L_X2Y119_SLICE_X0Y119_C2 = CLBLL_L_X2Y121_SLICE_X0Y121_AO6;
  assign CLBLL_L_X2Y119_SLICE_X0Y119_C3 = CLBLL_L_X2Y117_SLICE_X1Y117_AQ;
  assign CLBLL_L_X2Y119_SLICE_X0Y119_C4 = CLBLM_R_X3Y121_SLICE_X2Y121_AO6;
  assign CLBLL_L_X2Y119_SLICE_X0Y119_C5 = 1'b1;
  assign CLBLL_L_X2Y119_SLICE_X0Y119_C6 = LIOB33_X0Y67_IOB_X0Y68_I;
  assign CLBLL_L_X2Y119_SLICE_X0Y119_D1 = CLBLL_L_X4Y117_SLICE_X4Y117_AQ;
  assign CLBLL_L_X2Y119_SLICE_X0Y119_D2 = CLBLM_R_X3Y117_SLICE_X2Y117_CO6;
  assign CLBLL_L_X2Y119_SLICE_X0Y119_D3 = CLBLL_L_X2Y122_SLICE_X0Y122_AO6;
  assign CLBLL_L_X2Y119_SLICE_X0Y119_D4 = RIOB33_X105Y113_IOB_X1Y113_I;
  assign CLBLL_L_X2Y119_SLICE_X0Y119_D5 = 1'b1;
  assign CLBLL_L_X2Y119_SLICE_X0Y119_D6 = CLBLL_L_X2Y120_SLICE_X0Y120_AO6;
  assign LIOB33_X0Y107_IOB_X0Y108_O = CLBLL_L_X2Y111_SLICE_X0Y111_BO5;
  assign LIOB33_X0Y107_IOB_X0Y107_O = CLBLL_L_X2Y109_SLICE_X0Y109_AO6;
  assign CLBLM_R_X7Y122_SLICE_X9Y122_D5 = CLBLM_R_X5Y120_SLICE_X6Y120_A5Q;
  assign LIOI3_X0Y73_ILOGIC_X0Y74_D = LIOB33_X0Y73_IOB_X0Y74_I;
  assign CLBLL_L_X2Y119_SLICE_X1Y119_A1 = CLBLM_R_X3Y124_SLICE_X2Y124_AO6;
  assign CLBLL_L_X2Y119_SLICE_X1Y119_A2 = RIOB33_X105Y131_IOB_X1Y132_I;
  assign CLBLL_L_X2Y119_SLICE_X1Y119_A3 = RIOB33_X105Y133_IOB_X1Y133_I;
  assign CLBLL_L_X2Y119_SLICE_X1Y119_A4 = RIOB33_X105Y133_IOB_X1Y134_I;
  assign CLBLL_L_X2Y119_SLICE_X1Y119_A5 = RIOB33_X105Y131_IOB_X1Y131_I;
  assign CLBLL_L_X2Y119_SLICE_X1Y119_A6 = 1'b1;
  assign LIOI3_X0Y73_ILOGIC_X0Y73_D = LIOB33_X0Y73_IOB_X0Y73_I;
  assign CLBLL_L_X2Y119_SLICE_X1Y119_B1 = CLBLL_L_X4Y120_SLICE_X5Y120_DO6;
  assign CLBLL_L_X2Y119_SLICE_X1Y119_B2 = CLBLM_R_X3Y120_SLICE_X3Y120_BO6;
  assign CLBLL_L_X2Y119_SLICE_X1Y119_B3 = CLBLM_R_X3Y121_SLICE_X2Y121_CO6;
  assign CLBLL_L_X2Y119_SLICE_X1Y119_B4 = CLBLL_L_X4Y120_SLICE_X4Y120_AO6;
  assign CLBLL_L_X2Y119_SLICE_X1Y119_B5 = CLBLL_L_X4Y120_SLICE_X4Y120_BO6;
  assign CLBLL_L_X2Y119_SLICE_X1Y119_B6 = CLBLL_L_X2Y119_SLICE_X1Y119_CO6;
  assign CLBLM_R_X7Y122_SLICE_X9Y122_D6 = CLBLM_R_X7Y120_SLICE_X9Y120_A5Q;
  assign RIOI3_X105Y117_ILOGIC_X1Y118_D = RIOB33_X105Y117_IOB_X1Y118_I;
  assign RIOB33_X105Y193_IOB_X1Y194_O = CLBLM_R_X11Y128_SLICE_X15Y128_AQ;
  assign CLBLL_L_X2Y119_SLICE_X1Y119_C1 = CLBLL_L_X2Y118_SLICE_X1Y118_BO6;
  assign CLBLL_L_X2Y119_SLICE_X1Y119_C2 = CLBLL_L_X2Y122_SLICE_X0Y122_BO6;
  assign CLBLL_L_X2Y119_SLICE_X1Y119_C3 = CLBLL_L_X2Y118_SLICE_X0Y118_DO6;
  assign CLBLL_L_X2Y119_SLICE_X1Y119_C4 = CLBLL_L_X2Y120_SLICE_X1Y120_BO6;
  assign CLBLL_L_X2Y119_SLICE_X1Y119_C5 = CLBLL_L_X2Y121_SLICE_X1Y121_CO6;
  assign CLBLL_L_X2Y119_SLICE_X1Y119_C6 = CLBLL_L_X4Y118_SLICE_X4Y118_CO6;
  assign RIOB33_X105Y193_IOB_X1Y193_O = CLBLM_L_X10Y124_SLICE_X13Y124_AQ;
  assign CLBLL_L_X2Y119_SLICE_X1Y119_D1 = CLBLL_L_X2Y121_SLICE_X1Y121_AO6;
  assign CLBLL_L_X2Y119_SLICE_X1Y119_D2 = RIOB33_X105Y105_IOB_X1Y106_I;
  assign CLBLL_L_X2Y119_SLICE_X1Y119_D3 = CLBLM_R_X3Y122_SLICE_X2Y122_BO5;
  assign CLBLL_L_X2Y119_SLICE_X1Y119_D4 = CLBLM_R_X5Y116_SLICE_X7Y116_AQ;
  assign CLBLL_L_X2Y119_SLICE_X1Y119_D5 = CLBLL_L_X2Y122_SLICE_X0Y122_AO6;
  assign CLBLL_L_X2Y119_SLICE_X1Y119_D6 = CLBLL_L_X4Y118_SLICE_X5Y118_BQ;
  assign CLBLM_R_X11Y120_SLICE_X14Y120_C4 = CLBLM_L_X12Y119_SLICE_X17Y119_AO5;
  assign CLBLM_R_X7Y121_SLICE_X9Y121_A1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y121_SLICE_X9Y121_A2 = CLBLM_L_X8Y133_SLICE_X11Y133_AO6;
  assign CLBLM_R_X7Y121_SLICE_X9Y121_A3 = CLBLM_R_X7Y121_SLICE_X9Y121_AQ;
  assign CLBLM_R_X7Y121_SLICE_X9Y121_A4 = CLBLM_R_X7Y121_SLICE_X8Y121_BQ;
  assign CLBLM_R_X7Y121_SLICE_X9Y121_A5 = CLBLM_R_X7Y121_SLICE_X9Y121_CO5;
  assign CLBLM_R_X7Y121_SLICE_X9Y121_A6 = CLBLL_L_X4Y115_SLICE_X4Y115_CQ;
  assign LIOI3_X0Y175_OLOGIC_X0Y176_T1 = 1'b1;
  assign CLBLM_R_X7Y121_SLICE_X9Y121_AX = CLBLM_R_X7Y121_SLICE_X9Y121_CO6;
  assign CLBLM_R_X11Y120_SLICE_X14Y120_C5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y121_SLICE_X9Y121_B1 = CLBLM_L_X8Y115_SLICE_X11Y115_CQ;
  assign CLBLM_R_X7Y121_SLICE_X9Y121_B2 = CLBLM_R_X7Y121_SLICE_X9Y121_BQ;
  assign CLBLM_R_X7Y121_SLICE_X9Y121_B3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y121_SLICE_X9Y121_B4 = CLBLM_R_X7Y121_SLICE_X9Y121_DO5;
  assign CLBLM_R_X7Y121_SLICE_X9Y121_B5 = CLBLM_R_X7Y121_SLICE_X8Y121_AQ;
  assign CLBLM_R_X7Y121_SLICE_X9Y121_B6 = CLBLM_L_X8Y133_SLICE_X11Y133_AO6;
  assign CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_I = CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_O;
  assign CLBLM_R_X5Y111_SLICE_X7Y111_A1 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_R_X5Y111_SLICE_X7Y111_A2 = CLBLM_R_X3Y118_SLICE_X2Y118_AQ;
  assign CLBLM_R_X5Y111_SLICE_X7Y111_A3 = CLBLM_R_X5Y111_SLICE_X7Y111_AQ;
  assign CLBLM_R_X5Y111_SLICE_X7Y111_A4 = CLBLM_R_X7Y110_SLICE_X8Y110_AQ;
  assign CLBLM_R_X5Y111_SLICE_X7Y111_A5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X5Y111_SLICE_X7Y111_A6 = CLBLM_R_X5Y112_SLICE_X7Y112_CO6;
  assign CLBLM_R_X7Y121_SLICE_X9Y121_C1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y121_SLICE_X9Y121_C2 = CLBLM_L_X8Y133_SLICE_X11Y133_AO6;
  assign CLBLM_R_X7Y121_SLICE_X9Y121_C3 = CLBLM_R_X7Y121_SLICE_X9Y121_A5Q;
  assign CLBLM_R_X5Y111_SLICE_X7Y111_B1 = CLBLM_R_X5Y113_SLICE_X7Y113_CO6;
  assign CLBLM_R_X5Y111_SLICE_X7Y111_B2 = CLBLM_R_X5Y111_SLICE_X7Y111_BQ;
  assign CLBLM_R_X5Y111_SLICE_X7Y111_B3 = CLBLM_R_X5Y110_SLICE_X6Y110_BO6;
  assign CLBLM_R_X5Y111_SLICE_X7Y111_B4 = CLBLL_L_X4Y110_SLICE_X4Y110_CQ;
  assign CLBLM_R_X5Y111_SLICE_X7Y111_B5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X5Y111_SLICE_X7Y111_B6 = CLBLM_R_X5Y110_SLICE_X7Y110_AO5;
  assign CLBLM_R_X7Y121_SLICE_X9Y121_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X7Y121_SLICE_X9Y121_D1 = CLBLM_L_X8Y120_SLICE_X10Y120_CQ;
  assign CLBLM_R_X5Y111_SLICE_X7Y111_C1 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X5Y111_SLICE_X7Y111_C2 = CLBLL_L_X2Y120_SLICE_X0Y120_CO6;
  assign CLBLM_R_X5Y111_SLICE_X7Y111_C3 = CLBLL_L_X4Y120_SLICE_X5Y120_DO6;
  assign CLBLM_R_X5Y111_SLICE_X7Y111_C4 = CLBLL_L_X2Y119_SLICE_X0Y119_BO6;
  assign CLBLM_R_X5Y111_SLICE_X7Y111_C5 = CLBLM_R_X3Y120_SLICE_X3Y120_BO6;
  assign CLBLM_R_X5Y111_SLICE_X7Y111_C6 = 1'b1;
  assign CLBLM_R_X7Y121_SLICE_X9Y121_D3 = CLBLM_R_X5Y121_SLICE_X7Y121_DO6;
  assign CLBLM_R_X7Y121_SLICE_X9Y121_D4 = CLBLM_R_X7Y121_SLICE_X9Y121_A5Q;
  assign CLBLM_R_X5Y111_SLICE_X7Y111_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X7Y121_SLICE_X8Y121_A1 = 1'b1;
  assign CLBLM_R_X7Y121_SLICE_X8Y121_A2 = CLBLM_R_X7Y121_SLICE_X9Y121_DO5;
  assign CLBLM_R_X7Y121_SLICE_X8Y121_A3 = CLBLM_R_X7Y121_SLICE_X8Y121_AQ;
  assign CLBLM_R_X7Y121_SLICE_X8Y121_A4 = CLBLM_R_X7Y122_SLICE_X9Y122_BO6;
  assign CLBLM_R_X7Y121_SLICE_X8Y121_A5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X5Y111_SLICE_X7Y111_D1 = CLBLL_L_X4Y120_SLICE_X5Y120_AO6;
  assign CLBLM_R_X5Y111_SLICE_X7Y111_D2 = CLBLM_R_X5Y119_SLICE_X7Y119_CO6;
  assign CLBLM_R_X5Y111_SLICE_X7Y111_D3 = 1'b1;
  assign CLBLM_R_X5Y111_SLICE_X7Y111_D4 = CLBLM_R_X5Y111_SLICE_X7Y111_CO6;
  assign CLBLM_R_X5Y111_SLICE_X7Y111_D5 = CLBLL_L_X2Y120_SLICE_X1Y120_DO6;
  assign CLBLM_R_X5Y111_SLICE_X7Y111_D6 = CLBLM_R_X3Y119_SLICE_X2Y119_AO6;
  assign CLBLM_R_X7Y121_SLICE_X8Y121_A6 = CLBLL_L_X4Y121_SLICE_X5Y121_AQ;
  assign CLBLM_R_X7Y121_SLICE_X8Y121_B1 = CLBLM_R_X7Y121_SLICE_X9Y121_A5Q;
  assign CLBLM_R_X7Y121_SLICE_X8Y121_B2 = CLBLM_R_X7Y121_SLICE_X8Y121_BQ;
  assign CLBLM_R_X7Y121_SLICE_X8Y121_B3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y121_SLICE_X8Y121_B4 = CLBLM_R_X7Y122_SLICE_X9Y122_BO6;
  assign CLBLM_R_X5Y111_SLICE_X6Y111_A1 = CLBLM_R_X5Y115_SLICE_X6Y115_DO6;
  assign CLBLM_R_X5Y111_SLICE_X6Y111_A2 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X5Y111_SLICE_X6Y111_A3 = CLBLM_R_X5Y111_SLICE_X6Y111_AQ;
  assign CLBLM_R_X5Y111_SLICE_X6Y111_A4 = CLBLL_L_X4Y111_SLICE_X5Y111_CO6;
  assign CLBLM_R_X5Y111_SLICE_X6Y111_A5 = CLBLM_L_X10Y110_SLICE_X13Y110_AQ;
  assign CLBLM_R_X5Y111_SLICE_X6Y111_A6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y121_SLICE_X8Y121_C1 = CLBLM_R_X7Y127_SLICE_X8Y127_AQ;
  assign CLBLM_R_X7Y121_SLICE_X8Y121_C2 = CLBLM_L_X8Y121_SLICE_X10Y121_AQ;
  assign CLBLM_R_X7Y121_SLICE_X8Y121_C3 = CLBLL_L_X2Y117_SLICE_X0Y117_A5Q;
  assign CLBLM_R_X5Y111_SLICE_X6Y111_B1 = CLBLM_R_X5Y112_SLICE_X6Y112_CO6;
  assign CLBLM_R_X5Y111_SLICE_X6Y111_B2 = CLBLM_R_X7Y117_SLICE_X8Y117_CQ;
  assign CLBLM_R_X5Y111_SLICE_X6Y111_B3 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X5Y111_SLICE_X6Y111_B4 = CLBLM_R_X7Y110_SLICE_X9Y110_AQ;
  assign CLBLM_R_X5Y111_SLICE_X6Y111_B5 = 1'b1;
  assign CLBLM_R_X5Y111_SLICE_X6Y111_B6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y121_SLICE_X8Y121_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X7Y121_SLICE_X8Y121_D1 = CLBLM_R_X7Y121_SLICE_X9Y121_AQ;
  assign CLBLM_R_X5Y111_SLICE_X6Y111_C1 = CLBLM_R_X5Y110_SLICE_X6Y110_AQ;
  assign CLBLM_R_X5Y111_SLICE_X6Y111_C2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X5Y111_SLICE_X6Y111_C3 = CLBLM_R_X5Y111_SLICE_X6Y111_BQ;
  assign CLBLM_R_X5Y111_SLICE_X6Y111_C4 = CLBLL_L_X4Y110_SLICE_X4Y110_A5Q;
  assign CLBLM_R_X5Y111_SLICE_X6Y111_C5 = CLBLM_R_X5Y111_SLICE_X6Y111_DO6;
  assign CLBLM_R_X5Y111_SLICE_X6Y111_C6 = 1'b1;
  assign CLBLM_R_X7Y121_SLICE_X8Y121_D2 = CLBLM_R_X7Y121_SLICE_X9Y121_A5Q;
  assign CLBLM_R_X7Y121_SLICE_X8Y121_D3 = CLBLM_R_X7Y121_SLICE_X8Y121_BQ;
  assign CLBLM_R_X7Y121_SLICE_X8Y121_D4 = CLBLM_L_X8Y120_SLICE_X10Y120_CQ;
  assign CLBLM_R_X5Y111_SLICE_X6Y111_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X7Y121_SLICE_X8Y121_D6 = CLBLM_R_X7Y121_SLICE_X9Y121_BQ;
  assign CLBLM_R_X5Y111_SLICE_X6Y111_D1 = CLBLL_L_X4Y115_SLICE_X4Y115_BQ;
  assign CLBLM_R_X5Y111_SLICE_X6Y111_D2 = CLBLM_R_X5Y111_SLICE_X6Y111_CQ;
  assign CLBLM_R_X5Y111_SLICE_X6Y111_D3 = 1'b1;
  assign CLBLM_R_X5Y111_SLICE_X6Y111_D4 = CLBLM_R_X5Y115_SLICE_X6Y115_BQ;
  assign CLBLM_R_X5Y111_SLICE_X6Y111_D5 = CLBLM_R_X7Y113_SLICE_X8Y113_AQ;
  assign CLBLM_R_X5Y111_SLICE_X6Y111_D6 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign LIOI3_X0Y133_OLOGIC_X0Y133_D1 = CLBLM_R_X7Y124_SLICE_X8Y124_A5Q;
  assign CLBLM_L_X10Y118_SLICE_X12Y118_B6 = 1'b1;
  assign LIOI3_X0Y175_OLOGIC_X0Y175_T1 = 1'b1;
  assign CLBLM_L_X10Y118_SLICE_X12Y118_C1 = CLBLM_R_X7Y119_SLICE_X8Y119_BQ;
  assign CLBLM_L_X10Y118_SLICE_X12Y118_C2 = CLBLM_L_X10Y121_SLICE_X12Y121_DO6;
  assign CLBLM_L_X10Y118_SLICE_X12Y118_C4 = CLBLL_L_X4Y110_SLICE_X4Y110_CQ;
  assign CLBLM_L_X8Y128_SLICE_X11Y128_A1 = 1'b1;
  assign CLBLM_L_X8Y128_SLICE_X11Y128_A2 = 1'b1;
  assign CLBLM_L_X8Y128_SLICE_X11Y128_A3 = 1'b1;
  assign CLBLM_L_X8Y128_SLICE_X11Y128_A4 = 1'b1;
  assign CLBLM_L_X8Y128_SLICE_X11Y128_A5 = 1'b1;
  assign CLBLM_L_X8Y128_SLICE_X11Y128_A6 = 1'b1;
  assign CLBLL_L_X2Y120_SLICE_X0Y120_A1 = RIOB33_X105Y133_IOB_X1Y133_I;
  assign CLBLL_L_X2Y120_SLICE_X0Y120_A2 = CLBLM_R_X3Y122_SLICE_X3Y122_AO6;
  assign CLBLL_L_X2Y120_SLICE_X0Y120_A3 = RIOB33_X105Y131_IOB_X1Y132_I;
  assign CLBLL_L_X2Y120_SLICE_X0Y120_A4 = RIOB33_X105Y133_IOB_X1Y134_I;
  assign CLBLL_L_X2Y120_SLICE_X0Y120_A5 = RIOB33_X105Y131_IOB_X1Y131_I;
  assign CLBLL_L_X2Y120_SLICE_X0Y120_A6 = 1'b1;
  assign CLBLM_L_X8Y128_SLICE_X11Y128_B1 = 1'b1;
  assign CLBLM_L_X8Y128_SLICE_X11Y128_B2 = 1'b1;
  assign CLBLL_L_X2Y120_SLICE_X0Y120_B1 = CLBLL_L_X4Y122_SLICE_X5Y122_DO6;
  assign CLBLL_L_X2Y120_SLICE_X0Y120_B2 = CLBLM_R_X3Y124_SLICE_X2Y124_AO6;
  assign CLBLL_L_X2Y120_SLICE_X0Y120_B3 = RIOB33_X105Y131_IOB_X1Y132_I;
  assign CLBLL_L_X2Y120_SLICE_X0Y120_B4 = RIOB33_X105Y133_IOB_X1Y134_I;
  assign CLBLL_L_X2Y120_SLICE_X0Y120_B5 = RIOB33_X105Y131_IOB_X1Y131_I;
  assign CLBLL_L_X2Y120_SLICE_X0Y120_B6 = RIOB33_X105Y133_IOB_X1Y133_I;
  assign CLBLM_L_X8Y128_SLICE_X11Y128_B4 = 1'b1;
  assign CLBLM_L_X8Y128_SLICE_X11Y128_B5 = 1'b1;
  assign CLBLL_L_X2Y120_SLICE_X0Y120_C1 = CLBLM_R_X5Y122_SLICE_X6Y122_CO6;
  assign CLBLL_L_X2Y120_SLICE_X0Y120_C2 = CLBLL_L_X4Y118_SLICE_X4Y118_CO6;
  assign CLBLL_L_X2Y120_SLICE_X0Y120_C3 = CLBLL_L_X2Y122_SLICE_X0Y122_CO6;
  assign CLBLL_L_X2Y120_SLICE_X0Y120_C4 = CLBLM_R_X3Y118_SLICE_X2Y118_DO6;
  assign CLBLL_L_X2Y120_SLICE_X0Y120_C5 = CLBLL_L_X2Y119_SLICE_X1Y119_DO6;
  assign CLBLL_L_X2Y120_SLICE_X0Y120_C6 = CLBLL_L_X2Y121_SLICE_X1Y121_CO6;
  assign CLBLM_L_X8Y128_SLICE_X11Y128_C4 = 1'b1;
  assign CLBLM_L_X8Y128_SLICE_X11Y128_C5 = 1'b1;
  assign CLBLM_L_X8Y128_SLICE_X11Y128_C6 = 1'b1;
  assign CLBLM_L_X8Y128_SLICE_X11Y128_D1 = 1'b1;
  assign CLBLM_L_X8Y128_SLICE_X11Y128_D2 = 1'b1;
  assign CLBLM_L_X8Y128_SLICE_X11Y128_D4 = 1'b1;
  assign CLBLM_L_X8Y128_SLICE_X11Y128_D5 = 1'b1;
  assign CLBLL_L_X2Y120_SLICE_X0Y120_D1 = 1'b1;
  assign CLBLL_L_X2Y120_SLICE_X0Y120_D2 = 1'b1;
  assign CLBLL_L_X2Y120_SLICE_X0Y120_D3 = 1'b1;
  assign CLBLL_L_X2Y120_SLICE_X0Y120_D4 = 1'b1;
  assign CLBLL_L_X2Y120_SLICE_X0Y120_D5 = 1'b1;
  assign CLBLL_L_X2Y120_SLICE_X0Y120_D6 = 1'b1;
  assign CLBLM_L_X8Y128_SLICE_X11Y128_D6 = 1'b1;
  assign CLBLM_L_X8Y128_SLICE_X10Y128_A1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y128_SLICE_X10Y128_A2 = RIOB33_X105Y143_IOB_X1Y143_I;
  assign CLBLM_L_X8Y128_SLICE_X10Y128_A3 = 1'b1;
  assign CLBLM_L_X8Y120_SLICE_X10Y120_A3 = CLBLM_L_X8Y119_SLICE_X10Y119_CQ;
  assign CLBLM_L_X8Y128_SLICE_X10Y128_A4 = CLBLL_L_X4Y121_SLICE_X5Y121_BO5;
  assign CLBLM_L_X8Y128_SLICE_X10Y128_A5 = CLBLM_L_X8Y122_SLICE_X10Y122_AQ;
  assign CLBLM_L_X8Y128_SLICE_X10Y128_A6 = 1'b1;
  assign CLBLM_L_X8Y120_SLICE_X10Y120_A4 = CLBLM_R_X7Y121_SLICE_X8Y121_CQ;
  assign CLBLM_L_X8Y128_SLICE_X10Y128_B1 = 1'b1;
  assign CLBLM_L_X8Y128_SLICE_X10Y128_B2 = 1'b1;
  assign CLBLM_L_X8Y128_SLICE_X10Y128_B3 = 1'b1;
  assign CLBLM_L_X8Y120_SLICE_X10Y120_A5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y128_SLICE_X10Y128_B4 = 1'b1;
  assign CLBLM_L_X8Y128_SLICE_X10Y128_B5 = 1'b1;
  assign CLBLM_L_X8Y128_SLICE_X10Y128_B6 = 1'b1;
  assign RIOB33_X105Y195_IOB_X1Y196_O = CLBLM_R_X11Y120_SLICE_X14Y120_AQ;
  assign CLBLM_L_X8Y128_SLICE_X10Y128_C1 = 1'b1;
  assign CLBLM_L_X8Y128_SLICE_X10Y128_C2 = 1'b1;
  assign CLBLM_L_X8Y128_SLICE_X10Y128_C3 = 1'b1;
  assign CLBLM_L_X8Y128_SLICE_X10Y128_C4 = 1'b1;
  assign CLBLM_L_X8Y128_SLICE_X10Y128_C5 = 1'b1;
  assign CLBLM_L_X8Y128_SLICE_X10Y128_C6 = 1'b1;
  assign CLBLL_L_X2Y120_SLICE_X1Y120_A1 = RIOB33_X105Y133_IOB_X1Y134_I;
  assign CLBLL_L_X2Y120_SLICE_X1Y120_A2 = RIOB33_X105Y133_IOB_X1Y133_I;
  assign CLBLL_L_X2Y120_SLICE_X1Y120_A3 = RIOB33_X105Y131_IOB_X1Y131_I;
  assign CLBLL_L_X2Y120_SLICE_X1Y120_A4 = RIOB33_X105Y131_IOB_X1Y132_I;
  assign CLBLL_L_X2Y120_SLICE_X1Y120_A5 = CLBLM_R_X3Y124_SLICE_X2Y124_AO6;
  assign CLBLL_L_X2Y120_SLICE_X1Y120_A6 = 1'b1;
  assign CLBLL_L_X2Y120_SLICE_X1Y120_B1 = CLBLL_L_X4Y121_SLICE_X4Y121_CO5;
  assign CLBLL_L_X2Y120_SLICE_X1Y120_B2 = CLBLM_R_X3Y122_SLICE_X2Y122_AO6;
  assign CLBLL_L_X2Y120_SLICE_X1Y120_B3 = CLBLL_L_X2Y120_SLICE_X0Y120_AO6;
  assign CLBLM_L_X8Y128_SLICE_X10Y128_D4 = 1'b1;
  assign CLBLL_L_X2Y120_SLICE_X1Y120_B4 = CLBLL_L_X4Y122_SLICE_X5Y122_DO6;
  assign CLBLL_L_X2Y120_SLICE_X1Y120_B5 = CLBLL_L_X2Y119_SLICE_X1Y119_AO6;
  assign CLBLL_L_X2Y120_SLICE_X1Y120_B6 = CLBLM_R_X3Y122_SLICE_X2Y122_CO6;
  assign CLBLM_L_X8Y128_SLICE_X10Y128_D1 = 1'b1;
  assign CLBLM_L_X8Y128_SLICE_X10Y128_D2 = 1'b1;
  assign CLBLM_L_X8Y128_SLICE_X10Y128_D3 = 1'b1;
  assign CLBLL_L_X2Y120_SLICE_X1Y120_C1 = CLBLL_L_X2Y121_SLICE_X1Y121_AO6;
  assign CLBLL_L_X2Y120_SLICE_X1Y120_C2 = CLBLM_R_X3Y122_SLICE_X2Y122_AO6;
  assign CLBLL_L_X2Y120_SLICE_X1Y120_C3 = CLBLM_R_X3Y121_SLICE_X2Y121_AO5;
  assign CLBLL_L_X2Y120_SLICE_X1Y120_C4 = CLBLL_L_X4Y121_SLICE_X4Y121_CO5;
  assign CLBLL_L_X2Y120_SLICE_X1Y120_C5 = CLBLL_L_X2Y120_SLICE_X0Y120_AO6;
  assign CLBLL_L_X2Y120_SLICE_X1Y120_C6 = CLBLM_R_X3Y122_SLICE_X2Y122_CO6;
  assign CLBLM_L_X8Y120_SLICE_X10Y120_B3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLL_L_X2Y120_SLICE_X1Y120_D1 = CLBLL_L_X2Y120_SLICE_X1Y120_CO6;
  assign CLBLL_L_X2Y120_SLICE_X1Y120_D2 = CLBLM_R_X3Y119_SLICE_X3Y119_CO6;
  assign CLBLL_L_X2Y120_SLICE_X1Y120_D3 = CLBLM_R_X3Y120_SLICE_X2Y120_DO6;
  assign CLBLL_L_X2Y120_SLICE_X1Y120_D4 = CLBLL_L_X2Y120_SLICE_X1Y120_AO5;
  assign CLBLL_L_X2Y120_SLICE_X1Y120_D5 = CLBLL_L_X4Y122_SLICE_X5Y122_DO6;
  assign CLBLL_L_X2Y120_SLICE_X1Y120_D6 = CLBLM_R_X3Y121_SLICE_X3Y121_DO6;
  assign CLBLM_L_X8Y120_SLICE_X10Y120_B4 = CLBLM_R_X7Y122_SLICE_X9Y122_BQ;
  assign LIOB33_X0Y193_IOB_X0Y194_O = LIOB33_X0Y59_IOB_X0Y60_I;
  assign RIOI3_X105Y177_OLOGIC_X1Y177_D1 = CLBLM_R_X103Y177_SLICE_X163Y177_AO6;
  assign CLBLM_R_X7Y122_SLICE_X9Y122_A1 = CLBLL_L_X2Y117_SLICE_X0Y117_CQ;
  assign CLBLM_R_X7Y122_SLICE_X9Y122_A2 = 1'b1;
  assign CLBLM_R_X7Y122_SLICE_X9Y122_A3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y122_SLICE_X9Y122_A4 = CLBLM_L_X10Y122_SLICE_X13Y122_AQ;
  assign CLBLM_R_X7Y122_SLICE_X9Y122_A5 = RIOB33_X105Y143_IOB_X1Y144_I;
  assign CLBLM_R_X7Y122_SLICE_X9Y122_A6 = 1'b1;
  assign CLBLM_R_X7Y122_SLICE_X9Y122_B1 = CLBLM_L_X8Y120_SLICE_X10Y120_A5Q;
  assign CLBLM_R_X7Y122_SLICE_X9Y122_B2 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X7Y122_SLICE_X9Y122_B3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y122_SLICE_X9Y122_B4 = CLBLM_R_X3Y112_SLICE_X3Y112_BQ;
  assign CLBLM_R_X7Y122_SLICE_X9Y122_B5 = CLBLM_L_X8Y120_SLICE_X11Y120_C5Q;
  assign CLBLM_R_X7Y122_SLICE_X9Y122_B6 = 1'b1;
  assign CLBLM_R_X7Y123_SLICE_X9Y123_D2 = CLBLM_R_X7Y122_SLICE_X8Y122_AQ;
  assign CLBLM_R_X5Y112_SLICE_X7Y112_A1 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X5Y112_SLICE_X7Y112_A2 = CLBLM_R_X3Y119_SLICE_X2Y119_AO6;
  assign CLBLM_R_X5Y112_SLICE_X7Y112_A3 = CLBLM_R_X5Y116_SLICE_X7Y116_CQ;
  assign CLBLM_R_X5Y112_SLICE_X7Y112_A4 = CLBLM_R_X7Y109_SLICE_X8Y109_AQ;
  assign CLBLM_R_X5Y112_SLICE_X7Y112_A5 = CLBLM_R_X7Y113_SLICE_X8Y113_BO6;
  assign CLBLM_R_X5Y112_SLICE_X7Y112_A6 = 1'b1;
  assign CLBLM_R_X7Y122_SLICE_X9Y122_C1 = CLBLM_L_X10Y118_SLICE_X12Y118_B5Q;
  assign CLBLM_R_X7Y122_SLICE_X9Y122_C2 = CLBLM_R_X5Y122_SLICE_X6Y122_AO5;
  assign CLBLM_R_X7Y122_SLICE_X9Y122_C3 = CLBLM_L_X10Y123_SLICE_X13Y123_DO6;
  assign CLBLM_R_X5Y112_SLICE_X7Y112_B1 = CLBLM_R_X5Y112_SLICE_X7Y112_DO6;
  assign CLBLM_R_X5Y112_SLICE_X7Y112_B2 = CLBLM_L_X8Y115_SLICE_X10Y115_CQ;
  assign CLBLM_L_X8Y120_SLICE_X10Y120_C6 = CLBLM_L_X8Y120_SLICE_X11Y120_C5Q;
  assign CLBLM_R_X5Y112_SLICE_X7Y112_B3 = CLBLM_R_X5Y111_SLICE_X7Y111_AQ;
  assign CLBLM_R_X5Y112_SLICE_X7Y112_B4 = RIOB33_X105Y121_IOB_X1Y121_I;
  assign CLBLM_R_X5Y112_SLICE_X7Y112_B5 = CLBLM_R_X5Y110_SLICE_X7Y110_DO5;
  assign CLBLM_R_X5Y112_SLICE_X7Y112_B6 = CLBLM_R_X5Y112_SLICE_X7Y112_AO5;
  assign CLBLM_R_X7Y122_SLICE_X9Y122_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X5Y112_SLICE_X7Y112_C1 = CLBLM_R_X5Y114_SLICE_X7Y114_AQ;
  assign CLBLM_R_X5Y112_SLICE_X7Y112_C2 = CLBLM_R_X7Y118_SLICE_X9Y118_CQ;
  assign CLBLM_R_X5Y112_SLICE_X7Y112_C3 = CLBLM_R_X7Y120_SLICE_X9Y120_CQ;
  assign CLBLM_R_X5Y112_SLICE_X7Y112_C4 = CLBLM_R_X5Y115_SLICE_X7Y115_A5Q;
  assign CLBLM_R_X5Y112_SLICE_X7Y112_C5 = RIOB33_X105Y121_IOB_X1Y121_I;
  assign CLBLM_R_X5Y112_SLICE_X7Y112_C6 = CLBLM_R_X5Y114_SLICE_X7Y114_BO6;
  assign CLBLM_R_X7Y122_SLICE_X9Y122_D3 = CLBLM_L_X10Y123_SLICE_X13Y123_DO6;
  assign CLBLM_R_X7Y122_SLICE_X9Y122_D4 = CLBLM_R_X5Y122_SLICE_X6Y122_AO5;
  assign CLBLM_R_X7Y122_SLICE_X8Y122_A1 = 1'b1;
  assign CLBLM_R_X7Y122_SLICE_X8Y122_A2 = CLBLM_L_X10Y122_SLICE_X12Y122_AQ;
  assign CLBLM_R_X7Y122_SLICE_X8Y122_A3 = CLBLM_L_X10Y124_SLICE_X13Y124_BO6;
  assign CLBLM_R_X7Y122_SLICE_X8Y122_A4 = CLBLM_R_X5Y122_SLICE_X6Y122_BQ;
  assign CLBLM_L_X8Y120_SLICE_X10Y120_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X7Y122_SLICE_X8Y122_A5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X5Y112_SLICE_X7Y112_D1 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_R_X5Y112_SLICE_X7Y112_D2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X5Y112_SLICE_X7Y112_D3 = CLBLM_R_X7Y109_SLICE_X8Y109_AQ;
  assign CLBLM_R_X5Y112_SLICE_X7Y112_D4 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X5Y112_SLICE_X7Y112_D5 = CLBLM_R_X3Y118_SLICE_X2Y118_AQ;
  assign CLBLM_R_X5Y112_SLICE_X7Y112_D6 = CLBLM_R_X5Y116_SLICE_X7Y116_CQ;
  assign CLBLM_R_X7Y122_SLICE_X8Y122_A6 = 1'b1;
  assign CLBLM_R_X7Y122_SLICE_X8Y122_B1 = 1'b1;
  assign CLBLM_R_X7Y122_SLICE_X8Y122_B2 = CLBLM_R_X7Y123_SLICE_X8Y123_BQ;
  assign CLBLM_R_X7Y122_SLICE_X8Y122_B3 = CLBLM_L_X10Y124_SLICE_X13Y124_BO6;
  assign CLBLM_R_X7Y122_SLICE_X8Y122_B4 = 1'b1;
  assign CLBLM_R_X5Y112_SLICE_X6Y112_A1 = CLBLM_R_X3Y118_SLICE_X2Y118_AQ;
  assign CLBLM_R_X5Y112_SLICE_X6Y112_A2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X5Y112_SLICE_X6Y112_A3 = CLBLM_R_X5Y112_SLICE_X6Y112_AQ;
  assign CLBLM_R_X5Y112_SLICE_X6Y112_A4 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_R_X5Y112_SLICE_X6Y112_A5 = CLBLM_R_X5Y112_SLICE_X6Y112_CO6;
  assign CLBLM_R_X5Y112_SLICE_X6Y112_A6 = CLBLM_R_X5Y125_SLICE_X6Y125_A5Q;
  assign CLBLM_R_X7Y122_SLICE_X8Y122_C1 = CLBLM_L_X10Y124_SLICE_X13Y124_BO6;
  assign CLBLM_R_X7Y122_SLICE_X8Y122_C2 = 1'b1;
  assign CLBLM_R_X7Y122_SLICE_X8Y122_C3 = CLBLM_L_X8Y118_SLICE_X10Y118_BQ;
  assign CLBLM_R_X5Y112_SLICE_X6Y112_B1 = RIOB33_X105Y121_IOB_X1Y121_I;
  assign CLBLM_R_X5Y112_SLICE_X6Y112_B2 = CLBLM_R_X5Y119_SLICE_X6Y119_BQ;
  assign CLBLM_R_X5Y112_SLICE_X6Y112_B3 = CLBLM_R_X5Y112_SLICE_X6Y112_AQ;
  assign CLBLM_R_X5Y112_SLICE_X6Y112_B4 = CLBLM_L_X8Y115_SLICE_X10Y115_CQ;
  assign CLBLM_R_X5Y112_SLICE_X6Y112_B5 = CLBLM_R_X5Y111_SLICE_X7Y111_AQ;
  assign CLBLM_R_X5Y112_SLICE_X6Y112_B6 = 1'b1;
  assign CLBLM_R_X7Y122_SLICE_X8Y122_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X7Y122_SLICE_X8Y122_D1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y122_SLICE_X8Y122_D2 = CLBLM_R_X7Y122_SLICE_X8Y122_AQ;
  assign CLBLM_R_X5Y112_SLICE_X6Y112_C1 = CLBLL_L_X4Y111_SLICE_X5Y111_AQ;
  assign CLBLM_R_X5Y112_SLICE_X6Y112_C2 = CLBLM_R_X5Y114_SLICE_X7Y114_AQ;
  assign CLBLM_R_X5Y112_SLICE_X6Y112_C3 = RIOB33_X105Y121_IOB_X1Y121_I;
  assign CLBLM_R_X5Y112_SLICE_X6Y112_C4 = CLBLM_R_X7Y120_SLICE_X9Y120_CQ;
  assign CLBLM_R_X5Y112_SLICE_X6Y112_C5 = CLBLM_R_X5Y114_SLICE_X7Y114_BO5;
  assign CLBLM_R_X5Y112_SLICE_X6Y112_C6 = CLBLM_L_X8Y115_SLICE_X10Y115_CQ;
  assign CLBLM_R_X7Y122_SLICE_X8Y122_D3 = CLBLM_R_X7Y122_SLICE_X8Y122_DQ;
  assign CLBLM_R_X7Y122_SLICE_X8Y122_D4 = 1'b1;
  assign CLBLM_R_X7Y122_SLICE_X8Y122_D5 = 1'b1;
  assign CLBLM_R_X5Y112_SLICE_X6Y112_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X7Y122_SLICE_X8Y122_D6 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X5Y112_SLICE_X6Y112_D1 = CLBLM_R_X7Y110_SLICE_X9Y110_CQ;
  assign CLBLM_R_X5Y112_SLICE_X6Y112_D2 = CLBLM_R_X5Y113_SLICE_X6Y113_DO5;
  assign CLBLM_R_X5Y112_SLICE_X6Y112_D3 = CLBLL_L_X4Y121_SLICE_X4Y121_AQ;
  assign CLBLM_R_X5Y112_SLICE_X6Y112_D4 = 1'b1;
  assign CLBLM_R_X5Y112_SLICE_X6Y112_D5 = RIOB33_X105Y121_IOB_X1Y121_I;
  assign CLBLM_R_X5Y112_SLICE_X6Y112_D6 = CLBLM_R_X5Y119_SLICE_X6Y119_BQ;
  assign LIOI3_X0Y197_OLOGIC_X0Y198_D1 = LIOB33_X0Y73_IOB_X0Y73_I;
  assign LIOI3_X0Y197_OLOGIC_X0Y198_T1 = 1'b1;
  assign LIOI3_X0Y135_OLOGIC_X0Y136_D1 = CLBLM_R_X7Y124_SLICE_X8Y124_CQ;
  assign LIOI3_X0Y197_OLOGIC_X0Y197_D1 = LIOB33_X0Y71_IOB_X0Y72_I;
  assign LIOI3_X0Y135_OLOGIC_X0Y136_T1 = 1'b1;
  assign RIOI3_X105Y179_OLOGIC_X1Y180_D1 = CLBLM_R_X11Y113_SLICE_X15Y113_DO6;
  assign LIOI3_X0Y197_OLOGIC_X0Y197_T1 = 1'b1;
  assign LIOI3_X0Y135_OLOGIC_X0Y135_D1 = CLBLL_L_X4Y123_SLICE_X4Y123_AQ;
  assign LIOB33_X0Y111_IOB_X0Y112_O = CLBLM_R_X11Y114_SLICE_X14Y114_D5Q;
  assign LIOB33_X0Y111_IOB_X0Y111_O = 1'b0;
  assign CLBLL_L_X2Y121_SLICE_X0Y121_A1 = CLBLM_R_X3Y124_SLICE_X2Y124_AO5;
  assign CLBLL_L_X2Y121_SLICE_X0Y121_A2 = RIOB33_X105Y133_IOB_X1Y133_I;
  assign CLBLL_L_X2Y121_SLICE_X0Y121_A3 = RIOB33_X105Y131_IOB_X1Y131_I;
  assign CLBLL_L_X2Y121_SLICE_X0Y121_A4 = RIOB33_X105Y133_IOB_X1Y134_I;
  assign CLBLL_L_X2Y121_SLICE_X0Y121_A5 = RIOB33_X105Y131_IOB_X1Y132_I;
  assign CLBLL_L_X2Y121_SLICE_X0Y121_A6 = 1'b1;
  assign RIOI3_X105Y179_OLOGIC_X1Y180_T1 = 1'b1;
  assign LIOI3_X0Y135_OLOGIC_X0Y135_T1 = 1'b1;
  assign CLBLL_L_X2Y121_SLICE_X0Y121_B1 = 1'b1;
  assign CLBLL_L_X2Y121_SLICE_X0Y121_B2 = RIOB33_X105Y133_IOB_X1Y133_I;
  assign CLBLL_L_X2Y121_SLICE_X0Y121_B3 = RIOB33_X105Y131_IOB_X1Y131_I;
  assign CLBLL_L_X2Y121_SLICE_X0Y121_B4 = RIOB33_X105Y133_IOB_X1Y134_I;
  assign CLBLL_L_X2Y121_SLICE_X0Y121_B5 = RIOB33_X105Y131_IOB_X1Y132_I;
  assign CLBLL_L_X2Y121_SLICE_X0Y121_B6 = 1'b1;
  assign RIOI3_X105Y179_OLOGIC_X1Y179_D1 = CLBLM_R_X11Y128_SLICE_X14Y128_AO5;
  assign CLBLL_L_X2Y121_SLICE_X0Y121_C1 = RIOB33_X105Y131_IOB_X1Y132_I;
  assign CLBLL_L_X2Y121_SLICE_X0Y121_C2 = CLBLL_L_X2Y121_SLICE_X0Y121_BO5;
  assign CLBLL_L_X2Y121_SLICE_X0Y121_C3 = CLBLM_R_X5Y121_SLICE_X6Y121_B5Q;
  assign CLBLL_L_X2Y121_SLICE_X0Y121_C4 = CLBLL_L_X2Y121_SLICE_X0Y121_AO5;
  assign CLBLL_L_X2Y121_SLICE_X0Y121_C5 = CLBLM_R_X3Y124_SLICE_X2Y124_AO5;
  assign CLBLL_L_X2Y121_SLICE_X0Y121_C6 = LIOB33_X0Y53_IOB_X0Y54_I;
  assign LIOI3_TBYTESRC_X0Y169_OLOGIC_X0Y170_D1 = RIOB33_SING_X105Y149_IOB_X1Y149_I;
  assign RIOI3_X105Y179_OLOGIC_X1Y179_T1 = 1'b1;
  assign LIOI3_TBYTESRC_X0Y169_OLOGIC_X0Y170_T1 = 1'b1;
  assign CLBLL_L_X2Y121_SLICE_X0Y121_D1 = RIOB33_X105Y131_IOB_X1Y132_I;
  assign CLBLL_L_X2Y121_SLICE_X0Y121_D2 = CLBLL_L_X2Y120_SLICE_X1Y120_AO6;
  assign CLBLL_L_X2Y121_SLICE_X0Y121_D3 = CLBLM_R_X3Y124_SLICE_X2Y124_AO5;
  assign CLBLL_L_X2Y121_SLICE_X0Y121_D4 = CLBLL_L_X4Y117_SLICE_X4Y117_BQ;
  assign CLBLL_L_X2Y121_SLICE_X0Y121_D5 = CLBLL_L_X2Y121_SLICE_X0Y121_BO5;
  assign CLBLL_L_X2Y121_SLICE_X0Y121_D6 = CLBLL_L_X2Y117_SLICE_X0Y117_BQ;
  assign RIOB33_X105Y197_IOB_X1Y197_O = CLBLM_L_X8Y122_SLICE_X10Y122_BO5;
  assign RIOB33_X105Y197_IOB_X1Y198_O = CLBLM_L_X8Y122_SLICE_X10Y122_BO5;
  assign LIOI3_TBYTESRC_X0Y169_OLOGIC_X0Y169_D1 = RIOB33_X105Y121_IOB_X1Y122_I;
  assign CLBLM_R_X37Y119_SLICE_X57Y119_B1 = 1'b1;
  assign LIOI3_TBYTESRC_X0Y169_OLOGIC_X0Y169_T1 = 1'b1;
  assign CLBLL_L_X2Y121_SLICE_X1Y121_A1 = CLBLM_R_X3Y124_SLICE_X2Y124_AO6;
  assign CLBLL_L_X2Y121_SLICE_X1Y121_A2 = RIOB33_X105Y133_IOB_X1Y134_I;
  assign CLBLL_L_X2Y121_SLICE_X1Y121_A3 = RIOB33_X105Y131_IOB_X1Y132_I;
  assign CLBLL_L_X2Y121_SLICE_X1Y121_A4 = RIOB33_X105Y133_IOB_X1Y133_I;
  assign CLBLL_L_X2Y121_SLICE_X1Y121_A5 = RIOB33_X105Y131_IOB_X1Y131_I;
  assign CLBLL_L_X2Y121_SLICE_X1Y121_A6 = 1'b1;
  assign CLBLL_L_X2Y121_SLICE_X1Y121_B1 = 1'b1;
  assign CLBLL_L_X2Y121_SLICE_X1Y121_B2 = RIOB33_X105Y133_IOB_X1Y134_I;
  assign CLBLL_L_X2Y121_SLICE_X1Y121_B3 = RIOB33_X105Y131_IOB_X1Y132_I;
  assign CLBLL_L_X2Y121_SLICE_X1Y121_B4 = RIOB33_X105Y131_IOB_X1Y131_I;
  assign CLBLL_L_X2Y121_SLICE_X1Y121_B5 = RIOB33_X105Y133_IOB_X1Y133_I;
  assign CLBLL_L_X2Y121_SLICE_X1Y121_B6 = 1'b1;
  assign CLBLL_L_X2Y121_SLICE_X1Y121_C1 = CLBLM_R_X3Y122_SLICE_X2Y122_AO6;
  assign CLBLL_L_X2Y121_SLICE_X1Y121_C2 = CLBLM_R_X3Y122_SLICE_X2Y122_CO6;
  assign CLBLL_L_X2Y121_SLICE_X1Y121_C3 = CLBLL_L_X2Y121_SLICE_X1Y121_AO5;
  assign CLBLL_L_X2Y121_SLICE_X1Y121_C4 = CLBLL_L_X4Y121_SLICE_X4Y121_DO6;
  assign CLBLL_L_X2Y121_SLICE_X1Y121_C5 = CLBLL_L_X4Y122_SLICE_X5Y122_AO6;
  assign CLBLL_L_X2Y121_SLICE_X1Y121_C6 = CLBLL_L_X2Y119_SLICE_X1Y119_AO6;
  assign CLBLL_L_X2Y121_SLICE_X1Y121_D1 = CLBLM_R_X3Y122_SLICE_X2Y122_AO6;
  assign CLBLL_L_X2Y121_SLICE_X1Y121_D2 = CLBLM_R_X3Y122_SLICE_X2Y122_CO6;
  assign CLBLL_L_X2Y121_SLICE_X1Y121_D3 = CLBLL_L_X2Y121_SLICE_X1Y121_AO6;
  assign CLBLL_L_X2Y121_SLICE_X1Y121_D4 = CLBLL_L_X4Y121_SLICE_X4Y121_DO6;
  assign CLBLL_L_X2Y121_SLICE_X1Y121_D5 = CLBLM_R_X3Y121_SLICE_X2Y121_AO5;
  assign CLBLL_L_X2Y121_SLICE_X1Y121_D6 = CLBLL_L_X2Y120_SLICE_X1Y120_AO5;
  assign CLBLM_R_X37Y119_SLICE_X57Y119_B3 = 1'b1;
  assign LIOI3_TBYTESRC_X0Y131_OLOGIC_X0Y132_T1 = 1'b1;
  assign CLBLM_R_X37Y119_SLICE_X57Y119_B4 = 1'b1;
  assign CLBLM_L_X8Y110_SLICE_X11Y110_C4 = 1'b1;
  assign CLBLM_L_X8Y110_SLICE_X11Y110_C5 = 1'b1;
  assign CLBLM_R_X7Y123_SLICE_X9Y123_A1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y123_SLICE_X9Y123_A2 = CLBLM_R_X7Y122_SLICE_X8Y122_AQ;
  assign CLBLM_R_X7Y123_SLICE_X9Y123_A3 = CLBLM_R_X7Y123_SLICE_X9Y123_AQ;
  assign CLBLM_R_X7Y123_SLICE_X9Y123_A4 = CLBLM_R_X7Y123_SLICE_X9Y123_BO6;
  assign CLBLM_R_X7Y123_SLICE_X9Y123_A5 = CLBLM_R_X7Y118_SLICE_X8Y118_BQ;
  assign CLBLM_R_X7Y123_SLICE_X9Y123_A6 = 1'b1;
  assign CLBLM_R_X7Y123_SLICE_X9Y123_B1 = CLBLM_R_X7Y122_SLICE_X8Y122_AQ;
  assign CLBLM_R_X7Y123_SLICE_X9Y123_B2 = CLBLM_R_X7Y124_SLICE_X9Y124_AQ;
  assign CLBLM_R_X7Y123_SLICE_X9Y123_B3 = CLBLM_R_X7Y123_SLICE_X9Y123_AQ;
  assign CLBLM_R_X7Y123_SLICE_X9Y123_B4 = CLBLM_L_X10Y123_SLICE_X12Y123_AO6;
  assign CLBLM_R_X7Y123_SLICE_X9Y123_B5 = CLBLM_R_X7Y123_SLICE_X8Y123_AQ;
  assign CLBLM_R_X7Y123_SLICE_X9Y123_B6 = 1'b1;
  assign CLBLM_R_X5Y113_SLICE_X7Y113_A1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X5Y113_SLICE_X7Y113_A2 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X5Y113_SLICE_X7Y113_A3 = CLBLM_R_X5Y113_SLICE_X7Y113_AQ;
  assign CLBLM_R_X5Y113_SLICE_X7Y113_A4 = CLBLM_L_X8Y112_SLICE_X10Y112_AQ;
  assign CLBLM_R_X5Y113_SLICE_X7Y113_A5 = CLBLM_R_X3Y114_SLICE_X3Y114_BQ;
  assign CLBLM_R_X5Y113_SLICE_X7Y113_A6 = 1'b1;
  assign CLBLM_R_X7Y123_SLICE_X9Y123_C1 = CLBLM_R_X7Y123_SLICE_X8Y123_AQ;
  assign CLBLM_R_X7Y123_SLICE_X9Y123_C2 = CLBLM_R_X7Y123_SLICE_X9Y123_AQ;
  assign CLBLM_R_X7Y123_SLICE_X9Y123_C3 = CLBLM_R_X7Y122_SLICE_X8Y122_AQ;
  assign CLBLM_R_X5Y113_SLICE_X7Y113_B1 = CLBLM_R_X7Y122_SLICE_X8Y122_DQ;
  assign CLBLM_R_X5Y113_SLICE_X7Y113_B2 = CLBLM_R_X7Y109_SLICE_X8Y109_CQ;
  assign CLBLM_R_X5Y113_SLICE_X7Y113_B3 = CLBLM_R_X5Y113_SLICE_X7Y113_AQ;
  assign CLBLM_R_X5Y113_SLICE_X7Y113_B4 = CLBLM_R_X5Y121_SLICE_X7Y121_AQ;
  assign CLBLM_R_X5Y113_SLICE_X7Y113_B5 = CLBLL_L_X4Y111_SLICE_X5Y111_AQ;
  assign CLBLM_R_X5Y113_SLICE_X7Y113_B6 = CLBLL_L_X4Y111_SLICE_X4Y111_DQ;
  assign CLBLM_R_X7Y123_SLICE_X9Y123_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X7Y123_SLICE_X9Y123_D1 = CLBLM_R_X7Y123_SLICE_X8Y123_AQ;
  assign CLBLM_R_X5Y113_SLICE_X7Y113_C1 = CLBLL_L_X4Y112_SLICE_X4Y112_DO6;
  assign CLBLM_R_X5Y113_SLICE_X7Y113_C2 = CLBLM_R_X5Y117_SLICE_X7Y117_BQ;
  assign CLBLM_R_X5Y113_SLICE_X7Y113_C3 = CLBLM_L_X8Y112_SLICE_X10Y112_CQ;
  assign CLBLM_R_X5Y113_SLICE_X7Y113_C4 = CLBLM_R_X7Y119_SLICE_X8Y119_CQ;
  assign CLBLM_R_X5Y113_SLICE_X7Y113_C5 = CLBLM_R_X5Y113_SLICE_X7Y113_DO6;
  assign CLBLM_R_X5Y113_SLICE_X7Y113_C6 = CLBLM_R_X5Y114_SLICE_X7Y114_BO6;
  assign CLBLM_R_X7Y123_SLICE_X9Y123_D3 = 1'b1;
  assign CLBLM_R_X7Y123_SLICE_X9Y123_D4 = 1'b1;
  assign CLBLM_R_X5Y113_SLICE_X7Y113_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X7Y123_SLICE_X8Y123_A1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y123_SLICE_X8Y123_A2 = CLBLM_R_X7Y123_SLICE_X9Y123_BO6;
  assign CLBLM_R_X7Y123_SLICE_X8Y123_A3 = CLBLM_R_X7Y123_SLICE_X8Y123_AQ;
  assign CLBLM_R_X7Y123_SLICE_X8Y123_A4 = CLBLM_R_X7Y122_SLICE_X8Y122_AQ;
  assign CLBLM_R_X7Y123_SLICE_X8Y123_A5 = CLBLM_R_X7Y123_SLICE_X9Y123_AQ;
  assign CLBLM_R_X5Y113_SLICE_X7Y113_D1 = CLBLM_R_X3Y111_SLICE_X3Y111_AQ;
  assign CLBLM_R_X5Y113_SLICE_X7Y113_D2 = CLBLM_R_X5Y117_SLICE_X7Y117_BQ;
  assign CLBLM_R_X5Y113_SLICE_X7Y113_D3 = CLBLM_R_X7Y119_SLICE_X8Y119_DQ;
  assign CLBLM_R_X5Y113_SLICE_X7Y113_D4 = CLBLM_R_X7Y111_SLICE_X8Y111_DO6;
  assign CLBLM_R_X5Y113_SLICE_X7Y113_D5 = CLBLM_R_X5Y113_SLICE_X7Y113_BO6;
  assign CLBLM_R_X5Y113_SLICE_X7Y113_D6 = CLBLL_L_X4Y116_SLICE_X4Y116_BQ;
  assign CLBLM_R_X7Y123_SLICE_X8Y123_A6 = CLBLM_R_X7Y120_SLICE_X8Y120_BQ;
  assign CLBLM_R_X7Y123_SLICE_X8Y123_B1 = 1'b1;
  assign CLBLM_R_X7Y123_SLICE_X8Y123_B2 = 1'b1;
  assign CLBLM_R_X7Y123_SLICE_X8Y123_B3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y123_SLICE_X8Y123_B4 = CLBLM_R_X7Y119_SLICE_X8Y119_C5Q;
  assign CLBLM_R_X5Y113_SLICE_X6Y113_A1 = CLBLM_R_X5Y114_SLICE_X7Y114_DO6;
  assign CLBLM_R_X5Y113_SLICE_X6Y113_A2 = CLBLM_L_X8Y121_SLICE_X11Y121_BQ;
  assign CLBLM_R_X5Y113_SLICE_X6Y113_A3 = CLBLM_R_X5Y113_SLICE_X6Y113_AQ;
  assign CLBLM_R_X5Y113_SLICE_X6Y113_A4 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_R_X5Y113_SLICE_X6Y113_A5 = CLBLM_R_X3Y118_SLICE_X2Y118_AQ;
  assign CLBLM_R_X5Y113_SLICE_X6Y113_A6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y123_SLICE_X8Y123_C1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y123_SLICE_X8Y123_C2 = CLBLM_R_X7Y123_SLICE_X8Y123_CQ;
  assign CLBLM_R_X7Y123_SLICE_X8Y123_C3 = CLBLM_R_X7Y123_SLICE_X8Y123_BQ;
  assign CLBLM_R_X5Y113_SLICE_X6Y113_B1 = CLBLL_L_X4Y113_SLICE_X4Y113_CO6;
  assign CLBLM_R_X5Y113_SLICE_X6Y113_B2 = CLBLM_R_X5Y113_SLICE_X6Y113_BQ;
  assign CLBLM_R_X5Y113_SLICE_X6Y113_B3 = CLBLM_R_X5Y110_SLICE_X7Y110_BQ;
  assign CLBLM_R_X5Y113_SLICE_X6Y113_B4 = CLBLL_L_X4Y113_SLICE_X4Y113_AQ;
  assign CLBLM_R_X5Y113_SLICE_X6Y113_B5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X5Y113_SLICE_X6Y113_B6 = CLBLM_R_X7Y113_SLICE_X9Y113_BQ;
  assign CLBLM_R_X7Y123_SLICE_X8Y123_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X7Y123_SLICE_X8Y123_D1 = 1'b1;
  assign CLBLM_R_X7Y123_SLICE_X8Y123_D4 = 1'b1;
  assign CLBLM_R_X5Y113_SLICE_X6Y113_C1 = CLBLM_R_X3Y118_SLICE_X2Y118_AQ;
  assign CLBLM_R_X5Y113_SLICE_X6Y113_C2 = CLBLM_R_X5Y113_SLICE_X6Y113_CQ;
  assign CLBLM_R_X5Y113_SLICE_X6Y113_C3 = CLBLM_R_X5Y113_SLICE_X6Y113_AQ;
  assign CLBLM_R_X5Y113_SLICE_X6Y113_C4 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_R_X5Y113_SLICE_X6Y113_C5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X5Y113_SLICE_X6Y113_C6 = CLBLM_L_X8Y113_SLICE_X11Y113_CQ;
  assign CLBLM_R_X7Y123_SLICE_X8Y123_D5 = 1'b1;
  assign CLBLM_R_X7Y123_SLICE_X8Y123_D6 = 1'b1;
  assign CLBLM_R_X5Y113_SLICE_X6Y113_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X5Y113_SLICE_X6Y113_D1 = CLBLL_L_X4Y121_SLICE_X4Y121_AQ;
  assign CLBLM_R_X5Y113_SLICE_X6Y113_D2 = CLBLM_R_X7Y120_SLICE_X9Y120_CQ;
  assign CLBLM_R_X5Y113_SLICE_X6Y113_D3 = CLBLL_L_X4Y114_SLICE_X4Y114_BQ;
  assign CLBLM_R_X5Y113_SLICE_X6Y113_D4 = CLBLM_R_X5Y114_SLICE_X7Y114_AQ;
  assign CLBLM_R_X5Y113_SLICE_X6Y113_D5 = CLBLM_R_X7Y119_SLICE_X8Y119_DQ;
  assign CLBLM_R_X5Y113_SLICE_X6Y113_D6 = 1'b1;
  assign CLBLM_L_X8Y110_SLICE_X10Y110_A1 = CLBLM_R_X5Y111_SLICE_X7Y111_DO6;
  assign LIOB33_X0Y101_IOB_X0Y101_O = CLBLL_L_X2Y111_SLICE_X0Y111_CO6;
  assign LIOB33_X0Y113_IOB_X0Y114_O = CLBLM_R_X5Y117_SLICE_X6Y117_DQ;
  assign LIOB33_X0Y113_IOB_X0Y113_O = RIOB33_X105Y121_IOB_X1Y121_I;
  assign CLBLL_L_X2Y122_SLICE_X0Y122_A1 = RIOB33_X105Y133_IOB_X1Y133_I;
  assign CLBLL_L_X2Y122_SLICE_X0Y122_A2 = RIOB33_X105Y131_IOB_X1Y131_I;
  assign CLBLL_L_X2Y122_SLICE_X0Y122_A3 = RIOB33_X105Y133_IOB_X1Y134_I;
  assign CLBLL_L_X2Y122_SLICE_X0Y122_A4 = CLBLM_R_X3Y124_SLICE_X2Y124_AO6;
  assign CLBLL_L_X2Y122_SLICE_X0Y122_A5 = RIOB33_X105Y131_IOB_X1Y132_I;
  assign CLBLL_L_X2Y122_SLICE_X0Y122_A6 = 1'b1;
  assign CLBLL_L_X2Y122_SLICE_X0Y122_B1 = CLBLL_L_X2Y122_SLICE_X0Y122_DO6;
  assign CLBLL_L_X2Y122_SLICE_X0Y122_B2 = CLBLL_L_X2Y122_SLICE_X1Y122_BO6;
  assign CLBLL_L_X2Y122_SLICE_X0Y122_B3 = CLBLL_L_X2Y123_SLICE_X0Y123_AO6;
  assign CLBLL_L_X2Y122_SLICE_X0Y122_B4 = CLBLL_L_X4Y122_SLICE_X5Y122_BO6;
  assign CLBLL_L_X2Y122_SLICE_X0Y122_B5 = CLBLM_R_X5Y122_SLICE_X6Y122_CO6;
  assign CLBLL_L_X2Y122_SLICE_X0Y122_B6 = CLBLL_L_X2Y121_SLICE_X0Y121_CO6;
  assign CLBLM_R_X103Y169_SLICE_X163Y169_A6 = 1'b1;
  assign CLBLM_L_X8Y110_SLICE_X10Y110_B3 = CLBLM_L_X8Y118_SLICE_X10Y118_DQ;
  assign RIOI3_X105Y117_ILOGIC_X1Y117_D = RIOB33_X105Y117_IOB_X1Y117_I;
  assign CLBLL_L_X2Y122_SLICE_X0Y122_C1 = RIOB33_X105Y113_IOB_X1Y114_I;
  assign CLBLL_L_X2Y122_SLICE_X0Y122_C2 = CLBLL_L_X2Y121_SLICE_X0Y121_CO6;
  assign CLBLL_L_X2Y122_SLICE_X0Y122_C3 = CLBLL_L_X2Y122_SLICE_X1Y122_BO6;
  assign CLBLL_L_X2Y122_SLICE_X0Y122_C4 = CLBLL_L_X2Y122_SLICE_X0Y122_AO5;
  assign CLBLL_L_X2Y122_SLICE_X0Y122_C5 = CLBLL_L_X2Y122_SLICE_X0Y122_DO6;
  assign CLBLL_L_X2Y122_SLICE_X0Y122_C6 = CLBLL_L_X4Y122_SLICE_X5Y122_BO6;
  assign CLBLL_L_X2Y122_SLICE_X0Y122_D1 = CLBLL_L_X2Y121_SLICE_X0Y121_BO6;
  assign CLBLL_L_X2Y122_SLICE_X0Y122_D2 = LIOB33_X0Y69_IOB_X0Y70_I;
  assign CLBLL_L_X2Y122_SLICE_X0Y122_D3 = CLBLL_L_X2Y117_SLICE_X0Y117_CQ;
  assign CLBLL_L_X2Y122_SLICE_X0Y122_D4 = CLBLM_R_X3Y124_SLICE_X2Y124_AO5;
  assign CLBLL_L_X2Y122_SLICE_X0Y122_D5 = CLBLL_L_X2Y120_SLICE_X1Y120_AO6;
  assign CLBLL_L_X2Y122_SLICE_X0Y122_D6 = 1'b1;
  assign LIOB33_X0Y191_IOB_X0Y192_O = LIOB33_X0Y51_IOB_X0Y52_I;
  assign LIOB33_X0Y191_IOB_X0Y191_O = RIOB33_X105Y147_IOB_X1Y148_I;
  assign RIOB33_X105Y195_IOB_X1Y195_O = CLBLM_R_X11Y119_SLICE_X14Y119_AQ;
  assign RIOB33_X105Y173_IOB_X1Y174_O = CLBLM_R_X103Y174_SLICE_X163Y174_AO6;
  assign CLBLL_L_X2Y122_SLICE_X1Y122_A1 = CLBLL_L_X2Y122_SLICE_X1Y122_DO6;
  assign CLBLL_L_X2Y122_SLICE_X1Y122_A2 = LIOB33_X0Y71_IOB_X0Y71_I;
  assign CLBLL_L_X2Y122_SLICE_X1Y122_A3 = RIOB33_X105Y131_IOB_X1Y132_I;
  assign CLBLL_L_X2Y122_SLICE_X1Y122_A4 = RIOB33_X105Y131_IOB_X1Y131_I;
  assign CLBLL_L_X2Y122_SLICE_X1Y122_A5 = LIOB33_X0Y61_IOB_X0Y61_I;
  assign CLBLL_L_X2Y122_SLICE_X1Y122_A6 = CLBLM_R_X3Y124_SLICE_X2Y124_AO5;
  assign RIOI3_X105Y177_OLOGIC_X1Y178_D1 = CLBLM_R_X103Y177_SLICE_X163Y177_AO5;
  assign CLBLM_R_X103Y169_SLICE_X163Y169_A1 = CLBLM_L_X10Y114_SLICE_X12Y114_AQ;
  assign CLBLM_R_X103Y169_SLICE_X163Y169_A2 = 1'b1;
  assign CLBLL_L_X2Y122_SLICE_X1Y122_B1 = CLBLM_R_X3Y124_SLICE_X2Y124_AO5;
  assign CLBLL_L_X2Y122_SLICE_X1Y122_B2 = CLBLL_L_X2Y121_SLICE_X1Y121_BO5;
  assign CLBLL_L_X2Y122_SLICE_X1Y122_B3 = 1'b1;
  assign CLBLL_L_X2Y122_SLICE_X1Y122_B4 = CLBLL_L_X2Y121_SLICE_X1Y121_BO6;
  assign CLBLL_L_X2Y122_SLICE_X1Y122_B5 = CLBLM_R_X5Y122_SLICE_X7Y122_DQ;
  assign CLBLL_L_X2Y122_SLICE_X1Y122_B6 = LIOB33_X0Y59_IOB_X0Y59_I;
  assign CLBLM_R_X103Y169_SLICE_X163Y169_A3 = RIOB33_X105Y143_IOB_X1Y143_I;
  assign CLBLM_R_X103Y169_SLICE_X163Y169_A4 = 1'b1;
  assign CLBLM_R_X103Y169_SLICE_X163Y169_A5 = CLBLM_R_X11Y122_SLICE_X14Y122_AQ;
  assign CLBLL_L_X2Y122_SLICE_X1Y122_C1 = 1'b1;
  assign CLBLL_L_X2Y122_SLICE_X1Y122_C2 = CLBLL_L_X2Y121_SLICE_X1Y121_BO5;
  assign CLBLL_L_X2Y122_SLICE_X1Y122_C3 = LIOB33_X0Y63_IOB_X0Y63_I;
  assign CLBLL_L_X2Y122_SLICE_X1Y122_C4 = CLBLM_R_X3Y124_SLICE_X2Y124_AO5;
  assign CLBLL_L_X2Y122_SLICE_X1Y122_C5 = CLBLM_R_X3Y116_SLICE_X3Y116_CQ;
  assign CLBLL_L_X2Y122_SLICE_X1Y122_C6 = CLBLL_L_X2Y121_SLICE_X1Y121_BO6;
  assign CLBLM_R_X103Y169_SLICE_X163Y169_B2 = 1'b1;
  assign CLBLM_R_X103Y169_SLICE_X163Y169_B3 = 1'b1;
  assign CLBLM_R_X103Y169_SLICE_X163Y169_B4 = 1'b1;
  assign CLBLM_R_X103Y169_SLICE_X163Y169_B5 = 1'b1;
  assign CLBLM_R_X103Y169_SLICE_X163Y169_B6 = 1'b1;
  assign CLBLM_R_X103Y169_SLICE_X163Y169_C1 = 1'b1;
  assign CLBLL_L_X2Y122_SLICE_X1Y122_D1 = 1'b1;
  assign CLBLL_L_X2Y122_SLICE_X1Y122_D2 = RIOB33_X105Y133_IOB_X1Y133_I;
  assign CLBLL_L_X2Y122_SLICE_X1Y122_D3 = 1'b1;
  assign CLBLL_L_X2Y122_SLICE_X1Y122_D4 = RIOB33_X105Y133_IOB_X1Y134_I;
  assign CLBLL_L_X2Y122_SLICE_X1Y122_D5 = 1'b1;
  assign CLBLL_L_X2Y122_SLICE_X1Y122_D6 = 1'b1;
  assign CLBLM_R_X103Y169_SLICE_X163Y169_C6 = 1'b1;
  assign CLBLM_R_X103Y169_SLICE_X163Y169_D1 = 1'b1;
  assign CLBLM_R_X103Y169_SLICE_X163Y169_D2 = 1'b1;
  assign CLBLM_R_X103Y169_SLICE_X163Y169_D3 = 1'b1;
  assign CLBLM_R_X103Y169_SLICE_X163Y169_D4 = 1'b1;
  assign CLBLM_R_X103Y169_SLICE_X163Y169_D5 = 1'b1;
  assign CLBLM_R_X103Y169_SLICE_X163Y169_D6 = 1'b1;
  assign CLBLM_R_X103Y169_SLICE_X162Y169_A1 = 1'b1;
  assign CLBLM_R_X103Y169_SLICE_X162Y169_A2 = 1'b1;
  assign CLBLM_R_X103Y169_SLICE_X162Y169_A3 = 1'b1;
  assign CLBLM_R_X103Y169_SLICE_X162Y169_A4 = 1'b1;
  assign CLBLM_R_X103Y169_SLICE_X162Y169_A5 = 1'b1;
  assign CLBLM_R_X103Y169_SLICE_X162Y169_A6 = 1'b1;
  assign CLBLM_R_X103Y169_SLICE_X162Y169_B1 = 1'b1;
  assign CLBLM_R_X103Y169_SLICE_X162Y169_B2 = 1'b1;
  assign CLBLM_R_X103Y169_SLICE_X162Y169_B3 = 1'b1;
  assign CLBLM_R_X103Y169_SLICE_X162Y169_B4 = 1'b1;
  assign CLBLM_R_X103Y169_SLICE_X162Y169_B5 = 1'b1;
  assign CLBLM_R_X103Y169_SLICE_X162Y169_B6 = 1'b1;
  assign CLBLM_R_X103Y169_SLICE_X163Y169_B1 = 1'b1;
  assign CLBLM_R_X103Y169_SLICE_X162Y169_C1 = 1'b1;
  assign CLBLM_R_X103Y169_SLICE_X162Y169_C2 = 1'b1;
  assign CLBLM_R_X103Y169_SLICE_X162Y169_C3 = 1'b1;
  assign CLBLM_R_X7Y124_SLICE_X9Y124_A1 = CLBLM_R_X7Y123_SLICE_X9Y123_DO6;
  assign CLBLM_R_X7Y124_SLICE_X9Y124_A2 = 1'b1;
  assign CLBLM_R_X7Y124_SLICE_X9Y124_A3 = CLBLM_R_X7Y124_SLICE_X9Y124_AQ;
  assign CLBLM_R_X7Y124_SLICE_X9Y124_A4 = CLBLM_R_X5Y114_SLICE_X6Y114_BQ;
  assign CLBLM_R_X7Y124_SLICE_X9Y124_A5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y124_SLICE_X9Y124_A6 = CLBLM_L_X10Y123_SLICE_X12Y123_AO6;
  assign CLBLM_R_X103Y169_SLICE_X162Y169_C4 = 1'b1;
  assign CLBLM_R_X103Y169_SLICE_X162Y169_C5 = 1'b1;
  assign CLBLM_R_X103Y169_SLICE_X162Y169_C6 = 1'b1;
  assign CLBLM_R_X7Y124_SLICE_X9Y124_B1 = 1'b1;
  assign CLBLM_R_X7Y124_SLICE_X9Y124_B2 = 1'b1;
  assign CLBLM_R_X7Y124_SLICE_X9Y124_B3 = 1'b1;
  assign CLBLM_R_X7Y124_SLICE_X9Y124_B4 = 1'b1;
  assign CLBLM_R_X7Y124_SLICE_X9Y124_B5 = 1'b1;
  assign CLBLM_R_X7Y124_SLICE_X9Y124_B6 = 1'b1;
  assign CLBLM_R_X103Y169_SLICE_X162Y169_D1 = 1'b1;
  assign CLBLM_R_X103Y169_SLICE_X162Y169_D2 = 1'b1;
  assign CLBLM_R_X5Y114_SLICE_X7Y114_A1 = CLBLM_R_X5Y114_SLICE_X7Y114_AQ;
  assign CLBLM_R_X5Y114_SLICE_X7Y114_A2 = CLBLL_L_X4Y111_SLICE_X4Y111_DQ;
  assign CLBLM_R_X5Y114_SLICE_X7Y114_A3 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X5Y114_SLICE_X7Y114_A4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X5Y114_SLICE_X7Y114_A5 = 1'b1;
  assign CLBLM_R_X5Y114_SLICE_X7Y114_A6 = CLBLL_L_X4Y115_SLICE_X4Y115_CQ;
  assign CLBLM_R_X7Y124_SLICE_X9Y124_C1 = 1'b1;
  assign CLBLM_R_X7Y124_SLICE_X9Y124_C2 = 1'b1;
  assign CLBLM_R_X7Y124_SLICE_X9Y124_C3 = 1'b1;
  assign CLBLM_R_X5Y114_SLICE_X7Y114_B1 = 1'b1;
  assign CLBLM_R_X5Y114_SLICE_X7Y114_B2 = CLBLL_L_X4Y114_SLICE_X4Y114_BQ;
  assign CLBLM_R_X5Y114_SLICE_X7Y114_B3 = 1'b1;
  assign CLBLM_R_X5Y114_SLICE_X7Y114_B4 = 1'b1;
  assign CLBLM_R_X5Y114_SLICE_X7Y114_B5 = CLBLL_L_X4Y121_SLICE_X4Y121_AQ;
  assign CLBLM_R_X5Y114_SLICE_X7Y114_B6 = 1'b1;
  assign CLBLM_R_X7Y124_SLICE_X9Y124_D1 = 1'b1;
  assign CLBLM_R_X5Y114_SLICE_X7Y114_C1 = CLBLL_L_X4Y120_SLICE_X4Y120_BO6;
  assign CLBLM_R_X5Y114_SLICE_X7Y114_C2 = CLBLM_R_X5Y112_SLICE_X7Y112_AO5;
  assign CLBLM_R_X5Y114_SLICE_X7Y114_C3 = CLBLM_R_X5Y112_SLICE_X7Y112_DO6;
  assign CLBLM_R_X5Y114_SLICE_X7Y114_C4 = CLBLM_R_X7Y115_SLICE_X8Y115_CQ;
  assign CLBLM_R_X5Y114_SLICE_X7Y114_C5 = CLBLM_R_X3Y114_SLICE_X3Y114_AQ;
  assign CLBLM_R_X5Y114_SLICE_X7Y114_C6 = RIOB33_X105Y121_IOB_X1Y121_I;
  assign CLBLM_R_X7Y124_SLICE_X9Y124_D3 = 1'b1;
  assign CLBLM_R_X7Y124_SLICE_X9Y124_D4 = 1'b1;
  assign CLBLM_R_X5Y114_SLICE_X7Y114_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X7Y124_SLICE_X8Y124_A1 = CLBLM_R_X5Y124_SLICE_X6Y124_AQ;
  assign CLBLM_R_X7Y124_SLICE_X8Y124_A2 = RIOB33_X105Y121_IOB_X1Y121_I;
  assign CLBLM_R_X7Y124_SLICE_X8Y124_A3 = CLBLM_R_X7Y124_SLICE_X8Y124_AQ;
  assign CLBLM_R_X7Y124_SLICE_X8Y124_A4 = CLBLM_R_X7Y120_SLICE_X9Y120_A5Q;
  assign CLBLM_R_X7Y124_SLICE_X8Y124_A5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X5Y114_SLICE_X7Y114_D1 = CLBLM_R_X5Y121_SLICE_X7Y121_AQ;
  assign CLBLM_R_X5Y114_SLICE_X7Y114_D2 = CLBLM_R_X7Y120_SLICE_X9Y120_CQ;
  assign CLBLM_R_X5Y114_SLICE_X7Y114_D3 = RIOB33_X105Y121_IOB_X1Y121_I;
  assign CLBLM_R_X5Y114_SLICE_X7Y114_D4 = CLBLM_R_X7Y115_SLICE_X8Y115_CQ;
  assign CLBLM_R_X5Y114_SLICE_X7Y114_D5 = CLBLM_R_X5Y114_SLICE_X7Y114_AQ;
  assign CLBLM_R_X5Y114_SLICE_X7Y114_D6 = CLBLM_R_X5Y114_SLICE_X7Y114_BO6;
  assign CLBLM_R_X7Y124_SLICE_X8Y124_A6 = CLBLM_L_X10Y123_SLICE_X13Y123_DO6;
  assign CLBLM_R_X7Y124_SLICE_X8Y124_AX = CLBLM_R_X7Y124_SLICE_X8Y124_DO6;
  assign CLBLM_R_X7Y124_SLICE_X8Y124_B1 = CLBLL_L_X4Y119_SLICE_X4Y119_C5Q;
  assign CLBLM_R_X7Y124_SLICE_X8Y124_B2 = CLBLM_R_X7Y124_SLICE_X8Y124_BQ;
  assign CLBLM_R_X7Y124_SLICE_X8Y124_B3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y124_SLICE_X8Y124_B4 = CLBLM_R_X7Y116_SLICE_X8Y116_CQ;
  assign CLBLM_R_X5Y114_SLICE_X6Y114_A1 = CLBLL_L_X4Y119_SLICE_X4Y119_B5Q;
  assign CLBLM_R_X5Y114_SLICE_X6Y114_A2 = CLBLM_R_X5Y113_SLICE_X6Y113_CQ;
  assign CLBLM_R_X5Y114_SLICE_X6Y114_A3 = CLBLM_R_X5Y114_SLICE_X6Y114_AQ;
  assign CLBLM_R_X5Y114_SLICE_X6Y114_A4 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_R_X5Y114_SLICE_X6Y114_A5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X5Y114_SLICE_X6Y114_A6 = CLBLM_R_X3Y118_SLICE_X2Y118_AQ;
  assign CLBLM_R_X7Y124_SLICE_X8Y124_C1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y124_SLICE_X8Y124_C2 = CLBLM_R_X7Y124_SLICE_X8Y124_CQ;
  assign CLBLM_R_X7Y124_SLICE_X8Y124_C3 = CLBLL_L_X4Y119_SLICE_X4Y119_C5Q;
  assign CLBLM_R_X5Y114_SLICE_X6Y114_B1 = 1'b1;
  assign CLBLM_R_X5Y114_SLICE_X6Y114_B2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X5Y114_SLICE_X6Y114_B3 = CLBLL_L_X4Y111_SLICE_X4Y111_CQ;
  assign CLBLM_R_X5Y114_SLICE_X6Y114_B4 = CLBLM_R_X5Y118_SLICE_X6Y118_BQ;
  assign CLBLM_R_X5Y114_SLICE_X6Y114_B5 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X5Y114_SLICE_X6Y114_B6 = CLBLL_L_X4Y114_SLICE_X4Y114_DO6;
  assign CLBLM_R_X7Y124_SLICE_X8Y124_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X7Y124_SLICE_X8Y124_D1 = CLBLM_R_X7Y124_SLICE_X9Y124_AQ;
  assign CLBLM_R_X7Y124_SLICE_X8Y124_D2 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X5Y114_SLICE_X6Y114_C1 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X5Y114_SLICE_X6Y114_C2 = CLBLM_R_X7Y115_SLICE_X8Y115_BQ;
  assign CLBLL_L_X4Y122_SLICE_X5Y122_C1 = CLBLM_R_X3Y124_SLICE_X2Y124_BO6;
  assign CLBLM_R_X5Y114_SLICE_X6Y114_C3 = 1'b1;
  assign CLBLM_R_X5Y114_SLICE_X6Y114_C4 = CLBLM_R_X5Y112_SLICE_X6Y112_BO5;
  assign CLBLM_R_X5Y114_SLICE_X6Y114_C5 = CLBLM_R_X5Y117_SLICE_X6Y117_CQ;
  assign CLBLM_R_X5Y114_SLICE_X6Y114_C6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y124_SLICE_X8Y124_D3 = CLBLL_L_X4Y119_SLICE_X4Y119_C5Q;
  assign CLBLM_R_X7Y124_SLICE_X8Y124_D4 = CLBLM_R_X7Y124_SLICE_X8Y124_A5Q;
  assign CLBLM_R_X5Y114_SLICE_X6Y114_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X7Y124_SLICE_X8Y124_D6 = 1'b1;
  assign CLBLM_R_X5Y114_SLICE_X6Y114_D1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X5Y114_SLICE_X6Y114_D2 = CLBLM_L_X10Y115_SLICE_X12Y115_BQ;
  assign CLBLM_R_X5Y114_SLICE_X6Y114_D3 = CLBLM_R_X5Y114_SLICE_X6Y114_DQ;
  assign CLBLM_R_X5Y114_SLICE_X6Y114_D4 = 1'b1;
  assign CLBLM_R_X5Y114_SLICE_X6Y114_D5 = CLBLL_L_X4Y114_SLICE_X4Y114_CQ;
  assign CLBLM_R_X5Y114_SLICE_X6Y114_D6 = CLBLM_R_X5Y111_SLICE_X7Y111_DO6;
  assign LIOB33_X0Y115_IOB_X0Y115_O = CLBLM_R_X11Y114_SLICE_X14Y114_DQ;
  assign LIOB33_X0Y115_IOB_X0Y116_O = CLBLM_L_X8Y123_SLICE_X11Y123_AQ;
  assign LIOB33_SING_X0Y149_IOB_X0Y149_O = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLL_L_X2Y123_SLICE_X0Y123_A1 = RIOB33_X105Y113_IOB_X1Y114_I;
  assign CLBLL_L_X2Y123_SLICE_X0Y123_A2 = CLBLM_R_X3Y124_SLICE_X2Y124_AO6;
  assign CLBLL_L_X2Y123_SLICE_X0Y123_A3 = RIOB33_X105Y133_IOB_X1Y133_I;
  assign CLBLL_L_X2Y123_SLICE_X0Y123_A4 = RIOB33_X105Y133_IOB_X1Y134_I;
  assign CLBLL_L_X2Y123_SLICE_X0Y123_A5 = RIOB33_X105Y131_IOB_X1Y131_I;
  assign CLBLL_L_X2Y123_SLICE_X0Y123_A6 = RIOB33_X105Y131_IOB_X1Y132_I;
  assign CLBLL_L_X2Y123_SLICE_X0Y123_B1 = 1'b1;
  assign CLBLL_L_X2Y123_SLICE_X0Y123_B2 = 1'b1;
  assign CLBLL_L_X2Y123_SLICE_X0Y123_B3 = 1'b1;
  assign CLBLL_L_X2Y123_SLICE_X0Y123_B4 = 1'b1;
  assign CLBLL_L_X2Y123_SLICE_X0Y123_B5 = 1'b1;
  assign CLBLL_L_X2Y123_SLICE_X0Y123_B6 = 1'b1;
  assign CLBLL_L_X2Y123_SLICE_X0Y123_C1 = 1'b1;
  assign CLBLL_L_X2Y123_SLICE_X0Y123_C2 = 1'b1;
  assign CLBLL_L_X2Y123_SLICE_X0Y123_C3 = 1'b1;
  assign CLBLL_L_X2Y123_SLICE_X0Y123_C4 = 1'b1;
  assign CLBLL_L_X2Y123_SLICE_X0Y123_C5 = 1'b1;
  assign CLBLL_L_X2Y123_SLICE_X0Y123_C6 = 1'b1;
  assign CLBLL_L_X2Y123_SLICE_X0Y123_D1 = 1'b1;
  assign CLBLL_L_X2Y123_SLICE_X0Y123_D2 = 1'b1;
  assign CLBLL_L_X2Y123_SLICE_X0Y123_D3 = 1'b1;
  assign CLBLL_L_X2Y123_SLICE_X0Y123_D4 = 1'b1;
  assign CLBLL_L_X2Y123_SLICE_X0Y123_D5 = 1'b1;
  assign CLBLL_L_X2Y123_SLICE_X0Y123_D6 = 1'b1;
  assign RIOI3_X105Y177_OLOGIC_X1Y178_T1 = 1'b1;
  assign CLBLL_L_X2Y123_SLICE_X1Y123_A1 = 1'b1;
  assign CLBLL_L_X2Y123_SLICE_X1Y123_A2 = 1'b1;
  assign CLBLL_L_X2Y123_SLICE_X1Y123_A3 = 1'b1;
  assign CLBLL_L_X2Y123_SLICE_X1Y123_A4 = 1'b1;
  assign CLBLL_L_X2Y123_SLICE_X1Y123_A5 = 1'b1;
  assign CLBLL_L_X2Y123_SLICE_X1Y123_A6 = 1'b1;
  assign CLBLL_L_X2Y123_SLICE_X1Y123_B1 = 1'b1;
  assign CLBLL_L_X2Y123_SLICE_X1Y123_B2 = 1'b1;
  assign CLBLL_L_X2Y123_SLICE_X1Y123_B3 = 1'b1;
  assign CLBLL_L_X2Y123_SLICE_X1Y123_B4 = 1'b1;
  assign CLBLL_L_X2Y123_SLICE_X1Y123_B5 = 1'b1;
  assign CLBLL_L_X2Y123_SLICE_X1Y123_B6 = 1'b1;
  assign CLBLL_L_X2Y123_SLICE_X1Y123_C1 = 1'b1;
  assign CLBLL_L_X2Y123_SLICE_X1Y123_C2 = 1'b1;
  assign CLBLL_L_X2Y123_SLICE_X1Y123_C3 = 1'b1;
  assign CLBLL_L_X2Y123_SLICE_X1Y123_C4 = 1'b1;
  assign CLBLL_L_X2Y123_SLICE_X1Y123_C5 = 1'b1;
  assign CLBLL_L_X2Y123_SLICE_X1Y123_C6 = 1'b1;
  assign LIOI3_X0Y139_OLOGIC_X0Y140_D1 = CLBLL_L_X4Y123_SLICE_X4Y123_BQ;
  assign LIOI3_X0Y175_OLOGIC_X0Y175_D1 = RIOB33_X105Y127_IOB_X1Y127_I;
  assign CLBLL_L_X2Y123_SLICE_X1Y123_D1 = 1'b1;
  assign CLBLL_L_X2Y123_SLICE_X1Y123_D2 = 1'b1;
  assign CLBLL_L_X2Y123_SLICE_X1Y123_D3 = 1'b1;
  assign CLBLL_L_X2Y123_SLICE_X1Y123_D4 = 1'b1;
  assign CLBLL_L_X2Y123_SLICE_X1Y123_D5 = 1'b1;
  assign CLBLL_L_X2Y123_SLICE_X1Y123_D6 = 1'b1;
  assign CLBLM_R_X103Y169_SLICE_X163Y169_C2 = 1'b1;
  assign LIOI3_X0Y139_OLOGIC_X0Y140_T1 = 1'b1;
  assign RIOI3_X105Y183_OLOGIC_X1Y184_D1 = CLBLM_R_X11Y117_SLICE_X14Y117_DO5;
  assign LIOI3_X0Y139_OLOGIC_X0Y139_D1 = CLBLM_R_X5Y124_SLICE_X6Y124_AQ;
  assign RIOI3_X105Y183_OLOGIC_X1Y184_T1 = 1'b1;
  assign LIOI3_X0Y139_OLOGIC_X0Y139_T1 = 1'b1;
  assign CLBLM_R_X103Y169_SLICE_X163Y169_C3 = 1'b1;
  assign RIOI3_X105Y183_OLOGIC_X1Y183_D1 = CLBLM_R_X11Y117_SLICE_X14Y117_DO6;
  assign LIOB33_SING_X0Y150_IOB_X0Y150_O = LIOB33_X0Y63_IOB_X0Y63_I;
  assign LIOI3_TBYTESRC_X0Y181_OLOGIC_X0Y182_D1 = RIOB33_X105Y133_IOB_X1Y134_I;
  assign RIOI3_X105Y183_OLOGIC_X1Y183_T1 = 1'b1;
  assign LIOI3_TBYTESRC_X0Y107_OLOGIC_X0Y108_T1 = 1'b1;
  assign CLBLM_R_X7Y125_SLICE_X9Y125_A1 = 1'b1;
  assign CLBLM_R_X7Y125_SLICE_X9Y125_A2 = 1'b1;
  assign CLBLM_R_X7Y125_SLICE_X9Y125_A3 = 1'b1;
  assign CLBLM_R_X7Y125_SLICE_X9Y125_A4 = 1'b1;
  assign CLBLM_R_X7Y125_SLICE_X9Y125_A5 = 1'b1;
  assign CLBLM_R_X7Y125_SLICE_X9Y125_A6 = 1'b1;
  assign CLBLM_R_X103Y169_SLICE_X163Y169_C4 = 1'b1;
  assign LIOI3_TBYTESRC_X0Y181_OLOGIC_X0Y182_T1 = 1'b1;
  assign CLBLM_R_X7Y125_SLICE_X9Y125_B1 = 1'b1;
  assign CLBLM_R_X7Y125_SLICE_X9Y125_B2 = 1'b1;
  assign CLBLM_R_X7Y125_SLICE_X9Y125_B3 = 1'b1;
  assign CLBLM_R_X7Y125_SLICE_X9Y125_B4 = 1'b1;
  assign CLBLM_R_X7Y125_SLICE_X9Y125_B5 = 1'b1;
  assign CLBLM_R_X7Y125_SLICE_X9Y125_B6 = 1'b1;
  assign LIOI3_TBYTESRC_X0Y181_OLOGIC_X0Y181_D1 = RIOB33_X105Y133_IOB_X1Y133_I;
  assign CLBLM_R_X5Y115_SLICE_X7Y115_A1 = CLBLM_R_X7Y115_SLICE_X9Y115_CQ;
  assign CLBLM_R_X5Y115_SLICE_X7Y115_A2 = CLBLM_L_X8Y117_SLICE_X11Y117_AQ;
  assign CLBLM_R_X5Y115_SLICE_X7Y115_A3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X5Y115_SLICE_X7Y115_A4 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X5Y115_SLICE_X7Y115_A5 = CLBLM_R_X5Y115_SLICE_X7Y115_A5Q;
  assign CLBLM_R_X5Y115_SLICE_X7Y115_A6 = 1'b1;
  assign CLBLM_R_X7Y125_SLICE_X9Y125_C1 = 1'b1;
  assign CLBLM_R_X7Y125_SLICE_X9Y125_C2 = 1'b1;
  assign CLBLM_R_X7Y125_SLICE_X9Y125_C3 = 1'b1;
  assign CLBLM_R_X5Y115_SLICE_X7Y115_B1 = CLBLM_R_X5Y110_SLICE_X7Y110_AQ;
  assign CLBLM_R_X5Y115_SLICE_X7Y115_B2 = 1'b1;
  assign CLBLM_R_X5Y115_SLICE_X7Y115_B3 = CLBLM_R_X5Y119_SLICE_X6Y119_BQ;
  assign CLBLM_R_X5Y115_SLICE_X7Y115_B4 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X5Y115_SLICE_X7Y115_B5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X5Y115_SLICE_X7Y115_B6 = 1'b1;
  assign CLBLM_R_X7Y125_SLICE_X9Y125_D1 = 1'b1;
  assign CLBLM_R_X7Y125_SLICE_X9Y125_D2 = 1'b1;
  assign CLBLM_R_X5Y115_SLICE_X7Y115_C1 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X5Y115_SLICE_X7Y115_C2 = CLBLM_R_X5Y116_SLICE_X7Y116_CQ;
  assign CLBLM_R_X5Y115_SLICE_X7Y115_C3 = CLBLM_R_X7Y109_SLICE_X8Y109_AQ;
  assign CLBLM_R_X5Y115_SLICE_X7Y115_C4 = CLBLL_L_X4Y113_SLICE_X5Y113_DO6;
  assign CLBLM_R_X5Y115_SLICE_X7Y115_C5 = CLBLL_L_X2Y119_SLICE_X0Y119_BO6;
  assign CLBLM_R_X5Y115_SLICE_X7Y115_C6 = 1'b1;
  assign CLBLM_R_X7Y125_SLICE_X9Y125_D3 = 1'b1;
  assign CLBLM_R_X7Y125_SLICE_X9Y125_D4 = 1'b1;
  assign CLBLM_R_X5Y115_SLICE_X7Y115_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X7Y125_SLICE_X8Y125_A1 = 1'b1;
  assign CLBLM_R_X7Y125_SLICE_X8Y125_A2 = CLBLM_R_X7Y124_SLICE_X8Y124_A5Q;
  assign CLBLM_R_X7Y125_SLICE_X8Y125_A3 = 1'b1;
  assign CLBLM_R_X7Y125_SLICE_X8Y125_A4 = CLBLL_L_X4Y123_SLICE_X4Y123_AQ;
  assign CLBLM_R_X7Y125_SLICE_X8Y125_A5 = CLBLM_R_X7Y124_SLICE_X8Y124_BQ;
  assign CLBLM_R_X5Y115_SLICE_X7Y115_D1 = CLBLM_R_X5Y115_SLICE_X7Y115_CO5;
  assign CLBLM_R_X5Y115_SLICE_X7Y115_D2 = CLBLM_L_X8Y114_SLICE_X10Y114_C5Q;
  assign CLBLM_R_X5Y115_SLICE_X7Y115_D3 = CLBLL_L_X4Y115_SLICE_X5Y115_AQ;
  assign CLBLM_R_X5Y115_SLICE_X7Y115_D4 = RIOB33_X105Y121_IOB_X1Y121_I;
  assign CLBLM_R_X5Y115_SLICE_X7Y115_D5 = CLBLM_R_X5Y112_SLICE_X7Y112_AO5;
  assign CLBLM_R_X5Y115_SLICE_X7Y115_D6 = CLBLL_L_X2Y120_SLICE_X0Y120_CO6;
  assign CLBLM_R_X7Y125_SLICE_X8Y125_A6 = 1'b1;
  assign CLBLM_R_X7Y125_SLICE_X8Y125_B1 = 1'b1;
  assign CLBLM_R_X7Y125_SLICE_X8Y125_B2 = 1'b1;
  assign CLBLM_R_X7Y125_SLICE_X8Y125_B3 = 1'b1;
  assign CLBLM_R_X7Y125_SLICE_X8Y125_B4 = 1'b1;
  assign CLBLM_R_X5Y115_SLICE_X6Y115_A1 = CLBLM_R_X7Y115_SLICE_X9Y115_DQ;
  assign CLBLM_R_X5Y115_SLICE_X6Y115_A2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X5Y115_SLICE_X6Y115_A3 = CLBLM_R_X5Y115_SLICE_X6Y115_AQ;
  assign CLBLM_R_X5Y115_SLICE_X6Y115_A4 = CLBLM_R_X7Y115_SLICE_X8Y115_BQ;
  assign CLBLM_R_X5Y115_SLICE_X6Y115_A5 = CLBLM_R_X5Y115_SLICE_X6Y115_CO5;
  assign CLBLM_R_X5Y115_SLICE_X6Y115_A6 = 1'b1;
  assign CLBLM_R_X7Y125_SLICE_X8Y125_C1 = 1'b1;
  assign CLBLM_R_X7Y125_SLICE_X8Y125_C2 = 1'b1;
  assign CLBLM_R_X7Y125_SLICE_X8Y125_C3 = 1'b1;
  assign CLBLM_R_X5Y115_SLICE_X6Y115_B1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X5Y115_SLICE_X6Y115_B2 = CLBLM_L_X8Y115_SLICE_X11Y115_C5Q;
  assign CLBLM_R_X5Y115_SLICE_X6Y115_B3 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X5Y115_SLICE_X6Y115_B4 = 1'b1;
  assign CLBLM_R_X5Y115_SLICE_X6Y115_B5 = CLBLM_R_X7Y113_SLICE_X8Y113_AQ;
  assign CLBLM_R_X5Y115_SLICE_X6Y115_B6 = CLBLM_R_X7Y115_SLICE_X8Y115_DO6;
  assign CLBLM_R_X7Y125_SLICE_X8Y125_D1 = 1'b1;
  assign CLBLM_R_X7Y125_SLICE_X8Y125_D2 = 1'b1;
  assign CLBLM_R_X7Y125_SLICE_X8Y125_D3 = 1'b1;
  assign CLBLM_R_X5Y115_SLICE_X6Y115_C1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X5Y115_SLICE_X6Y115_C2 = CLBLM_R_X5Y121_SLICE_X6Y121_AQ;
  assign CLBLM_R_X5Y115_SLICE_X6Y115_C3 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X5Y115_SLICE_X6Y115_C4 = CLBLM_R_X7Y114_SLICE_X8Y114_BQ;
  assign CLBLM_R_X5Y115_SLICE_X6Y115_C5 = RIOB33_X105Y121_IOB_X1Y121_I;
  assign CLBLM_R_X5Y115_SLICE_X6Y115_C6 = 1'b1;
  assign CLBLM_R_X7Y125_SLICE_X8Y125_D4 = 1'b1;
  assign CLBLM_R_X7Y125_SLICE_X8Y125_D5 = 1'b1;
  assign CLBLM_R_X7Y125_SLICE_X8Y125_D6 = 1'b1;
  assign CLBLM_R_X5Y115_SLICE_X6Y115_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign RIOI3_TBYTETERM_X105Y113_ILOGIC_X1Y113_D = RIOB33_X105Y113_IOB_X1Y113_I;
  assign CLBLM_R_X5Y115_SLICE_X6Y115_D1 = CLBLL_L_X4Y115_SLICE_X4Y115_DQ;
  assign CLBLM_R_X5Y115_SLICE_X6Y115_D2 = CLBLM_R_X5Y114_SLICE_X6Y114_CQ;
  assign CLBLM_R_X5Y115_SLICE_X6Y115_D3 = CLBLM_R_X7Y116_SLICE_X8Y116_BQ;
  assign CLBLM_R_X5Y115_SLICE_X6Y115_D4 = CLBLL_L_X4Y115_SLICE_X5Y115_BQ;
  assign CLBLM_R_X5Y115_SLICE_X6Y115_D5 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X5Y115_SLICE_X6Y115_D6 = CLBLM_R_X7Y115_SLICE_X8Y115_BQ;
  assign LIOB33_SING_X0Y199_IOB_X0Y199_O = LIOB33_X0Y73_IOB_X0Y74_I;
  assign LIOB33_X0Y121_IOB_X0Y122_O = CLBLM_R_X5Y121_SLICE_X6Y121_A5Q;
  assign LIOB33_X0Y121_IOB_X0Y121_O = CLBLM_L_X8Y123_SLICE_X11Y123_A5Q;
  assign LIOI3_X0Y77_ILOGIC_X0Y78_D = LIOB33_X0Y77_IOB_X0Y78_I;
  assign LIOI3_X0Y77_ILOGIC_X0Y77_D = LIOB33_X0Y77_IOB_X0Y77_I;
  assign RIOI3_X105Y123_ILOGIC_X1Y124_D = RIOB33_X105Y123_IOB_X1Y124_I;
  assign RIOI3_X105Y123_ILOGIC_X1Y123_D = RIOB33_X105Y123_IOB_X1Y123_I;
  assign CLBLM_R_X7Y127_SLICE_X9Y127_C4 = 1'b1;
  assign CLBLM_R_X7Y127_SLICE_X9Y127_C5 = 1'b1;
  assign CLBLM_R_X7Y127_SLICE_X9Y127_C6 = 1'b1;
  assign RIOI3_TBYTESRC_X105Y107_ILOGIC_X1Y108_D = RIOB33_X105Y107_IOB_X1Y108_I;
  assign RIOI3_TBYTESRC_X105Y107_ILOGIC_X1Y107_D = RIOB33_X105Y107_IOB_X1Y107_I;
  assign CLBLM_R_X7Y127_SLICE_X9Y127_D5 = 1'b1;
  assign CLBLM_R_X7Y127_SLICE_X9Y127_D6 = 1'b1;
  assign CLBLM_R_X103Y172_SLICE_X163Y172_B4 = 1'b1;
  assign CLBLM_R_X5Y116_SLICE_X7Y116_A1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X5Y116_SLICE_X7Y116_A2 = CLBLM_R_X7Y113_SLICE_X8Y113_AQ;
  assign CLBLM_R_X5Y116_SLICE_X7Y116_A3 = CLBLM_R_X5Y116_SLICE_X7Y116_AQ;
  assign CLBLM_R_X5Y116_SLICE_X7Y116_A4 = CLBLM_L_X10Y116_SLICE_X13Y116_AQ;
  assign CLBLM_R_X5Y116_SLICE_X7Y116_A5 = 1'b1;
  assign CLBLM_R_X5Y116_SLICE_X7Y116_A6 = CLBLM_R_X5Y115_SLICE_X6Y115_CO5;
  assign RIOI3_X105Y167_OLOGIC_X1Y168_D1 = CLBLM_R_X7Y151_SLICE_X8Y151_AO6;
  assign CLBLM_R_X5Y116_SLICE_X7Y116_AX = CLBLM_R_X5Y116_SLICE_X7Y116_BO6;
  assign CLBLM_R_X5Y116_SLICE_X7Y116_B1 = CLBLM_R_X5Y116_SLICE_X7Y116_DO6;
  assign CLBLM_R_X5Y116_SLICE_X7Y116_B2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X5Y116_SLICE_X7Y116_B3 = CLBLM_R_X5Y123_SLICE_X6Y123_AQ;
  assign CLBLM_R_X5Y116_SLICE_X7Y116_B4 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_R_X5Y116_SLICE_X7Y116_B5 = CLBLM_R_X3Y118_SLICE_X2Y118_AQ;
  assign CLBLM_R_X5Y116_SLICE_X7Y116_B6 = 1'b1;
  assign CLBLM_R_X5Y116_SLICE_X7Y116_C1 = CLBLM_R_X3Y118_SLICE_X2Y118_AQ;
  assign CLBLM_R_X5Y116_SLICE_X7Y116_C2 = CLBLM_R_X5Y116_SLICE_X7Y116_CQ;
  assign CLBLM_R_X5Y116_SLICE_X7Y116_C3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X5Y116_SLICE_X7Y116_C4 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_R_X5Y116_SLICE_X7Y116_C5 = CLBLM_R_X7Y124_SLICE_X8Y124_A5Q;
  assign CLBLM_R_X5Y116_SLICE_X7Y116_C6 = CLBLM_R_X5Y110_SLICE_X7Y110_BQ;
  assign LIOB33_X0Y119_IOB_X0Y119_O = CLBLM_L_X8Y114_SLICE_X10Y114_CQ;
  assign LIOB33_X0Y119_IOB_X0Y120_O = CLBLM_R_X3Y116_SLICE_X3Y116_A5Q;
  assign CLBLM_R_X5Y116_SLICE_X7Y116_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X5Y116_SLICE_X7Y116_D1 = CLBLL_L_X4Y121_SLICE_X4Y121_AQ;
  assign CLBLM_R_X5Y116_SLICE_X7Y116_D2 = CLBLM_R_X7Y120_SLICE_X9Y120_CQ;
  assign CLBLM_R_X5Y116_SLICE_X7Y116_D3 = CLBLM_R_X7Y111_SLICE_X8Y111_AQ;
  assign CLBLM_R_X5Y116_SLICE_X7Y116_D4 = CLBLM_R_X5Y116_SLICE_X7Y116_A5Q;
  assign CLBLM_R_X5Y116_SLICE_X7Y116_D5 = CLBLM_R_X5Y114_SLICE_X7Y114_AQ;
  assign CLBLM_R_X5Y116_SLICE_X7Y116_D6 = CLBLL_L_X4Y114_SLICE_X4Y114_BQ;
  assign CLBLM_L_X10Y119_SLICE_X12Y119_A5 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_R_X5Y116_SLICE_X6Y116_A1 = 1'b1;
  assign CLBLM_R_X5Y116_SLICE_X6Y116_A2 = CLBLM_L_X8Y119_SLICE_X10Y119_AQ;
  assign CLBLM_R_X5Y116_SLICE_X6Y116_A3 = CLBLM_R_X5Y116_SLICE_X6Y116_AQ;
  assign CLBLM_R_X5Y116_SLICE_X6Y116_A4 = CLBLL_L_X4Y111_SLICE_X4Y111_CQ;
  assign CLBLM_R_X5Y116_SLICE_X6Y116_A5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X5Y116_SLICE_X6Y116_A6 = CLBLM_R_X5Y115_SLICE_X6Y115_CO5;
  assign CLBLM_R_X5Y116_SLICE_X6Y116_AX = CLBLM_R_X5Y116_SLICE_X6Y116_CO6;
  assign CLBLM_R_X5Y116_SLICE_X6Y116_B1 = CLBLM_R_X5Y110_SLICE_X7Y110_BQ;
  assign CLBLM_R_X5Y116_SLICE_X6Y116_B2 = CLBLM_R_X5Y116_SLICE_X6Y116_BQ;
  assign CLBLM_R_X5Y116_SLICE_X6Y116_B3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X5Y116_SLICE_X6Y116_B4 = CLBLL_L_X4Y118_SLICE_X5Y118_AQ;
  assign CLBLM_R_X5Y116_SLICE_X6Y116_B5 = CLBLM_L_X10Y114_SLICE_X13Y114_D5Q;
  assign CLBLM_R_X5Y116_SLICE_X6Y116_B6 = CLBLM_R_X5Y116_SLICE_X7Y116_BO5;
  assign CLBLM_R_X7Y127_SLICE_X8Y127_B5 = 1'b1;
  assign CLBLM_R_X7Y127_SLICE_X8Y127_B6 = 1'b1;
  assign RIOI3_X105Y167_OLOGIC_X1Y168_T1 = 1'b1;
  assign CLBLM_R_X5Y116_SLICE_X6Y116_C1 = CLBLL_L_X4Y115_SLICE_X5Y115_AQ;
  assign CLBLM_R_X5Y116_SLICE_X6Y116_C2 = CLBLM_L_X8Y114_SLICE_X10Y114_C5Q;
  assign CLBLM_R_X5Y116_SLICE_X6Y116_C3 = RIOB33_X105Y121_IOB_X1Y121_I;
  assign CLBLM_R_X5Y116_SLICE_X6Y116_C4 = CLBLM_R_X5Y123_SLICE_X7Y123_AQ;
  assign CLBLM_R_X5Y116_SLICE_X6Y116_C5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X5Y116_SLICE_X6Y116_C6 = 1'b1;
  assign CLBLM_R_X5Y116_SLICE_X6Y116_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X5Y116_SLICE_X6Y116_D1 = CLBLM_R_X5Y116_SLICE_X6Y116_CO5;
  assign CLBLM_R_X5Y116_SLICE_X6Y116_D2 = CLBLM_R_X5Y116_SLICE_X6Y116_AQ;
  assign CLBLM_R_X5Y116_SLICE_X6Y116_D3 = 1'b1;
  assign CLBLM_R_X5Y116_SLICE_X6Y116_D4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X5Y116_SLICE_X6Y116_D5 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X5Y116_SLICE_X6Y116_D6 = CLBLM_R_X7Y116_SLICE_X8Y116_BQ;
  assign CLBLM_L_X10Y119_SLICE_X12Y119_B3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y119_SLICE_X12Y119_B4 = 1'b1;
  assign CLBLM_L_X10Y119_SLICE_X12Y119_B5 = CLBLM_R_X5Y119_SLICE_X7Y119_AO6;
  assign CLBLM_L_X10Y119_SLICE_X12Y119_B6 = CLBLM_L_X10Y117_SLICE_X13Y117_BQ;
  assign CLBLM_R_X7Y127_SLICE_X8Y127_C4 = 1'b1;
  assign CLBLM_R_X7Y127_SLICE_X8Y127_C5 = 1'b1;
  assign CLBLM_R_X7Y127_SLICE_X8Y127_C6 = 1'b1;
  assign RIOI3_X105Y167_OLOGIC_X1Y167_D1 = LIOB33_SING_X0Y50_IOB_X0Y50_I;
  assign CLBLM_L_X8Y133_SLICE_X11Y133_A1 = CLBLM_L_X8Y120_SLICE_X10Y120_A5Q;
  assign CLBLM_L_X8Y133_SLICE_X11Y133_A2 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X8Y133_SLICE_X11Y133_A3 = RIOB33_X105Y139_IOB_X1Y140_I;
  assign CLBLM_L_X8Y133_SLICE_X11Y133_A4 = RIOB33_X105Y141_IOB_X1Y141_I;
  assign CLBLM_L_X8Y133_SLICE_X11Y133_A5 = CLBLM_L_X8Y120_SLICE_X11Y120_C5Q;
  assign CLBLM_L_X8Y133_SLICE_X11Y133_A6 = 1'b1;
  assign CLBLM_L_X10Y119_SLICE_X12Y119_C4 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X8Y133_SLICE_X11Y133_B1 = 1'b1;
  assign CLBLM_L_X8Y133_SLICE_X11Y133_B2 = 1'b1;
  assign CLBLM_L_X8Y133_SLICE_X11Y133_B3 = 1'b1;
  assign CLBLM_L_X8Y133_SLICE_X11Y133_B4 = 1'b1;
  assign CLBLM_L_X8Y133_SLICE_X11Y133_B5 = 1'b1;
  assign CLBLM_L_X8Y133_SLICE_X11Y133_B6 = 1'b1;
  assign CLBLM_L_X8Y133_SLICE_X11Y133_C1 = 1'b1;
  assign CLBLM_L_X8Y133_SLICE_X11Y133_C2 = 1'b1;
  assign CLBLM_L_X8Y133_SLICE_X11Y133_C3 = 1'b1;
  assign CLBLM_L_X8Y133_SLICE_X11Y133_C4 = 1'b1;
  assign CLBLM_L_X8Y133_SLICE_X11Y133_C5 = 1'b1;
  assign CLBLM_L_X8Y133_SLICE_X11Y133_C6 = 1'b1;
  assign RIOI3_X105Y177_OLOGIC_X1Y177_T1 = 1'b1;
  assign CLBLM_L_X8Y133_SLICE_X11Y133_D1 = 1'b1;
  assign CLBLM_L_X8Y133_SLICE_X11Y133_D2 = 1'b1;
  assign CLBLM_L_X8Y133_SLICE_X11Y133_D3 = 1'b1;
  assign CLBLM_L_X8Y133_SLICE_X11Y133_D4 = 1'b1;
  assign CLBLM_L_X8Y133_SLICE_X11Y133_D5 = 1'b1;
  assign CLBLM_L_X8Y133_SLICE_X11Y133_D6 = 1'b1;
  assign RIOI3_X105Y167_OLOGIC_X1Y167_T1 = 1'b1;
  assign CLBLM_L_X8Y133_SLICE_X10Y133_A1 = 1'b1;
  assign CLBLM_L_X8Y133_SLICE_X10Y133_A2 = 1'b1;
  assign CLBLM_L_X8Y133_SLICE_X10Y133_A3 = 1'b1;
  assign CLBLM_L_X8Y133_SLICE_X10Y133_A4 = 1'b1;
  assign CLBLM_L_X8Y133_SLICE_X10Y133_A5 = 1'b1;
  assign CLBLM_L_X8Y133_SLICE_X10Y133_A6 = 1'b1;
  assign CLBLM_L_X8Y133_SLICE_X10Y133_B1 = 1'b1;
  assign CLBLM_L_X8Y133_SLICE_X10Y133_B2 = 1'b1;
  assign CLBLM_L_X8Y133_SLICE_X10Y133_B3 = 1'b1;
  assign CLBLM_L_X8Y133_SLICE_X10Y133_B4 = 1'b1;
  assign CLBLM_L_X8Y133_SLICE_X10Y133_B5 = 1'b1;
  assign CLBLM_L_X8Y133_SLICE_X10Y133_B6 = 1'b1;
  assign CLBLM_L_X8Y121_SLICE_X10Y121_A4 = CLBLM_L_X10Y123_SLICE_X12Y123_AO6;
  assign CLBLM_L_X8Y133_SLICE_X10Y133_C1 = 1'b1;
  assign CLBLM_L_X8Y133_SLICE_X10Y133_C2 = 1'b1;
  assign CLBLM_L_X8Y121_SLICE_X10Y121_A5 = CLBLM_L_X8Y122_SLICE_X11Y122_AQ;
  assign CLBLM_L_X8Y133_SLICE_X10Y133_C3 = 1'b1;
  assign CLBLM_L_X8Y133_SLICE_X10Y133_C4 = 1'b1;
  assign CLBLM_L_X8Y133_SLICE_X10Y133_C5 = 1'b1;
  assign CLBLM_L_X8Y133_SLICE_X10Y133_C6 = 1'b1;
  assign CLBLM_L_X8Y121_SLICE_X10Y121_A6 = CLBLM_R_X7Y123_SLICE_X9Y123_CO6;
  assign CLBLM_R_X103Y172_SLICE_X163Y172_A1 = RIOB33_X105Y143_IOB_X1Y143_I;
  assign CLBLM_R_X103Y172_SLICE_X163Y172_A2 = CLBLM_L_X8Y116_SLICE_X10Y116_AQ;
  assign CLBLM_R_X103Y172_SLICE_X163Y172_A3 = 1'b1;
  assign CLBLM_R_X103Y172_SLICE_X163Y172_A4 = CLBLM_R_X13Y119_SLICE_X18Y119_AQ;
  assign CLBLM_R_X103Y172_SLICE_X163Y172_A5 = 1'b1;
  assign CLBLM_R_X103Y172_SLICE_X163Y172_A6 = 1'b1;
  assign CLBLM_L_X8Y133_SLICE_X10Y133_D1 = 1'b1;
  assign CLBLM_L_X8Y133_SLICE_X10Y133_D2 = 1'b1;
  assign CLBLM_L_X8Y133_SLICE_X10Y133_D3 = 1'b1;
  assign CLBLM_L_X8Y133_SLICE_X10Y133_D4 = 1'b1;
  assign CLBLM_L_X8Y133_SLICE_X10Y133_D5 = 1'b1;
  assign CLBLM_L_X8Y133_SLICE_X10Y133_D6 = 1'b1;
  assign CLBLM_R_X103Y172_SLICE_X163Y172_B1 = 1'b1;
  assign CLBLM_R_X103Y172_SLICE_X163Y172_B2 = 1'b1;
  assign CLBLM_R_X103Y172_SLICE_X163Y172_B3 = 1'b1;
  assign CLBLM_R_X103Y172_SLICE_X163Y172_B5 = 1'b1;
  assign CLBLM_R_X103Y172_SLICE_X163Y172_B6 = 1'b1;
  assign CLBLM_R_X103Y172_SLICE_X163Y172_C1 = 1'b1;
  assign CLBLM_R_X103Y172_SLICE_X163Y172_C2 = 1'b1;
  assign CLBLM_R_X103Y172_SLICE_X163Y172_C3 = 1'b1;
  assign CLBLM_R_X103Y172_SLICE_X163Y172_C4 = 1'b1;
  assign CLBLM_R_X103Y172_SLICE_X163Y172_C5 = 1'b1;
  assign CLBLM_R_X103Y172_SLICE_X163Y172_C6 = 1'b1;
  assign CLBLM_R_X103Y172_SLICE_X163Y172_D1 = 1'b1;
  assign CLBLM_R_X103Y172_SLICE_X163Y172_D2 = 1'b1;
  assign CLBLM_R_X103Y172_SLICE_X163Y172_D3 = 1'b1;
  assign CLBLM_R_X103Y172_SLICE_X163Y172_D4 = 1'b1;
  assign CLBLM_R_X103Y172_SLICE_X163Y172_D5 = 1'b1;
  assign CLBLM_R_X103Y172_SLICE_X163Y172_D6 = 1'b1;
  assign CLBLM_L_X8Y121_SLICE_X10Y121_B3 = CLBLM_R_X7Y114_SLICE_X8Y114_BQ;
  assign CLBLM_R_X103Y172_SLICE_X162Y172_A1 = 1'b1;
  assign CLBLM_L_X8Y121_SLICE_X10Y121_B4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X103Y172_SLICE_X162Y172_A2 = 1'b1;
  assign CLBLM_R_X103Y172_SLICE_X162Y172_A3 = 1'b1;
  assign CLBLM_R_X103Y172_SLICE_X162Y172_A4 = 1'b1;
  assign CLBLM_R_X103Y172_SLICE_X162Y172_A5 = 1'b1;
  assign CLBLM_R_X103Y172_SLICE_X162Y172_A6 = 1'b1;
  assign CLBLM_L_X8Y121_SLICE_X10Y121_B6 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X103Y172_SLICE_X162Y172_B1 = 1'b1;
  assign CLBLM_R_X103Y172_SLICE_X162Y172_B2 = 1'b1;
  assign CLBLM_R_X103Y172_SLICE_X162Y172_B3 = 1'b1;
  assign CLBLM_R_X103Y172_SLICE_X162Y172_B4 = 1'b1;
  assign CLBLM_R_X103Y172_SLICE_X162Y172_B5 = 1'b1;
  assign CLBLM_R_X103Y172_SLICE_X162Y172_B6 = 1'b1;
  assign CLBLM_R_X103Y172_SLICE_X162Y172_C1 = 1'b1;
  assign CLBLM_R_X103Y172_SLICE_X162Y172_C2 = 1'b1;
  assign CLBLM_R_X103Y172_SLICE_X162Y172_C3 = 1'b1;
  assign CLBLM_R_X7Y127_SLICE_X9Y127_A1 = 1'b1;
  assign CLBLM_R_X7Y127_SLICE_X9Y127_A2 = 1'b1;
  assign CLBLM_R_X7Y127_SLICE_X9Y127_A3 = 1'b1;
  assign CLBLM_R_X7Y127_SLICE_X9Y127_A4 = 1'b1;
  assign CLBLM_R_X7Y127_SLICE_X9Y127_A5 = 1'b1;
  assign CLBLM_R_X7Y127_SLICE_X9Y127_A6 = 1'b1;
  assign CLBLM_R_X103Y172_SLICE_X162Y172_C4 = 1'b1;
  assign CLBLM_R_X103Y172_SLICE_X162Y172_C5 = 1'b1;
  assign CLBLM_R_X103Y172_SLICE_X162Y172_C6 = 1'b1;
  assign CLBLM_R_X7Y127_SLICE_X9Y127_B1 = 1'b1;
  assign CLBLM_R_X7Y127_SLICE_X9Y127_B2 = 1'b1;
  assign CLBLM_R_X7Y127_SLICE_X9Y127_B3 = 1'b1;
  assign CLBLM_R_X7Y127_SLICE_X9Y127_B4 = 1'b1;
  assign CLBLM_R_X7Y127_SLICE_X9Y127_B5 = 1'b1;
  assign CLBLM_R_X7Y127_SLICE_X9Y127_B6 = 1'b1;
  assign CLBLM_R_X103Y172_SLICE_X162Y172_D1 = 1'b1;
  assign CLBLM_R_X103Y172_SLICE_X162Y172_D2 = 1'b1;
  assign CLBLM_R_X5Y117_SLICE_X7Y117_A1 = CLBLM_R_X5Y117_SLICE_X7Y117_AQ;
  assign CLBLM_R_X5Y117_SLICE_X7Y117_A2 = CLBLL_L_X2Y112_SLICE_X1Y112_BQ;
  assign CLBLM_R_X5Y117_SLICE_X7Y117_A3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X5Y117_SLICE_X7Y117_A4 = CLBLM_R_X3Y112_SLICE_X3Y112_AQ;
  assign CLBLM_R_X5Y117_SLICE_X7Y117_A5 = CLBLM_R_X5Y123_SLICE_X7Y123_AQ;
  assign CLBLM_R_X5Y117_SLICE_X7Y117_A6 = CLBLM_L_X8Y112_SLICE_X10Y112_CQ;
  assign CLBLM_R_X7Y127_SLICE_X9Y127_C1 = 1'b1;
  assign CLBLM_R_X7Y127_SLICE_X9Y127_C2 = 1'b1;
  assign CLBLM_R_X7Y127_SLICE_X9Y127_C3 = 1'b1;
  assign CLBLM_R_X5Y117_SLICE_X7Y117_B1 = 1'b1;
  assign CLBLM_R_X5Y117_SLICE_X7Y117_B2 = CLBLM_R_X5Y117_SLICE_X7Y117_BQ;
  assign CLBLM_R_X5Y117_SLICE_X7Y117_B3 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X5Y117_SLICE_X7Y117_B4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X5Y117_SLICE_X7Y117_B5 = CLBLM_L_X12Y118_SLICE_X16Y118_BQ;
  assign CLBLM_R_X5Y117_SLICE_X7Y117_B6 = 1'b1;
  assign CLBLM_R_X7Y127_SLICE_X9Y127_D1 = 1'b1;
  assign CLBLM_R_X7Y127_SLICE_X9Y127_D2 = 1'b1;
  assign CLBLM_R_X5Y117_SLICE_X7Y117_C1 = CLBLL_L_X4Y120_SLICE_X5Y120_AO6;
  assign CLBLM_R_X5Y117_SLICE_X7Y117_C2 = CLBLM_R_X5Y111_SLICE_X7Y111_CO6;
  assign CLBLM_R_X5Y117_SLICE_X7Y117_C3 = CLBLL_L_X2Y120_SLICE_X1Y120_DO6;
  assign CLBLM_R_X5Y117_SLICE_X7Y117_C4 = CLBLM_R_X3Y119_SLICE_X2Y119_AO6;
  assign CLBLM_R_X5Y117_SLICE_X7Y117_C5 = CLBLM_R_X7Y120_SLICE_X9Y120_D5Q;
  assign CLBLM_R_X5Y117_SLICE_X7Y117_C6 = CLBLM_R_X5Y118_SLICE_X7Y118_DO6;
  assign CLBLM_R_X7Y127_SLICE_X9Y127_D3 = 1'b1;
  assign CLBLM_R_X7Y127_SLICE_X9Y127_D4 = 1'b1;
  assign CLBLM_R_X5Y117_SLICE_X7Y117_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X7Y127_SLICE_X8Y127_A1 = 1'b1;
  assign CLBLM_R_X7Y127_SLICE_X8Y127_A2 = 1'b1;
  assign CLBLM_R_X7Y127_SLICE_X8Y127_A3 = 1'b1;
  assign CLBLM_R_X7Y127_SLICE_X8Y127_A4 = 1'b1;
  assign CLBLM_R_X7Y127_SLICE_X8Y127_A5 = 1'b1;
  assign CLBLM_R_X5Y117_SLICE_X7Y117_D1 = 1'b1;
  assign CLBLM_R_X5Y117_SLICE_X7Y117_D2 = RIOB33_X105Y135_IOB_X1Y135_I;
  assign CLBLM_R_X5Y117_SLICE_X7Y117_D3 = RIOB33_X105Y135_IOB_X1Y136_I;
  assign CLBLM_R_X5Y117_SLICE_X7Y117_D4 = RIOB33_X105Y131_IOB_X1Y131_I;
  assign CLBLM_R_X5Y117_SLICE_X7Y117_D5 = CLBLM_L_X8Y121_SLICE_X10Y121_DO6;
  assign CLBLM_R_X5Y117_SLICE_X7Y117_D6 = 1'b1;
  assign CLBLM_R_X7Y127_SLICE_X8Y127_A6 = 1'b1;
  assign CLBLM_R_X7Y127_SLICE_X8Y127_AX = CLBLM_L_X8Y128_SLICE_X10Y128_AO6;
  assign CLBLM_R_X7Y127_SLICE_X8Y127_B1 = 1'b1;
  assign CLBLM_R_X7Y127_SLICE_X8Y127_B2 = 1'b1;
  assign CLBLM_R_X7Y127_SLICE_X8Y127_B3 = 1'b1;
  assign CLBLM_R_X7Y127_SLICE_X8Y127_B4 = 1'b1;
  assign CLBLM_R_X5Y117_SLICE_X6Y117_A1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X5Y117_SLICE_X6Y117_A2 = CLBLL_L_X4Y111_SLICE_X4Y111_AO5;
  assign CLBLM_R_X5Y117_SLICE_X6Y117_A3 = CLBLM_R_X5Y117_SLICE_X6Y117_AQ;
  assign CLBLM_R_X5Y117_SLICE_X6Y117_A4 = CLBLL_L_X4Y110_SLICE_X5Y110_BQ;
  assign CLBLM_R_X5Y117_SLICE_X6Y117_A5 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X5Y117_SLICE_X6Y117_A6 = CLBLL_L_X4Y120_SLICE_X4Y120_AO6;
  assign CLBLM_R_X7Y127_SLICE_X8Y127_C1 = 1'b1;
  assign CLBLM_R_X7Y127_SLICE_X8Y127_C2 = 1'b1;
  assign CLBLM_R_X7Y127_SLICE_X8Y127_C3 = 1'b1;
  assign CLBLM_R_X5Y117_SLICE_X6Y117_B1 = RIOB33_X105Y135_IOB_X1Y136_I;
  assign CLBLM_R_X5Y117_SLICE_X6Y117_B2 = CLBLM_L_X8Y121_SLICE_X10Y121_DO6;
  assign CLBLM_R_X5Y117_SLICE_X6Y117_B3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X5Y117_SLICE_X6Y117_B4 = RIOB33_X105Y135_IOB_X1Y135_I;
  assign CLBLM_R_X5Y117_SLICE_X6Y117_B5 = CLBLM_R_X3Y111_SLICE_X3Y111_AQ;
  assign CLBLM_R_X5Y117_SLICE_X6Y117_B6 = RIOB33_X105Y131_IOB_X1Y131_I;
  assign CLBLM_R_X7Y127_SLICE_X8Y127_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X7Y127_SLICE_X8Y127_D1 = 1'b1;
  assign CLBLM_R_X7Y127_SLICE_X8Y127_D2 = 1'b1;
  assign CLBLM_R_X5Y117_SLICE_X6Y117_C1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X5Y117_SLICE_X6Y117_C2 = CLBLM_R_X5Y117_SLICE_X6Y117_CQ;
  assign CLBLM_R_X5Y117_SLICE_X6Y117_C3 = CLBLL_L_X4Y118_SLICE_X5Y118_AQ;
  assign CLBLM_R_X5Y117_SLICE_X6Y117_C4 = CLBLM_L_X10Y123_SLICE_X13Y123_AQ;
  assign CLBLM_R_X5Y117_SLICE_X6Y117_C5 = CLBLM_L_X8Y112_SLICE_X10Y112_CQ;
  assign CLBLM_R_X5Y117_SLICE_X6Y117_C6 = CLBLL_L_X2Y112_SLICE_X1Y112_BQ;
  assign CLBLM_R_X7Y127_SLICE_X8Y127_D3 = 1'b1;
  assign CLBLM_R_X7Y127_SLICE_X8Y127_D4 = 1'b1;
  assign CLBLM_R_X7Y127_SLICE_X8Y127_D5 = 1'b1;
  assign CLBLM_R_X5Y117_SLICE_X6Y117_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X7Y127_SLICE_X8Y127_D6 = 1'b1;
  assign RIOI3_X105Y185_OLOGIC_X1Y185_D1 = CLBLM_R_X7Y119_SLICE_X9Y119_DO5;
  assign LIOI3_TBYTESRC_X0Y193_OLOGIC_X0Y194_D1 = LIOB33_X0Y59_IOB_X0Y60_I;
  assign CLBLM_R_X5Y117_SLICE_X6Y117_D1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X5Y117_SLICE_X6Y117_D2 = 1'b1;
  assign CLBLM_R_X5Y117_SLICE_X6Y117_D3 = CLBLM_R_X5Y113_SLICE_X6Y113_CQ;
  assign CLBLM_R_X5Y117_SLICE_X6Y117_D4 = CLBLM_R_X5Y121_SLICE_X6Y121_BQ;
  assign CLBLM_R_X5Y117_SLICE_X6Y117_D5 = RIOB33_X105Y101_IOB_X1Y101_I;
  assign CLBLM_R_X5Y117_SLICE_X6Y117_D6 = 1'b1;
  assign RIOI3_X105Y185_OLOGIC_X1Y185_T1 = 1'b1;
  assign LIOI3_TBYTESRC_X0Y193_OLOGIC_X0Y194_T1 = 1'b1;
  assign LIOI3_TBYTESRC_X0Y193_OLOGIC_X0Y193_D1 = LIOB33_X0Y55_IOB_X0Y56_I;
  assign LIOI3_TBYTESRC_X0Y193_OLOGIC_X0Y193_T1 = 1'b1;
  assign CLBLM_R_X11Y123_SLICE_X14Y123_C4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign RIOB33_X105Y175_IOB_X1Y176_O = CLBLM_R_X103Y174_SLICE_X163Y174_AO5;
  assign RIOI3_SING_X105Y199_OLOGIC_X1Y199_T1 = 1'b1;
  assign CLBLM_L_X8Y111_SLICE_X11Y111_B2 = CLBLL_L_X2Y119_SLICE_X1Y119_BO6;
  assign LIOI3_X0Y79_ILOGIC_X0Y79_D = LIOB33_X0Y79_IOB_X0Y79_I;
  assign RIOI3_X105Y125_ILOGIC_X1Y126_D = RIOB33_X105Y125_IOB_X1Y126_I;
  assign RIOI3_X105Y125_ILOGIC_X1Y125_D = RIOB33_X105Y125_IOB_X1Y125_I;
  assign LIOB33_X0Y123_IOB_X0Y124_O = CLBLL_L_X4Y116_SLICE_X4Y116_C5Q;
  assign LIOB33_X0Y123_IOB_X0Y123_O = CLBLM_R_X5Y117_SLICE_X6Y117_D5Q;
  assign CLBLM_L_X8Y111_SLICE_X11Y111_C1 = CLBLM_R_X7Y111_SLICE_X9Y111_AO5;
  assign CLBLM_R_X7Y128_SLICE_X9Y128_A1 = 1'b1;
  assign CLBLM_R_X7Y128_SLICE_X9Y128_A2 = 1'b1;
  assign CLBLM_R_X7Y128_SLICE_X9Y128_A3 = 1'b1;
  assign CLBLM_R_X7Y128_SLICE_X9Y128_A4 = 1'b1;
  assign CLBLM_R_X7Y128_SLICE_X9Y128_A5 = 1'b1;
  assign CLBLM_R_X7Y128_SLICE_X9Y128_A6 = 1'b1;
  assign CLBLM_R_X7Y128_SLICE_X9Y128_B1 = 1'b1;
  assign CLBLM_R_X7Y128_SLICE_X9Y128_B2 = 1'b1;
  assign CLBLM_R_X7Y128_SLICE_X9Y128_B3 = 1'b1;
  assign CLBLM_R_X7Y128_SLICE_X9Y128_B4 = 1'b1;
  assign CLBLM_R_X7Y128_SLICE_X9Y128_B5 = 1'b1;
  assign CLBLM_R_X7Y128_SLICE_X9Y128_B6 = 1'b1;
  assign CLBLM_R_X5Y118_SLICE_X7Y118_A1 = 1'b1;
  assign CLBLM_R_X5Y118_SLICE_X7Y118_A2 = CLBLM_R_X5Y114_SLICE_X6Y114_BQ;
  assign CLBLM_R_X5Y118_SLICE_X7Y118_A3 = CLBLM_R_X5Y118_SLICE_X7Y118_AQ;
  assign CLBLM_R_X5Y118_SLICE_X7Y118_A4 = CLBLM_R_X7Y118_SLICE_X8Y118_DQ;
  assign CLBLM_R_X5Y118_SLICE_X7Y118_A5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X5Y118_SLICE_X7Y118_A6 = CLBLM_R_X5Y115_SLICE_X6Y115_CO6;
  assign CLBLM_R_X7Y128_SLICE_X9Y128_C1 = 1'b1;
  assign CLBLM_R_X7Y128_SLICE_X9Y128_C2 = 1'b1;
  assign CLBLM_R_X7Y128_SLICE_X9Y128_C3 = 1'b1;
  assign CLBLM_R_X5Y118_SLICE_X7Y118_B1 = CLBLL_L_X4Y119_SLICE_X4Y119_B5Q;
  assign CLBLM_R_X5Y118_SLICE_X7Y118_B2 = CLBLM_R_X5Y116_SLICE_X6Y116_A5Q;
  assign CLBLM_R_X5Y118_SLICE_X7Y118_B3 = CLBLM_R_X5Y119_SLICE_X6Y119_B5Q;
  assign CLBLM_R_X5Y118_SLICE_X7Y118_B4 = CLBLM_R_X5Y125_SLICE_X6Y125_A5Q;
  assign CLBLM_R_X5Y118_SLICE_X7Y118_B5 = CLBLM_R_X3Y117_SLICE_X3Y117_AQ;
  assign CLBLM_R_X5Y118_SLICE_X7Y118_B6 = 1'b1;
  assign CLBLM_R_X7Y128_SLICE_X9Y128_D1 = 1'b1;
  assign CLBLM_R_X7Y128_SLICE_X9Y128_D2 = 1'b1;
  assign CLBLM_R_X5Y118_SLICE_X7Y118_C1 = CLBLL_L_X4Y120_SLICE_X4Y120_AO6;
  assign CLBLM_R_X5Y118_SLICE_X7Y118_C2 = CLBLM_R_X3Y113_SLICE_X3Y113_DO6;
  assign CLBLM_R_X5Y118_SLICE_X7Y118_C3 = CLBLM_R_X5Y120_SLICE_X7Y120_DO6;
  assign CLBLM_R_X5Y118_SLICE_X7Y118_C4 = CLBLL_L_X4Y120_SLICE_X4Y120_BO6;
  assign CLBLM_R_X5Y118_SLICE_X7Y118_C5 = CLBLM_R_X3Y120_SLICE_X3Y120_BO6;
  assign CLBLM_R_X5Y118_SLICE_X7Y118_C6 = CLBLL_L_X2Y120_SLICE_X0Y120_CO6;
  assign CLBLM_R_X7Y128_SLICE_X9Y128_D3 = 1'b1;
  assign CLBLM_R_X7Y128_SLICE_X9Y128_D4 = 1'b1;
  assign CLBLM_L_X10Y127_SLICE_X13Y127_B1 = 1'b1;
  assign CLBLM_R_X5Y118_SLICE_X7Y118_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X7Y128_SLICE_X8Y128_A3 = CLBLM_R_X7Y128_SLICE_X8Y128_AQ;
  assign CLBLM_R_X7Y128_SLICE_X8Y128_A4 = RIOB33_X105Y141_IOB_X1Y142_I;
  assign CLBLM_R_X7Y128_SLICE_X8Y128_A5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y128_SLICE_X8Y128_A6 = 1'b1;
  assign CLBLM_R_X5Y118_SLICE_X7Y118_D1 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X5Y118_SLICE_X7Y118_D2 = CLBLM_R_X5Y122_SLICE_X7Y122_A5Q;
  assign CLBLM_R_X5Y118_SLICE_X7Y118_D3 = CLBLM_L_X8Y119_SLICE_X11Y119_C5Q;
  assign CLBLM_R_X5Y118_SLICE_X7Y118_D4 = CLBLM_R_X5Y121_SLICE_X7Y121_A5Q;
  assign CLBLM_R_X5Y118_SLICE_X7Y118_D5 = CLBLM_R_X5Y118_SLICE_X7Y118_BO5;
  assign CLBLM_R_X5Y118_SLICE_X7Y118_D6 = CLBLM_R_X3Y117_SLICE_X3Y117_AQ;
  assign CLBLM_R_X7Y128_SLICE_X8Y128_B1 = 1'b1;
  assign CLBLM_R_X7Y128_SLICE_X8Y128_B2 = 1'b1;
  assign CLBLM_R_X7Y128_SLICE_X8Y128_B3 = 1'b1;
  assign CLBLM_R_X7Y128_SLICE_X8Y128_B4 = 1'b1;
  assign CLBLM_R_X7Y128_SLICE_X8Y128_B5 = 1'b1;
  assign CLBLM_R_X5Y118_SLICE_X6Y118_A1 = CLBLL_L_X4Y111_SLICE_X4Y111_AO5;
  assign CLBLM_R_X5Y118_SLICE_X6Y118_A2 = CLBLL_L_X4Y120_SLICE_X4Y120_BO6;
  assign CLBLM_R_X5Y118_SLICE_X6Y118_A3 = CLBLM_R_X5Y118_SLICE_X6Y118_AQ;
  assign CLBLM_R_X5Y118_SLICE_X6Y118_A4 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X5Y118_SLICE_X6Y118_A5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X5Y118_SLICE_X6Y118_A6 = CLBLM_R_X7Y120_SLICE_X9Y120_A5Q;
  assign CLBLM_R_X7Y128_SLICE_X8Y128_C1 = 1'b1;
  assign CLBLM_R_X7Y128_SLICE_X8Y128_C2 = 1'b1;
  assign CLBLM_R_X7Y128_SLICE_X8Y128_C3 = 1'b1;
  assign CLBLM_R_X5Y118_SLICE_X6Y118_B1 = CLBLM_R_X5Y118_SLICE_X6Y118_CQ;
  assign CLBLM_R_X5Y118_SLICE_X6Y118_B2 = CLBLM_R_X5Y118_SLICE_X6Y118_BQ;
  assign CLBLM_R_X5Y118_SLICE_X6Y118_B3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X5Y118_SLICE_X6Y118_B4 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_R_X5Y118_SLICE_X6Y118_B5 = CLBLM_R_X3Y118_SLICE_X2Y118_AQ;
  assign CLBLM_R_X5Y118_SLICE_X6Y118_B6 = CLBLM_R_X3Y116_SLICE_X3Y116_CQ;
  assign CLBLM_R_X7Y128_SLICE_X8Y128_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X7Y128_SLICE_X8Y128_D1 = 1'b1;
  assign CLBLM_R_X7Y128_SLICE_X8Y128_D2 = 1'b1;
  assign CLBLM_R_X5Y118_SLICE_X6Y118_C1 = CLBLM_R_X3Y118_SLICE_X2Y118_AQ;
  assign CLBLM_R_X5Y118_SLICE_X6Y118_C2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X5Y118_SLICE_X6Y118_C3 = CLBLM_R_X5Y110_SLICE_X6Y110_AQ;
  assign CLBLM_R_X5Y118_SLICE_X6Y118_C4 = CLBLM_R_X5Y122_SLICE_X7Y122_A5Q;
  assign CLBLM_R_X5Y118_SLICE_X6Y118_C5 = CLBLM_R_X5Y118_SLICE_X6Y118_CQ;
  assign CLBLM_R_X5Y118_SLICE_X6Y118_C6 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_R_X7Y128_SLICE_X8Y128_D3 = 1'b1;
  assign CLBLM_R_X7Y128_SLICE_X8Y128_D4 = 1'b1;
  assign CLBLM_R_X7Y128_SLICE_X8Y128_D5 = 1'b1;
  assign CLBLM_R_X5Y118_SLICE_X6Y118_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X7Y128_SLICE_X8Y128_D6 = 1'b1;
  assign CLBLM_R_X5Y118_SLICE_X6Y118_D1 = CLBLM_R_X7Y117_SLICE_X9Y117_CQ;
  assign CLBLM_R_X5Y118_SLICE_X6Y118_D2 = CLBLM_R_X5Y117_SLICE_X6Y117_CQ;
  assign CLBLM_R_X5Y118_SLICE_X6Y118_D3 = CLBLM_R_X3Y121_SLICE_X2Y121_AO5;
  assign CLBLM_R_X5Y118_SLICE_X6Y118_D4 = CLBLM_R_X3Y121_SLICE_X2Y121_AO6;
  assign CLBLM_R_X5Y118_SLICE_X6Y118_D5 = CLBLL_L_X2Y120_SLICE_X0Y120_AO5;
  assign CLBLM_R_X5Y118_SLICE_X6Y118_D6 = CLBLL_L_X4Y117_SLICE_X5Y117_CQ;
  assign CLBLM_R_X103Y174_SLICE_X163Y174_A1 = RIOB33_X105Y143_IOB_X1Y143_I;
  assign CLBLM_R_X103Y174_SLICE_X163Y174_A2 = 1'b1;
  assign CLBLM_R_X103Y174_SLICE_X163Y174_A3 = CLBLM_R_X11Y128_SLICE_X15Y128_AQ;
  assign CLBLM_R_X103Y174_SLICE_X163Y174_A4 = 1'b1;
  assign CLBLM_R_X103Y174_SLICE_X163Y174_A5 = CLBLM_L_X12Y115_SLICE_X16Y115_AQ;
  assign CLBLM_R_X103Y174_SLICE_X163Y174_A6 = 1'b1;
  assign CLBLM_R_X103Y174_SLICE_X163Y174_B1 = 1'b1;
  assign CLBLM_R_X103Y174_SLICE_X163Y174_B2 = 1'b1;
  assign CLBLM_R_X103Y174_SLICE_X163Y174_B3 = 1'b1;
  assign CLBLM_R_X103Y174_SLICE_X163Y174_B4 = 1'b1;
  assign CLBLM_R_X103Y174_SLICE_X163Y174_B5 = 1'b1;
  assign CLBLM_R_X103Y174_SLICE_X163Y174_B6 = 1'b1;
  assign CLBLM_R_X103Y174_SLICE_X163Y174_C1 = 1'b1;
  assign CLBLM_R_X103Y174_SLICE_X163Y174_C2 = 1'b1;
  assign CLBLM_R_X103Y174_SLICE_X163Y174_C3 = 1'b1;
  assign CLBLM_R_X103Y174_SLICE_X163Y174_C4 = 1'b1;
  assign CLBLM_R_X103Y174_SLICE_X163Y174_C5 = 1'b1;
  assign CLBLM_R_X103Y174_SLICE_X163Y174_C6 = 1'b1;
  assign LIOB33_X0Y125_IOB_X0Y125_O = CLBLM_R_X7Y115_SLICE_X9Y115_CQ;
  assign LIOB33_X0Y125_IOB_X0Y126_O = CLBLM_R_X5Y124_SLICE_X6Y124_CQ;
  assign CLBLM_R_X103Y174_SLICE_X163Y174_D1 = 1'b1;
  assign CLBLM_R_X103Y174_SLICE_X163Y174_D2 = 1'b1;
  assign CLBLM_R_X103Y174_SLICE_X163Y174_D3 = 1'b1;
  assign CLBLM_R_X103Y174_SLICE_X163Y174_D4 = 1'b1;
  assign CLBLM_R_X103Y174_SLICE_X163Y174_D5 = 1'b1;
  assign CLBLM_R_X103Y174_SLICE_X163Y174_D6 = 1'b1;
  assign CLBLM_R_X103Y174_SLICE_X162Y174_A1 = 1'b1;
  assign CLBLM_R_X103Y174_SLICE_X162Y174_A2 = 1'b1;
  assign CLBLM_R_X103Y174_SLICE_X162Y174_A3 = 1'b1;
  assign CLBLM_R_X103Y174_SLICE_X162Y174_A4 = 1'b1;
  assign CLBLM_R_X103Y174_SLICE_X162Y174_A5 = 1'b1;
  assign CLBLM_R_X103Y174_SLICE_X162Y174_A6 = 1'b1;
  assign CLBLM_R_X103Y174_SLICE_X162Y174_B1 = 1'b1;
  assign CLBLM_R_X103Y174_SLICE_X162Y174_B2 = 1'b1;
  assign CLBLM_R_X103Y174_SLICE_X162Y174_B3 = 1'b1;
  assign CLBLM_R_X103Y174_SLICE_X162Y174_B4 = 1'b1;
  assign CLBLM_R_X103Y174_SLICE_X162Y174_B5 = 1'b1;
  assign CLBLM_R_X103Y174_SLICE_X162Y174_B6 = 1'b1;
  assign CLBLM_R_X103Y174_SLICE_X162Y174_C1 = 1'b1;
  assign CLBLM_R_X103Y174_SLICE_X162Y174_C2 = 1'b1;
  assign CLBLM_R_X103Y174_SLICE_X162Y174_C3 = 1'b1;
  assign CLBLM_R_X103Y174_SLICE_X162Y174_C4 = 1'b1;
  assign CLBLM_R_X103Y174_SLICE_X162Y174_C5 = 1'b1;
  assign CLBLM_R_X103Y174_SLICE_X162Y174_C6 = 1'b1;
  assign CLBLM_R_X103Y174_SLICE_X162Y174_D1 = 1'b1;
  assign CLBLM_R_X103Y174_SLICE_X162Y174_D2 = 1'b1;
  assign CLBLM_R_X103Y174_SLICE_X162Y174_D3 = 1'b1;
  assign CLBLM_R_X103Y174_SLICE_X162Y174_D4 = 1'b1;
  assign CLBLM_R_X103Y174_SLICE_X162Y174_D5 = 1'b1;
  assign CLBLM_R_X103Y174_SLICE_X162Y174_D6 = 1'b1;
  assign LIOI3_X0Y55_ILOGIC_X0Y56_D = LIOB33_X0Y55_IOB_X0Y56_I;
  assign CLBLM_R_X5Y119_SLICE_X7Y119_A1 = CLBLM_R_X5Y119_SLICE_X7Y119_DO6;
  assign CLBLM_R_X5Y119_SLICE_X7Y119_A2 = CLBLM_R_X5Y118_SLICE_X7Y118_BO6;
  assign CLBLM_R_X5Y119_SLICE_X7Y119_A3 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X5Y119_SLICE_X7Y119_A4 = CLBLM_R_X7Y120_SLICE_X9Y120_D5Q;
  assign CLBLM_R_X5Y119_SLICE_X7Y119_A5 = CLBLL_L_X2Y119_SLICE_X1Y119_BO6;
  assign CLBLM_R_X5Y119_SLICE_X7Y119_A6 = CLBLM_L_X8Y119_SLICE_X11Y119_C5Q;
  assign CLBLM_R_X5Y119_SLICE_X7Y119_B1 = CLBLL_L_X4Y119_SLICE_X4Y119_B5Q;
  assign CLBLM_R_X5Y119_SLICE_X7Y119_B2 = CLBLM_R_X5Y122_SLICE_X7Y122_A5Q;
  assign CLBLM_R_X5Y119_SLICE_X7Y119_B3 = CLBLM_R_X3Y117_SLICE_X3Y117_AQ;
  assign CLBLM_R_X5Y119_SLICE_X7Y119_B4 = CLBLM_R_X5Y125_SLICE_X6Y125_A5Q;
  assign CLBLM_R_X5Y119_SLICE_X7Y119_B5 = CLBLM_R_X5Y116_SLICE_X6Y116_A5Q;
  assign CLBLM_R_X5Y119_SLICE_X7Y119_B6 = CLBLM_L_X8Y119_SLICE_X11Y119_C5Q;
  assign CLBLM_R_X5Y119_SLICE_X7Y119_C1 = CLBLM_R_X7Y120_SLICE_X9Y120_D5Q;
  assign CLBLM_R_X5Y119_SLICE_X7Y119_C2 = 1'b1;
  assign CLBLM_R_X5Y119_SLICE_X7Y119_C3 = CLBLM_R_X5Y119_SLICE_X6Y119_B5Q;
  assign CLBLM_R_X5Y119_SLICE_X7Y119_C4 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X5Y119_SLICE_X7Y119_C5 = CLBLM_R_X5Y121_SLICE_X7Y121_A5Q;
  assign CLBLM_R_X5Y119_SLICE_X7Y119_C6 = CLBLM_R_X5Y119_SLICE_X7Y119_BO6;
  assign CLBLM_R_X5Y119_SLICE_X7Y119_D1 = 1'b1;
  assign CLBLM_R_X5Y119_SLICE_X7Y119_D2 = 1'b1;
  assign CLBLM_R_X5Y119_SLICE_X7Y119_D3 = CLBLM_R_X5Y122_SLICE_X7Y122_A5Q;
  assign CLBLM_R_X5Y119_SLICE_X7Y119_D4 = 1'b1;
  assign CLBLM_R_X5Y119_SLICE_X7Y119_D5 = CLBLM_R_X5Y121_SLICE_X7Y121_A5Q;
  assign CLBLM_R_X5Y119_SLICE_X7Y119_D6 = 1'b1;
  assign CLBLM_R_X5Y119_SLICE_X6Y119_A1 = CLBLM_R_X5Y114_SLICE_X7Y114_CO6;
  assign CLBLM_R_X5Y119_SLICE_X6Y119_A2 = CLBLM_R_X5Y121_SLICE_X6Y121_A5Q;
  assign CLBLM_R_X5Y119_SLICE_X6Y119_A3 = CLBLM_R_X5Y119_SLICE_X6Y119_AQ;
  assign CLBLM_R_X5Y119_SLICE_X6Y119_A4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X5Y119_SLICE_X6Y119_A5 = CLBLM_R_X3Y118_SLICE_X2Y118_AQ;
  assign CLBLM_R_X5Y119_SLICE_X6Y119_A6 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_R_X5Y119_SLICE_X6Y119_B1 = CLBLM_R_X7Y120_SLICE_X8Y120_DQ;
  assign CLBLM_R_X5Y119_SLICE_X6Y119_B2 = CLBLL_L_X4Y118_SLICE_X5Y118_BQ;
  assign CLBLM_R_X5Y119_SLICE_X6Y119_B3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X5Y119_SLICE_X6Y119_B4 = CLBLM_R_X7Y121_SLICE_X9Y121_BQ;
  assign CLBLM_R_X5Y119_SLICE_X6Y119_B5 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X5Y119_SLICE_X6Y119_B6 = 1'b1;
  assign CLBLM_R_X5Y119_SLICE_X6Y119_C1 = 1'b1;
  assign CLBLM_R_X5Y119_SLICE_X6Y119_C2 = CLBLM_R_X5Y119_SLICE_X6Y119_CQ;
  assign CLBLM_R_X5Y119_SLICE_X6Y119_C3 = CLBLM_R_X5Y115_SLICE_X6Y115_AQ;
  assign CLBLM_R_X5Y119_SLICE_X6Y119_C4 = CLBLM_L_X8Y119_SLICE_X11Y119_C5Q;
  assign CLBLM_R_X5Y119_SLICE_X6Y119_C5 = CLBLM_R_X3Y116_SLICE_X2Y116_DO6;
  assign CLBLM_R_X5Y119_SLICE_X6Y119_C6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X5Y119_SLICE_X6Y119_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X5Y119_SLICE_X6Y119_D1 = RIOB33_X105Y131_IOB_X1Y132_I;
  assign CLBLM_R_X5Y119_SLICE_X6Y119_D2 = RIOB33_X105Y131_IOB_X1Y131_I;
  assign CLBLM_R_X5Y119_SLICE_X6Y119_D3 = RIOB33_X105Y133_IOB_X1Y134_I;
  assign CLBLM_R_X5Y119_SLICE_X6Y119_D4 = CLBLM_L_X8Y118_SLICE_X10Y118_D5Q;
  assign CLBLM_R_X5Y119_SLICE_X6Y119_D5 = RIOB33_X105Y133_IOB_X1Y133_I;
  assign CLBLM_R_X5Y119_SLICE_X6Y119_D6 = CLBLM_R_X3Y122_SLICE_X3Y122_AO6;
  assign LIOI3_X0Y55_ILOGIC_X0Y55_D = LIOB33_X0Y55_IOB_X0Y55_I;
  assign LIOI3_X0Y177_OLOGIC_X0Y177_T1 = 1'b1;
  assign LIOI3_X0Y145_OLOGIC_X0Y146_D1 = LIOB33_X0Y59_IOB_X0Y59_I;
  assign LIOI3_X0Y145_OLOGIC_X0Y146_T1 = 1'b1;
  assign RIOI3_X105Y189_OLOGIC_X1Y190_D1 = CLBLM_R_X13Y119_SLICE_X18Y119_AQ;
  assign LIOI3_X0Y145_OLOGIC_X0Y145_D1 = LIOB33_X0Y57_IOB_X0Y58_I;
  assign RIOI3_X105Y189_OLOGIC_X1Y190_T1 = 1'b1;
  assign CLBLL_L_X4Y117_SLICE_X4Y117_B3 = CLBLM_L_X10Y112_SLICE_X13Y112_CQ;
  assign CLBLM_R_X13Y120_SLICE_X19Y120_A5 = 1'b1;
  assign CLBLL_L_X4Y117_SLICE_X4Y117_B4 = CLBLM_R_X3Y116_SLICE_X2Y116_CO6;
  assign LIOI3_X0Y145_OLOGIC_X0Y145_T1 = 1'b1;
  assign RIOI3_X105Y189_OLOGIC_X1Y189_D1 = CLBLM_L_X8Y122_SLICE_X10Y122_AQ;
  assign RIOI3_X105Y189_OLOGIC_X1Y189_T1 = 1'b1;
  assign LIOB33_X0Y127_IOB_X0Y128_O = CLBLL_L_X2Y117_SLICE_X0Y117_A5Q;
  assign LIOB33_X0Y127_IOB_X0Y127_O = CLBLL_L_X4Y121_SLICE_X4Y121_BQ;
  assign CLBLL_L_X4Y117_SLICE_X4Y117_C3 = 1'b1;
  assign CLBLL_L_X4Y117_SLICE_X4Y117_C5 = CLBLM_R_X3Y122_SLICE_X3Y122_AO6;
  assign CLBLM_R_X5Y120_SLICE_X7Y120_A1 = CLBLM_R_X7Y121_SLICE_X8Y121_BQ;
  assign CLBLM_R_X5Y120_SLICE_X7Y120_A2 = CLBLM_R_X11Y121_SLICE_X14Y121_CO6;
  assign CLBLM_R_X5Y120_SLICE_X7Y120_A3 = CLBLM_R_X5Y120_SLICE_X7Y120_AQ;
  assign CLBLM_R_X5Y120_SLICE_X7Y120_A4 = 1'b1;
  assign CLBLM_R_X5Y120_SLICE_X7Y120_A5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X5Y120_SLICE_X7Y120_A6 = CLBLM_L_X8Y115_SLICE_X10Y115_AQ;
  assign CLBLM_R_X5Y120_SLICE_X7Y120_B1 = 1'b1;
  assign CLBLM_R_X5Y120_SLICE_X7Y120_B2 = CLBLM_R_X5Y120_SLICE_X7Y120_BQ;
  assign CLBLM_R_X5Y120_SLICE_X7Y120_B3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X5Y120_SLICE_X7Y120_B4 = CLBLM_R_X7Y113_SLICE_X8Y113_AQ;
  assign CLBLM_R_X5Y120_SLICE_X7Y120_B5 = CLBLM_R_X5Y115_SLICE_X6Y115_CO5;
  assign CLBLM_R_X5Y120_SLICE_X7Y120_B6 = CLBLL_L_X4Y119_SLICE_X4Y119_CQ;
  assign CLBLM_R_X3Y110_SLICE_X3Y110_A1 = CLBLL_L_X4Y111_SLICE_X4Y111_AO5;
  assign CLBLM_R_X3Y110_SLICE_X3Y110_A2 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X3Y110_SLICE_X3Y110_A3 = CLBLM_R_X3Y110_SLICE_X3Y110_AQ;
  assign CLBLM_R_X3Y110_SLICE_X3Y110_A4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X3Y110_SLICE_X3Y110_A5 = CLBLM_L_X10Y110_SLICE_X13Y110_BQ;
  assign CLBLM_R_X3Y110_SLICE_X3Y110_A6 = CLBLL_L_X2Y120_SLICE_X0Y120_CO6;
  assign CLBLM_R_X5Y120_SLICE_X7Y120_C1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X5Y120_SLICE_X7Y120_C2 = CLBLM_R_X5Y120_SLICE_X7Y120_CQ;
  assign CLBLM_R_X5Y120_SLICE_X7Y120_C3 = CLBLM_R_X5Y121_SLICE_X7Y121_A5Q;
  assign CLBLM_R_X3Y110_SLICE_X3Y110_B1 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_R_X3Y110_SLICE_X3Y110_B2 = CLBLM_R_X3Y110_SLICE_X3Y110_BQ;
  assign CLBLM_R_X3Y110_SLICE_X3Y110_B3 = 1'b1;
  assign CLBLM_R_X3Y110_SLICE_X3Y110_B4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X3Y110_SLICE_X3Y110_B5 = CLBLM_R_X3Y118_SLICE_X2Y118_AQ;
  assign CLBLM_R_X3Y110_SLICE_X3Y110_B6 = CLBLM_R_X3Y112_SLICE_X3Y112_CQ;
  assign CLBLM_R_X5Y120_SLICE_X7Y120_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X5Y120_SLICE_X7Y120_D1 = CLBLM_R_X3Y119_SLICE_X2Y119_AO6;
  assign CLBLM_R_X3Y110_SLICE_X3Y110_C1 = 1'b1;
  assign CLBLM_R_X3Y110_SLICE_X3Y110_C2 = 1'b1;
  assign CLBLM_R_X3Y110_SLICE_X3Y110_C3 = 1'b1;
  assign CLBLM_R_X3Y110_SLICE_X3Y110_C4 = 1'b1;
  assign CLBLM_R_X3Y110_SLICE_X3Y110_C5 = 1'b1;
  assign CLBLM_R_X3Y110_SLICE_X3Y110_C6 = 1'b1;
  assign CLBLM_R_X5Y120_SLICE_X7Y120_D6 = 1'b1;
  assign CLBLM_R_X3Y110_SLICE_X3Y110_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X5Y120_SLICE_X6Y120_A1 = CLBLM_R_X7Y122_SLICE_X9Y122_CO6;
  assign CLBLM_R_X5Y120_SLICE_X6Y120_A2 = CLBLM_R_X5Y119_SLICE_X6Y119_CQ;
  assign CLBLM_R_X5Y120_SLICE_X6Y120_A3 = CLBLL_L_X4Y120_SLICE_X4Y120_BO6;
  assign CLBLM_R_X5Y120_SLICE_X6Y120_A4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X5Y120_SLICE_X6Y120_A5 = CLBLM_R_X7Y109_SLICE_X8Y109_AQ;
  assign CLBLM_R_X3Y110_SLICE_X3Y110_D1 = 1'b1;
  assign CLBLM_R_X3Y110_SLICE_X3Y110_D2 = 1'b1;
  assign CLBLM_R_X3Y110_SLICE_X3Y110_D3 = 1'b1;
  assign CLBLM_R_X3Y110_SLICE_X3Y110_D4 = 1'b1;
  assign CLBLM_R_X3Y110_SLICE_X3Y110_D5 = 1'b1;
  assign CLBLM_R_X3Y110_SLICE_X3Y110_D6 = 1'b1;
  assign CLBLM_R_X5Y120_SLICE_X6Y120_A6 = 1'b1;
  assign CLBLM_R_X5Y120_SLICE_X6Y120_B1 = 1'b1;
  assign CLBLM_R_X5Y120_SLICE_X6Y120_B2 = CLBLM_R_X5Y120_SLICE_X6Y120_BQ;
  assign CLBLM_R_X5Y120_SLICE_X6Y120_B3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X5Y120_SLICE_X6Y120_B4 = CLBLM_R_X7Y116_SLICE_X8Y116_BQ;
  assign CLBLM_R_X3Y110_SLICE_X2Y110_A1 = 1'b1;
  assign CLBLM_R_X3Y110_SLICE_X2Y110_A2 = 1'b1;
  assign CLBLM_R_X3Y110_SLICE_X2Y110_A3 = 1'b1;
  assign CLBLM_R_X3Y110_SLICE_X2Y110_A4 = 1'b1;
  assign CLBLM_R_X3Y110_SLICE_X2Y110_A5 = 1'b1;
  assign CLBLM_R_X3Y110_SLICE_X2Y110_A6 = 1'b1;
  assign CLBLL_L_X52Y126_SLICE_X78Y126_D1 = 1'b1;
  assign CLBLM_R_X5Y120_SLICE_X6Y120_C1 = CLBLM_R_X3Y121_SLICE_X2Y121_AO5;
  assign CLBLM_R_X3Y110_SLICE_X2Y110_AX = CLBLM_R_X3Y111_SLICE_X2Y111_BO6;
  assign CLBLM_R_X5Y120_SLICE_X6Y120_C2 = 1'b1;
  assign CLBLM_R_X3Y110_SLICE_X2Y110_B1 = 1'b1;
  assign CLBLM_R_X3Y110_SLICE_X2Y110_B2 = 1'b1;
  assign CLBLM_R_X3Y110_SLICE_X2Y110_B3 = 1'b1;
  assign CLBLM_R_X3Y110_SLICE_X2Y110_B4 = 1'b1;
  assign CLBLM_R_X3Y110_SLICE_X2Y110_B5 = 1'b1;
  assign CLBLM_R_X3Y110_SLICE_X2Y110_B6 = 1'b1;
  assign CLBLM_R_X5Y120_SLICE_X6Y120_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X5Y120_SLICE_X6Y120_D1 = CLBLM_R_X5Y120_SLICE_X7Y120_AQ;
  assign CLBLM_R_X5Y120_SLICE_X6Y120_D2 = 1'b1;
  assign CLBLM_R_X3Y110_SLICE_X2Y110_C1 = 1'b1;
  assign CLBLM_R_X3Y110_SLICE_X2Y110_C2 = 1'b1;
  assign CLBLM_R_X3Y110_SLICE_X2Y110_C3 = 1'b1;
  assign CLBLM_R_X3Y110_SLICE_X2Y110_C4 = 1'b1;
  assign CLBLM_R_X3Y110_SLICE_X2Y110_C5 = 1'b1;
  assign CLBLM_R_X3Y110_SLICE_X2Y110_C6 = 1'b1;
  assign CLBLM_R_X5Y120_SLICE_X6Y120_D3 = CLBLL_L_X2Y120_SLICE_X0Y120_AO5;
  assign CLBLM_R_X5Y120_SLICE_X6Y120_D4 = CLBLM_R_X7Y112_SLICE_X8Y112_CQ;
  assign CLBLM_R_X5Y120_SLICE_X6Y120_D5 = 1'b1;
  assign CLBLM_R_X3Y110_SLICE_X2Y110_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLL_L_X52Y126_SLICE_X78Y126_D2 = 1'b1;
  assign CLBLM_R_X103Y169_SLICE_X162Y169_D5 = 1'b1;
  assign CLBLM_R_X3Y110_SLICE_X2Y110_D1 = 1'b1;
  assign CLBLM_R_X3Y110_SLICE_X2Y110_D2 = 1'b1;
  assign CLBLM_R_X3Y110_SLICE_X2Y110_D3 = 1'b1;
  assign CLBLM_R_X3Y110_SLICE_X2Y110_D4 = 1'b1;
  assign CLBLM_R_X3Y110_SLICE_X2Y110_D5 = 1'b1;
  assign CLBLM_R_X3Y110_SLICE_X2Y110_D6 = 1'b1;
  assign RIOI3_TBYTESRC_X105Y131_ILOGIC_X1Y132_D = RIOB33_X105Y131_IOB_X1Y132_I;
  assign CLBLM_R_X103Y169_SLICE_X162Y169_D6 = 1'b1;
  assign RIOI3_TBYTESRC_X105Y131_ILOGIC_X1Y131_D = RIOB33_X105Y131_IOB_X1Y131_I;
  assign LIOB33_X0Y129_IOB_X0Y130_O = CLBLL_L_X52Y126_SLICE_X78Y126_AO6;
  assign CLBLM_R_X7Y128_SLICE_X9Y128_C4 = 1'b1;
  assign LIOB33_X0Y129_IOB_X0Y129_O = CLBLM_R_X3Y115_SLICE_X3Y115_CQ;
  assign CLBLM_R_X7Y128_SLICE_X9Y128_C5 = 1'b1;
  assign CLBLM_R_X7Y128_SLICE_X9Y128_C6 = 1'b1;
  assign CLBLL_L_X52Y126_SLICE_X78Y126_D6 = 1'b1;
  assign LIOI3_X0Y151_OLOGIC_X0Y152_T1 = 1'b1;
  assign CLBLM_L_X10Y120_SLICE_X13Y120_C4 = CLBLM_L_X10Y120_SLICE_X13Y120_AQ;
  assign CLBLM_L_X10Y120_SLICE_X13Y120_C5 = CLBLM_R_X7Y120_SLICE_X9Y120_A5Q;
  assign CLBLM_L_X10Y120_SLICE_X13Y120_C6 = CLBLM_R_X7Y124_SLICE_X8Y124_AQ;
  assign CLBLM_L_X10Y120_SLICE_X13Y120_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X7Y128_SLICE_X9Y128_D5 = 1'b1;
  assign CLBLM_R_X7Y128_SLICE_X9Y128_D6 = 1'b1;
  assign CLBLM_L_X10Y120_SLICE_X13Y120_D1 = CLBLM_L_X10Y120_SLICE_X13Y120_BQ;
  assign CLBLM_L_X10Y120_SLICE_X13Y120_D2 = CLBLM_L_X10Y123_SLICE_X12Y123_CO6;
  assign CLBLM_L_X10Y120_SLICE_X13Y120_D3 = 1'b1;
  assign CLBLM_L_X10Y120_SLICE_X13Y120_D4 = CLBLM_L_X10Y120_SLICE_X13Y120_CO6;
  assign CLBLM_L_X10Y120_SLICE_X13Y120_D5 = CLBLM_L_X10Y121_SLICE_X12Y121_BQ;
  assign CLBLM_R_X7Y128_SLICE_X8Y128_A1 = CLBLM_L_X8Y120_SLICE_X10Y120_A5Q;
  assign CLBLM_L_X10Y120_SLICE_X13Y120_D6 = CLBLM_L_X8Y122_SLICE_X11Y122_DO6;
  assign CLBLM_R_X5Y121_SLICE_X7Y121_A1 = CLBLM_R_X5Y122_SLICE_X7Y122_DQ;
  assign CLBLM_R_X5Y121_SLICE_X7Y121_A2 = CLBLM_R_X5Y123_SLICE_X6Y123_BQ;
  assign CLBLM_R_X5Y121_SLICE_X7Y121_A3 = CLBLM_R_X5Y121_SLICE_X7Y121_AQ;
  assign CLBLM_R_X5Y121_SLICE_X7Y121_A4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X5Y121_SLICE_X7Y121_A5 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X5Y121_SLICE_X7Y121_A6 = 1'b1;
  assign CLBLM_L_X12Y121_SLICE_X17Y121_D2 = 1'b1;
  assign CLBLM_R_X7Y128_SLICE_X8Y128_A2 = CLBLM_L_X8Y117_SLICE_X11Y117_BQ;
  assign CLBLM_R_X5Y121_SLICE_X7Y121_B1 = RIOB33_X105Y131_IOB_X1Y131_I;
  assign CLBLM_R_X5Y121_SLICE_X7Y121_B2 = RIOB33_X105Y133_IOB_X1Y133_I;
  assign CLBLM_R_X5Y121_SLICE_X7Y121_B3 = RIOB33_X105Y133_IOB_X1Y134_I;
  assign CLBLM_R_X5Y121_SLICE_X7Y121_B4 = RIOB33_X105Y131_IOB_X1Y132_I;
  assign CLBLM_R_X5Y121_SLICE_X7Y121_B5 = CLBLM_L_X8Y118_SLICE_X10Y118_BQ;
  assign CLBLM_R_X5Y121_SLICE_X7Y121_B6 = CLBLM_R_X3Y122_SLICE_X3Y122_AO6;
  assign CLBLM_R_X3Y111_SLICE_X3Y111_A1 = CLBLL_L_X2Y113_SLICE_X1Y113_C5Q;
  assign CLBLM_R_X3Y111_SLICE_X3Y111_A2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X3Y111_SLICE_X3Y111_A3 = CLBLM_R_X3Y111_SLICE_X3Y111_AQ;
  assign CLBLM_R_X3Y111_SLICE_X3Y111_A4 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X3Y111_SLICE_X3Y111_A5 = CLBLL_L_X4Y110_SLICE_X4Y110_DQ;
  assign CLBLM_R_X3Y111_SLICE_X3Y111_A6 = 1'b1;
  assign CLBLM_R_X5Y121_SLICE_X7Y121_C1 = CLBLM_R_X5Y121_SLICE_X6Y121_AQ;
  assign CLBLM_R_X5Y121_SLICE_X7Y121_C2 = RIOB33_X105Y133_IOB_X1Y133_I;
  assign CLBLM_R_X5Y121_SLICE_X7Y121_C3 = RIOB33_X105Y133_IOB_X1Y134_I;
  assign CLBLM_R_X3Y111_SLICE_X3Y111_B1 = 1'b1;
  assign CLBLM_L_X12Y121_SLICE_X17Y121_D3 = 1'b1;
  assign CLBLM_R_X3Y111_SLICE_X3Y111_B2 = CLBLM_R_X3Y111_SLICE_X3Y111_BQ;
  assign CLBLM_R_X3Y111_SLICE_X3Y111_B3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X3Y111_SLICE_X3Y111_B4 = CLBLM_R_X3Y113_SLICE_X3Y113_BO6;
  assign CLBLM_R_X3Y111_SLICE_X3Y111_B5 = CLBLM_L_X10Y117_SLICE_X13Y117_BQ;
  assign CLBLM_L_X10Y120_SLICE_X12Y120_A1 = CLBLM_R_X3Y118_SLICE_X2Y118_AQ;
  assign CLBLM_R_X3Y111_SLICE_X3Y111_B6 = CLBLM_R_X5Y110_SLICE_X7Y110_BQ;
  assign CLBLM_R_X3Y111_SLICE_X3Y111_C1 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X10Y120_SLICE_X12Y120_A2 = CLBLM_L_X10Y121_SLICE_X13Y121_BQ;
  assign CLBLM_R_X3Y111_SLICE_X3Y111_C2 = CLBLM_L_X8Y112_SLICE_X10Y112_CQ;
  assign CLBLM_R_X3Y111_SLICE_X3Y111_C3 = CLBLM_R_X3Y116_SLICE_X3Y116_DO6;
  assign CLBLM_R_X3Y111_SLICE_X3Y111_C4 = CLBLM_R_X3Y119_SLICE_X2Y119_AO6;
  assign CLBLM_R_X3Y111_SLICE_X3Y111_C5 = CLBLM_R_X3Y111_SLICE_X3Y111_DO6;
  assign CLBLM_L_X10Y120_SLICE_X12Y120_A3 = CLBLM_L_X10Y120_SLICE_X12Y120_AQ;
  assign CLBLM_R_X3Y111_SLICE_X3Y111_C6 = CLBLL_L_X2Y112_SLICE_X1Y112_BQ;
  assign CLBLM_R_X3Y111_SLICE_X3Y111_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X5Y121_SLICE_X6Y121_A1 = CLBLM_R_X5Y117_SLICE_X6Y117_AQ;
  assign CLBLM_R_X5Y121_SLICE_X6Y121_A2 = CLBLM_R_X7Y114_SLICE_X8Y114_BQ;
  assign CLBLM_L_X10Y120_SLICE_X12Y120_A4 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_R_X5Y121_SLICE_X6Y121_A3 = CLBLM_R_X5Y121_SLICE_X6Y121_AQ;
  assign CLBLM_R_X5Y121_SLICE_X6Y121_A4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X3Y111_SLICE_X3Y111_D1 = CLBLM_R_X3Y115_SLICE_X3Y115_CQ;
  assign CLBLM_L_X12Y121_SLICE_X17Y121_D4 = 1'b1;
  assign CLBLM_L_X10Y120_SLICE_X12Y120_A5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X3Y111_SLICE_X3Y111_D2 = CLBLM_L_X8Y112_SLICE_X11Y112_AQ;
  assign CLBLM_R_X3Y111_SLICE_X3Y111_D3 = CLBLL_L_X4Y120_SLICE_X5Y120_DO6;
  assign CLBLM_R_X3Y111_SLICE_X3Y111_D4 = CLBLM_R_X7Y115_SLICE_X9Y115_C5Q;
  assign CLBLM_L_X10Y120_SLICE_X12Y120_A6 = CLBLM_R_X5Y115_SLICE_X7Y115_DO6;
  assign CLBLM_R_X3Y111_SLICE_X3Y111_D5 = CLBLL_L_X2Y120_SLICE_X1Y120_DO6;
  assign CLBLM_R_X3Y111_SLICE_X3Y111_D6 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X5Y121_SLICE_X6Y121_AX = CLBLM_R_X5Y123_SLICE_X6Y123_DO6;
  assign CLBLM_R_X5Y121_SLICE_X6Y121_B1 = CLBLM_R_X7Y122_SLICE_X9Y122_A5Q;
  assign CLBLM_R_X5Y121_SLICE_X6Y121_B2 = CLBLM_R_X5Y121_SLICE_X6Y121_BQ;
  assign CLBLM_R_X3Y111_SLICE_X2Y111_A1 = CLBLM_R_X5Y115_SLICE_X6Y115_CO6;
  assign CLBLM_R_X3Y111_SLICE_X2Y111_A2 = 1'b1;
  assign CLBLM_R_X3Y111_SLICE_X2Y111_A3 = CLBLM_R_X3Y111_SLICE_X2Y111_AQ;
  assign CLBLM_R_X3Y111_SLICE_X2Y111_A4 = CLBLM_R_X7Y124_SLICE_X8Y124_CQ;
  assign CLBLM_R_X3Y111_SLICE_X2Y111_A5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X3Y111_SLICE_X2Y111_A6 = CLBLL_L_X4Y111_SLICE_X5Y111_A5Q;
  assign CLBLM_R_X5Y121_SLICE_X6Y121_BX = CLBLM_R_X5Y121_SLICE_X6Y121_CO6;
  assign CLBLM_R_X5Y121_SLICE_X6Y121_C1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X5Y121_SLICE_X6Y121_C2 = CLBLM_R_X11Y121_SLICE_X14Y121_AQ;
  assign CLBLM_R_X5Y121_SLICE_X6Y121_C3 = CLBLM_R_X3Y116_SLICE_X2Y116_CO6;
  assign CLBLM_R_X3Y111_SLICE_X2Y111_B1 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X3Y111_SLICE_X2Y111_B2 = CLBLL_L_X4Y121_SLICE_X4Y121_BQ;
  assign CLBLM_R_X3Y111_SLICE_X2Y111_B3 = CLBLM_R_X3Y110_SLICE_X2Y110_AQ;
  assign CLBLM_R_X3Y111_SLICE_X2Y111_B4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X3Y111_SLICE_X2Y111_B5 = CLBLM_R_X3Y110_SLICE_X3Y110_AQ;
  assign CLBLM_R_X3Y111_SLICE_X2Y111_B6 = 1'b1;
  assign CLBLM_R_X5Y121_SLICE_X6Y121_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X5Y121_SLICE_X6Y121_D1 = CLBLM_R_X5Y117_SLICE_X6Y117_AQ;
  assign CLBLM_R_X3Y111_SLICE_X2Y111_C1 = CLBLM_R_X3Y120_SLICE_X3Y120_BO6;
  assign CLBLM_L_X10Y120_SLICE_X12Y120_B1 = CLBLM_R_X3Y118_SLICE_X2Y118_AQ;
  assign CLBLM_R_X3Y111_SLICE_X2Y111_C2 = CLBLM_R_X3Y111_SLICE_X3Y111_AO5;
  assign CLBLM_R_X3Y111_SLICE_X2Y111_C3 = CLBLM_R_X3Y117_SLICE_X2Y117_BO5;
  assign CLBLM_R_X3Y111_SLICE_X2Y111_C4 = CLBLL_L_X4Y120_SLICE_X4Y120_BO6;
  assign CLBLM_R_X3Y111_SLICE_X2Y111_C5 = CLBLM_R_X3Y111_SLICE_X2Y111_BO5;
  assign CLBLM_L_X10Y120_SLICE_X12Y120_B2 = CLBLM_L_X10Y120_SLICE_X12Y120_BQ;
  assign CLBLM_R_X3Y111_SLICE_X2Y111_C6 = CLBLL_L_X4Y120_SLICE_X5Y120_DO6;
  assign CLBLM_R_X5Y121_SLICE_X6Y121_D4 = CLBLM_R_X3Y121_SLICE_X2Y121_AO6;
  assign CLBLM_R_X3Y111_SLICE_X2Y111_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X5Y121_SLICE_X6Y121_D6 = CLBLL_L_X4Y121_SLICE_X4Y121_CO6;
  assign CLBLM_L_X10Y120_SLICE_X12Y120_B3 = CLBLM_L_X10Y120_SLICE_X12Y120_DQ;
  assign CLBLM_L_X10Y120_SLICE_X12Y120_B4 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_R_X3Y111_SLICE_X2Y111_D2 = 1'b1;
  assign CLBLM_R_X3Y111_SLICE_X2Y111_D3 = 1'b1;
  assign CLBLM_R_X3Y111_SLICE_X2Y111_D1 = 1'b1;
  assign CLBLM_R_X3Y111_SLICE_X2Y111_D4 = 1'b1;
  assign CLBLM_R_X3Y111_SLICE_X2Y111_D5 = 1'b1;
  assign CLBLM_L_X10Y120_SLICE_X12Y120_B5 = CLBLM_R_X7Y120_SLICE_X9Y120_BQ;
  assign CLBLM_L_X12Y121_SLICE_X17Y121_D6 = 1'b1;
  assign CLBLM_R_X3Y111_SLICE_X2Y111_D6 = 1'b1;
  assign CLBLM_L_X10Y120_SLICE_X12Y120_B6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y128_SLICE_X8Y128_C4 = 1'b1;
  assign CLBLM_R_X7Y128_SLICE_X8Y128_C5 = 1'b1;
  assign CLBLM_R_X7Y128_SLICE_X8Y128_C6 = 1'b1;
  assign CLBLM_L_X10Y120_SLICE_X12Y120_C1 = CLBLM_R_X11Y119_SLICE_X14Y119_AO6;
  assign LIOB33_X0Y131_IOB_X0Y132_O = CLBLM_R_X7Y128_SLICE_X8Y128_AQ;
  assign LIOB33_X0Y131_IOB_X0Y131_O = CLBLM_R_X7Y128_SLICE_X8Y128_AO5;
  assign CLBLM_L_X8Y122_SLICE_X11Y122_D4 = CLBLM_R_X7Y123_SLICE_X9Y123_BO5;
  assign CLBLM_L_X10Y120_SLICE_X12Y120_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X8Y122_SLICE_X10Y122_A3 = CLBLM_L_X10Y124_SLICE_X12Y124_AQ;
  assign CLBLM_R_X103Y177_SLICE_X163Y177_A1 = 1'b1;
  assign CLBLM_R_X103Y177_SLICE_X163Y177_A2 = RIOB33_X105Y143_IOB_X1Y143_I;
  assign CLBLM_R_X103Y177_SLICE_X163Y177_A3 = CLBLM_R_X11Y119_SLICE_X14Y119_AQ;
  assign CLBLM_R_X103Y177_SLICE_X163Y177_A4 = 1'b1;
  assign CLBLM_R_X103Y177_SLICE_X163Y177_A5 = CLBLM_L_X12Y115_SLICE_X16Y115_BQ;
  assign CLBLM_R_X103Y177_SLICE_X163Y177_A6 = 1'b1;
  assign CLBLM_L_X8Y122_SLICE_X10Y122_A5 = CLBLM_R_X5Y120_SLICE_X6Y120_A5Q;
  assign CLBLM_R_X103Y177_SLICE_X163Y177_B1 = 1'b1;
  assign CLBLM_R_X103Y177_SLICE_X163Y177_B2 = 1'b1;
  assign CLBLM_R_X103Y177_SLICE_X163Y177_B3 = 1'b1;
  assign CLBLM_R_X103Y177_SLICE_X163Y177_B4 = 1'b1;
  assign CLBLM_R_X103Y177_SLICE_X163Y177_B5 = 1'b1;
  assign CLBLM_L_X10Y120_SLICE_X12Y120_D3 = CLBLM_L_X10Y120_SLICE_X12Y120_DQ;
  assign CLBLM_R_X103Y177_SLICE_X163Y177_B6 = 1'b1;
  assign CLBLM_L_X10Y120_SLICE_X12Y120_D4 = CLBLM_L_X12Y119_SLICE_X17Y119_AO5;
  assign CLBLM_R_X103Y177_SLICE_X163Y177_C1 = 1'b1;
  assign CLBLM_R_X103Y177_SLICE_X163Y177_C2 = 1'b1;
  assign CLBLM_R_X103Y177_SLICE_X163Y177_C3 = 1'b1;
  assign CLBLM_R_X103Y177_SLICE_X163Y177_C4 = 1'b1;
  assign CLBLM_R_X103Y177_SLICE_X163Y177_C5 = 1'b1;
  assign CLBLM_R_X103Y177_SLICE_X163Y177_C6 = 1'b1;
  assign CLBLM_L_X10Y120_SLICE_X12Y120_D6 = CLBLM_L_X10Y121_SLICE_X12Y121_AQ;
  assign CLBLM_R_X103Y177_SLICE_X163Y177_D1 = 1'b1;
  assign CLBLM_R_X103Y177_SLICE_X163Y177_D2 = 1'b1;
  assign CLBLM_R_X103Y177_SLICE_X163Y177_D3 = 1'b1;
  assign CLBLM_R_X103Y177_SLICE_X163Y177_D4 = 1'b1;
  assign CLBLM_R_X103Y177_SLICE_X163Y177_D5 = 1'b1;
  assign CLBLM_R_X103Y177_SLICE_X163Y177_D6 = 1'b1;
  assign LIOI3_X0Y147_OLOGIC_X0Y148_D1 = LIOB33_X0Y61_IOB_X0Y61_I;
  assign CLBLM_R_X103Y177_SLICE_X162Y177_A1 = 1'b1;
  assign CLBLM_R_X103Y177_SLICE_X162Y177_A2 = 1'b1;
  assign CLBLM_R_X103Y177_SLICE_X162Y177_A3 = 1'b1;
  assign CLBLM_R_X103Y177_SLICE_X162Y177_A4 = 1'b1;
  assign CLBLM_R_X103Y177_SLICE_X162Y177_A5 = 1'b1;
  assign CLBLM_R_X103Y177_SLICE_X162Y177_A6 = 1'b1;
  assign CLBLM_L_X8Y122_SLICE_X10Y122_B3 = RIOB33_X105Y129_IOB_X1Y130_I;
  assign LIOI3_X0Y147_OLOGIC_X0Y148_T1 = 1'b1;
  assign RIOI3_X105Y191_OLOGIC_X1Y192_D1 = CLBLM_L_X12Y115_SLICE_X16Y115_AQ;
  assign CLBLM_R_X103Y177_SLICE_X162Y177_B1 = 1'b1;
  assign CLBLM_R_X103Y177_SLICE_X162Y177_B2 = 1'b1;
  assign CLBLM_R_X103Y177_SLICE_X162Y177_B3 = 1'b1;
  assign CLBLM_R_X103Y177_SLICE_X162Y177_B4 = 1'b1;
  assign CLBLM_R_X103Y177_SLICE_X162Y177_B5 = 1'b1;
  assign CLBLM_R_X103Y177_SLICE_X162Y177_B6 = 1'b1;
  assign LIOI3_X0Y147_OLOGIC_X0Y147_D1 = LIOB33_X0Y71_IOB_X0Y71_I;
  assign RIOI3_X105Y191_OLOGIC_X1Y192_T1 = 1'b1;
  assign CLBLM_R_X103Y177_SLICE_X162Y177_C1 = 1'b1;
  assign CLBLM_R_X103Y177_SLICE_X162Y177_C2 = 1'b1;
  assign CLBLM_R_X103Y177_SLICE_X162Y177_C3 = 1'b1;
  assign CLBLM_R_X103Y177_SLICE_X162Y177_C4 = 1'b1;
  assign CLBLM_R_X103Y177_SLICE_X162Y177_C5 = 1'b1;
  assign CLBLM_R_X103Y177_SLICE_X162Y177_C6 = 1'b1;
  assign LIOI3_X0Y147_OLOGIC_X0Y147_T1 = 1'b1;
  assign RIOI3_X105Y191_OLOGIC_X1Y191_D1 = CLBLM_L_X8Y116_SLICE_X10Y116_AQ;
  assign CLBLM_R_X103Y177_SLICE_X162Y177_D1 = 1'b1;
  assign CLBLM_R_X103Y177_SLICE_X162Y177_D2 = 1'b1;
  assign CLBLM_R_X103Y177_SLICE_X162Y177_D3 = 1'b1;
  assign CLBLM_R_X103Y177_SLICE_X162Y177_D4 = 1'b1;
  assign CLBLM_R_X103Y177_SLICE_X162Y177_D5 = 1'b1;
  assign CLBLM_R_X103Y177_SLICE_X162Y177_D6 = 1'b1;
  assign RIOI3_X105Y191_OLOGIC_X1Y191_T1 = 1'b1;
  assign CLBLM_R_X5Y122_SLICE_X7Y122_A1 = 1'b1;
  assign CLBLM_R_X5Y122_SLICE_X7Y122_A2 = CLBLM_R_X3Y120_SLICE_X3Y120_BO6;
  assign CLBLM_R_X5Y122_SLICE_X7Y122_A3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X5Y122_SLICE_X7Y122_A4 = CLBLM_L_X8Y120_SLICE_X10Y120_CQ;
  assign CLBLM_R_X5Y122_SLICE_X7Y122_A5 = CLBLL_L_X4Y119_SLICE_X4Y119_C5Q;
  assign CLBLM_R_X5Y122_SLICE_X7Y122_A6 = 1'b1;
  assign CLBLM_R_X5Y122_SLICE_X7Y122_B1 = CLBLM_L_X8Y121_SLICE_X11Y121_DQ;
  assign CLBLM_R_X5Y122_SLICE_X7Y122_B2 = CLBLM_R_X5Y122_SLICE_X7Y122_BQ;
  assign CLBLM_R_X5Y122_SLICE_X7Y122_B3 = CLBLM_R_X5Y122_SLICE_X7Y122_AQ;
  assign CLBLM_R_X5Y122_SLICE_X7Y122_B4 = 1'b1;
  assign CLBLM_R_X5Y122_SLICE_X7Y122_B5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X5Y122_SLICE_X7Y122_B6 = CLBLM_R_X11Y121_SLICE_X14Y121_CO6;
  assign LIOB33_X0Y101_IOB_X0Y102_O = CLBLL_L_X2Y111_SLICE_X0Y111_AO5;
  assign CLBLM_R_X3Y112_SLICE_X3Y112_A1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X3Y112_SLICE_X3Y112_A2 = CLBLM_R_X3Y113_SLICE_X3Y113_BO6;
  assign CLBLM_L_X8Y122_SLICE_X10Y122_C4 = CLBLM_L_X10Y124_SLICE_X13Y124_BO6;
  assign CLBLM_R_X3Y112_SLICE_X3Y112_A3 = CLBLM_R_X3Y112_SLICE_X3Y112_AQ;
  assign CLBLM_R_X3Y112_SLICE_X3Y112_A4 = CLBLM_R_X3Y111_SLICE_X3Y111_BQ;
  assign CLBLM_R_X3Y112_SLICE_X3Y112_A5 = CLBLM_R_X5Y110_SLICE_X7Y110_BQ;
  assign CLBLM_R_X3Y112_SLICE_X3Y112_A6 = CLBLM_R_X7Y115_SLICE_X8Y115_CQ;
  assign CLBLM_L_X8Y122_SLICE_X10Y122_C5 = CLBLM_L_X8Y122_SLICE_X10Y122_DO6;
  assign CLBLM_R_X5Y122_SLICE_X7Y122_C1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X3Y112_SLICE_X3Y112_B1 = CLBLL_L_X4Y111_SLICE_X5Y111_A5Q;
  assign CLBLM_R_X3Y112_SLICE_X3Y112_B2 = CLBLL_L_X2Y112_SLICE_X1Y112_AQ;
  assign CLBLM_R_X3Y112_SLICE_X3Y112_B3 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X3Y112_SLICE_X3Y112_B4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X3Y112_SLICE_X3Y112_B5 = CLBLM_R_X7Y113_SLICE_X9Y113_AQ;
  assign CLBLM_R_X3Y112_SLICE_X3Y112_B6 = 1'b1;
  assign CLBLM_R_X5Y122_SLICE_X7Y122_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X5Y122_SLICE_X7Y122_D1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X3Y112_SLICE_X3Y112_C1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X3Y112_SLICE_X3Y112_C2 = CLBLM_R_X3Y119_SLICE_X2Y119_AO6;
  assign CLBLM_R_X3Y112_SLICE_X3Y112_C3 = CLBLL_L_X4Y115_SLICE_X4Y115_AQ;
  assign CLBLM_R_X3Y112_SLICE_X3Y112_C4 = CLBLL_L_X2Y112_SLICE_X1Y112_AQ;
  assign CLBLM_R_X3Y112_SLICE_X3Y112_C5 = CLBLM_R_X3Y112_SLICE_X3Y112_DO6;
  assign CLBLM_R_X3Y112_SLICE_X3Y112_C6 = 1'b1;
  assign CLBLM_R_X5Y122_SLICE_X7Y122_D3 = CLBLM_R_X5Y122_SLICE_X7Y122_DQ;
  assign CLBLM_R_X5Y122_SLICE_X7Y122_D4 = CLBLM_R_X3Y116_SLICE_X2Y116_DO6;
  assign CLBLM_R_X3Y112_SLICE_X3Y112_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X5Y122_SLICE_X6Y122_A1 = RIOB33_X105Y121_IOB_X1Y121_I;
  assign CLBLM_R_X5Y122_SLICE_X6Y122_A3 = CLBLM_R_X5Y122_SLICE_X6Y122_AQ;
  assign CLBLM_R_X5Y122_SLICE_X6Y122_A4 = CLBLM_R_X3Y116_SLICE_X2Y116_CO6;
  assign CLBLM_R_X5Y122_SLICE_X6Y122_A5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X5Y122_SLICE_X6Y122_A6 = 1'b1;
  assign CLBLM_R_X3Y112_SLICE_X3Y112_D1 = CLBLM_R_X3Y112_SLICE_X3Y112_C5Q;
  assign CLBLM_R_X3Y112_SLICE_X3Y112_D2 = CLBLM_R_X3Y112_SLICE_X2Y112_CO6;
  assign CLBLM_R_X3Y112_SLICE_X3Y112_D3 = CLBLM_R_X3Y112_SLICE_X2Y112_BQ;
  assign CLBLM_R_X3Y112_SLICE_X3Y112_D4 = CLBLM_R_X3Y112_SLICE_X2Y112_AQ;
  assign CLBLM_R_X3Y112_SLICE_X3Y112_D5 = CLBLL_L_X2Y112_SLICE_X1Y112_A5Q;
  assign CLBLM_R_X3Y112_SLICE_X3Y112_D6 = CLBLM_L_X10Y113_SLICE_X13Y113_BO6;
  assign CLBLM_R_X5Y122_SLICE_X6Y122_B1 = CLBLM_R_X3Y116_SLICE_X2Y116_DO6;
  assign CLBLM_R_X5Y122_SLICE_X6Y122_B2 = CLBLM_R_X5Y122_SLICE_X6Y122_BQ;
  assign CLBLM_R_X5Y122_SLICE_X6Y122_B3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X5Y122_SLICE_X6Y122_B4 = CLBLM_L_X8Y120_SLICE_X10Y120_D5Q;
  assign CLBLM_R_X5Y122_SLICE_X6Y122_B5 = 1'b1;
  assign CLBLM_R_X3Y112_SLICE_X2Y112_A1 = CLBLM_R_X3Y112_SLICE_X2Y112_DO6;
  assign CLBLM_R_X3Y112_SLICE_X2Y112_A2 = CLBLM_R_X7Y110_SLICE_X9Y110_CQ;
  assign CLBLM_R_X3Y112_SLICE_X2Y112_A3 = CLBLM_R_X3Y112_SLICE_X2Y112_AQ;
  assign CLBLM_R_X3Y112_SLICE_X2Y112_A4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X3Y112_SLICE_X2Y112_A5 = 1'b1;
  assign CLBLM_R_X3Y112_SLICE_X2Y112_A6 = CLBLL_L_X2Y112_SLICE_X1Y112_CO5;
  assign CLBLM_R_X5Y122_SLICE_X6Y122_C1 = CLBLM_R_X3Y122_SLICE_X3Y122_AO6;
  assign CLBLM_R_X5Y122_SLICE_X6Y122_C2 = CLBLL_L_X4Y123_SLICE_X5Y123_AO6;
  assign CLBLM_R_X5Y122_SLICE_X6Y122_C3 = RIOB33_X105Y131_IOB_X1Y131_I;
  assign CLBLM_R_X3Y112_SLICE_X2Y112_B1 = CLBLM_R_X3Y112_SLICE_X2Y112_DO6;
  assign CLBLM_R_X3Y112_SLICE_X2Y112_B2 = CLBLM_R_X3Y112_SLICE_X2Y112_BQ;
  assign CLBLM_R_X3Y112_SLICE_X2Y112_B3 = CLBLM_R_X3Y112_SLICE_X2Y112_AQ;
  assign CLBLM_R_X3Y112_SLICE_X2Y112_B4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X3Y112_SLICE_X2Y112_B5 = CLBLM_R_X11Y116_SLICE_X14Y116_AQ;
  assign CLBLM_R_X3Y112_SLICE_X2Y112_B6 = CLBLL_L_X2Y112_SLICE_X1Y112_CO5;
  assign CLBLM_R_X5Y122_SLICE_X6Y122_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X5Y122_SLICE_X6Y122_D1 = CLBLM_R_X3Y122_SLICE_X3Y122_AO6;
  assign CLBLM_R_X5Y122_SLICE_X6Y122_D2 = CLBLM_R_X7Y118_SLICE_X8Y118_AQ;
  assign CLBLM_R_X3Y112_SLICE_X2Y112_C1 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X3Y112_SLICE_X2Y112_C2 = CLBLM_R_X7Y113_SLICE_X9Y113_A5Q;
  assign CLBLM_R_X3Y112_SLICE_X2Y112_C3 = CLBLM_R_X7Y115_SLICE_X9Y115_C5Q;
  assign CLBLM_R_X3Y112_SLICE_X2Y112_C4 = CLBLM_R_X7Y120_SLICE_X9Y120_DQ;
  assign CLBLM_R_X3Y112_SLICE_X2Y112_C5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X3Y112_SLICE_X2Y112_C6 = CLBLM_R_X3Y115_SLICE_X3Y115_CQ;
  assign CLBLM_R_X5Y122_SLICE_X6Y122_D3 = CLBLL_L_X4Y123_SLICE_X5Y123_AO6;
  assign CLBLM_R_X5Y122_SLICE_X6Y122_D4 = CLBLM_R_X11Y121_SLICE_X14Y121_AQ;
  assign CLBLM_R_X5Y122_SLICE_X6Y122_D5 = RIOB33_X105Y131_IOB_X1Y131_I;
  assign CLBLM_R_X3Y112_SLICE_X2Y112_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X5Y122_SLICE_X6Y122_D6 = CLBLM_R_X3Y124_SLICE_X2Y124_BO6;
  assign CLBLM_R_X3Y112_SLICE_X2Y112_D1 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X3Y112_SLICE_X2Y112_D2 = CLBLM_R_X7Y120_SLICE_X9Y120_DQ;
  assign CLBLM_R_X3Y112_SLICE_X2Y112_D3 = CLBLM_R_X7Y113_SLICE_X9Y113_A5Q;
  assign CLBLM_R_X3Y112_SLICE_X2Y112_D4 = CLBLM_R_X3Y115_SLICE_X3Y115_CQ;
  assign CLBLM_R_X3Y112_SLICE_X2Y112_D5 = CLBLM_R_X7Y115_SLICE_X9Y115_C5Q;
  assign CLBLM_R_X3Y112_SLICE_X2Y112_D6 = 1'b1;
  assign LIOB33_X0Y133_IOB_X0Y134_O = CLBLM_R_X7Y124_SLICE_X8Y124_BQ;
  assign LIOB33_X0Y133_IOB_X0Y133_O = CLBLM_R_X7Y124_SLICE_X8Y124_A5Q;
  assign RIOI3_X105Y129_ILOGIC_X1Y130_D = RIOB33_X105Y129_IOB_X1Y130_I;
  assign RIOI3_X105Y129_ILOGIC_X1Y129_D = RIOB33_X105Y129_IOB_X1Y129_I;
  assign LIOI3_X0Y177_OLOGIC_X0Y178_D1 = RIOB33_X105Y129_IOB_X1Y130_I;
  assign CLBLM_L_X10Y110_SLICE_X13Y110_D6 = 1'b1;
  assign RIOI3_TBYTESRC_X105Y143_ILOGIC_X1Y144_D = RIOB33_X105Y143_IOB_X1Y144_I;
  assign RIOB33_X105Y177_IOB_X1Y178_O = CLBLM_R_X103Y177_SLICE_X163Y177_AO5;
  assign RIOI3_TBYTESRC_X105Y143_ILOGIC_X1Y143_D = RIOB33_X105Y143_IOB_X1Y143_I;
  assign CLBLM_L_X8Y112_SLICE_X11Y112_B1 = CLBLL_L_X4Y110_SLICE_X5Y110_AQ;
  assign CLBLM_L_X8Y112_SLICE_X11Y112_B2 = CLBLL_L_X4Y110_SLICE_X5Y110_BQ;
  assign CLBLM_L_X8Y112_SLICE_X11Y112_B3 = CLBLM_L_X8Y110_SLICE_X10Y110_BQ;
  assign CLBLM_L_X8Y112_SLICE_X11Y112_B4 = CLBLM_L_X10Y112_SLICE_X13Y112_CQ;
  assign LIOI3_X0Y79_OLOGIC_X0Y80_D1 = CLBLL_L_X2Y111_SLICE_X0Y111_AO6;
  assign CLBLM_L_X8Y112_SLICE_X11Y112_B5 = CLBLM_R_X7Y110_SLICE_X8Y110_CQ;
  assign CLBLM_L_X8Y112_SLICE_X11Y112_B6 = 1'b1;
  assign CLBLM_R_X5Y120_SLICE_X7Y120_C4 = 1'b1;
  assign CLBLM_R_X5Y120_SLICE_X7Y120_C5 = CLBLM_R_X3Y116_SLICE_X2Y116_DO6;
  assign CLBLM_R_X5Y120_SLICE_X7Y120_C6 = CLBLM_L_X10Y120_SLICE_X12Y120_CQ;
  assign CLBLM_L_X8Y112_SLICE_X11Y112_C1 = CLBLM_L_X10Y111_SLICE_X12Y111_AO5;
  assign CLBLM_L_X8Y112_SLICE_X11Y112_C2 = CLBLM_R_X5Y111_SLICE_X7Y111_DO6;
  assign CLBLM_L_X8Y112_SLICE_X11Y112_C3 = CLBLM_L_X8Y115_SLICE_X11Y115_CQ;
  assign CLBLM_L_X8Y112_SLICE_X11Y112_C4 = CLBLM_R_X7Y112_SLICE_X9Y112_BQ;
  assign CLBLM_L_X8Y112_SLICE_X11Y112_C5 = CLBLM_L_X8Y110_SLICE_X10Y110_AQ;
  assign CLBLM_R_X5Y123_SLICE_X7Y123_A1 = CLBLM_R_X7Y123_SLICE_X8Y123_CQ;
  assign CLBLM_L_X8Y112_SLICE_X11Y112_C6 = CLBLM_L_X8Y112_SLICE_X11Y112_BO6;
  assign CLBLM_R_X5Y123_SLICE_X7Y123_A2 = 1'b1;
  assign CLBLM_R_X5Y123_SLICE_X7Y123_A3 = CLBLM_R_X5Y123_SLICE_X7Y123_AQ;
  assign CLBLM_R_X5Y123_SLICE_X7Y123_A4 = CLBLM_R_X7Y122_SLICE_X9Y122_BO6;
  assign CLBLM_R_X5Y123_SLICE_X7Y123_A5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X5Y123_SLICE_X7Y123_A6 = CLBLM_R_X7Y121_SLICE_X8Y121_DO6;
  assign LIOI3_X0Y79_OLOGIC_X0Y80_T1 = 1'b1;
  assign CLBLM_R_X5Y123_SLICE_X7Y123_B1 = 1'b1;
  assign CLBLM_R_X5Y123_SLICE_X7Y123_B2 = 1'b1;
  assign CLBLM_R_X5Y123_SLICE_X7Y123_B3 = 1'b1;
  assign CLBLM_R_X5Y123_SLICE_X7Y123_B4 = 1'b1;
  assign CLBLM_R_X5Y123_SLICE_X7Y123_B5 = 1'b1;
  assign CLBLM_R_X5Y120_SLICE_X7Y120_D2 = CLBLL_L_X4Y120_SLICE_X5Y120_DO6;
  assign CLBLM_L_X8Y112_SLICE_X11Y112_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X10Y110_SLICE_X12Y110_B5 = 1'b1;
  assign CLBLM_R_X5Y123_SLICE_X7Y123_B6 = 1'b1;
  assign CLBLM_R_X3Y113_SLICE_X3Y113_A1 = CLBLM_R_X3Y114_SLICE_X2Y114_DQ;
  assign CLBLM_R_X3Y113_SLICE_X3Y113_A2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y110_SLICE_X12Y110_B6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X3Y113_SLICE_X3Y113_A3 = CLBLM_R_X3Y113_SLICE_X3Y113_AQ;
  assign CLBLM_R_X3Y113_SLICE_X3Y113_A4 = CLBLL_L_X2Y112_SLICE_X1Y112_BQ;
  assign CLBLM_R_X3Y113_SLICE_X3Y113_A5 = CLBLM_R_X3Y117_SLICE_X3Y117_C5Q;
  assign CLBLM_R_X3Y113_SLICE_X3Y113_A6 = CLBLM_L_X8Y112_SLICE_X10Y112_CQ;
  assign CLBLM_R_X5Y120_SLICE_X7Y120_D3 = CLBLL_L_X2Y119_SLICE_X0Y119_BO6;
  assign CLBLM_R_X5Y120_SLICE_X7Y120_D4 = CLBLL_L_X2Y120_SLICE_X1Y120_DO6;
  assign CLBLM_R_X3Y113_SLICE_X3Y113_B1 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_R_X3Y113_SLICE_X3Y113_B2 = CLBLM_R_X3Y118_SLICE_X2Y118_AQ;
  assign CLBLM_R_X3Y113_SLICE_X3Y113_B3 = CLBLL_L_X4Y118_SLICE_X5Y118_AQ;
  assign CLBLM_R_X3Y113_SLICE_X3Y113_B4 = 1'b1;
  assign CLBLM_R_X3Y113_SLICE_X3Y113_B5 = CLBLM_R_X5Y116_SLICE_X6Y116_BQ;
  assign CLBLM_R_X3Y113_SLICE_X3Y113_B6 = 1'b1;
  assign CLBLM_R_X5Y120_SLICE_X7Y120_D5 = CLBLM_R_X3Y120_SLICE_X3Y120_BO6;
  assign CLBLM_R_X5Y123_SLICE_X7Y123_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X3Y113_SLICE_X3Y113_C1 = CLBLM_R_X3Y112_SLICE_X3Y112_AQ;
  assign CLBLM_R_X3Y113_SLICE_X3Y113_C2 = CLBLM_R_X3Y117_SLICE_X3Y117_C5Q;
  assign CLBLM_R_X3Y113_SLICE_X3Y113_C3 = CLBLM_R_X3Y114_SLICE_X2Y114_DQ;
  assign CLBLM_R_X3Y113_SLICE_X3Y113_C4 = CLBLM_R_X3Y113_SLICE_X2Y113_DO5;
  assign CLBLM_R_X3Y113_SLICE_X3Y113_C5 = CLBLM_R_X3Y113_SLICE_X3Y113_BO5;
  assign CLBLM_R_X3Y113_SLICE_X3Y113_C6 = CLBLM_R_X3Y113_SLICE_X2Y113_BQ;
  assign CLBLM_R_X5Y123_SLICE_X7Y123_D3 = 1'b1;
  assign CLBLM_R_X5Y123_SLICE_X7Y123_D4 = 1'b1;
  assign CLBLM_R_X3Y113_SLICE_X3Y113_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X5Y123_SLICE_X6Y123_A1 = CLBLM_R_X5Y125_SLICE_X6Y125_BO5;
  assign CLBLM_R_X5Y123_SLICE_X6Y123_A2 = CLBLM_R_X7Y124_SLICE_X8Y124_DO5;
  assign CLBLM_L_X8Y112_SLICE_X11Y112_D1 = 1'b1;
  assign CLBLM_R_X5Y123_SLICE_X6Y123_A3 = CLBLM_R_X5Y123_SLICE_X6Y123_AQ;
  assign CLBLM_R_X5Y123_SLICE_X6Y123_A4 = CLBLM_R_X3Y117_SLICE_X3Y117_AQ;
  assign CLBLM_R_X3Y113_SLICE_X3Y113_D1 = CLBLM_R_X3Y111_SLICE_X3Y111_BQ;
  assign CLBLM_R_X3Y113_SLICE_X3Y113_D2 = CLBLM_R_X3Y112_SLICE_X3Y112_AQ;
  assign CLBLM_R_X3Y113_SLICE_X3Y113_D3 = CLBLM_R_X3Y114_SLICE_X2Y114_DQ;
  assign CLBLM_R_X3Y113_SLICE_X3Y113_D4 = CLBLM_R_X3Y113_SLICE_X2Y113_DO5;
  assign CLBLM_R_X3Y113_SLICE_X3Y113_D5 = CLBLM_R_X3Y113_SLICE_X3Y113_BO5;
  assign CLBLM_R_X3Y113_SLICE_X3Y113_D6 = CLBLM_R_X3Y113_SLICE_X2Y113_BQ;
  assign CLBLM_L_X8Y112_SLICE_X11Y112_D3 = CLBLM_L_X10Y120_SLICE_X12Y120_BQ;
  assign CLBLM_R_X5Y123_SLICE_X6Y123_A6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X5Y123_SLICE_X6Y123_B1 = CLBLM_R_X7Y121_SLICE_X8Y121_DO6;
  assign CLBLM_L_X8Y112_SLICE_X11Y112_D4 = CLBLM_L_X8Y111_SLICE_X10Y111_CO6;
  assign CLBLM_R_X5Y123_SLICE_X6Y123_B2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X3Y113_SLICE_X2Y113_A1 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_R_X3Y113_SLICE_X2Y113_A2 = CLBLM_R_X5Y112_SLICE_X6Y112_DO6;
  assign CLBLM_R_X3Y113_SLICE_X2Y113_A3 = CLBLM_R_X3Y113_SLICE_X2Y113_AQ;
  assign CLBLM_L_X8Y112_SLICE_X11Y112_D5 = CLBLM_L_X8Y113_SLICE_X10Y113_BO6;
  assign CLBLM_R_X3Y113_SLICE_X2Y113_A4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X3Y113_SLICE_X2Y113_A5 = CLBLM_R_X3Y112_SLICE_X2Y112_BQ;
  assign CLBLM_R_X3Y113_SLICE_X2Y113_A6 = CLBLM_R_X3Y118_SLICE_X2Y118_AQ;
  assign CLBLM_L_X8Y112_SLICE_X11Y112_D6 = CLBLM_L_X8Y112_SLICE_X11Y112_AQ;
  assign CLBLM_R_X5Y123_SLICE_X6Y123_C1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X3Y113_SLICE_X2Y113_B1 = CLBLM_R_X3Y113_SLICE_X2Y113_DO6;
  assign CLBLM_R_X3Y113_SLICE_X2Y113_B2 = CLBLM_R_X3Y113_SLICE_X2Y113_BQ;
  assign CLBLM_R_X3Y113_SLICE_X2Y113_B3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X3Y113_SLICE_X2Y113_B4 = CLBLM_R_X5Y110_SLICE_X7Y110_BQ;
  assign CLBLM_R_X3Y113_SLICE_X2Y113_B5 = CLBLM_R_X3Y113_SLICE_X2Y113_CO5;
  assign CLBLM_R_X3Y113_SLICE_X2Y113_B6 = CLBLM_L_X8Y112_SLICE_X10Y112_CQ;
  assign CLBLM_R_X5Y123_SLICE_X6Y123_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X5Y123_SLICE_X6Y123_D1 = CLBLM_R_X5Y123_SLICE_X7Y123_AQ;
  assign CLBLM_R_X5Y123_SLICE_X6Y123_D2 = CLBLM_R_X7Y121_SLICE_X8Y121_DO6;
  assign CLBLM_R_X3Y113_SLICE_X2Y113_C1 = CLBLM_R_X5Y113_SLICE_X6Y113_BQ;
  assign CLBLM_R_X3Y113_SLICE_X2Y113_C2 = CLBLL_L_X4Y113_SLICE_X4Y113_CO6;
  assign CLBLM_R_X3Y113_SLICE_X2Y113_C3 = CLBLM_R_X3Y114_SLICE_X2Y114_DQ;
  assign CLBLM_R_X3Y113_SLICE_X2Y113_C4 = CLBLM_R_X3Y113_SLICE_X2Y113_BQ;
  assign CLBLM_R_X3Y113_SLICE_X2Y113_C5 = CLBLL_L_X4Y113_SLICE_X4Y113_AQ;
  assign CLBLM_R_X3Y113_SLICE_X2Y113_C6 = 1'b1;
  assign CLBLM_R_X5Y123_SLICE_X6Y123_D3 = CLBLM_R_X5Y123_SLICE_X6Y123_BQ;
  assign CLBLM_R_X5Y123_SLICE_X6Y123_D4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X3Y113_SLICE_X2Y113_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X5Y123_SLICE_X6Y123_D6 = 1'b1;
  assign CLBLM_R_X3Y113_SLICE_X2Y113_D1 = CLBLM_R_X5Y113_SLICE_X6Y113_BQ;
  assign CLBLM_R_X3Y113_SLICE_X2Y113_D2 = 1'b1;
  assign CLBLM_R_X3Y113_SLICE_X2Y113_D3 = CLBLL_L_X4Y113_SLICE_X4Y113_CO6;
  assign CLBLM_R_X3Y113_SLICE_X2Y113_D4 = 1'b1;
  assign CLBLM_R_X3Y113_SLICE_X2Y113_D5 = CLBLL_L_X4Y113_SLICE_X4Y113_AQ;
  assign CLBLM_R_X3Y113_SLICE_X2Y113_D6 = 1'b1;
  assign CLBLM_R_X5Y120_SLICE_X6Y120_B5 = CLBLL_L_X4Y117_SLICE_X5Y117_AQ;
  assign CLBLM_R_X5Y120_SLICE_X6Y120_B6 = CLBLM_R_X5Y115_SLICE_X6Y115_CO5;
  assign CLBLM_R_X5Y120_SLICE_X6Y120_C3 = CLBLL_L_X2Y120_SLICE_X0Y120_AO5;
  assign CLBLM_R_X5Y120_SLICE_X6Y120_C4 = CLBLM_R_X5Y117_SLICE_X7Y117_AQ;
  assign CLBLM_R_X5Y120_SLICE_X6Y120_C5 = CLBLM_L_X8Y118_SLICE_X10Y118_AQ;
  assign CLBLM_R_X5Y120_SLICE_X6Y120_C6 = 1'b1;
  assign CLBLM_L_X8Y112_SLICE_X10Y112_C6 = CLBLM_R_X3Y118_SLICE_X2Y118_AQ;
  assign CLBLM_R_X5Y120_SLICE_X6Y120_D6 = CLBLM_R_X3Y121_SLICE_X2Y121_AO6;
  assign CLBLM_L_X8Y112_SLICE_X10Y112_D1 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X8Y112_SLICE_X10Y112_D2 = 1'b1;
  assign CLBLM_R_X5Y124_SLICE_X7Y124_A1 = 1'b1;
  assign CLBLM_R_X5Y124_SLICE_X7Y124_A2 = 1'b1;
  assign CLBLM_R_X5Y124_SLICE_X7Y124_A3 = 1'b1;
  assign CLBLM_R_X5Y124_SLICE_X7Y124_A4 = 1'b1;
  assign CLBLM_R_X5Y124_SLICE_X7Y124_A5 = 1'b1;
  assign CLBLM_R_X5Y124_SLICE_X7Y124_A6 = 1'b1;
  assign CLBLM_R_X5Y124_SLICE_X7Y124_B1 = 1'b1;
  assign CLBLM_R_X5Y124_SLICE_X7Y124_B2 = 1'b1;
  assign CLBLM_R_X5Y124_SLICE_X7Y124_B3 = 1'b1;
  assign CLBLM_R_X5Y124_SLICE_X7Y124_B4 = 1'b1;
  assign CLBLM_R_X5Y124_SLICE_X7Y124_B5 = 1'b1;
  assign CLBLM_R_X5Y124_SLICE_X7Y124_B6 = 1'b1;
  assign CLBLM_R_X3Y114_SLICE_X3Y114_A1 = CLBLM_R_X3Y114_SLICE_X3Y114_CQ;
  assign CLBLM_R_X3Y114_SLICE_X3Y114_A2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X3Y114_SLICE_X3Y114_A3 = CLBLL_L_X4Y114_SLICE_X4Y114_DO6;
  assign CLBLM_R_X3Y114_SLICE_X3Y114_A4 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_R_X3Y114_SLICE_X3Y114_A5 = CLBLM_R_X3Y118_SLICE_X2Y118_AQ;
  assign CLBLM_R_X3Y114_SLICE_X3Y114_A6 = CLBLM_R_X3Y114_SLICE_X3Y114_AQ;
  assign CLBLM_R_X5Y124_SLICE_X7Y124_C1 = 1'b1;
  assign CLBLM_R_X5Y124_SLICE_X7Y124_C2 = 1'b1;
  assign CLBLM_R_X5Y124_SLICE_X7Y124_C3 = 1'b1;
  assign CLBLM_R_X3Y114_SLICE_X3Y114_B1 = CLBLL_L_X4Y119_SLICE_X4Y119_DQ;
  assign CLBLM_R_X3Y114_SLICE_X3Y114_B2 = CLBLM_R_X3Y117_SLICE_X3Y117_BQ;
  assign CLBLM_R_X3Y114_SLICE_X3Y114_B3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X3Y114_SLICE_X3Y114_B4 = CLBLM_R_X3Y115_SLICE_X2Y115_BQ;
  assign CLBLM_R_X3Y114_SLICE_X3Y114_B5 = CLBLM_R_X3Y113_SLICE_X3Y113_CO6;
  assign CLBLM_R_X3Y114_SLICE_X3Y114_B6 = CLBLM_R_X3Y111_SLICE_X3Y111_BQ;
  assign CLBLM_R_X5Y124_SLICE_X7Y124_D1 = 1'b1;
  assign CLBLM_R_X5Y124_SLICE_X7Y124_D2 = 1'b1;
  assign CLBLM_R_X3Y114_SLICE_X3Y114_C1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X3Y114_SLICE_X3Y114_C2 = CLBLM_L_X10Y113_SLICE_X13Y113_BO6;
  assign CLBLM_R_X3Y114_SLICE_X3Y114_C3 = CLBLM_R_X7Y119_SLICE_X8Y119_D5Q;
  assign CLBLM_R_X3Y114_SLICE_X3Y114_C4 = CLBLM_R_X11Y113_SLICE_X15Y113_BQ;
  assign CLBLM_R_X3Y114_SLICE_X3Y114_C5 = CLBLM_R_X3Y114_SLICE_X3Y114_CQ;
  assign CLBLM_R_X3Y114_SLICE_X3Y114_C6 = CLBLM_R_X5Y116_SLICE_X6Y116_BQ;
  assign CLBLM_R_X5Y124_SLICE_X7Y124_D3 = 1'b1;
  assign CLBLM_R_X5Y124_SLICE_X7Y124_D4 = 1'b1;
  assign CLBLM_R_X3Y114_SLICE_X3Y114_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X5Y124_SLICE_X6Y124_A1 = CLBLL_L_X4Y119_SLICE_X4Y119_C5Q;
  assign CLBLM_R_X5Y124_SLICE_X6Y124_A2 = CLBLM_L_X10Y122_SLICE_X13Y122_BQ;
  assign CLBLM_R_X5Y124_SLICE_X6Y124_A3 = CLBLM_R_X5Y124_SLICE_X6Y124_AQ;
  assign CLBLM_R_X5Y124_SLICE_X6Y124_A4 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X5Y124_SLICE_X6Y124_A5 = CLBLM_R_X5Y125_SLICE_X6Y125_DO6;
  assign CLBLM_R_X3Y114_SLICE_X3Y114_D1 = 1'b1;
  assign CLBLM_R_X3Y114_SLICE_X3Y114_D2 = 1'b1;
  assign CLBLM_R_X3Y114_SLICE_X3Y114_D3 = RIOB33_X105Y121_IOB_X1Y121_I;
  assign CLBLM_R_X3Y114_SLICE_X3Y114_D4 = CLBLM_R_X3Y114_SLICE_X3Y114_AQ;
  assign CLBLM_R_X3Y114_SLICE_X3Y114_D5 = CLBLM_R_X7Y115_SLICE_X8Y115_CQ;
  assign CLBLM_R_X3Y114_SLICE_X3Y114_D6 = 1'b1;
  assign CLBLM_R_X5Y124_SLICE_X6Y124_B2 = CLBLM_R_X5Y124_SLICE_X6Y124_BQ;
  assign CLBLM_R_X5Y124_SLICE_X6Y124_B3 = CLBLL_L_X4Y119_SLICE_X4Y119_C5Q;
  assign CLBLM_R_X5Y124_SLICE_X6Y124_B4 = CLBLM_R_X5Y125_SLICE_X6Y125_CO5;
  assign CLBLM_R_X5Y124_SLICE_X6Y124_B5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X5Y124_SLICE_X6Y124_B6 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X5Y124_SLICE_X6Y124_B1 = CLBLM_R_X5Y111_SLICE_X6Y111_AQ;
  assign CLBLM_R_X3Y114_SLICE_X2Y114_A1 = CLBLM_R_X5Y115_SLICE_X7Y115_AQ;
  assign CLBLM_R_X3Y114_SLICE_X2Y114_A2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X3Y114_SLICE_X2Y114_A3 = CLBLM_R_X11Y115_SLICE_X15Y115_AQ;
  assign CLBLM_R_X3Y114_SLICE_X2Y114_A4 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X3Y114_SLICE_X2Y114_A5 = CLBLL_L_X2Y114_SLICE_X1Y114_BO6;
  assign CLBLM_R_X3Y114_SLICE_X2Y114_A6 = 1'b1;
  assign CLBLM_R_X5Y124_SLICE_X6Y124_C1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X5Y124_SLICE_X6Y124_C2 = CLBLL_L_X4Y123_SLICE_X4Y123_BQ;
  assign CLBLM_R_X5Y124_SLICE_X6Y124_C3 = CLBLL_L_X4Y119_SLICE_X4Y119_C5Q;
  assign CLBLM_R_X3Y114_SLICE_X2Y114_B1 = 1'b1;
  assign CLBLM_R_X3Y114_SLICE_X2Y114_B2 = CLBLM_R_X3Y114_SLICE_X2Y114_BQ;
  assign CLBLM_R_X3Y114_SLICE_X2Y114_B3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X3Y114_SLICE_X2Y114_B4 = CLBLM_R_X3Y114_SLICE_X2Y114_CQ;
  assign CLBLM_R_X3Y114_SLICE_X2Y114_B5 = CLBLM_R_X3Y112_SLICE_X3Y112_BQ;
  assign CLBLM_R_X3Y114_SLICE_X2Y114_B6 = CLBLM_R_X5Y115_SLICE_X6Y115_CO6;
  assign CLBLM_R_X5Y124_SLICE_X6Y124_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X5Y124_SLICE_X6Y124_D1 = 1'b1;
  assign CLBLM_R_X5Y124_SLICE_X6Y124_D2 = 1'b1;
  assign CLBLM_R_X3Y114_SLICE_X2Y114_C1 = CLBLM_R_X7Y123_SLICE_X8Y123_AQ;
  assign CLBLM_R_X3Y114_SLICE_X2Y114_C2 = CLBLM_R_X3Y114_SLICE_X2Y114_CQ;
  assign CLBLM_R_X3Y114_SLICE_X2Y114_C3 = CLBLM_R_X5Y111_SLICE_X7Y111_DO6;
  assign CLBLM_R_X3Y114_SLICE_X2Y114_C4 = CLBLM_R_X3Y114_SLICE_X2Y114_AO5;
  assign CLBLM_R_X3Y114_SLICE_X2Y114_C5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X3Y114_SLICE_X2Y114_C6 = CLBLL_L_X2Y114_SLICE_X1Y114_BO5;
  assign CLBLM_R_X5Y124_SLICE_X6Y124_D3 = 1'b1;
  assign CLBLM_R_X5Y124_SLICE_X6Y124_D4 = 1'b1;
  assign CLBLM_R_X5Y124_SLICE_X6Y124_D5 = 1'b1;
  assign CLBLM_R_X3Y114_SLICE_X2Y114_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X5Y124_SLICE_X6Y124_D6 = 1'b1;
  assign LIOI3_X0Y151_OLOGIC_X0Y151_T1 = 1'b1;
  assign RIOI3_X105Y195_OLOGIC_X1Y195_D1 = CLBLM_R_X11Y119_SLICE_X14Y119_AQ;
  assign CLBLM_R_X3Y114_SLICE_X2Y114_D1 = CLBLM_R_X3Y113_SLICE_X2Y113_CO5;
  assign CLBLM_R_X3Y114_SLICE_X2Y114_D2 = CLBLM_R_X3Y113_SLICE_X2Y113_CO6;
  assign CLBLM_R_X3Y114_SLICE_X2Y114_D3 = CLBLM_R_X3Y114_SLICE_X2Y114_DQ;
  assign CLBLM_R_X3Y114_SLICE_X2Y114_D4 = CLBLM_R_X5Y110_SLICE_X7Y110_BQ;
  assign CLBLM_R_X3Y114_SLICE_X2Y114_D5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X3Y114_SLICE_X2Y114_D6 = CLBLL_L_X4Y118_SLICE_X5Y118_AQ;
  assign CLBLL_L_X4Y118_SLICE_X4Y118_A3 = CLBLL_L_X4Y118_SLICE_X4Y118_AQ;
  assign RIOI3_X105Y195_OLOGIC_X1Y195_T1 = 1'b1;
  assign CLBLL_L_X4Y118_SLICE_X4Y118_A4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign LIOI3_X0Y141_OLOGIC_X0Y142_T1 = 1'b1;
  assign CLBLL_L_X4Y118_SLICE_X4Y118_A5 = CLBLM_R_X5Y118_SLICE_X6Y118_AQ;
  assign CLBLL_L_X4Y118_SLICE_X4Y118_A6 = 1'b1;
  assign RIOI3_TBYTESRC_X105Y157_OLOGIC_X1Y158_D1 = CLBLM_R_X37Y119_SLICE_X56Y119_AO6;
  assign RIOI3_TBYTESRC_X105Y157_OLOGIC_X1Y158_T1 = 1'b1;
  assign RIOI3_TBYTESRC_X105Y157_OLOGIC_X1Y157_D1 = RIOB33_X105Y125_IOB_X1Y126_I;
  assign CLBLL_L_X4Y118_SLICE_X4Y118_B6 = CLBLM_R_X5Y121_SLICE_X6Y121_BQ;
  assign RIOI3_TBYTESRC_X105Y157_OLOGIC_X1Y157_T1 = 1'b1;
  assign LIOI3_X0Y141_OLOGIC_X0Y141_D1 = CLBLM_R_X5Y123_SLICE_X6Y123_AQ;
  assign CLBLL_L_X4Y118_SLICE_X4Y118_C1 = CLBLL_L_X4Y117_SLICE_X5Y117_BQ;
  assign CLBLL_L_X4Y118_SLICE_X4Y118_C4 = CLBLM_R_X7Y118_SLICE_X9Y118_BQ;
  assign CLBLL_L_X4Y118_SLICE_X4Y118_C6 = 1'b1;
  assign LIOI3_X0Y141_OLOGIC_X0Y141_T1 = 1'b1;
  assign CLBLL_L_X4Y118_SLICE_X4Y118_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign RIOB33_X105Y155_IOB_X1Y156_O = RIOB33_X105Y103_IOB_X1Y104_I;
  assign RIOB33_X105Y155_IOB_X1Y155_O = RIOB33_X105Y103_IOB_X1Y103_I;
  assign RIOI3_X105Y127_ILOGIC_X1Y127_D = RIOB33_X105Y127_IOB_X1Y127_I;
  assign CLBLL_L_X4Y118_SLICE_X4Y118_D4 = CLBLM_R_X3Y121_SLICE_X2Y121_AO5;
  assign RIOI3_X105Y133_ILOGIC_X1Y134_D = RIOB33_X105Y133_IOB_X1Y134_I;
  assign LIOI3_TBYTESRC_X0Y143_OLOGIC_X0Y143_D1 = LIOB33_X0Y55_IOB_X0Y55_I;
  assign RIOI3_X105Y133_ILOGIC_X1Y133_D = RIOB33_X105Y133_IOB_X1Y133_I;
  assign CLBLL_L_X4Y118_SLICE_X4Y118_D6 = CLBLM_R_X5Y118_SLICE_X6Y118_AQ;
  assign CLBLM_R_X5Y125_SLICE_X7Y125_A1 = 1'b1;
  assign CLBLM_R_X5Y125_SLICE_X7Y125_A2 = 1'b1;
  assign CLBLM_R_X5Y125_SLICE_X7Y125_A3 = 1'b1;
  assign CLBLM_R_X5Y125_SLICE_X7Y125_A4 = 1'b1;
  assign CLBLM_R_X5Y125_SLICE_X7Y125_A5 = 1'b1;
  assign CLBLM_R_X5Y125_SLICE_X7Y125_A6 = 1'b1;
  assign CLBLM_R_X5Y125_SLICE_X7Y125_B1 = 1'b1;
  assign CLBLM_R_X5Y125_SLICE_X7Y125_B2 = 1'b1;
  assign CLBLM_R_X5Y125_SLICE_X7Y125_B3 = 1'b1;
  assign CLBLM_R_X5Y125_SLICE_X7Y125_B4 = 1'b1;
  assign CLBLM_R_X5Y125_SLICE_X7Y125_B5 = 1'b1;
  assign CLBLM_R_X5Y125_SLICE_X7Y125_B6 = 1'b1;
  assign CLBLM_R_X3Y115_SLICE_X3Y115_A1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X3Y115_SLICE_X3Y115_A2 = CLBLL_L_X4Y111_SLICE_X4Y111_AO5;
  assign CLBLM_R_X3Y115_SLICE_X3Y115_A3 = CLBLM_R_X3Y120_SLICE_X3Y120_BO6;
  assign CLBLM_R_X3Y115_SLICE_X3Y115_A4 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X3Y115_SLICE_X3Y115_A5 = CLBLL_L_X4Y112_SLICE_X4Y112_BQ;
  assign CLBLM_R_X3Y115_SLICE_X3Y115_A6 = CLBLM_R_X3Y115_SLICE_X3Y115_AQ;
  assign CLBLM_R_X5Y125_SLICE_X7Y125_C1 = 1'b1;
  assign CLBLM_R_X5Y125_SLICE_X7Y125_C2 = 1'b1;
  assign CLBLM_R_X5Y125_SLICE_X7Y125_C3 = 1'b1;
  assign CLBLM_R_X3Y115_SLICE_X3Y115_B1 = 1'b1;
  assign CLBLM_R_X3Y115_SLICE_X3Y115_B2 = CLBLM_R_X3Y115_SLICE_X3Y115_BQ;
  assign CLBLM_R_X3Y115_SLICE_X3Y115_B3 = CLBLL_L_X4Y111_SLICE_X5Y111_BQ;
  assign CLBLM_R_X3Y115_SLICE_X3Y115_B4 = CLBLM_R_X5Y115_SLICE_X6Y115_CO6;
  assign CLBLM_R_X3Y115_SLICE_X3Y115_B5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X3Y115_SLICE_X3Y115_B6 = CLBLM_R_X3Y116_SLICE_X3Y116_A5Q;
  assign CLBLM_L_X10Y126_SLICE_X12Y126_AX = CLBLM_R_X11Y128_SLICE_X14Y128_AO6;
  assign CLBLM_R_X5Y125_SLICE_X7Y125_D1 = 1'b1;
  assign CLBLM_R_X3Y115_SLICE_X3Y115_C1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X3Y115_SLICE_X3Y115_C2 = CLBLM_R_X3Y112_SLICE_X2Y112_BQ;
  assign CLBLM_R_X3Y115_SLICE_X3Y115_C3 = CLBLL_L_X4Y115_SLICE_X4Y115_C5Q;
  assign CLBLM_R_X3Y115_SLICE_X3Y115_C4 = CLBLM_R_X3Y112_SLICE_X3Y112_C5Q;
  assign CLBLM_R_X3Y115_SLICE_X3Y115_C5 = CLBLL_L_X2Y112_SLICE_X1Y112_A5Q;
  assign CLBLM_R_X3Y115_SLICE_X3Y115_C6 = CLBLM_R_X3Y112_SLICE_X2Y112_AQ;
  assign CLBLM_R_X5Y125_SLICE_X7Y125_D3 = 1'b1;
  assign CLBLM_R_X5Y125_SLICE_X7Y125_D4 = 1'b1;
  assign CLBLM_R_X3Y115_SLICE_X3Y115_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X5Y125_SLICE_X6Y125_A1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X5Y125_SLICE_X6Y125_A2 = CLBLM_L_X8Y119_SLICE_X10Y119_A5Q;
  assign CLBLM_R_X5Y125_SLICE_X6Y125_A3 = CLBLM_R_X5Y125_SLICE_X6Y125_AQ;
  assign CLBLM_R_X5Y125_SLICE_X6Y125_A4 = CLBLL_L_X4Y119_SLICE_X4Y119_C5Q;
  assign CLBLM_R_X5Y125_SLICE_X6Y125_A5 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X3Y115_SLICE_X3Y115_D1 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X3Y115_SLICE_X3Y115_D2 = CLBLM_R_X3Y117_SLICE_X3Y117_A5Q;
  assign CLBLM_R_X3Y115_SLICE_X3Y115_D3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X3Y115_SLICE_X3Y115_D4 = 1'b1;
  assign CLBLM_R_X3Y115_SLICE_X3Y115_D5 = CLBLM_R_X3Y114_SLICE_X3Y114_DO6;
  assign CLBLM_R_X3Y115_SLICE_X3Y115_D6 = CLBLL_L_X4Y112_SLICE_X4Y112_BQ;
  assign CLBLM_R_X5Y125_SLICE_X6Y125_A6 = CLBLM_R_X5Y125_SLICE_X6Y125_CO6;
  assign CLBLM_R_X5Y125_SLICE_X6Y125_AX = CLBLM_R_X5Y125_SLICE_X6Y125_BO6;
  assign CLBLM_R_X5Y125_SLICE_X6Y125_B1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X5Y125_SLICE_X6Y125_B2 = CLBLM_R_X5Y124_SLICE_X6Y124_AQ;
  assign CLBLM_R_X5Y125_SLICE_X6Y125_B3 = CLBLM_R_X5Y125_SLICE_X6Y125_AQ;
  assign CLBLM_R_X5Y125_SLICE_X6Y125_B4 = CLBLM_R_X5Y123_SLICE_X6Y123_CQ;
  assign CLBLM_R_X3Y115_SLICE_X2Y115_A1 = 1'b1;
  assign CLBLM_R_X3Y115_SLICE_X2Y115_A2 = CLBLL_L_X4Y112_SLICE_X4Y112_BQ;
  assign CLBLM_R_X3Y115_SLICE_X2Y115_A3 = CLBLM_R_X3Y115_SLICE_X2Y115_AQ;
  assign CLBLM_R_X3Y115_SLICE_X2Y115_A4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X3Y115_SLICE_X2Y115_A5 = CLBLM_R_X5Y115_SLICE_X6Y115_CO5;
  assign CLBLM_R_X3Y115_SLICE_X2Y115_A6 = CLBLM_R_X3Y115_SLICE_X2Y115_DQ;
  assign CLBLM_R_X5Y125_SLICE_X6Y125_C1 = CLBLL_L_X4Y123_SLICE_X4Y123_AQ;
  assign CLBLM_R_X5Y125_SLICE_X6Y125_C2 = CLBLM_R_X7Y124_SLICE_X8Y124_A5Q;
  assign CLBLM_R_X5Y125_SLICE_X6Y125_C3 = CLBLM_R_X5Y124_SLICE_X6Y124_BQ;
  assign CLBLM_R_X3Y115_SLICE_X2Y115_B1 = 1'b1;
  assign CLBLM_R_X3Y115_SLICE_X2Y115_B2 = CLBLM_R_X3Y115_SLICE_X2Y115_BQ;
  assign CLBLM_R_X3Y115_SLICE_X2Y115_B3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X3Y115_SLICE_X2Y115_B4 = CLBLM_R_X5Y110_SLICE_X7Y110_BQ;
  assign CLBLM_R_X3Y115_SLICE_X2Y115_B5 = CLBLM_R_X3Y118_SLICE_X3Y118_AQ;
  assign CLBLM_R_X3Y115_SLICE_X2Y115_B6 = CLBLM_R_X3Y113_SLICE_X2Y113_CO6;
  assign CLBLM_R_X5Y125_SLICE_X6Y125_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X5Y125_SLICE_X6Y125_D1 = CLBLL_L_X4Y123_SLICE_X4Y123_AQ;
  assign CLBLM_R_X5Y125_SLICE_X6Y125_D2 = CLBLM_R_X5Y125_SLICE_X6Y125_AQ;
  assign CLBLM_R_X3Y115_SLICE_X2Y115_C1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X3Y115_SLICE_X2Y115_C2 = CLBLM_R_X3Y115_SLICE_X2Y115_CQ;
  assign CLBLM_R_X3Y115_SLICE_X2Y115_C3 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_R_X3Y115_SLICE_X2Y115_C4 = CLBLM_R_X3Y118_SLICE_X2Y118_AQ;
  assign CLBLM_R_X3Y115_SLICE_X2Y115_C5 = CLBLM_R_X7Y121_SLICE_X8Y121_C5Q;
  assign CLBLM_R_X3Y115_SLICE_X2Y115_C6 = CLBLM_R_X11Y115_SLICE_X14Y115_BQ;
  assign CLBLM_R_X5Y125_SLICE_X6Y125_D3 = CLBLM_R_X7Y124_SLICE_X8Y124_A5Q;
  assign CLBLM_R_X5Y125_SLICE_X6Y125_D4 = CLBLM_R_X7Y124_SLICE_X8Y124_CQ;
  assign CLBLM_R_X5Y125_SLICE_X6Y125_D5 = CLBLM_R_X7Y124_SLICE_X8Y124_BQ;
  assign CLBLM_R_X3Y115_SLICE_X2Y115_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X5Y125_SLICE_X6Y125_D6 = CLBLM_R_X5Y124_SLICE_X6Y124_BQ;
  assign RIOI3_X105Y121_ILOGIC_X1Y122_D = RIOB33_X105Y121_IOB_X1Y122_I;
  assign CLBLM_R_X3Y115_SLICE_X2Y115_D1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X3Y115_SLICE_X2Y115_D2 = CLBLM_R_X3Y113_SLICE_X2Y113_BQ;
  assign CLBLM_R_X3Y115_SLICE_X2Y115_D3 = CLBLM_L_X10Y113_SLICE_X13Y113_BO6;
  assign CLBLM_R_X3Y115_SLICE_X2Y115_D4 = CLBLM_R_X3Y115_SLICE_X2Y115_DQ;
  assign CLBLM_R_X3Y115_SLICE_X2Y115_D5 = CLBLM_R_X7Y119_SLICE_X8Y119_D5Q;
  assign CLBLM_R_X3Y115_SLICE_X2Y115_D6 = CLBLM_R_X5Y113_SLICE_X6Y113_BQ;
  assign RIOI3_X105Y121_ILOGIC_X1Y121_D = RIOB33_X105Y121_IOB_X1Y121_I;
  assign CLBLM_L_X10Y121_SLICE_X13Y121_C4 = CLBLM_R_X11Y121_SLICE_X14Y121_DO6;
  assign CLBLM_L_X10Y121_SLICE_X13Y121_C5 = 1'b1;
  assign CLBLM_L_X10Y121_SLICE_X13Y121_C6 = CLBLM_L_X10Y117_SLICE_X13Y117_CQ;
  assign CLBLM_L_X10Y121_SLICE_X13Y121_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X10Y121_SLICE_X13Y121_D1 = CLBLM_L_X8Y122_SLICE_X11Y122_BQ;
  assign CLBLM_L_X10Y121_SLICE_X13Y121_D2 = CLBLM_L_X10Y120_SLICE_X13Y120_AQ;
  assign CLBLM_L_X10Y121_SLICE_X13Y121_D3 = CLBLM_L_X10Y122_SLICE_X12Y122_CO6;
  assign CLBLM_L_X10Y121_SLICE_X13Y121_D4 = CLBLM_L_X10Y123_SLICE_X12Y123_CO6;
  assign LIOB33_X0Y141_IOB_X0Y142_O = LIOB33_X0Y53_IOB_X0Y54_I;
  assign CLBLL_L_X52Y126_SLICE_X79Y126_D3 = 1'b1;
  assign LIOB33_X0Y141_IOB_X0Y141_O = CLBLM_R_X5Y123_SLICE_X6Y123_AQ;
  assign CLBLM_L_X10Y121_SLICE_X13Y121_D5 = CLBLM_L_X10Y121_SLICE_X13Y121_CQ;
  assign CLBLM_L_X10Y121_SLICE_X13Y121_D6 = CLBLM_L_X8Y122_SLICE_X11Y122_DO6;
  assign CLBLM_R_X3Y116_SLICE_X3Y116_A1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X3Y116_SLICE_X3Y116_A2 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_R_X3Y116_SLICE_X3Y116_A3 = CLBLM_R_X3Y116_SLICE_X3Y116_AQ;
  assign CLBLM_R_X3Y116_SLICE_X3Y116_A4 = CLBLL_L_X4Y121_SLICE_X4Y121_BQ;
  assign CLBLM_R_X3Y116_SLICE_X3Y116_A5 = CLBLM_R_X3Y118_SLICE_X2Y118_AQ;
  assign CLBLM_R_X3Y116_SLICE_X3Y116_A6 = CLBLM_R_X11Y113_SLICE_X14Y113_BQ;
  assign CLBLM_R_X3Y116_SLICE_X3Y116_AX = CLBLM_L_X10Y116_SLICE_X13Y116_AO6;
  assign CLBLM_R_X3Y116_SLICE_X3Y116_B1 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X3Y116_SLICE_X3Y116_B2 = 1'b1;
  assign CLBLM_R_X3Y116_SLICE_X3Y116_B3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X3Y116_SLICE_X3Y116_B4 = 1'b1;
  assign CLBLM_R_X3Y116_SLICE_X3Y116_B5 = CLBLL_L_X2Y117_SLICE_X1Y117_AQ;
  assign CLBLM_R_X3Y116_SLICE_X3Y116_B6 = CLBLM_R_X5Y115_SLICE_X7Y115_BQ;
  assign CLBLM_R_X3Y116_SLICE_X3Y116_C1 = CLBLL_L_X4Y114_SLICE_X5Y114_AQ;
  assign CLBLM_R_X3Y116_SLICE_X3Y116_C2 = CLBLM_R_X3Y116_SLICE_X3Y116_CQ;
  assign CLBLM_R_X3Y116_SLICE_X3Y116_C3 = CLBLM_R_X3Y116_SLICE_X2Y116_DO6;
  assign CLBLM_R_X3Y116_SLICE_X3Y116_C4 = CLBLM_R_X5Y119_SLICE_X6Y119_B5Q;
  assign CLBLM_R_X3Y116_SLICE_X3Y116_C5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X3Y116_SLICE_X3Y116_C6 = 1'b1;
  assign CLBLM_L_X10Y121_SLICE_X12Y121_A1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign LIOI3_SING_X0Y100_OLOGIC_X0Y100_D1 = CLBLL_L_X2Y111_SLICE_X0Y111_BO6;
  assign CLBLM_R_X3Y116_SLICE_X3Y116_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X10Y121_SLICE_X12Y121_A2 = CLBLM_L_X8Y122_SLICE_X11Y122_BQ;
  assign CLBLM_R_X3Y116_SLICE_X3Y116_D1 = CLBLL_L_X2Y119_SLICE_X0Y119_BO6;
  assign CLBLM_L_X10Y121_SLICE_X12Y121_A3 = CLBLM_L_X10Y121_SLICE_X12Y121_AQ;
  assign CLBLM_R_X3Y116_SLICE_X3Y116_D2 = CLBLM_R_X7Y113_SLICE_X9Y113_A5Q;
  assign CLBLM_R_X3Y116_SLICE_X3Y116_D3 = CLBLM_R_X3Y120_SLICE_X3Y120_BO6;
  assign CLBLM_R_X3Y116_SLICE_X3Y116_D4 = CLBLM_R_X5Y124_SLICE_X6Y124_CQ;
  assign CLBLM_R_X3Y116_SLICE_X3Y116_D5 = 1'b1;
  assign CLBLM_L_X10Y121_SLICE_X12Y121_A4 = CLBLM_R_X7Y123_SLICE_X9Y123_CO6;
  assign CLBLM_R_X3Y116_SLICE_X3Y116_D6 = 1'b1;
  assign LIOI3_SING_X0Y100_OLOGIC_X0Y100_T1 = 1'b1;
  assign CLBLM_L_X10Y121_SLICE_X12Y121_A5 = CLBLM_L_X10Y123_SLICE_X12Y123_AO6;
  assign CLBLM_R_X3Y116_SLICE_X2Y116_A1 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X3Y116_SLICE_X2Y116_A2 = LIOB33_X0Y53_IOB_X0Y53_I;
  assign CLBLM_R_X3Y116_SLICE_X2Y116_A3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y121_SLICE_X12Y121_A6 = CLBLM_R_X7Y120_SLICE_X8Y120_CQ;
  assign CLBLM_R_X3Y116_SLICE_X2Y116_A4 = CLBLL_L_X4Y121_SLICE_X4Y121_BQ;
  assign CLBLM_R_X3Y116_SLICE_X2Y116_A5 = CLBLM_R_X3Y110_SLICE_X2Y110_AQ;
  assign CLBLM_R_X3Y116_SLICE_X2Y116_A6 = CLBLM_R_X11Y115_SLICE_X14Y115_BQ;
  assign CLBLM_R_X3Y116_SLICE_X2Y116_B1 = CLBLL_L_X4Y116_SLICE_X4Y116_CQ;
  assign CLBLM_R_X3Y116_SLICE_X2Y116_B2 = CLBLM_R_X3Y116_SLICE_X2Y116_BQ;
  assign CLBLM_R_X3Y116_SLICE_X2Y116_B3 = CLBLM_R_X5Y111_SLICE_X6Y111_CQ;
  assign CLBLM_R_X3Y116_SLICE_X2Y116_B4 = 1'b1;
  assign CLBLM_R_X3Y116_SLICE_X2Y116_B5 = CLBLM_R_X5Y115_SLICE_X6Y115_CO6;
  assign CLBLM_R_X3Y116_SLICE_X2Y116_B6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y123_SLICE_X12Y123_C1 = CLBLM_L_X10Y124_SLICE_X12Y124_AQ;
  assign CLBLM_R_X3Y116_SLICE_X2Y116_C1 = CLBLM_R_X3Y110_SLICE_X2Y110_AQ;
  assign CLBLM_R_X3Y116_SLICE_X2Y116_C2 = LIOB33_X0Y53_IOB_X0Y53_I;
  assign CLBLM_R_X3Y116_SLICE_X2Y116_C3 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X3Y116_SLICE_X2Y116_C4 = CLBLM_R_X3Y117_SLICE_X3Y117_A5Q;
  assign CLBLM_R_X3Y116_SLICE_X2Y116_C5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X3Y116_SLICE_X2Y116_C6 = CLBLL_L_X4Y121_SLICE_X4Y121_BQ;
  assign CLBLM_R_X3Y116_SLICE_X2Y116_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X10Y121_SLICE_X12Y121_B1 = CLBLM_L_X8Y116_SLICE_X11Y116_DQ;
  assign CLBLM_L_X10Y121_SLICE_X12Y121_B2 = CLBLM_L_X10Y121_SLICE_X12Y121_BQ;
  assign CLBLM_R_X3Y116_SLICE_X2Y116_D1 = CLBLL_L_X2Y113_SLICE_X1Y113_C5Q;
  assign CLBLM_R_X3Y116_SLICE_X2Y116_D2 = CLBLL_L_X2Y114_SLICE_X1Y114_BO5;
  assign CLBLM_R_X3Y116_SLICE_X2Y116_D3 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X10Y123_SLICE_X12Y123_C2 = CLBLM_R_X7Y123_SLICE_X9Y123_BO5;
  assign CLBLM_L_X10Y121_SLICE_X12Y121_B3 = CLBLM_L_X10Y121_SLICE_X12Y121_AQ;
  assign CLBLM_R_X3Y116_SLICE_X2Y116_D4 = CLBLM_L_X8Y116_SLICE_X10Y116_AO6;
  assign CLBLM_R_X3Y116_SLICE_X2Y116_D5 = CLBLM_R_X3Y117_SLICE_X2Y117_BO5;
  assign CLBLM_R_X3Y116_SLICE_X2Y116_D6 = CLBLM_R_X5Y111_SLICE_X7Y111_DO6;
  assign CLBLM_L_X10Y121_SLICE_X12Y121_B4 = CLBLM_L_X10Y123_SLICE_X12Y123_AO6;
  assign CLBLM_L_X10Y121_SLICE_X12Y121_B5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y121_SLICE_X12Y121_B6 = CLBLM_R_X7Y123_SLICE_X9Y123_CO6;
  assign CLBLM_L_X10Y123_SLICE_X12Y123_C3 = CLBLM_R_X5Y120_SLICE_X6Y120_A5Q;
  assign CLBLM_L_X10Y121_SLICE_X12Y121_C1 = CLBLM_L_X10Y121_SLICE_X13Y121_CQ;
  assign CLBLM_L_X10Y121_SLICE_X12Y121_C2 = CLBLM_L_X10Y121_SLICE_X12Y121_AQ;
  assign CLBLM_L_X8Y123_SLICE_X11Y123_D3 = 1'b1;
  assign CLBLM_L_X10Y121_SLICE_X12Y121_C3 = CLBLM_L_X10Y123_SLICE_X12Y123_CO6;
  assign CLBLM_L_X10Y121_SLICE_X12Y121_C4 = CLBLM_L_X10Y120_SLICE_X13Y120_AQ;
  assign CLBLM_L_X8Y123_SLICE_X11Y123_D5 = 1'b1;
  assign LIOI3_X0Y153_OLOGIC_X0Y154_D1 = LIOB33_X0Y67_IOB_X0Y68_I;
  assign CLBLM_L_X10Y121_SLICE_X12Y121_C5 = CLBLM_L_X10Y122_SLICE_X12Y122_CO6;
  assign CLBLM_L_X8Y123_SLICE_X11Y123_D6 = 1'b1;
  assign CLBLM_L_X10Y121_SLICE_X12Y121_C6 = CLBLM_L_X8Y122_SLICE_X11Y122_DO6;
  assign CLBLM_L_X10Y123_SLICE_X12Y123_C5 = CLBLM_L_X10Y118_SLICE_X12Y118_B5Q;
  assign LIOI3_X0Y153_OLOGIC_X0Y154_T1 = 1'b1;
  assign RIOI3_X105Y197_OLOGIC_X1Y198_D1 = CLBLM_L_X8Y122_SLICE_X10Y122_BO5;
  assign LIOI3_X0Y153_OLOGIC_X0Y153_D1 = LIOB33_X0Y67_IOB_X0Y67_I;
  assign RIOI3_X105Y197_OLOGIC_X1Y198_T1 = 1'b1;
  assign LIOI3_X0Y153_OLOGIC_X0Y153_T1 = 1'b1;
  assign RIOI3_X105Y197_OLOGIC_X1Y197_D1 = CLBLM_L_X8Y122_SLICE_X10Y122_BO5;
  assign RIOI3_X105Y197_OLOGIC_X1Y197_T1 = 1'b1;
  assign RIOI3_TBYTESRC_X105Y169_OLOGIC_X1Y170_D1 = CLBLM_R_X103Y169_SLICE_X163Y169_AO5;
  assign CLBLM_L_X10Y121_SLICE_X12Y121_D5 = CLBLM_L_X8Y121_SLICE_X11Y121_DQ;
  assign RIOI3_TBYTESRC_X105Y169_OLOGIC_X1Y170_T1 = 1'b1;
  assign RIOI3_TBYTESRC_X105Y169_OLOGIC_X1Y169_D1 = CLBLM_R_X103Y169_SLICE_X163Y169_AO6;
  assign LIOB33_X0Y143_IOB_X0Y143_O = LIOB33_X0Y55_IOB_X0Y55_I;
  assign CLBLM_L_X8Y123_SLICE_X10Y123_B4 = 1'b1;
  assign RIOI3_TBYTESRC_X105Y169_OLOGIC_X1Y169_T1 = 1'b1;
  assign CLBLM_R_X3Y117_SLICE_X3Y117_A1 = CLBLM_R_X5Y116_SLICE_X7Y116_A5Q;
  assign CLBLM_R_X3Y117_SLICE_X3Y117_A2 = CLBLM_R_X3Y116_SLICE_X2Y116_AQ;
  assign CLBLM_R_X3Y117_SLICE_X3Y117_A3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X3Y117_SLICE_X3Y117_A4 = CLBLM_R_X7Y121_SLICE_X8Y121_AQ;
  assign CLBLM_R_X3Y117_SLICE_X3Y117_A5 = CLBLM_R_X3Y117_SLICE_X2Y117_AQ;
  assign CLBLM_R_X3Y117_SLICE_X3Y117_A6 = 1'b1;
  assign CLBLM_R_X3Y117_SLICE_X3Y117_B1 = RIOB33_X105Y119_IOB_X1Y119_I;
  assign CLBLM_R_X3Y117_SLICE_X3Y117_B2 = CLBLM_R_X3Y117_SLICE_X3Y117_BQ;
  assign CLBLM_R_X3Y117_SLICE_X3Y117_B3 = CLBLM_R_X3Y117_SLICE_X3Y117_CQ;
  assign CLBLM_R_X3Y117_SLICE_X3Y117_B4 = CLBLM_R_X3Y112_SLICE_X2Y112_AQ;
  assign CLBLM_R_X3Y117_SLICE_X3Y117_B5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X3Y117_SLICE_X3Y117_B6 = 1'b1;
  assign CLBLM_R_X3Y117_SLICE_X3Y117_C1 = CLBLM_R_X3Y117_SLICE_X3Y117_C5Q;
  assign CLBLM_R_X3Y117_SLICE_X3Y117_C2 = RIOB33_X105Y119_IOB_X1Y119_I;
  assign CLBLM_R_X3Y117_SLICE_X3Y117_C3 = CLBLM_L_X8Y114_SLICE_X10Y114_C5Q;
  assign CLBLM_R_X3Y117_SLICE_X3Y117_C4 = CLBLM_R_X5Y114_SLICE_X6Y114_CQ;
  assign CLBLM_R_X3Y117_SLICE_X3Y117_C5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X3Y117_SLICE_X3Y117_C6 = 1'b1;
  assign CLBLM_R_X3Y117_SLICE_X3Y117_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X3Y117_SLICE_X3Y117_D1 = CLBLM_R_X3Y115_SLICE_X3Y115_BQ;
  assign CLBLM_R_X3Y117_SLICE_X3Y117_D2 = CLBLM_R_X3Y122_SLICE_X3Y122_AO5;
  assign CLBLM_R_X3Y117_SLICE_X3Y117_D3 = RIOB33_X105Y135_IOB_X1Y136_I;
  assign CLBLM_R_X3Y117_SLICE_X3Y117_D4 = CLBLM_R_X3Y117_SLICE_X2Y117_AQ;
  assign CLBLM_R_X3Y117_SLICE_X3Y117_D5 = CLBLL_L_X2Y121_SLICE_X1Y121_BO5;
  assign CLBLM_R_X3Y117_SLICE_X3Y117_D6 = RIOB33_X105Y135_IOB_X1Y135_I;
  assign CLBLM_R_X3Y117_SLICE_X2Y117_A1 = CLBLM_L_X10Y113_SLICE_X13Y113_BO6;
  assign CLBLM_R_X3Y117_SLICE_X2Y117_A2 = CLBLM_R_X7Y128_SLICE_X8Y128_AQ;
  assign CLBLM_R_X3Y117_SLICE_X2Y117_A3 = CLBLM_R_X3Y117_SLICE_X2Y117_AQ;
  assign CLBLM_R_X3Y117_SLICE_X2Y117_A4 = CLBLM_R_X7Y119_SLICE_X8Y119_D5Q;
  assign CLBLM_R_X3Y117_SLICE_X2Y117_A5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X3Y117_SLICE_X2Y117_A6 = CLBLM_R_X3Y114_SLICE_X2Y114_DQ;
  assign CLBLM_R_X3Y117_SLICE_X2Y117_B1 = CLBLL_L_X2Y113_SLICE_X1Y113_C5Q;
  assign CLBLM_R_X3Y117_SLICE_X2Y117_B2 = CLBLL_L_X2Y117_SLICE_X0Y117_A5Q;
  assign CLBLM_R_X3Y117_SLICE_X2Y117_B3 = CLBLM_R_X7Y121_SLICE_X8Y121_C5Q;
  assign CLBLM_R_X3Y117_SLICE_X2Y117_B4 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X3Y117_SLICE_X2Y117_B5 = CLBLM_R_X5Y115_SLICE_X7Y115_AQ;
  assign CLBLM_R_X3Y117_SLICE_X2Y117_B6 = 1'b1;
  assign RIOB33_X105Y179_IOB_X1Y180_O = CLBLM_R_X11Y113_SLICE_X15Y113_DO6;
  assign CLBLM_R_X3Y117_SLICE_X2Y117_C1 = CLBLM_R_X5Y116_SLICE_X6Y116_AQ;
  assign CLBLM_R_X3Y117_SLICE_X2Y117_C2 = CLBLM_R_X3Y114_SLICE_X3Y114_CQ;
  assign CLBLM_R_X3Y117_SLICE_X2Y117_C3 = CLBLM_R_X3Y122_SLICE_X3Y122_AO5;
  assign CLBLM_R_X3Y117_SLICE_X2Y117_C4 = CLBLL_L_X2Y120_SLICE_X1Y120_AO6;
  assign CLBLM_R_X3Y117_SLICE_X2Y117_C5 = RIOB33_X105Y135_IOB_X1Y136_I;
  assign CLBLM_R_X3Y117_SLICE_X2Y117_C6 = RIOB33_X105Y135_IOB_X1Y135_I;
  assign LIOI3_X0Y123_OLOGIC_X0Y123_T1 = 1'b1;
  assign LIOI3_SING_X0Y149_OLOGIC_X0Y149_D1 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign RIOI3_X105Y135_ILOGIC_X1Y136_D = RIOB33_X105Y135_IOB_X1Y136_I;
  assign CLBLM_R_X3Y117_SLICE_X2Y117_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X7Y119_SLICE_X9Y119_C4 = 1'b1;
  assign RIOI3_X105Y135_ILOGIC_X1Y135_D = RIOB33_X105Y135_IOB_X1Y135_I;
  assign CLBLM_R_X7Y119_SLICE_X9Y119_C5 = 1'b1;
  assign CLBLM_R_X3Y117_SLICE_X2Y117_D1 = CLBLL_L_X2Y120_SLICE_X1Y120_AO6;
  assign CLBLM_R_X3Y117_SLICE_X2Y117_D2 = CLBLL_L_X4Y114_SLICE_X4Y114_AQ;
  assign CLBLM_R_X3Y117_SLICE_X2Y117_D3 = CLBLM_R_X3Y122_SLICE_X3Y122_AO6;
  assign CLBLM_R_X3Y117_SLICE_X2Y117_D4 = CLBLL_L_X2Y121_SLICE_X1Y121_BO6;
  assign CLBLM_R_X3Y117_SLICE_X2Y117_D5 = 1'b1;
  assign CLBLM_R_X3Y117_SLICE_X2Y117_D6 = CLBLM_R_X3Y114_SLICE_X2Y114_BQ;
  assign CLBLM_R_X7Y119_SLICE_X9Y119_C6 = CLBLM_R_X5Y120_SLICE_X7Y120_CQ;
  assign LIOI3_SING_X0Y149_OLOGIC_X0Y149_T1 = 1'b1;
  assign CLBLM_R_X7Y119_SLICE_X9Y119_D2 = CLBLM_R_X7Y118_SLICE_X8Y118_DQ;
  assign CLBLM_R_X7Y119_SLICE_X9Y119_D5 = CLBLM_R_X3Y117_SLICE_X3Y117_BQ;
  assign CLBLM_R_X7Y119_SLICE_X9Y119_D6 = 1'b1;
  assign CLBLM_L_X8Y113_SLICE_X11Y113_A2 = CLBLM_L_X8Y112_SLICE_X10Y112_BQ;
  assign CLBLM_L_X8Y113_SLICE_X11Y113_A3 = CLBLM_L_X8Y113_SLICE_X11Y113_AQ;
  assign CLBLM_L_X8Y113_SLICE_X11Y113_B1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign LIOB33_X0Y145_IOB_X0Y146_O = LIOB33_X0Y59_IOB_X0Y59_I;
  assign LIOB33_X0Y145_IOB_X0Y145_O = LIOB33_X0Y57_IOB_X0Y58_I;
  assign CLBLM_L_X8Y113_SLICE_X11Y113_B2 = CLBLM_L_X8Y113_SLICE_X11Y113_BQ;
  assign CLBLM_L_X8Y113_SLICE_X11Y113_B3 = CLBLM_L_X8Y111_SLICE_X10Y111_AQ;
  assign CLBLM_L_X8Y113_SLICE_X11Y113_B4 = CLBLM_L_X10Y113_SLICE_X12Y113_DO6;
  assign CLBLM_L_X8Y113_SLICE_X11Y113_B5 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X5Y121_SLICE_X7Y121_C4 = CLBLM_R_X3Y122_SLICE_X3Y122_AO6;
  assign CLBLM_R_X5Y121_SLICE_X7Y121_C5 = RIOB33_X105Y131_IOB_X1Y131_I;
  assign RIOI3_X105Y171_OLOGIC_X1Y172_D1 = CLBLM_R_X103Y172_SLICE_X163Y172_AO6;
  assign CLBLM_R_X5Y121_SLICE_X7Y121_C6 = RIOB33_X105Y131_IOB_X1Y132_I;
  assign CLBLM_R_X5Y121_SLICE_X7Y121_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X7Y119_SLICE_X8Y119_B5 = 1'b1;
  assign CLBLM_L_X8Y113_SLICE_X11Y113_C2 = CLBLM_L_X8Y113_SLICE_X11Y113_CQ;
  assign CLBLM_R_X7Y119_SLICE_X8Y119_B6 = CLBLM_L_X10Y122_SLICE_X12Y122_AQ;
  assign CLBLM_L_X8Y113_SLICE_X11Y113_C3 = CLBLM_L_X8Y111_SLICE_X11Y111_AO6;
  assign CLBLM_L_X8Y113_SLICE_X11Y113_C4 = CLBLM_R_X11Y123_SLICE_X14Y123_CO6;
  assign CLBLM_L_X8Y113_SLICE_X11Y113_C5 = CLBLM_L_X10Y113_SLICE_X12Y113_CO6;
  assign CLBLM_L_X8Y113_SLICE_X11Y113_C6 = CLBLM_R_X5Y121_SLICE_X6Y121_CO5;
  assign CLBLM_L_X10Y111_SLICE_X12Y111_B3 = CLBLM_L_X8Y110_SLICE_X10Y110_BQ;
  assign CLBLM_R_X3Y118_SLICE_X3Y118_A1 = CLBLL_L_X4Y117_SLICE_X5Y117_DQ;
  assign CLBLM_R_X3Y118_SLICE_X3Y118_A2 = CLBLM_R_X11Y121_SLICE_X14Y121_CO6;
  assign CLBLM_L_X10Y111_SLICE_X12Y111_B4 = CLBLM_L_X10Y115_SLICE_X12Y115_BQ;
  assign CLBLM_R_X3Y118_SLICE_X3Y118_A3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X3Y118_SLICE_X3Y118_A4 = CLBLM_R_X3Y118_SLICE_X3Y118_AQ;
  assign CLBLM_R_X3Y118_SLICE_X3Y118_A5 = 1'b1;
  assign CLBLM_L_X8Y113_SLICE_X11Y113_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X3Y118_SLICE_X3Y118_A6 = CLBLL_L_X2Y112_SLICE_X1Y112_A5Q;
  assign CLBLM_L_X10Y111_SLICE_X12Y111_B5 = CLBLM_R_X7Y110_SLICE_X8Y110_CQ;
  assign CLBLM_R_X3Y118_SLICE_X3Y118_B1 = CLBLM_R_X3Y121_SLICE_X3Y121_CO6;
  assign CLBLM_R_X3Y118_SLICE_X3Y118_B2 = RIOB33_X105Y133_IOB_X1Y133_I;
  assign CLBLM_R_X3Y118_SLICE_X3Y118_B3 = CLBLL_L_X4Y117_SLICE_X5Y117_AQ;
  assign CLBLM_R_X3Y118_SLICE_X3Y118_B4 = CLBLM_R_X3Y110_SLICE_X3Y110_AQ;
  assign CLBLM_R_X3Y118_SLICE_X3Y118_B5 = RIOB33_X105Y131_IOB_X1Y131_I;
  assign CLBLM_R_X3Y118_SLICE_X3Y118_B6 = RIOB33_X105Y133_IOB_X1Y134_I;
  assign CLBLM_R_X5Y121_SLICE_X7Y121_D3 = CLBLM_R_X7Y121_SLICE_X8Y121_AQ;
  assign CLBLM_R_X5Y121_SLICE_X7Y121_D4 = CLBLM_R_X5Y123_SLICE_X6Y123_CQ;
  assign CLBLM_R_X3Y118_SLICE_X3Y118_C1 = CLBLM_R_X3Y115_SLICE_X3Y115_AQ;
  assign CLBLM_R_X3Y118_SLICE_X3Y118_C2 = 1'b1;
  assign CLBLM_R_X3Y118_SLICE_X3Y118_C3 = CLBLL_L_X2Y120_SLICE_X0Y120_AO5;
  assign CLBLM_R_X3Y118_SLICE_X3Y118_C4 = CLBLM_R_X3Y121_SLICE_X2Y121_AO6;
  assign CLBLM_R_X3Y118_SLICE_X3Y118_C5 = 1'b1;
  assign CLBLM_R_X3Y118_SLICE_X3Y118_C6 = CLBLM_R_X3Y118_SLICE_X3Y118_AQ;
  assign CLBLM_R_X5Y121_SLICE_X7Y121_D5 = 1'b1;
  assign CLBLM_R_X5Y121_SLICE_X7Y121_D6 = CLBLM_R_X5Y123_SLICE_X6Y123_BQ;
  assign CLBLM_R_X3Y118_SLICE_X3Y118_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X7Y119_SLICE_X8Y119_C5 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X7Y119_SLICE_X8Y119_C6 = 1'b1;
  assign CLBLM_R_X3Y118_SLICE_X3Y118_D1 = CLBLL_L_X2Y115_SLICE_X1Y115_AQ;
  assign CLBLM_R_X3Y118_SLICE_X3Y118_D2 = CLBLM_L_X10Y114_SLICE_X13Y114_D5Q;
  assign CLBLM_R_X3Y118_SLICE_X3Y118_D3 = 1'b1;
  assign CLBLM_R_X3Y118_SLICE_X3Y118_D4 = CLBLL_L_X4Y121_SLICE_X4Y121_CO6;
  assign CLBLM_R_X3Y118_SLICE_X3Y118_D5 = 1'b1;
  assign CLBLM_R_X3Y118_SLICE_X3Y118_D6 = CLBLM_R_X3Y121_SLICE_X2Y121_AO5;
  assign CLBLM_L_X8Y113_SLICE_X11Y113_D1 = CLBLM_L_X10Y113_SLICE_X12Y113_AO6;
  assign CLBLM_L_X8Y113_SLICE_X11Y113_D2 = CLBLM_L_X10Y114_SLICE_X12Y114_AO6;
  assign CLBLM_R_X3Y118_SLICE_X2Y118_A1 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_R_X3Y118_SLICE_X2Y118_A2 = RIOB33_X105Y119_IOB_X1Y119_I;
  assign CLBLM_R_X3Y118_SLICE_X2Y118_A3 = CLBLM_R_X3Y118_SLICE_X2Y118_AQ;
  assign CLBLM_L_X8Y113_SLICE_X11Y113_D3 = CLBLM_R_X7Y115_SLICE_X9Y115_B5Q;
  assign CLBLM_R_X3Y118_SLICE_X2Y118_A4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X3Y118_SLICE_X2Y118_A5 = CLBLL_L_X4Y118_SLICE_X4Y118_AQ;
  assign CLBLM_R_X3Y118_SLICE_X2Y118_A6 = CLBLM_R_X3Y117_SLICE_X3Y117_CQ;
  assign CLBLM_L_X8Y113_SLICE_X11Y113_D4 = CLBLM_L_X8Y115_SLICE_X11Y115_CQ;
  assign CLBLM_R_X3Y118_SLICE_X2Y118_B1 = CLBLM_R_X3Y122_SLICE_X3Y122_AO5;
  assign CLBLM_R_X3Y118_SLICE_X2Y118_B2 = CLBLM_R_X5Y118_SLICE_X7Y118_AQ;
  assign CLBLM_L_X8Y113_SLICE_X11Y113_D5 = CLBLM_R_X5Y119_SLICE_X7Y119_CO6;
  assign CLBLM_R_X3Y118_SLICE_X2Y118_B3 = RIOB33_X105Y135_IOB_X1Y135_I;
  assign CLBLM_R_X3Y118_SLICE_X2Y118_B4 = CLBLL_L_X4Y118_SLICE_X5Y118_CQ;
  assign CLBLM_R_X3Y118_SLICE_X2Y118_B5 = RIOB33_X105Y135_IOB_X1Y136_I;
  assign CLBLM_R_X3Y118_SLICE_X2Y118_B6 = CLBLL_L_X2Y120_SLICE_X1Y120_AO6;
  assign CLBLM_L_X8Y113_SLICE_X11Y113_D6 = CLBLL_L_X2Y119_SLICE_X1Y119_BO6;
  assign CLBLM_R_X3Y118_SLICE_X2Y118_C1 = CLBLL_L_X2Y121_SLICE_X1Y121_BO5;
  assign CLBLM_R_X3Y118_SLICE_X2Y118_C2 = 1'b1;
  assign CLBLM_R_X3Y118_SLICE_X2Y118_C3 = CLBLL_L_X4Y118_SLICE_X4Y118_AQ;
  assign CLBLM_R_X3Y118_SLICE_X2Y118_C4 = CLBLM_R_X3Y122_SLICE_X3Y122_AO6;
  assign CLBLM_R_X3Y118_SLICE_X2Y118_C5 = CLBLL_L_X4Y119_SLICE_X4Y119_AQ;
  assign CLBLM_R_X3Y118_SLICE_X2Y118_C6 = CLBLL_L_X2Y121_SLICE_X1Y121_BO6;
  assign RIOI3_X105Y145_ILOGIC_X1Y145_D = RIOB33_X105Y145_IOB_X1Y145_I;
  assign RIOI3_X105Y171_OLOGIC_X1Y171_D1 = CLBLM_L_X8Y128_SLICE_X10Y128_AO5;
  assign CLBLM_R_X3Y118_SLICE_X2Y118_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X3Y118_SLICE_X2Y118_D1 = CLBLL_L_X4Y120_SLICE_X5Y120_BO6;
  assign CLBLM_R_X3Y118_SLICE_X2Y118_D2 = CLBLL_L_X2Y119_SLICE_X1Y119_AO5;
  assign CLBLM_R_X3Y118_SLICE_X2Y118_D3 = 1'b1;
  assign CLBLM_R_X3Y118_SLICE_X2Y118_D4 = CLBLM_R_X3Y118_SLICE_X2Y118_CO6;
  assign CLBLM_R_X3Y118_SLICE_X2Y118_D5 = CLBLM_R_X5Y115_SLICE_X6Y115_AQ;
  assign CLBLM_R_X3Y118_SLICE_X2Y118_D6 = CLBLL_L_X2Y112_SLICE_X1Y112_A5Q;
  assign CLBLM_R_X5Y121_SLICE_X6Y121_A5 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X5Y121_SLICE_X6Y121_A6 = RIOB33_X105Y121_IOB_X1Y121_I;
  assign LIOI3_SING_X0Y150_OLOGIC_X0Y150_D1 = LIOB33_X0Y63_IOB_X0Y63_I;
  assign LIOI3_TBYTETERM_X0Y137_OLOGIC_X0Y137_T1 = 1'b1;
  assign RIOI3_X105Y171_OLOGIC_X1Y171_T1 = 1'b1;
  assign CLBLM_R_X5Y121_SLICE_X6Y121_B3 = CLBLM_R_X5Y115_SLICE_X6Y115_CO5;
  assign LIOI3_SING_X0Y150_OLOGIC_X0Y150_T1 = 1'b1;
  assign CLBLM_R_X5Y121_SLICE_X6Y121_B4 = 1'b1;
  assign CLBLM_R_X5Y121_SLICE_X6Y121_B5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X5Y121_SLICE_X6Y121_B6 = CLBLL_L_X4Y115_SLICE_X5Y115_BQ;
endmodule
