module top(
  input LIOB33_SING_X0Y100_IOB_X0Y100_IPAD,
  input LIOB33_SING_X0Y149_IOB_X0Y149_IPAD,
  input LIOB33_SING_X0Y150_IOB_X0Y150_IPAD,
  input LIOB33_SING_X0Y50_IOB_X0Y50_IPAD,
  input LIOB33_SING_X0Y99_IOB_X0Y99_IPAD,
  input LIOB33_X0Y101_IOB_X0Y101_IPAD,
  input LIOB33_X0Y101_IOB_X0Y102_IPAD,
  input LIOB33_X0Y103_IOB_X0Y103_IPAD,
  input LIOB33_X0Y103_IOB_X0Y104_IPAD,
  input LIOB33_X0Y105_IOB_X0Y105_IPAD,
  input LIOB33_X0Y105_IOB_X0Y106_IPAD,
  input LIOB33_X0Y107_IOB_X0Y107_IPAD,
  input LIOB33_X0Y107_IOB_X0Y108_IPAD,
  input LIOB33_X0Y109_IOB_X0Y109_IPAD,
  input LIOB33_X0Y109_IOB_X0Y110_IPAD,
  input LIOB33_X0Y111_IOB_X0Y111_IPAD,
  input LIOB33_X0Y111_IOB_X0Y112_IPAD,
  input LIOB33_X0Y113_IOB_X0Y113_IPAD,
  input LIOB33_X0Y113_IOB_X0Y114_IPAD,
  input LIOB33_X0Y115_IOB_X0Y115_IPAD,
  input LIOB33_X0Y115_IOB_X0Y116_IPAD,
  input LIOB33_X0Y117_IOB_X0Y117_IPAD,
  input LIOB33_X0Y117_IOB_X0Y118_IPAD,
  input LIOB33_X0Y119_IOB_X0Y119_IPAD,
  input LIOB33_X0Y119_IOB_X0Y120_IPAD,
  input LIOB33_X0Y121_IOB_X0Y121_IPAD,
  input LIOB33_X0Y121_IOB_X0Y122_IPAD,
  input LIOB33_X0Y123_IOB_X0Y123_IPAD,
  input LIOB33_X0Y123_IOB_X0Y124_IPAD,
  input LIOB33_X0Y125_IOB_X0Y125_IPAD,
  input LIOB33_X0Y125_IOB_X0Y126_IPAD,
  input LIOB33_X0Y127_IOB_X0Y127_IPAD,
  input LIOB33_X0Y127_IOB_X0Y128_IPAD,
  input LIOB33_X0Y129_IOB_X0Y129_IPAD,
  input LIOB33_X0Y129_IOB_X0Y130_IPAD,
  input LIOB33_X0Y131_IOB_X0Y131_IPAD,
  input LIOB33_X0Y131_IOB_X0Y132_IPAD,
  input LIOB33_X0Y133_IOB_X0Y133_IPAD,
  input LIOB33_X0Y133_IOB_X0Y134_IPAD,
  input LIOB33_X0Y135_IOB_X0Y135_IPAD,
  input LIOB33_X0Y135_IOB_X0Y136_IPAD,
  input LIOB33_X0Y137_IOB_X0Y137_IPAD,
  input LIOB33_X0Y137_IOB_X0Y138_IPAD,
  input LIOB33_X0Y139_IOB_X0Y139_IPAD,
  input LIOB33_X0Y139_IOB_X0Y140_IPAD,
  input LIOB33_X0Y141_IOB_X0Y141_IPAD,
  input LIOB33_X0Y141_IOB_X0Y142_IPAD,
  input LIOB33_X0Y143_IOB_X0Y143_IPAD,
  input LIOB33_X0Y145_IOB_X0Y145_IPAD,
  input LIOB33_X0Y145_IOB_X0Y146_IPAD,
  input LIOB33_X0Y147_IOB_X0Y147_IPAD,
  input LIOB33_X0Y147_IOB_X0Y148_IPAD,
  input LIOB33_X0Y151_IOB_X0Y151_IPAD,
  input LIOB33_X0Y151_IOB_X0Y152_IPAD,
  input LIOB33_X0Y153_IOB_X0Y153_IPAD,
  input LIOB33_X0Y153_IOB_X0Y154_IPAD,
  input LIOB33_X0Y155_IOB_X0Y155_IPAD,
  input LIOB33_X0Y155_IOB_X0Y156_IPAD,
  input LIOB33_X0Y157_IOB_X0Y157_IPAD,
  input LIOB33_X0Y157_IOB_X0Y158_IPAD,
  input LIOB33_X0Y159_IOB_X0Y159_IPAD,
  input LIOB33_X0Y159_IOB_X0Y160_IPAD,
  input LIOB33_X0Y161_IOB_X0Y161_IPAD,
  input LIOB33_X0Y161_IOB_X0Y162_IPAD,
  input LIOB33_X0Y163_IOB_X0Y163_IPAD,
  input LIOB33_X0Y163_IOB_X0Y164_IPAD,
  input LIOB33_X0Y165_IOB_X0Y165_IPAD,
  input LIOB33_X0Y165_IOB_X0Y166_IPAD,
  input LIOB33_X0Y167_IOB_X0Y167_IPAD,
  input LIOB33_X0Y167_IOB_X0Y168_IPAD,
  input LIOB33_X0Y169_IOB_X0Y169_IPAD,
  input LIOB33_X0Y169_IOB_X0Y170_IPAD,
  input LIOB33_X0Y171_IOB_X0Y171_IPAD,
  input LIOB33_X0Y171_IOB_X0Y172_IPAD,
  input LIOB33_X0Y173_IOB_X0Y173_IPAD,
  input LIOB33_X0Y173_IOB_X0Y174_IPAD,
  input LIOB33_X0Y175_IOB_X0Y175_IPAD,
  input LIOB33_X0Y175_IOB_X0Y176_IPAD,
  input LIOB33_X0Y177_IOB_X0Y177_IPAD,
  input LIOB33_X0Y51_IOB_X0Y51_IPAD,
  input LIOB33_X0Y51_IOB_X0Y52_IPAD,
  input LIOB33_X0Y53_IOB_X0Y53_IPAD,
  input LIOB33_X0Y53_IOB_X0Y54_IPAD,
  input LIOB33_X0Y55_IOB_X0Y55_IPAD,
  input LIOB33_X0Y55_IOB_X0Y56_IPAD,
  input LIOB33_X0Y57_IOB_X0Y57_IPAD,
  input LIOB33_X0Y57_IOB_X0Y58_IPAD,
  input LIOB33_X0Y59_IOB_X0Y59_IPAD,
  input LIOB33_X0Y59_IOB_X0Y60_IPAD,
  input LIOB33_X0Y61_IOB_X0Y61_IPAD,
  input LIOB33_X0Y61_IOB_X0Y62_IPAD,
  input LIOB33_X0Y63_IOB_X0Y63_IPAD,
  input LIOB33_X0Y63_IOB_X0Y64_IPAD,
  input LIOB33_X0Y65_IOB_X0Y65_IPAD,
  input LIOB33_X0Y65_IOB_X0Y66_IPAD,
  input LIOB33_X0Y67_IOB_X0Y67_IPAD,
  input LIOB33_X0Y67_IOB_X0Y68_IPAD,
  input LIOB33_X0Y69_IOB_X0Y69_IPAD,
  input LIOB33_X0Y69_IOB_X0Y70_IPAD,
  input LIOB33_X0Y71_IOB_X0Y71_IPAD,
  input LIOB33_X0Y71_IOB_X0Y72_IPAD,
  input LIOB33_X0Y73_IOB_X0Y73_IPAD,
  input LIOB33_X0Y73_IOB_X0Y74_IPAD,
  input LIOB33_X0Y75_IOB_X0Y75_IPAD,
  input LIOB33_X0Y75_IOB_X0Y76_IPAD,
  input LIOB33_X0Y77_IOB_X0Y77_IPAD,
  input LIOB33_X0Y77_IOB_X0Y78_IPAD,
  input LIOB33_X0Y79_IOB_X0Y79_IPAD,
  input LIOB33_X0Y79_IOB_X0Y80_IPAD,
  input LIOB33_X0Y81_IOB_X0Y81_IPAD,
  input LIOB33_X0Y81_IOB_X0Y82_IPAD,
  input LIOB33_X0Y83_IOB_X0Y83_IPAD,
  input LIOB33_X0Y83_IOB_X0Y84_IPAD,
  input LIOB33_X0Y85_IOB_X0Y85_IPAD,
  input LIOB33_X0Y85_IOB_X0Y86_IPAD,
  input LIOB33_X0Y87_IOB_X0Y87_IPAD,
  input LIOB33_X0Y87_IOB_X0Y88_IPAD,
  input LIOB33_X0Y89_IOB_X0Y89_IPAD,
  input LIOB33_X0Y89_IOB_X0Y90_IPAD,
  input LIOB33_X0Y91_IOB_X0Y91_IPAD,
  input LIOB33_X0Y91_IOB_X0Y92_IPAD,
  input LIOB33_X0Y93_IOB_X0Y93_IPAD,
  input LIOB33_X0Y93_IOB_X0Y94_IPAD,
  input LIOB33_X0Y95_IOB_X0Y95_IPAD,
  input LIOB33_X0Y95_IOB_X0Y96_IPAD,
  input LIOB33_X0Y97_IOB_X0Y97_IPAD,
  input LIOB33_X0Y97_IOB_X0Y98_IPAD,
  input RIOB33_SING_X105Y100_IOB_X1Y100_IPAD,
  input RIOB33_SING_X105Y150_IOB_X1Y150_IPAD,
  input RIOB33_X105Y101_IOB_X1Y101_IPAD,
  input RIOB33_X105Y101_IOB_X1Y102_IPAD,
  input RIOB33_X105Y103_IOB_X1Y103_IPAD,
  input RIOB33_X105Y103_IOB_X1Y104_IPAD,
  input RIOB33_X105Y105_IOB_X1Y105_IPAD,
  input RIOB33_X105Y105_IOB_X1Y106_IPAD,
  input RIOB33_X105Y107_IOB_X1Y107_IPAD,
  input RIOB33_X105Y107_IOB_X1Y108_IPAD,
  input RIOB33_X105Y109_IOB_X1Y109_IPAD,
  input RIOB33_X105Y109_IOB_X1Y110_IPAD,
  input RIOB33_X105Y111_IOB_X1Y111_IPAD,
  input RIOB33_X105Y111_IOB_X1Y112_IPAD,
  input RIOB33_X105Y113_IOB_X1Y113_IPAD,
  input RIOB33_X105Y113_IOB_X1Y114_IPAD,
  input RIOB33_X105Y115_IOB_X1Y115_IPAD,
  input RIOB33_X105Y115_IOB_X1Y116_IPAD,
  input RIOB33_X105Y117_IOB_X1Y117_IPAD,
  input RIOB33_X105Y117_IOB_X1Y118_IPAD,
  input RIOB33_X105Y119_IOB_X1Y119_IPAD,
  input RIOB33_X105Y119_IOB_X1Y120_IPAD,
  input RIOB33_X105Y121_IOB_X1Y121_IPAD,
  input RIOB33_X105Y121_IOB_X1Y122_IPAD,
  input RIOB33_X105Y123_IOB_X1Y123_IPAD,
  input RIOB33_X105Y123_IOB_X1Y124_IPAD,
  input RIOB33_X105Y125_IOB_X1Y125_IPAD,
  input RIOB33_X105Y125_IOB_X1Y126_IPAD,
  input RIOB33_X105Y151_IOB_X1Y151_IPAD,
  input RIOB33_X105Y151_IOB_X1Y152_IPAD,
  input RIOB33_X105Y153_IOB_X1Y153_IPAD,
  input RIOB33_X105Y153_IOB_X1Y154_IPAD,
  input RIOB33_X105Y155_IOB_X1Y155_IPAD,
  input RIOB33_X105Y155_IOB_X1Y156_IPAD,
  input RIOB33_X105Y157_IOB_X1Y157_IPAD,
  input RIOB33_X105Y157_IOB_X1Y158_IPAD,
  input RIOB33_X105Y159_IOB_X1Y159_IPAD,
  input RIOB33_X105Y159_IOB_X1Y160_IPAD,
  input RIOB33_X105Y161_IOB_X1Y161_IPAD,
  input RIOB33_X105Y161_IOB_X1Y162_IPAD,
  input RIOB33_X105Y163_IOB_X1Y163_IPAD,
  input RIOB33_X105Y163_IOB_X1Y164_IPAD,
  input RIOB33_X105Y165_IOB_X1Y165_IPAD,
  input RIOB33_X105Y165_IOB_X1Y166_IPAD,
  input RIOB33_X105Y167_IOB_X1Y167_IPAD,
  input RIOB33_X105Y167_IOB_X1Y168_IPAD,
  input RIOB33_X105Y169_IOB_X1Y169_IPAD,
  input RIOB33_X105Y169_IOB_X1Y170_IPAD,
  input RIOB33_X105Y171_IOB_X1Y171_IPAD,
  input RIOB33_X105Y171_IOB_X1Y172_IPAD,
  output LIOB33_SING_X0Y199_IOB_X0Y199_OPAD,
  output LIOB33_SING_X0Y200_IOB_X0Y200_OPAD,
  output LIOB33_X0Y177_IOB_X0Y178_OPAD,
  output LIOB33_X0Y179_IOB_X0Y179_OPAD,
  output LIOB33_X0Y179_IOB_X0Y180_OPAD,
  output LIOB33_X0Y181_IOB_X0Y181_OPAD,
  output LIOB33_X0Y181_IOB_X0Y182_OPAD,
  output LIOB33_X0Y183_IOB_X0Y183_OPAD,
  output LIOB33_X0Y183_IOB_X0Y184_OPAD,
  output LIOB33_X0Y185_IOB_X0Y185_OPAD,
  output LIOB33_X0Y185_IOB_X0Y186_OPAD,
  output LIOB33_X0Y187_IOB_X0Y187_OPAD,
  output LIOB33_X0Y187_IOB_X0Y188_OPAD,
  output LIOB33_X0Y189_IOB_X0Y189_OPAD,
  output LIOB33_X0Y189_IOB_X0Y190_OPAD,
  output LIOB33_X0Y191_IOB_X0Y191_OPAD,
  output LIOB33_X0Y191_IOB_X0Y192_OPAD,
  output LIOB33_X0Y193_IOB_X0Y193_OPAD,
  output LIOB33_X0Y193_IOB_X0Y194_OPAD,
  output LIOB33_X0Y195_IOB_X0Y195_OPAD,
  output LIOB33_X0Y195_IOB_X0Y196_OPAD,
  output LIOB33_X0Y197_IOB_X0Y197_OPAD,
  output LIOB33_X0Y197_IOB_X0Y198_OPAD,
  output RIOB33_SING_X105Y149_IOB_X1Y149_OPAD,
  output RIOB33_SING_X105Y199_IOB_X1Y199_OPAD,
  output RIOB33_SING_X105Y50_IOB_X1Y50_OPAD,
  output RIOB33_SING_X105Y99_IOB_X1Y99_OPAD,
  output RIOB33_X105Y127_IOB_X1Y127_OPAD,
  output RIOB33_X105Y127_IOB_X1Y128_OPAD,
  output RIOB33_X105Y129_IOB_X1Y129_OPAD,
  output RIOB33_X105Y129_IOB_X1Y130_OPAD,
  output RIOB33_X105Y131_IOB_X1Y131_OPAD,
  output RIOB33_X105Y131_IOB_X1Y132_OPAD,
  output RIOB33_X105Y133_IOB_X1Y133_OPAD,
  output RIOB33_X105Y133_IOB_X1Y134_OPAD,
  output RIOB33_X105Y135_IOB_X1Y135_OPAD,
  output RIOB33_X105Y135_IOB_X1Y136_OPAD,
  output RIOB33_X105Y137_IOB_X1Y137_OPAD,
  output RIOB33_X105Y137_IOB_X1Y138_OPAD,
  output RIOB33_X105Y139_IOB_X1Y139_OPAD,
  output RIOB33_X105Y139_IOB_X1Y140_OPAD,
  output RIOB33_X105Y141_IOB_X1Y141_OPAD,
  output RIOB33_X105Y141_IOB_X1Y142_OPAD,
  output RIOB33_X105Y143_IOB_X1Y143_OPAD,
  output RIOB33_X105Y143_IOB_X1Y144_OPAD,
  output RIOB33_X105Y145_IOB_X1Y145_OPAD,
  output RIOB33_X105Y145_IOB_X1Y146_OPAD,
  output RIOB33_X105Y147_IOB_X1Y147_OPAD,
  output RIOB33_X105Y147_IOB_X1Y148_OPAD,
  output RIOB33_X105Y173_IOB_X1Y173_OPAD,
  output RIOB33_X105Y173_IOB_X1Y174_OPAD,
  output RIOB33_X105Y175_IOB_X1Y175_OPAD,
  output RIOB33_X105Y175_IOB_X1Y176_OPAD,
  output RIOB33_X105Y177_IOB_X1Y177_OPAD,
  output RIOB33_X105Y177_IOB_X1Y178_OPAD,
  output RIOB33_X105Y179_IOB_X1Y179_OPAD,
  output RIOB33_X105Y179_IOB_X1Y180_OPAD,
  output RIOB33_X105Y181_IOB_X1Y181_OPAD,
  output RIOB33_X105Y181_IOB_X1Y182_OPAD,
  output RIOB33_X105Y183_IOB_X1Y183_OPAD,
  output RIOB33_X105Y183_IOB_X1Y184_OPAD,
  output RIOB33_X105Y185_IOB_X1Y185_OPAD,
  output RIOB33_X105Y185_IOB_X1Y186_OPAD,
  output RIOB33_X105Y187_IOB_X1Y187_OPAD,
  output RIOB33_X105Y187_IOB_X1Y188_OPAD,
  output RIOB33_X105Y189_IOB_X1Y189_OPAD,
  output RIOB33_X105Y189_IOB_X1Y190_OPAD,
  output RIOB33_X105Y191_IOB_X1Y191_OPAD,
  output RIOB33_X105Y191_IOB_X1Y192_OPAD,
  output RIOB33_X105Y193_IOB_X1Y193_OPAD,
  output RIOB33_X105Y193_IOB_X1Y194_OPAD,
  output RIOB33_X105Y195_IOB_X1Y195_OPAD,
  output RIOB33_X105Y195_IOB_X1Y196_OPAD,
  output RIOB33_X105Y197_IOB_X1Y197_OPAD,
  output RIOB33_X105Y197_IOB_X1Y198_OPAD,
  output RIOB33_X105Y51_IOB_X1Y51_OPAD,
  output RIOB33_X105Y51_IOB_X1Y52_OPAD,
  output RIOB33_X105Y53_IOB_X1Y53_OPAD,
  output RIOB33_X105Y53_IOB_X1Y54_OPAD,
  output RIOB33_X105Y55_IOB_X1Y55_OPAD,
  output RIOB33_X105Y55_IOB_X1Y56_OPAD,
  output RIOB33_X105Y57_IOB_X1Y57_OPAD,
  output RIOB33_X105Y57_IOB_X1Y58_OPAD,
  output RIOB33_X105Y59_IOB_X1Y59_OPAD,
  output RIOB33_X105Y59_IOB_X1Y60_OPAD,
  output RIOB33_X105Y61_IOB_X1Y61_OPAD,
  output RIOB33_X105Y61_IOB_X1Y62_OPAD,
  output RIOB33_X105Y63_IOB_X1Y63_OPAD,
  output RIOB33_X105Y63_IOB_X1Y64_OPAD,
  output RIOB33_X105Y65_IOB_X1Y65_OPAD,
  output RIOB33_X105Y65_IOB_X1Y66_OPAD,
  output RIOB33_X105Y67_IOB_X1Y67_OPAD,
  output RIOB33_X105Y67_IOB_X1Y68_OPAD,
  output RIOB33_X105Y69_IOB_X1Y69_OPAD,
  output RIOB33_X105Y69_IOB_X1Y70_OPAD,
  output RIOB33_X105Y71_IOB_X1Y71_OPAD,
  output RIOB33_X105Y71_IOB_X1Y72_OPAD,
  output RIOB33_X105Y73_IOB_X1Y73_OPAD,
  output RIOB33_X105Y73_IOB_X1Y74_OPAD,
  output RIOB33_X105Y75_IOB_X1Y75_OPAD,
  output RIOB33_X105Y75_IOB_X1Y76_OPAD,
  output RIOB33_X105Y77_IOB_X1Y77_OPAD,
  output RIOB33_X105Y77_IOB_X1Y78_OPAD,
  output RIOB33_X105Y79_IOB_X1Y79_OPAD,
  output RIOB33_X105Y79_IOB_X1Y80_OPAD,
  output RIOB33_X105Y81_IOB_X1Y81_OPAD,
  output RIOB33_X105Y81_IOB_X1Y82_OPAD,
  output RIOB33_X105Y83_IOB_X1Y83_OPAD,
  output RIOB33_X105Y83_IOB_X1Y84_OPAD,
  output RIOB33_X105Y85_IOB_X1Y85_OPAD,
  output RIOB33_X105Y85_IOB_X1Y86_OPAD,
  output RIOB33_X105Y87_IOB_X1Y87_OPAD,
  output RIOB33_X105Y87_IOB_X1Y88_OPAD,
  output RIOB33_X105Y89_IOB_X1Y89_OPAD,
  output RIOB33_X105Y89_IOB_X1Y90_OPAD,
  output RIOB33_X105Y91_IOB_X1Y91_OPAD,
  output RIOB33_X105Y91_IOB_X1Y92_OPAD,
  output RIOB33_X105Y93_IOB_X1Y93_OPAD,
  output RIOB33_X105Y93_IOB_X1Y94_OPAD,
  output RIOB33_X105Y95_IOB_X1Y95_OPAD,
  output RIOB33_X105Y95_IOB_X1Y96_OPAD,
  output RIOB33_X105Y97_IOB_X1Y97_OPAD,
  output RIOB33_X105Y97_IOB_X1Y98_OPAD
  );
  wire [0:0] CLBLL_L_X100Y113_SLICE_X156Y113_A;
  wire [0:0] CLBLL_L_X100Y113_SLICE_X156Y113_A1;
  wire [0:0] CLBLL_L_X100Y113_SLICE_X156Y113_A2;
  wire [0:0] CLBLL_L_X100Y113_SLICE_X156Y113_A3;
  wire [0:0] CLBLL_L_X100Y113_SLICE_X156Y113_A4;
  wire [0:0] CLBLL_L_X100Y113_SLICE_X156Y113_A5;
  wire [0:0] CLBLL_L_X100Y113_SLICE_X156Y113_A6;
  wire [0:0] CLBLL_L_X100Y113_SLICE_X156Y113_AO5;
  wire [0:0] CLBLL_L_X100Y113_SLICE_X156Y113_AO6;
  wire [0:0] CLBLL_L_X100Y113_SLICE_X156Y113_A_CY;
  wire [0:0] CLBLL_L_X100Y113_SLICE_X156Y113_A_XOR;
  wire [0:0] CLBLL_L_X100Y113_SLICE_X156Y113_B;
  wire [0:0] CLBLL_L_X100Y113_SLICE_X156Y113_B1;
  wire [0:0] CLBLL_L_X100Y113_SLICE_X156Y113_B2;
  wire [0:0] CLBLL_L_X100Y113_SLICE_X156Y113_B3;
  wire [0:0] CLBLL_L_X100Y113_SLICE_X156Y113_B4;
  wire [0:0] CLBLL_L_X100Y113_SLICE_X156Y113_B5;
  wire [0:0] CLBLL_L_X100Y113_SLICE_X156Y113_B6;
  wire [0:0] CLBLL_L_X100Y113_SLICE_X156Y113_BO5;
  wire [0:0] CLBLL_L_X100Y113_SLICE_X156Y113_BO6;
  wire [0:0] CLBLL_L_X100Y113_SLICE_X156Y113_B_CY;
  wire [0:0] CLBLL_L_X100Y113_SLICE_X156Y113_B_XOR;
  wire [0:0] CLBLL_L_X100Y113_SLICE_X156Y113_C;
  wire [0:0] CLBLL_L_X100Y113_SLICE_X156Y113_C1;
  wire [0:0] CLBLL_L_X100Y113_SLICE_X156Y113_C2;
  wire [0:0] CLBLL_L_X100Y113_SLICE_X156Y113_C3;
  wire [0:0] CLBLL_L_X100Y113_SLICE_X156Y113_C4;
  wire [0:0] CLBLL_L_X100Y113_SLICE_X156Y113_C5;
  wire [0:0] CLBLL_L_X100Y113_SLICE_X156Y113_C6;
  wire [0:0] CLBLL_L_X100Y113_SLICE_X156Y113_CO5;
  wire [0:0] CLBLL_L_X100Y113_SLICE_X156Y113_CO6;
  wire [0:0] CLBLL_L_X100Y113_SLICE_X156Y113_C_CY;
  wire [0:0] CLBLL_L_X100Y113_SLICE_X156Y113_C_XOR;
  wire [0:0] CLBLL_L_X100Y113_SLICE_X156Y113_D;
  wire [0:0] CLBLL_L_X100Y113_SLICE_X156Y113_D1;
  wire [0:0] CLBLL_L_X100Y113_SLICE_X156Y113_D2;
  wire [0:0] CLBLL_L_X100Y113_SLICE_X156Y113_D3;
  wire [0:0] CLBLL_L_X100Y113_SLICE_X156Y113_D4;
  wire [0:0] CLBLL_L_X100Y113_SLICE_X156Y113_D5;
  wire [0:0] CLBLL_L_X100Y113_SLICE_X156Y113_D6;
  wire [0:0] CLBLL_L_X100Y113_SLICE_X156Y113_DO5;
  wire [0:0] CLBLL_L_X100Y113_SLICE_X156Y113_DO6;
  wire [0:0] CLBLL_L_X100Y113_SLICE_X156Y113_D_CY;
  wire [0:0] CLBLL_L_X100Y113_SLICE_X156Y113_D_XOR;
  wire [0:0] CLBLL_L_X100Y113_SLICE_X157Y113_A;
  wire [0:0] CLBLL_L_X100Y113_SLICE_X157Y113_A1;
  wire [0:0] CLBLL_L_X100Y113_SLICE_X157Y113_A2;
  wire [0:0] CLBLL_L_X100Y113_SLICE_X157Y113_A3;
  wire [0:0] CLBLL_L_X100Y113_SLICE_X157Y113_A4;
  wire [0:0] CLBLL_L_X100Y113_SLICE_X157Y113_A5;
  wire [0:0] CLBLL_L_X100Y113_SLICE_X157Y113_A6;
  wire [0:0] CLBLL_L_X100Y113_SLICE_X157Y113_AO5;
  wire [0:0] CLBLL_L_X100Y113_SLICE_X157Y113_AO6;
  wire [0:0] CLBLL_L_X100Y113_SLICE_X157Y113_A_CY;
  wire [0:0] CLBLL_L_X100Y113_SLICE_X157Y113_A_XOR;
  wire [0:0] CLBLL_L_X100Y113_SLICE_X157Y113_B;
  wire [0:0] CLBLL_L_X100Y113_SLICE_X157Y113_B1;
  wire [0:0] CLBLL_L_X100Y113_SLICE_X157Y113_B2;
  wire [0:0] CLBLL_L_X100Y113_SLICE_X157Y113_B3;
  wire [0:0] CLBLL_L_X100Y113_SLICE_X157Y113_B4;
  wire [0:0] CLBLL_L_X100Y113_SLICE_X157Y113_B5;
  wire [0:0] CLBLL_L_X100Y113_SLICE_X157Y113_B6;
  wire [0:0] CLBLL_L_X100Y113_SLICE_X157Y113_BO5;
  wire [0:0] CLBLL_L_X100Y113_SLICE_X157Y113_BO6;
  wire [0:0] CLBLL_L_X100Y113_SLICE_X157Y113_B_CY;
  wire [0:0] CLBLL_L_X100Y113_SLICE_X157Y113_B_XOR;
  wire [0:0] CLBLL_L_X100Y113_SLICE_X157Y113_C;
  wire [0:0] CLBLL_L_X100Y113_SLICE_X157Y113_C1;
  wire [0:0] CLBLL_L_X100Y113_SLICE_X157Y113_C2;
  wire [0:0] CLBLL_L_X100Y113_SLICE_X157Y113_C3;
  wire [0:0] CLBLL_L_X100Y113_SLICE_X157Y113_C4;
  wire [0:0] CLBLL_L_X100Y113_SLICE_X157Y113_C5;
  wire [0:0] CLBLL_L_X100Y113_SLICE_X157Y113_C6;
  wire [0:0] CLBLL_L_X100Y113_SLICE_X157Y113_CO5;
  wire [0:0] CLBLL_L_X100Y113_SLICE_X157Y113_CO6;
  wire [0:0] CLBLL_L_X100Y113_SLICE_X157Y113_C_CY;
  wire [0:0] CLBLL_L_X100Y113_SLICE_X157Y113_C_XOR;
  wire [0:0] CLBLL_L_X100Y113_SLICE_X157Y113_D;
  wire [0:0] CLBLL_L_X100Y113_SLICE_X157Y113_D1;
  wire [0:0] CLBLL_L_X100Y113_SLICE_X157Y113_D2;
  wire [0:0] CLBLL_L_X100Y113_SLICE_X157Y113_D3;
  wire [0:0] CLBLL_L_X100Y113_SLICE_X157Y113_D4;
  wire [0:0] CLBLL_L_X100Y113_SLICE_X157Y113_D5;
  wire [0:0] CLBLL_L_X100Y113_SLICE_X157Y113_D6;
  wire [0:0] CLBLL_L_X100Y113_SLICE_X157Y113_DO5;
  wire [0:0] CLBLL_L_X100Y113_SLICE_X157Y113_DO6;
  wire [0:0] CLBLL_L_X100Y113_SLICE_X157Y113_D_CY;
  wire [0:0] CLBLL_L_X100Y113_SLICE_X157Y113_D_XOR;
  wire [0:0] CLBLL_L_X100Y121_SLICE_X156Y121_A;
  wire [0:0] CLBLL_L_X100Y121_SLICE_X156Y121_A1;
  wire [0:0] CLBLL_L_X100Y121_SLICE_X156Y121_A2;
  wire [0:0] CLBLL_L_X100Y121_SLICE_X156Y121_A3;
  wire [0:0] CLBLL_L_X100Y121_SLICE_X156Y121_A4;
  wire [0:0] CLBLL_L_X100Y121_SLICE_X156Y121_A5;
  wire [0:0] CLBLL_L_X100Y121_SLICE_X156Y121_A6;
  wire [0:0] CLBLL_L_X100Y121_SLICE_X156Y121_AO5;
  wire [0:0] CLBLL_L_X100Y121_SLICE_X156Y121_AO6;
  wire [0:0] CLBLL_L_X100Y121_SLICE_X156Y121_A_CY;
  wire [0:0] CLBLL_L_X100Y121_SLICE_X156Y121_A_XOR;
  wire [0:0] CLBLL_L_X100Y121_SLICE_X156Y121_B;
  wire [0:0] CLBLL_L_X100Y121_SLICE_X156Y121_B1;
  wire [0:0] CLBLL_L_X100Y121_SLICE_X156Y121_B2;
  wire [0:0] CLBLL_L_X100Y121_SLICE_X156Y121_B3;
  wire [0:0] CLBLL_L_X100Y121_SLICE_X156Y121_B4;
  wire [0:0] CLBLL_L_X100Y121_SLICE_X156Y121_B5;
  wire [0:0] CLBLL_L_X100Y121_SLICE_X156Y121_B6;
  wire [0:0] CLBLL_L_X100Y121_SLICE_X156Y121_BO5;
  wire [0:0] CLBLL_L_X100Y121_SLICE_X156Y121_BO6;
  wire [0:0] CLBLL_L_X100Y121_SLICE_X156Y121_B_CY;
  wire [0:0] CLBLL_L_X100Y121_SLICE_X156Y121_B_XOR;
  wire [0:0] CLBLL_L_X100Y121_SLICE_X156Y121_C;
  wire [0:0] CLBLL_L_X100Y121_SLICE_X156Y121_C1;
  wire [0:0] CLBLL_L_X100Y121_SLICE_X156Y121_C2;
  wire [0:0] CLBLL_L_X100Y121_SLICE_X156Y121_C3;
  wire [0:0] CLBLL_L_X100Y121_SLICE_X156Y121_C4;
  wire [0:0] CLBLL_L_X100Y121_SLICE_X156Y121_C5;
  wire [0:0] CLBLL_L_X100Y121_SLICE_X156Y121_C6;
  wire [0:0] CLBLL_L_X100Y121_SLICE_X156Y121_CO5;
  wire [0:0] CLBLL_L_X100Y121_SLICE_X156Y121_CO6;
  wire [0:0] CLBLL_L_X100Y121_SLICE_X156Y121_C_CY;
  wire [0:0] CLBLL_L_X100Y121_SLICE_X156Y121_C_XOR;
  wire [0:0] CLBLL_L_X100Y121_SLICE_X156Y121_D;
  wire [0:0] CLBLL_L_X100Y121_SLICE_X156Y121_D1;
  wire [0:0] CLBLL_L_X100Y121_SLICE_X156Y121_D2;
  wire [0:0] CLBLL_L_X100Y121_SLICE_X156Y121_D3;
  wire [0:0] CLBLL_L_X100Y121_SLICE_X156Y121_D4;
  wire [0:0] CLBLL_L_X100Y121_SLICE_X156Y121_D5;
  wire [0:0] CLBLL_L_X100Y121_SLICE_X156Y121_D6;
  wire [0:0] CLBLL_L_X100Y121_SLICE_X156Y121_DO5;
  wire [0:0] CLBLL_L_X100Y121_SLICE_X156Y121_DO6;
  wire [0:0] CLBLL_L_X100Y121_SLICE_X156Y121_D_CY;
  wire [0:0] CLBLL_L_X100Y121_SLICE_X156Y121_D_XOR;
  wire [0:0] CLBLL_L_X100Y121_SLICE_X157Y121_A;
  wire [0:0] CLBLL_L_X100Y121_SLICE_X157Y121_A1;
  wire [0:0] CLBLL_L_X100Y121_SLICE_X157Y121_A2;
  wire [0:0] CLBLL_L_X100Y121_SLICE_X157Y121_A3;
  wire [0:0] CLBLL_L_X100Y121_SLICE_X157Y121_A4;
  wire [0:0] CLBLL_L_X100Y121_SLICE_X157Y121_A5;
  wire [0:0] CLBLL_L_X100Y121_SLICE_X157Y121_A6;
  wire [0:0] CLBLL_L_X100Y121_SLICE_X157Y121_AO5;
  wire [0:0] CLBLL_L_X100Y121_SLICE_X157Y121_AO6;
  wire [0:0] CLBLL_L_X100Y121_SLICE_X157Y121_A_CY;
  wire [0:0] CLBLL_L_X100Y121_SLICE_X157Y121_A_XOR;
  wire [0:0] CLBLL_L_X100Y121_SLICE_X157Y121_B;
  wire [0:0] CLBLL_L_X100Y121_SLICE_X157Y121_B1;
  wire [0:0] CLBLL_L_X100Y121_SLICE_X157Y121_B2;
  wire [0:0] CLBLL_L_X100Y121_SLICE_X157Y121_B3;
  wire [0:0] CLBLL_L_X100Y121_SLICE_X157Y121_B4;
  wire [0:0] CLBLL_L_X100Y121_SLICE_X157Y121_B5;
  wire [0:0] CLBLL_L_X100Y121_SLICE_X157Y121_B6;
  wire [0:0] CLBLL_L_X100Y121_SLICE_X157Y121_BO5;
  wire [0:0] CLBLL_L_X100Y121_SLICE_X157Y121_BO6;
  wire [0:0] CLBLL_L_X100Y121_SLICE_X157Y121_B_CY;
  wire [0:0] CLBLL_L_X100Y121_SLICE_X157Y121_B_XOR;
  wire [0:0] CLBLL_L_X100Y121_SLICE_X157Y121_C;
  wire [0:0] CLBLL_L_X100Y121_SLICE_X157Y121_C1;
  wire [0:0] CLBLL_L_X100Y121_SLICE_X157Y121_C2;
  wire [0:0] CLBLL_L_X100Y121_SLICE_X157Y121_C3;
  wire [0:0] CLBLL_L_X100Y121_SLICE_X157Y121_C4;
  wire [0:0] CLBLL_L_X100Y121_SLICE_X157Y121_C5;
  wire [0:0] CLBLL_L_X100Y121_SLICE_X157Y121_C6;
  wire [0:0] CLBLL_L_X100Y121_SLICE_X157Y121_CO5;
  wire [0:0] CLBLL_L_X100Y121_SLICE_X157Y121_CO6;
  wire [0:0] CLBLL_L_X100Y121_SLICE_X157Y121_C_CY;
  wire [0:0] CLBLL_L_X100Y121_SLICE_X157Y121_C_XOR;
  wire [0:0] CLBLL_L_X100Y121_SLICE_X157Y121_D;
  wire [0:0] CLBLL_L_X100Y121_SLICE_X157Y121_D1;
  wire [0:0] CLBLL_L_X100Y121_SLICE_X157Y121_D2;
  wire [0:0] CLBLL_L_X100Y121_SLICE_X157Y121_D3;
  wire [0:0] CLBLL_L_X100Y121_SLICE_X157Y121_D4;
  wire [0:0] CLBLL_L_X100Y121_SLICE_X157Y121_D5;
  wire [0:0] CLBLL_L_X100Y121_SLICE_X157Y121_D6;
  wire [0:0] CLBLL_L_X100Y121_SLICE_X157Y121_DO5;
  wire [0:0] CLBLL_L_X100Y121_SLICE_X157Y121_DO6;
  wire [0:0] CLBLL_L_X100Y121_SLICE_X157Y121_D_CY;
  wire [0:0] CLBLL_L_X100Y121_SLICE_X157Y121_D_XOR;
  wire [0:0] CLBLL_L_X100Y123_SLICE_X156Y123_A;
  wire [0:0] CLBLL_L_X100Y123_SLICE_X156Y123_A1;
  wire [0:0] CLBLL_L_X100Y123_SLICE_X156Y123_A2;
  wire [0:0] CLBLL_L_X100Y123_SLICE_X156Y123_A3;
  wire [0:0] CLBLL_L_X100Y123_SLICE_X156Y123_A4;
  wire [0:0] CLBLL_L_X100Y123_SLICE_X156Y123_A5;
  wire [0:0] CLBLL_L_X100Y123_SLICE_X156Y123_A6;
  wire [0:0] CLBLL_L_X100Y123_SLICE_X156Y123_AMUX;
  wire [0:0] CLBLL_L_X100Y123_SLICE_X156Y123_AO5;
  wire [0:0] CLBLL_L_X100Y123_SLICE_X156Y123_AO6;
  wire [0:0] CLBLL_L_X100Y123_SLICE_X156Y123_A_CY;
  wire [0:0] CLBLL_L_X100Y123_SLICE_X156Y123_A_XOR;
  wire [0:0] CLBLL_L_X100Y123_SLICE_X156Y123_B;
  wire [0:0] CLBLL_L_X100Y123_SLICE_X156Y123_B1;
  wire [0:0] CLBLL_L_X100Y123_SLICE_X156Y123_B2;
  wire [0:0] CLBLL_L_X100Y123_SLICE_X156Y123_B3;
  wire [0:0] CLBLL_L_X100Y123_SLICE_X156Y123_B4;
  wire [0:0] CLBLL_L_X100Y123_SLICE_X156Y123_B5;
  wire [0:0] CLBLL_L_X100Y123_SLICE_X156Y123_B6;
  wire [0:0] CLBLL_L_X100Y123_SLICE_X156Y123_BMUX;
  wire [0:0] CLBLL_L_X100Y123_SLICE_X156Y123_BO5;
  wire [0:0] CLBLL_L_X100Y123_SLICE_X156Y123_BO6;
  wire [0:0] CLBLL_L_X100Y123_SLICE_X156Y123_B_CY;
  wire [0:0] CLBLL_L_X100Y123_SLICE_X156Y123_B_XOR;
  wire [0:0] CLBLL_L_X100Y123_SLICE_X156Y123_C;
  wire [0:0] CLBLL_L_X100Y123_SLICE_X156Y123_C1;
  wire [0:0] CLBLL_L_X100Y123_SLICE_X156Y123_C2;
  wire [0:0] CLBLL_L_X100Y123_SLICE_X156Y123_C3;
  wire [0:0] CLBLL_L_X100Y123_SLICE_X156Y123_C4;
  wire [0:0] CLBLL_L_X100Y123_SLICE_X156Y123_C5;
  wire [0:0] CLBLL_L_X100Y123_SLICE_X156Y123_C6;
  wire [0:0] CLBLL_L_X100Y123_SLICE_X156Y123_CO5;
  wire [0:0] CLBLL_L_X100Y123_SLICE_X156Y123_CO6;
  wire [0:0] CLBLL_L_X100Y123_SLICE_X156Y123_C_CY;
  wire [0:0] CLBLL_L_X100Y123_SLICE_X156Y123_C_XOR;
  wire [0:0] CLBLL_L_X100Y123_SLICE_X156Y123_D;
  wire [0:0] CLBLL_L_X100Y123_SLICE_X156Y123_D1;
  wire [0:0] CLBLL_L_X100Y123_SLICE_X156Y123_D2;
  wire [0:0] CLBLL_L_X100Y123_SLICE_X156Y123_D3;
  wire [0:0] CLBLL_L_X100Y123_SLICE_X156Y123_D4;
  wire [0:0] CLBLL_L_X100Y123_SLICE_X156Y123_D5;
  wire [0:0] CLBLL_L_X100Y123_SLICE_X156Y123_D6;
  wire [0:0] CLBLL_L_X100Y123_SLICE_X156Y123_DO5;
  wire [0:0] CLBLL_L_X100Y123_SLICE_X156Y123_DO6;
  wire [0:0] CLBLL_L_X100Y123_SLICE_X156Y123_D_CY;
  wire [0:0] CLBLL_L_X100Y123_SLICE_X156Y123_D_XOR;
  wire [0:0] CLBLL_L_X100Y123_SLICE_X157Y123_A;
  wire [0:0] CLBLL_L_X100Y123_SLICE_X157Y123_A1;
  wire [0:0] CLBLL_L_X100Y123_SLICE_X157Y123_A2;
  wire [0:0] CLBLL_L_X100Y123_SLICE_X157Y123_A3;
  wire [0:0] CLBLL_L_X100Y123_SLICE_X157Y123_A4;
  wire [0:0] CLBLL_L_X100Y123_SLICE_X157Y123_A5;
  wire [0:0] CLBLL_L_X100Y123_SLICE_X157Y123_A6;
  wire [0:0] CLBLL_L_X100Y123_SLICE_X157Y123_AO5;
  wire [0:0] CLBLL_L_X100Y123_SLICE_X157Y123_AO6;
  wire [0:0] CLBLL_L_X100Y123_SLICE_X157Y123_A_CY;
  wire [0:0] CLBLL_L_X100Y123_SLICE_X157Y123_A_XOR;
  wire [0:0] CLBLL_L_X100Y123_SLICE_X157Y123_B;
  wire [0:0] CLBLL_L_X100Y123_SLICE_X157Y123_B1;
  wire [0:0] CLBLL_L_X100Y123_SLICE_X157Y123_B2;
  wire [0:0] CLBLL_L_X100Y123_SLICE_X157Y123_B3;
  wire [0:0] CLBLL_L_X100Y123_SLICE_X157Y123_B4;
  wire [0:0] CLBLL_L_X100Y123_SLICE_X157Y123_B5;
  wire [0:0] CLBLL_L_X100Y123_SLICE_X157Y123_B6;
  wire [0:0] CLBLL_L_X100Y123_SLICE_X157Y123_BO5;
  wire [0:0] CLBLL_L_X100Y123_SLICE_X157Y123_BO6;
  wire [0:0] CLBLL_L_X100Y123_SLICE_X157Y123_B_CY;
  wire [0:0] CLBLL_L_X100Y123_SLICE_X157Y123_B_XOR;
  wire [0:0] CLBLL_L_X100Y123_SLICE_X157Y123_C;
  wire [0:0] CLBLL_L_X100Y123_SLICE_X157Y123_C1;
  wire [0:0] CLBLL_L_X100Y123_SLICE_X157Y123_C2;
  wire [0:0] CLBLL_L_X100Y123_SLICE_X157Y123_C3;
  wire [0:0] CLBLL_L_X100Y123_SLICE_X157Y123_C4;
  wire [0:0] CLBLL_L_X100Y123_SLICE_X157Y123_C5;
  wire [0:0] CLBLL_L_X100Y123_SLICE_X157Y123_C6;
  wire [0:0] CLBLL_L_X100Y123_SLICE_X157Y123_CO5;
  wire [0:0] CLBLL_L_X100Y123_SLICE_X157Y123_CO6;
  wire [0:0] CLBLL_L_X100Y123_SLICE_X157Y123_C_CY;
  wire [0:0] CLBLL_L_X100Y123_SLICE_X157Y123_C_XOR;
  wire [0:0] CLBLL_L_X100Y123_SLICE_X157Y123_D;
  wire [0:0] CLBLL_L_X100Y123_SLICE_X157Y123_D1;
  wire [0:0] CLBLL_L_X100Y123_SLICE_X157Y123_D2;
  wire [0:0] CLBLL_L_X100Y123_SLICE_X157Y123_D3;
  wire [0:0] CLBLL_L_X100Y123_SLICE_X157Y123_D4;
  wire [0:0] CLBLL_L_X100Y123_SLICE_X157Y123_D5;
  wire [0:0] CLBLL_L_X100Y123_SLICE_X157Y123_D6;
  wire [0:0] CLBLL_L_X100Y123_SLICE_X157Y123_DO5;
  wire [0:0] CLBLL_L_X100Y123_SLICE_X157Y123_DO6;
  wire [0:0] CLBLL_L_X100Y123_SLICE_X157Y123_D_CY;
  wire [0:0] CLBLL_L_X100Y123_SLICE_X157Y123_D_XOR;
  wire [0:0] CLBLL_L_X2Y102_SLICE_X0Y102_A;
  wire [0:0] CLBLL_L_X2Y102_SLICE_X0Y102_A1;
  wire [0:0] CLBLL_L_X2Y102_SLICE_X0Y102_A2;
  wire [0:0] CLBLL_L_X2Y102_SLICE_X0Y102_A3;
  wire [0:0] CLBLL_L_X2Y102_SLICE_X0Y102_A4;
  wire [0:0] CLBLL_L_X2Y102_SLICE_X0Y102_A5;
  wire [0:0] CLBLL_L_X2Y102_SLICE_X0Y102_A6;
  wire [0:0] CLBLL_L_X2Y102_SLICE_X0Y102_AO5;
  wire [0:0] CLBLL_L_X2Y102_SLICE_X0Y102_AO6;
  wire [0:0] CLBLL_L_X2Y102_SLICE_X0Y102_A_CY;
  wire [0:0] CLBLL_L_X2Y102_SLICE_X0Y102_A_XOR;
  wire [0:0] CLBLL_L_X2Y102_SLICE_X0Y102_B;
  wire [0:0] CLBLL_L_X2Y102_SLICE_X0Y102_B1;
  wire [0:0] CLBLL_L_X2Y102_SLICE_X0Y102_B2;
  wire [0:0] CLBLL_L_X2Y102_SLICE_X0Y102_B3;
  wire [0:0] CLBLL_L_X2Y102_SLICE_X0Y102_B4;
  wire [0:0] CLBLL_L_X2Y102_SLICE_X0Y102_B5;
  wire [0:0] CLBLL_L_X2Y102_SLICE_X0Y102_B6;
  wire [0:0] CLBLL_L_X2Y102_SLICE_X0Y102_BO5;
  wire [0:0] CLBLL_L_X2Y102_SLICE_X0Y102_BO6;
  wire [0:0] CLBLL_L_X2Y102_SLICE_X0Y102_B_CY;
  wire [0:0] CLBLL_L_X2Y102_SLICE_X0Y102_B_XOR;
  wire [0:0] CLBLL_L_X2Y102_SLICE_X0Y102_C;
  wire [0:0] CLBLL_L_X2Y102_SLICE_X0Y102_C1;
  wire [0:0] CLBLL_L_X2Y102_SLICE_X0Y102_C2;
  wire [0:0] CLBLL_L_X2Y102_SLICE_X0Y102_C3;
  wire [0:0] CLBLL_L_X2Y102_SLICE_X0Y102_C4;
  wire [0:0] CLBLL_L_X2Y102_SLICE_X0Y102_C5;
  wire [0:0] CLBLL_L_X2Y102_SLICE_X0Y102_C6;
  wire [0:0] CLBLL_L_X2Y102_SLICE_X0Y102_CO5;
  wire [0:0] CLBLL_L_X2Y102_SLICE_X0Y102_CO6;
  wire [0:0] CLBLL_L_X2Y102_SLICE_X0Y102_C_CY;
  wire [0:0] CLBLL_L_X2Y102_SLICE_X0Y102_C_XOR;
  wire [0:0] CLBLL_L_X2Y102_SLICE_X0Y102_D;
  wire [0:0] CLBLL_L_X2Y102_SLICE_X0Y102_D1;
  wire [0:0] CLBLL_L_X2Y102_SLICE_X0Y102_D2;
  wire [0:0] CLBLL_L_X2Y102_SLICE_X0Y102_D3;
  wire [0:0] CLBLL_L_X2Y102_SLICE_X0Y102_D4;
  wire [0:0] CLBLL_L_X2Y102_SLICE_X0Y102_D5;
  wire [0:0] CLBLL_L_X2Y102_SLICE_X0Y102_D6;
  wire [0:0] CLBLL_L_X2Y102_SLICE_X0Y102_DO5;
  wire [0:0] CLBLL_L_X2Y102_SLICE_X0Y102_DO6;
  wire [0:0] CLBLL_L_X2Y102_SLICE_X0Y102_D_CY;
  wire [0:0] CLBLL_L_X2Y102_SLICE_X0Y102_D_XOR;
  wire [0:0] CLBLL_L_X2Y102_SLICE_X1Y102_A;
  wire [0:0] CLBLL_L_X2Y102_SLICE_X1Y102_A1;
  wire [0:0] CLBLL_L_X2Y102_SLICE_X1Y102_A2;
  wire [0:0] CLBLL_L_X2Y102_SLICE_X1Y102_A3;
  wire [0:0] CLBLL_L_X2Y102_SLICE_X1Y102_A4;
  wire [0:0] CLBLL_L_X2Y102_SLICE_X1Y102_A5;
  wire [0:0] CLBLL_L_X2Y102_SLICE_X1Y102_A6;
  wire [0:0] CLBLL_L_X2Y102_SLICE_X1Y102_AO5;
  wire [0:0] CLBLL_L_X2Y102_SLICE_X1Y102_AO6;
  wire [0:0] CLBLL_L_X2Y102_SLICE_X1Y102_A_CY;
  wire [0:0] CLBLL_L_X2Y102_SLICE_X1Y102_A_XOR;
  wire [0:0] CLBLL_L_X2Y102_SLICE_X1Y102_B;
  wire [0:0] CLBLL_L_X2Y102_SLICE_X1Y102_B1;
  wire [0:0] CLBLL_L_X2Y102_SLICE_X1Y102_B2;
  wire [0:0] CLBLL_L_X2Y102_SLICE_X1Y102_B3;
  wire [0:0] CLBLL_L_X2Y102_SLICE_X1Y102_B4;
  wire [0:0] CLBLL_L_X2Y102_SLICE_X1Y102_B5;
  wire [0:0] CLBLL_L_X2Y102_SLICE_X1Y102_B6;
  wire [0:0] CLBLL_L_X2Y102_SLICE_X1Y102_BO5;
  wire [0:0] CLBLL_L_X2Y102_SLICE_X1Y102_BO6;
  wire [0:0] CLBLL_L_X2Y102_SLICE_X1Y102_B_CY;
  wire [0:0] CLBLL_L_X2Y102_SLICE_X1Y102_B_XOR;
  wire [0:0] CLBLL_L_X2Y102_SLICE_X1Y102_C;
  wire [0:0] CLBLL_L_X2Y102_SLICE_X1Y102_C1;
  wire [0:0] CLBLL_L_X2Y102_SLICE_X1Y102_C2;
  wire [0:0] CLBLL_L_X2Y102_SLICE_X1Y102_C3;
  wire [0:0] CLBLL_L_X2Y102_SLICE_X1Y102_C4;
  wire [0:0] CLBLL_L_X2Y102_SLICE_X1Y102_C5;
  wire [0:0] CLBLL_L_X2Y102_SLICE_X1Y102_C6;
  wire [0:0] CLBLL_L_X2Y102_SLICE_X1Y102_CO5;
  wire [0:0] CLBLL_L_X2Y102_SLICE_X1Y102_CO6;
  wire [0:0] CLBLL_L_X2Y102_SLICE_X1Y102_C_CY;
  wire [0:0] CLBLL_L_X2Y102_SLICE_X1Y102_C_XOR;
  wire [0:0] CLBLL_L_X2Y102_SLICE_X1Y102_D;
  wire [0:0] CLBLL_L_X2Y102_SLICE_X1Y102_D1;
  wire [0:0] CLBLL_L_X2Y102_SLICE_X1Y102_D2;
  wire [0:0] CLBLL_L_X2Y102_SLICE_X1Y102_D3;
  wire [0:0] CLBLL_L_X2Y102_SLICE_X1Y102_D4;
  wire [0:0] CLBLL_L_X2Y102_SLICE_X1Y102_D5;
  wire [0:0] CLBLL_L_X2Y102_SLICE_X1Y102_D6;
  wire [0:0] CLBLL_L_X2Y102_SLICE_X1Y102_DO5;
  wire [0:0] CLBLL_L_X2Y102_SLICE_X1Y102_DO6;
  wire [0:0] CLBLL_L_X2Y102_SLICE_X1Y102_D_CY;
  wire [0:0] CLBLL_L_X2Y102_SLICE_X1Y102_D_XOR;
  wire [0:0] CLBLL_L_X2Y136_SLICE_X0Y136_A;
  wire [0:0] CLBLL_L_X2Y136_SLICE_X0Y136_A1;
  wire [0:0] CLBLL_L_X2Y136_SLICE_X0Y136_A2;
  wire [0:0] CLBLL_L_X2Y136_SLICE_X0Y136_A3;
  wire [0:0] CLBLL_L_X2Y136_SLICE_X0Y136_A4;
  wire [0:0] CLBLL_L_X2Y136_SLICE_X0Y136_A5;
  wire [0:0] CLBLL_L_X2Y136_SLICE_X0Y136_A6;
  wire [0:0] CLBLL_L_X2Y136_SLICE_X0Y136_AO5;
  wire [0:0] CLBLL_L_X2Y136_SLICE_X0Y136_AO6;
  wire [0:0] CLBLL_L_X2Y136_SLICE_X0Y136_A_CY;
  wire [0:0] CLBLL_L_X2Y136_SLICE_X0Y136_A_XOR;
  wire [0:0] CLBLL_L_X2Y136_SLICE_X0Y136_B;
  wire [0:0] CLBLL_L_X2Y136_SLICE_X0Y136_B1;
  wire [0:0] CLBLL_L_X2Y136_SLICE_X0Y136_B2;
  wire [0:0] CLBLL_L_X2Y136_SLICE_X0Y136_B3;
  wire [0:0] CLBLL_L_X2Y136_SLICE_X0Y136_B4;
  wire [0:0] CLBLL_L_X2Y136_SLICE_X0Y136_B5;
  wire [0:0] CLBLL_L_X2Y136_SLICE_X0Y136_B6;
  wire [0:0] CLBLL_L_X2Y136_SLICE_X0Y136_BO5;
  wire [0:0] CLBLL_L_X2Y136_SLICE_X0Y136_BO6;
  wire [0:0] CLBLL_L_X2Y136_SLICE_X0Y136_B_CY;
  wire [0:0] CLBLL_L_X2Y136_SLICE_X0Y136_B_XOR;
  wire [0:0] CLBLL_L_X2Y136_SLICE_X0Y136_C;
  wire [0:0] CLBLL_L_X2Y136_SLICE_X0Y136_C1;
  wire [0:0] CLBLL_L_X2Y136_SLICE_X0Y136_C2;
  wire [0:0] CLBLL_L_X2Y136_SLICE_X0Y136_C3;
  wire [0:0] CLBLL_L_X2Y136_SLICE_X0Y136_C4;
  wire [0:0] CLBLL_L_X2Y136_SLICE_X0Y136_C5;
  wire [0:0] CLBLL_L_X2Y136_SLICE_X0Y136_C6;
  wire [0:0] CLBLL_L_X2Y136_SLICE_X0Y136_CO5;
  wire [0:0] CLBLL_L_X2Y136_SLICE_X0Y136_CO6;
  wire [0:0] CLBLL_L_X2Y136_SLICE_X0Y136_C_CY;
  wire [0:0] CLBLL_L_X2Y136_SLICE_X0Y136_C_XOR;
  wire [0:0] CLBLL_L_X2Y136_SLICE_X0Y136_D;
  wire [0:0] CLBLL_L_X2Y136_SLICE_X0Y136_D1;
  wire [0:0] CLBLL_L_X2Y136_SLICE_X0Y136_D2;
  wire [0:0] CLBLL_L_X2Y136_SLICE_X0Y136_D3;
  wire [0:0] CLBLL_L_X2Y136_SLICE_X0Y136_D4;
  wire [0:0] CLBLL_L_X2Y136_SLICE_X0Y136_D5;
  wire [0:0] CLBLL_L_X2Y136_SLICE_X0Y136_D6;
  wire [0:0] CLBLL_L_X2Y136_SLICE_X0Y136_DO5;
  wire [0:0] CLBLL_L_X2Y136_SLICE_X0Y136_DO6;
  wire [0:0] CLBLL_L_X2Y136_SLICE_X0Y136_D_CY;
  wire [0:0] CLBLL_L_X2Y136_SLICE_X0Y136_D_XOR;
  wire [0:0] CLBLL_L_X2Y136_SLICE_X1Y136_A;
  wire [0:0] CLBLL_L_X2Y136_SLICE_X1Y136_A1;
  wire [0:0] CLBLL_L_X2Y136_SLICE_X1Y136_A2;
  wire [0:0] CLBLL_L_X2Y136_SLICE_X1Y136_A3;
  wire [0:0] CLBLL_L_X2Y136_SLICE_X1Y136_A4;
  wire [0:0] CLBLL_L_X2Y136_SLICE_X1Y136_A5;
  wire [0:0] CLBLL_L_X2Y136_SLICE_X1Y136_A6;
  wire [0:0] CLBLL_L_X2Y136_SLICE_X1Y136_AO5;
  wire [0:0] CLBLL_L_X2Y136_SLICE_X1Y136_AO6;
  wire [0:0] CLBLL_L_X2Y136_SLICE_X1Y136_A_CY;
  wire [0:0] CLBLL_L_X2Y136_SLICE_X1Y136_A_XOR;
  wire [0:0] CLBLL_L_X2Y136_SLICE_X1Y136_B;
  wire [0:0] CLBLL_L_X2Y136_SLICE_X1Y136_B1;
  wire [0:0] CLBLL_L_X2Y136_SLICE_X1Y136_B2;
  wire [0:0] CLBLL_L_X2Y136_SLICE_X1Y136_B3;
  wire [0:0] CLBLL_L_X2Y136_SLICE_X1Y136_B4;
  wire [0:0] CLBLL_L_X2Y136_SLICE_X1Y136_B5;
  wire [0:0] CLBLL_L_X2Y136_SLICE_X1Y136_B6;
  wire [0:0] CLBLL_L_X2Y136_SLICE_X1Y136_BO5;
  wire [0:0] CLBLL_L_X2Y136_SLICE_X1Y136_BO6;
  wire [0:0] CLBLL_L_X2Y136_SLICE_X1Y136_B_CY;
  wire [0:0] CLBLL_L_X2Y136_SLICE_X1Y136_B_XOR;
  wire [0:0] CLBLL_L_X2Y136_SLICE_X1Y136_C;
  wire [0:0] CLBLL_L_X2Y136_SLICE_X1Y136_C1;
  wire [0:0] CLBLL_L_X2Y136_SLICE_X1Y136_C2;
  wire [0:0] CLBLL_L_X2Y136_SLICE_X1Y136_C3;
  wire [0:0] CLBLL_L_X2Y136_SLICE_X1Y136_C4;
  wire [0:0] CLBLL_L_X2Y136_SLICE_X1Y136_C5;
  wire [0:0] CLBLL_L_X2Y136_SLICE_X1Y136_C6;
  wire [0:0] CLBLL_L_X2Y136_SLICE_X1Y136_CO5;
  wire [0:0] CLBLL_L_X2Y136_SLICE_X1Y136_CO6;
  wire [0:0] CLBLL_L_X2Y136_SLICE_X1Y136_C_CY;
  wire [0:0] CLBLL_L_X2Y136_SLICE_X1Y136_C_XOR;
  wire [0:0] CLBLL_L_X2Y136_SLICE_X1Y136_D;
  wire [0:0] CLBLL_L_X2Y136_SLICE_X1Y136_D1;
  wire [0:0] CLBLL_L_X2Y136_SLICE_X1Y136_D2;
  wire [0:0] CLBLL_L_X2Y136_SLICE_X1Y136_D3;
  wire [0:0] CLBLL_L_X2Y136_SLICE_X1Y136_D4;
  wire [0:0] CLBLL_L_X2Y136_SLICE_X1Y136_D5;
  wire [0:0] CLBLL_L_X2Y136_SLICE_X1Y136_D6;
  wire [0:0] CLBLL_L_X2Y136_SLICE_X1Y136_DO5;
  wire [0:0] CLBLL_L_X2Y136_SLICE_X1Y136_DO6;
  wire [0:0] CLBLL_L_X2Y136_SLICE_X1Y136_D_CY;
  wire [0:0] CLBLL_L_X2Y136_SLICE_X1Y136_D_XOR;
  wire [0:0] CLBLL_L_X2Y146_SLICE_X0Y146_A;
  wire [0:0] CLBLL_L_X2Y146_SLICE_X0Y146_A1;
  wire [0:0] CLBLL_L_X2Y146_SLICE_X0Y146_A2;
  wire [0:0] CLBLL_L_X2Y146_SLICE_X0Y146_A3;
  wire [0:0] CLBLL_L_X2Y146_SLICE_X0Y146_A4;
  wire [0:0] CLBLL_L_X2Y146_SLICE_X0Y146_A5;
  wire [0:0] CLBLL_L_X2Y146_SLICE_X0Y146_A6;
  wire [0:0] CLBLL_L_X2Y146_SLICE_X0Y146_AO5;
  wire [0:0] CLBLL_L_X2Y146_SLICE_X0Y146_AO6;
  wire [0:0] CLBLL_L_X2Y146_SLICE_X0Y146_A_CY;
  wire [0:0] CLBLL_L_X2Y146_SLICE_X0Y146_A_XOR;
  wire [0:0] CLBLL_L_X2Y146_SLICE_X0Y146_B;
  wire [0:0] CLBLL_L_X2Y146_SLICE_X0Y146_B1;
  wire [0:0] CLBLL_L_X2Y146_SLICE_X0Y146_B2;
  wire [0:0] CLBLL_L_X2Y146_SLICE_X0Y146_B3;
  wire [0:0] CLBLL_L_X2Y146_SLICE_X0Y146_B4;
  wire [0:0] CLBLL_L_X2Y146_SLICE_X0Y146_B5;
  wire [0:0] CLBLL_L_X2Y146_SLICE_X0Y146_B6;
  wire [0:0] CLBLL_L_X2Y146_SLICE_X0Y146_BO5;
  wire [0:0] CLBLL_L_X2Y146_SLICE_X0Y146_BO6;
  wire [0:0] CLBLL_L_X2Y146_SLICE_X0Y146_B_CY;
  wire [0:0] CLBLL_L_X2Y146_SLICE_X0Y146_B_XOR;
  wire [0:0] CLBLL_L_X2Y146_SLICE_X0Y146_C;
  wire [0:0] CLBLL_L_X2Y146_SLICE_X0Y146_C1;
  wire [0:0] CLBLL_L_X2Y146_SLICE_X0Y146_C2;
  wire [0:0] CLBLL_L_X2Y146_SLICE_X0Y146_C3;
  wire [0:0] CLBLL_L_X2Y146_SLICE_X0Y146_C4;
  wire [0:0] CLBLL_L_X2Y146_SLICE_X0Y146_C5;
  wire [0:0] CLBLL_L_X2Y146_SLICE_X0Y146_C6;
  wire [0:0] CLBLL_L_X2Y146_SLICE_X0Y146_CO5;
  wire [0:0] CLBLL_L_X2Y146_SLICE_X0Y146_CO6;
  wire [0:0] CLBLL_L_X2Y146_SLICE_X0Y146_C_CY;
  wire [0:0] CLBLL_L_X2Y146_SLICE_X0Y146_C_XOR;
  wire [0:0] CLBLL_L_X2Y146_SLICE_X0Y146_D;
  wire [0:0] CLBLL_L_X2Y146_SLICE_X0Y146_D1;
  wire [0:0] CLBLL_L_X2Y146_SLICE_X0Y146_D2;
  wire [0:0] CLBLL_L_X2Y146_SLICE_X0Y146_D3;
  wire [0:0] CLBLL_L_X2Y146_SLICE_X0Y146_D4;
  wire [0:0] CLBLL_L_X2Y146_SLICE_X0Y146_D5;
  wire [0:0] CLBLL_L_X2Y146_SLICE_X0Y146_D6;
  wire [0:0] CLBLL_L_X2Y146_SLICE_X0Y146_DO5;
  wire [0:0] CLBLL_L_X2Y146_SLICE_X0Y146_DO6;
  wire [0:0] CLBLL_L_X2Y146_SLICE_X0Y146_D_CY;
  wire [0:0] CLBLL_L_X2Y146_SLICE_X0Y146_D_XOR;
  wire [0:0] CLBLL_L_X2Y146_SLICE_X1Y146_A;
  wire [0:0] CLBLL_L_X2Y146_SLICE_X1Y146_A1;
  wire [0:0] CLBLL_L_X2Y146_SLICE_X1Y146_A2;
  wire [0:0] CLBLL_L_X2Y146_SLICE_X1Y146_A3;
  wire [0:0] CLBLL_L_X2Y146_SLICE_X1Y146_A4;
  wire [0:0] CLBLL_L_X2Y146_SLICE_X1Y146_A5;
  wire [0:0] CLBLL_L_X2Y146_SLICE_X1Y146_A6;
  wire [0:0] CLBLL_L_X2Y146_SLICE_X1Y146_AMUX;
  wire [0:0] CLBLL_L_X2Y146_SLICE_X1Y146_AO5;
  wire [0:0] CLBLL_L_X2Y146_SLICE_X1Y146_AO6;
  wire [0:0] CLBLL_L_X2Y146_SLICE_X1Y146_A_CY;
  wire [0:0] CLBLL_L_X2Y146_SLICE_X1Y146_A_XOR;
  wire [0:0] CLBLL_L_X2Y146_SLICE_X1Y146_B;
  wire [0:0] CLBLL_L_X2Y146_SLICE_X1Y146_B1;
  wire [0:0] CLBLL_L_X2Y146_SLICE_X1Y146_B2;
  wire [0:0] CLBLL_L_X2Y146_SLICE_X1Y146_B3;
  wire [0:0] CLBLL_L_X2Y146_SLICE_X1Y146_B4;
  wire [0:0] CLBLL_L_X2Y146_SLICE_X1Y146_B5;
  wire [0:0] CLBLL_L_X2Y146_SLICE_X1Y146_B6;
  wire [0:0] CLBLL_L_X2Y146_SLICE_X1Y146_BO5;
  wire [0:0] CLBLL_L_X2Y146_SLICE_X1Y146_BO6;
  wire [0:0] CLBLL_L_X2Y146_SLICE_X1Y146_B_CY;
  wire [0:0] CLBLL_L_X2Y146_SLICE_X1Y146_B_XOR;
  wire [0:0] CLBLL_L_X2Y146_SLICE_X1Y146_C;
  wire [0:0] CLBLL_L_X2Y146_SLICE_X1Y146_C1;
  wire [0:0] CLBLL_L_X2Y146_SLICE_X1Y146_C2;
  wire [0:0] CLBLL_L_X2Y146_SLICE_X1Y146_C3;
  wire [0:0] CLBLL_L_X2Y146_SLICE_X1Y146_C4;
  wire [0:0] CLBLL_L_X2Y146_SLICE_X1Y146_C5;
  wire [0:0] CLBLL_L_X2Y146_SLICE_X1Y146_C6;
  wire [0:0] CLBLL_L_X2Y146_SLICE_X1Y146_CO5;
  wire [0:0] CLBLL_L_X2Y146_SLICE_X1Y146_CO6;
  wire [0:0] CLBLL_L_X2Y146_SLICE_X1Y146_C_CY;
  wire [0:0] CLBLL_L_X2Y146_SLICE_X1Y146_C_XOR;
  wire [0:0] CLBLL_L_X2Y146_SLICE_X1Y146_D;
  wire [0:0] CLBLL_L_X2Y146_SLICE_X1Y146_D1;
  wire [0:0] CLBLL_L_X2Y146_SLICE_X1Y146_D2;
  wire [0:0] CLBLL_L_X2Y146_SLICE_X1Y146_D3;
  wire [0:0] CLBLL_L_X2Y146_SLICE_X1Y146_D4;
  wire [0:0] CLBLL_L_X2Y146_SLICE_X1Y146_D5;
  wire [0:0] CLBLL_L_X2Y146_SLICE_X1Y146_D6;
  wire [0:0] CLBLL_L_X2Y146_SLICE_X1Y146_DO5;
  wire [0:0] CLBLL_L_X2Y146_SLICE_X1Y146_DO6;
  wire [0:0] CLBLL_L_X2Y146_SLICE_X1Y146_D_CY;
  wire [0:0] CLBLL_L_X2Y146_SLICE_X1Y146_D_XOR;
  wire [0:0] CLBLL_L_X2Y173_SLICE_X0Y173_A;
  wire [0:0] CLBLL_L_X2Y173_SLICE_X0Y173_A1;
  wire [0:0] CLBLL_L_X2Y173_SLICE_X0Y173_A2;
  wire [0:0] CLBLL_L_X2Y173_SLICE_X0Y173_A3;
  wire [0:0] CLBLL_L_X2Y173_SLICE_X0Y173_A4;
  wire [0:0] CLBLL_L_X2Y173_SLICE_X0Y173_A5;
  wire [0:0] CLBLL_L_X2Y173_SLICE_X0Y173_A6;
  wire [0:0] CLBLL_L_X2Y173_SLICE_X0Y173_AO5;
  wire [0:0] CLBLL_L_X2Y173_SLICE_X0Y173_AO6;
  wire [0:0] CLBLL_L_X2Y173_SLICE_X0Y173_A_CY;
  wire [0:0] CLBLL_L_X2Y173_SLICE_X0Y173_A_XOR;
  wire [0:0] CLBLL_L_X2Y173_SLICE_X0Y173_B;
  wire [0:0] CLBLL_L_X2Y173_SLICE_X0Y173_B1;
  wire [0:0] CLBLL_L_X2Y173_SLICE_X0Y173_B2;
  wire [0:0] CLBLL_L_X2Y173_SLICE_X0Y173_B3;
  wire [0:0] CLBLL_L_X2Y173_SLICE_X0Y173_B4;
  wire [0:0] CLBLL_L_X2Y173_SLICE_X0Y173_B5;
  wire [0:0] CLBLL_L_X2Y173_SLICE_X0Y173_B6;
  wire [0:0] CLBLL_L_X2Y173_SLICE_X0Y173_BO5;
  wire [0:0] CLBLL_L_X2Y173_SLICE_X0Y173_BO6;
  wire [0:0] CLBLL_L_X2Y173_SLICE_X0Y173_B_CY;
  wire [0:0] CLBLL_L_X2Y173_SLICE_X0Y173_B_XOR;
  wire [0:0] CLBLL_L_X2Y173_SLICE_X0Y173_C;
  wire [0:0] CLBLL_L_X2Y173_SLICE_X0Y173_C1;
  wire [0:0] CLBLL_L_X2Y173_SLICE_X0Y173_C2;
  wire [0:0] CLBLL_L_X2Y173_SLICE_X0Y173_C3;
  wire [0:0] CLBLL_L_X2Y173_SLICE_X0Y173_C4;
  wire [0:0] CLBLL_L_X2Y173_SLICE_X0Y173_C5;
  wire [0:0] CLBLL_L_X2Y173_SLICE_X0Y173_C6;
  wire [0:0] CLBLL_L_X2Y173_SLICE_X0Y173_CO5;
  wire [0:0] CLBLL_L_X2Y173_SLICE_X0Y173_CO6;
  wire [0:0] CLBLL_L_X2Y173_SLICE_X0Y173_C_CY;
  wire [0:0] CLBLL_L_X2Y173_SLICE_X0Y173_C_XOR;
  wire [0:0] CLBLL_L_X2Y173_SLICE_X0Y173_D;
  wire [0:0] CLBLL_L_X2Y173_SLICE_X0Y173_D1;
  wire [0:0] CLBLL_L_X2Y173_SLICE_X0Y173_D2;
  wire [0:0] CLBLL_L_X2Y173_SLICE_X0Y173_D3;
  wire [0:0] CLBLL_L_X2Y173_SLICE_X0Y173_D4;
  wire [0:0] CLBLL_L_X2Y173_SLICE_X0Y173_D5;
  wire [0:0] CLBLL_L_X2Y173_SLICE_X0Y173_D6;
  wire [0:0] CLBLL_L_X2Y173_SLICE_X0Y173_DO5;
  wire [0:0] CLBLL_L_X2Y173_SLICE_X0Y173_DO6;
  wire [0:0] CLBLL_L_X2Y173_SLICE_X0Y173_D_CY;
  wire [0:0] CLBLL_L_X2Y173_SLICE_X0Y173_D_XOR;
  wire [0:0] CLBLL_L_X2Y173_SLICE_X1Y173_A;
  wire [0:0] CLBLL_L_X2Y173_SLICE_X1Y173_A1;
  wire [0:0] CLBLL_L_X2Y173_SLICE_X1Y173_A2;
  wire [0:0] CLBLL_L_X2Y173_SLICE_X1Y173_A3;
  wire [0:0] CLBLL_L_X2Y173_SLICE_X1Y173_A4;
  wire [0:0] CLBLL_L_X2Y173_SLICE_X1Y173_A5;
  wire [0:0] CLBLL_L_X2Y173_SLICE_X1Y173_A6;
  wire [0:0] CLBLL_L_X2Y173_SLICE_X1Y173_AMUX;
  wire [0:0] CLBLL_L_X2Y173_SLICE_X1Y173_AO5;
  wire [0:0] CLBLL_L_X2Y173_SLICE_X1Y173_AO6;
  wire [0:0] CLBLL_L_X2Y173_SLICE_X1Y173_A_CY;
  wire [0:0] CLBLL_L_X2Y173_SLICE_X1Y173_A_XOR;
  wire [0:0] CLBLL_L_X2Y173_SLICE_X1Y173_B;
  wire [0:0] CLBLL_L_X2Y173_SLICE_X1Y173_B1;
  wire [0:0] CLBLL_L_X2Y173_SLICE_X1Y173_B2;
  wire [0:0] CLBLL_L_X2Y173_SLICE_X1Y173_B3;
  wire [0:0] CLBLL_L_X2Y173_SLICE_X1Y173_B4;
  wire [0:0] CLBLL_L_X2Y173_SLICE_X1Y173_B5;
  wire [0:0] CLBLL_L_X2Y173_SLICE_X1Y173_B6;
  wire [0:0] CLBLL_L_X2Y173_SLICE_X1Y173_BMUX;
  wire [0:0] CLBLL_L_X2Y173_SLICE_X1Y173_BO5;
  wire [0:0] CLBLL_L_X2Y173_SLICE_X1Y173_BO6;
  wire [0:0] CLBLL_L_X2Y173_SLICE_X1Y173_B_CY;
  wire [0:0] CLBLL_L_X2Y173_SLICE_X1Y173_B_XOR;
  wire [0:0] CLBLL_L_X2Y173_SLICE_X1Y173_C;
  wire [0:0] CLBLL_L_X2Y173_SLICE_X1Y173_C1;
  wire [0:0] CLBLL_L_X2Y173_SLICE_X1Y173_C2;
  wire [0:0] CLBLL_L_X2Y173_SLICE_X1Y173_C3;
  wire [0:0] CLBLL_L_X2Y173_SLICE_X1Y173_C4;
  wire [0:0] CLBLL_L_X2Y173_SLICE_X1Y173_C5;
  wire [0:0] CLBLL_L_X2Y173_SLICE_X1Y173_C6;
  wire [0:0] CLBLL_L_X2Y173_SLICE_X1Y173_CO5;
  wire [0:0] CLBLL_L_X2Y173_SLICE_X1Y173_CO6;
  wire [0:0] CLBLL_L_X2Y173_SLICE_X1Y173_C_CY;
  wire [0:0] CLBLL_L_X2Y173_SLICE_X1Y173_C_XOR;
  wire [0:0] CLBLL_L_X2Y173_SLICE_X1Y173_D;
  wire [0:0] CLBLL_L_X2Y173_SLICE_X1Y173_D1;
  wire [0:0] CLBLL_L_X2Y173_SLICE_X1Y173_D2;
  wire [0:0] CLBLL_L_X2Y173_SLICE_X1Y173_D3;
  wire [0:0] CLBLL_L_X2Y173_SLICE_X1Y173_D4;
  wire [0:0] CLBLL_L_X2Y173_SLICE_X1Y173_D5;
  wire [0:0] CLBLL_L_X2Y173_SLICE_X1Y173_D6;
  wire [0:0] CLBLL_L_X2Y173_SLICE_X1Y173_DO5;
  wire [0:0] CLBLL_L_X2Y173_SLICE_X1Y173_DO6;
  wire [0:0] CLBLL_L_X2Y173_SLICE_X1Y173_D_CY;
  wire [0:0] CLBLL_L_X2Y173_SLICE_X1Y173_D_XOR;
  wire [0:0] CLBLL_L_X2Y175_SLICE_X0Y175_A;
  wire [0:0] CLBLL_L_X2Y175_SLICE_X0Y175_A1;
  wire [0:0] CLBLL_L_X2Y175_SLICE_X0Y175_A2;
  wire [0:0] CLBLL_L_X2Y175_SLICE_X0Y175_A3;
  wire [0:0] CLBLL_L_X2Y175_SLICE_X0Y175_A4;
  wire [0:0] CLBLL_L_X2Y175_SLICE_X0Y175_A5;
  wire [0:0] CLBLL_L_X2Y175_SLICE_X0Y175_A6;
  wire [0:0] CLBLL_L_X2Y175_SLICE_X0Y175_AO5;
  wire [0:0] CLBLL_L_X2Y175_SLICE_X0Y175_AO6;
  wire [0:0] CLBLL_L_X2Y175_SLICE_X0Y175_A_CY;
  wire [0:0] CLBLL_L_X2Y175_SLICE_X0Y175_A_XOR;
  wire [0:0] CLBLL_L_X2Y175_SLICE_X0Y175_B;
  wire [0:0] CLBLL_L_X2Y175_SLICE_X0Y175_B1;
  wire [0:0] CLBLL_L_X2Y175_SLICE_X0Y175_B2;
  wire [0:0] CLBLL_L_X2Y175_SLICE_X0Y175_B3;
  wire [0:0] CLBLL_L_X2Y175_SLICE_X0Y175_B4;
  wire [0:0] CLBLL_L_X2Y175_SLICE_X0Y175_B5;
  wire [0:0] CLBLL_L_X2Y175_SLICE_X0Y175_B6;
  wire [0:0] CLBLL_L_X2Y175_SLICE_X0Y175_BO5;
  wire [0:0] CLBLL_L_X2Y175_SLICE_X0Y175_BO6;
  wire [0:0] CLBLL_L_X2Y175_SLICE_X0Y175_B_CY;
  wire [0:0] CLBLL_L_X2Y175_SLICE_X0Y175_B_XOR;
  wire [0:0] CLBLL_L_X2Y175_SLICE_X0Y175_C;
  wire [0:0] CLBLL_L_X2Y175_SLICE_X0Y175_C1;
  wire [0:0] CLBLL_L_X2Y175_SLICE_X0Y175_C2;
  wire [0:0] CLBLL_L_X2Y175_SLICE_X0Y175_C3;
  wire [0:0] CLBLL_L_X2Y175_SLICE_X0Y175_C4;
  wire [0:0] CLBLL_L_X2Y175_SLICE_X0Y175_C5;
  wire [0:0] CLBLL_L_X2Y175_SLICE_X0Y175_C6;
  wire [0:0] CLBLL_L_X2Y175_SLICE_X0Y175_CO5;
  wire [0:0] CLBLL_L_X2Y175_SLICE_X0Y175_CO6;
  wire [0:0] CLBLL_L_X2Y175_SLICE_X0Y175_C_CY;
  wire [0:0] CLBLL_L_X2Y175_SLICE_X0Y175_C_XOR;
  wire [0:0] CLBLL_L_X2Y175_SLICE_X0Y175_D;
  wire [0:0] CLBLL_L_X2Y175_SLICE_X0Y175_D1;
  wire [0:0] CLBLL_L_X2Y175_SLICE_X0Y175_D2;
  wire [0:0] CLBLL_L_X2Y175_SLICE_X0Y175_D3;
  wire [0:0] CLBLL_L_X2Y175_SLICE_X0Y175_D4;
  wire [0:0] CLBLL_L_X2Y175_SLICE_X0Y175_D5;
  wire [0:0] CLBLL_L_X2Y175_SLICE_X0Y175_D6;
  wire [0:0] CLBLL_L_X2Y175_SLICE_X0Y175_DO5;
  wire [0:0] CLBLL_L_X2Y175_SLICE_X0Y175_DO6;
  wire [0:0] CLBLL_L_X2Y175_SLICE_X0Y175_D_CY;
  wire [0:0] CLBLL_L_X2Y175_SLICE_X0Y175_D_XOR;
  wire [0:0] CLBLL_L_X2Y175_SLICE_X1Y175_A;
  wire [0:0] CLBLL_L_X2Y175_SLICE_X1Y175_A1;
  wire [0:0] CLBLL_L_X2Y175_SLICE_X1Y175_A2;
  wire [0:0] CLBLL_L_X2Y175_SLICE_X1Y175_A3;
  wire [0:0] CLBLL_L_X2Y175_SLICE_X1Y175_A4;
  wire [0:0] CLBLL_L_X2Y175_SLICE_X1Y175_A5;
  wire [0:0] CLBLL_L_X2Y175_SLICE_X1Y175_A6;
  wire [0:0] CLBLL_L_X2Y175_SLICE_X1Y175_AO5;
  wire [0:0] CLBLL_L_X2Y175_SLICE_X1Y175_AO6;
  wire [0:0] CLBLL_L_X2Y175_SLICE_X1Y175_A_CY;
  wire [0:0] CLBLL_L_X2Y175_SLICE_X1Y175_A_XOR;
  wire [0:0] CLBLL_L_X2Y175_SLICE_X1Y175_B;
  wire [0:0] CLBLL_L_X2Y175_SLICE_X1Y175_B1;
  wire [0:0] CLBLL_L_X2Y175_SLICE_X1Y175_B2;
  wire [0:0] CLBLL_L_X2Y175_SLICE_X1Y175_B3;
  wire [0:0] CLBLL_L_X2Y175_SLICE_X1Y175_B4;
  wire [0:0] CLBLL_L_X2Y175_SLICE_X1Y175_B5;
  wire [0:0] CLBLL_L_X2Y175_SLICE_X1Y175_B6;
  wire [0:0] CLBLL_L_X2Y175_SLICE_X1Y175_BO5;
  wire [0:0] CLBLL_L_X2Y175_SLICE_X1Y175_BO6;
  wire [0:0] CLBLL_L_X2Y175_SLICE_X1Y175_B_CY;
  wire [0:0] CLBLL_L_X2Y175_SLICE_X1Y175_B_XOR;
  wire [0:0] CLBLL_L_X2Y175_SLICE_X1Y175_C;
  wire [0:0] CLBLL_L_X2Y175_SLICE_X1Y175_C1;
  wire [0:0] CLBLL_L_X2Y175_SLICE_X1Y175_C2;
  wire [0:0] CLBLL_L_X2Y175_SLICE_X1Y175_C3;
  wire [0:0] CLBLL_L_X2Y175_SLICE_X1Y175_C4;
  wire [0:0] CLBLL_L_X2Y175_SLICE_X1Y175_C5;
  wire [0:0] CLBLL_L_X2Y175_SLICE_X1Y175_C6;
  wire [0:0] CLBLL_L_X2Y175_SLICE_X1Y175_CO5;
  wire [0:0] CLBLL_L_X2Y175_SLICE_X1Y175_CO6;
  wire [0:0] CLBLL_L_X2Y175_SLICE_X1Y175_C_CY;
  wire [0:0] CLBLL_L_X2Y175_SLICE_X1Y175_C_XOR;
  wire [0:0] CLBLL_L_X2Y175_SLICE_X1Y175_D;
  wire [0:0] CLBLL_L_X2Y175_SLICE_X1Y175_D1;
  wire [0:0] CLBLL_L_X2Y175_SLICE_X1Y175_D2;
  wire [0:0] CLBLL_L_X2Y175_SLICE_X1Y175_D3;
  wire [0:0] CLBLL_L_X2Y175_SLICE_X1Y175_D4;
  wire [0:0] CLBLL_L_X2Y175_SLICE_X1Y175_D5;
  wire [0:0] CLBLL_L_X2Y175_SLICE_X1Y175_D6;
  wire [0:0] CLBLL_L_X2Y175_SLICE_X1Y175_DO5;
  wire [0:0] CLBLL_L_X2Y175_SLICE_X1Y175_DO6;
  wire [0:0] CLBLL_L_X2Y175_SLICE_X1Y175_D_CY;
  wire [0:0] CLBLL_L_X2Y175_SLICE_X1Y175_D_XOR;
  wire [0:0] CLBLL_L_X2Y98_SLICE_X0Y98_A;
  wire [0:0] CLBLL_L_X2Y98_SLICE_X0Y98_A1;
  wire [0:0] CLBLL_L_X2Y98_SLICE_X0Y98_A2;
  wire [0:0] CLBLL_L_X2Y98_SLICE_X0Y98_A3;
  wire [0:0] CLBLL_L_X2Y98_SLICE_X0Y98_A4;
  wire [0:0] CLBLL_L_X2Y98_SLICE_X0Y98_A5;
  wire [0:0] CLBLL_L_X2Y98_SLICE_X0Y98_A6;
  wire [0:0] CLBLL_L_X2Y98_SLICE_X0Y98_AO5;
  wire [0:0] CLBLL_L_X2Y98_SLICE_X0Y98_AO6;
  wire [0:0] CLBLL_L_X2Y98_SLICE_X0Y98_A_CY;
  wire [0:0] CLBLL_L_X2Y98_SLICE_X0Y98_A_XOR;
  wire [0:0] CLBLL_L_X2Y98_SLICE_X0Y98_B;
  wire [0:0] CLBLL_L_X2Y98_SLICE_X0Y98_B1;
  wire [0:0] CLBLL_L_X2Y98_SLICE_X0Y98_B2;
  wire [0:0] CLBLL_L_X2Y98_SLICE_X0Y98_B3;
  wire [0:0] CLBLL_L_X2Y98_SLICE_X0Y98_B4;
  wire [0:0] CLBLL_L_X2Y98_SLICE_X0Y98_B5;
  wire [0:0] CLBLL_L_X2Y98_SLICE_X0Y98_B6;
  wire [0:0] CLBLL_L_X2Y98_SLICE_X0Y98_BO5;
  wire [0:0] CLBLL_L_X2Y98_SLICE_X0Y98_BO6;
  wire [0:0] CLBLL_L_X2Y98_SLICE_X0Y98_B_CY;
  wire [0:0] CLBLL_L_X2Y98_SLICE_X0Y98_B_XOR;
  wire [0:0] CLBLL_L_X2Y98_SLICE_X0Y98_C;
  wire [0:0] CLBLL_L_X2Y98_SLICE_X0Y98_C1;
  wire [0:0] CLBLL_L_X2Y98_SLICE_X0Y98_C2;
  wire [0:0] CLBLL_L_X2Y98_SLICE_X0Y98_C3;
  wire [0:0] CLBLL_L_X2Y98_SLICE_X0Y98_C4;
  wire [0:0] CLBLL_L_X2Y98_SLICE_X0Y98_C5;
  wire [0:0] CLBLL_L_X2Y98_SLICE_X0Y98_C6;
  wire [0:0] CLBLL_L_X2Y98_SLICE_X0Y98_CO5;
  wire [0:0] CLBLL_L_X2Y98_SLICE_X0Y98_CO6;
  wire [0:0] CLBLL_L_X2Y98_SLICE_X0Y98_C_CY;
  wire [0:0] CLBLL_L_X2Y98_SLICE_X0Y98_C_XOR;
  wire [0:0] CLBLL_L_X2Y98_SLICE_X0Y98_D;
  wire [0:0] CLBLL_L_X2Y98_SLICE_X0Y98_D1;
  wire [0:0] CLBLL_L_X2Y98_SLICE_X0Y98_D2;
  wire [0:0] CLBLL_L_X2Y98_SLICE_X0Y98_D3;
  wire [0:0] CLBLL_L_X2Y98_SLICE_X0Y98_D4;
  wire [0:0] CLBLL_L_X2Y98_SLICE_X0Y98_D5;
  wire [0:0] CLBLL_L_X2Y98_SLICE_X0Y98_D6;
  wire [0:0] CLBLL_L_X2Y98_SLICE_X0Y98_DO5;
  wire [0:0] CLBLL_L_X2Y98_SLICE_X0Y98_DO6;
  wire [0:0] CLBLL_L_X2Y98_SLICE_X0Y98_D_CY;
  wire [0:0] CLBLL_L_X2Y98_SLICE_X0Y98_D_XOR;
  wire [0:0] CLBLL_L_X2Y98_SLICE_X1Y98_A;
  wire [0:0] CLBLL_L_X2Y98_SLICE_X1Y98_A1;
  wire [0:0] CLBLL_L_X2Y98_SLICE_X1Y98_A2;
  wire [0:0] CLBLL_L_X2Y98_SLICE_X1Y98_A3;
  wire [0:0] CLBLL_L_X2Y98_SLICE_X1Y98_A4;
  wire [0:0] CLBLL_L_X2Y98_SLICE_X1Y98_A5;
  wire [0:0] CLBLL_L_X2Y98_SLICE_X1Y98_A6;
  wire [0:0] CLBLL_L_X2Y98_SLICE_X1Y98_AO5;
  wire [0:0] CLBLL_L_X2Y98_SLICE_X1Y98_AO6;
  wire [0:0] CLBLL_L_X2Y98_SLICE_X1Y98_A_CY;
  wire [0:0] CLBLL_L_X2Y98_SLICE_X1Y98_A_XOR;
  wire [0:0] CLBLL_L_X2Y98_SLICE_X1Y98_B;
  wire [0:0] CLBLL_L_X2Y98_SLICE_X1Y98_B1;
  wire [0:0] CLBLL_L_X2Y98_SLICE_X1Y98_B2;
  wire [0:0] CLBLL_L_X2Y98_SLICE_X1Y98_B3;
  wire [0:0] CLBLL_L_X2Y98_SLICE_X1Y98_B4;
  wire [0:0] CLBLL_L_X2Y98_SLICE_X1Y98_B5;
  wire [0:0] CLBLL_L_X2Y98_SLICE_X1Y98_B6;
  wire [0:0] CLBLL_L_X2Y98_SLICE_X1Y98_BO5;
  wire [0:0] CLBLL_L_X2Y98_SLICE_X1Y98_BO6;
  wire [0:0] CLBLL_L_X2Y98_SLICE_X1Y98_B_CY;
  wire [0:0] CLBLL_L_X2Y98_SLICE_X1Y98_B_XOR;
  wire [0:0] CLBLL_L_X2Y98_SLICE_X1Y98_C;
  wire [0:0] CLBLL_L_X2Y98_SLICE_X1Y98_C1;
  wire [0:0] CLBLL_L_X2Y98_SLICE_X1Y98_C2;
  wire [0:0] CLBLL_L_X2Y98_SLICE_X1Y98_C3;
  wire [0:0] CLBLL_L_X2Y98_SLICE_X1Y98_C4;
  wire [0:0] CLBLL_L_X2Y98_SLICE_X1Y98_C5;
  wire [0:0] CLBLL_L_X2Y98_SLICE_X1Y98_C6;
  wire [0:0] CLBLL_L_X2Y98_SLICE_X1Y98_CO5;
  wire [0:0] CLBLL_L_X2Y98_SLICE_X1Y98_CO6;
  wire [0:0] CLBLL_L_X2Y98_SLICE_X1Y98_C_CY;
  wire [0:0] CLBLL_L_X2Y98_SLICE_X1Y98_C_XOR;
  wire [0:0] CLBLL_L_X2Y98_SLICE_X1Y98_D;
  wire [0:0] CLBLL_L_X2Y98_SLICE_X1Y98_D1;
  wire [0:0] CLBLL_L_X2Y98_SLICE_X1Y98_D2;
  wire [0:0] CLBLL_L_X2Y98_SLICE_X1Y98_D3;
  wire [0:0] CLBLL_L_X2Y98_SLICE_X1Y98_D4;
  wire [0:0] CLBLL_L_X2Y98_SLICE_X1Y98_D5;
  wire [0:0] CLBLL_L_X2Y98_SLICE_X1Y98_D6;
  wire [0:0] CLBLL_L_X2Y98_SLICE_X1Y98_DO5;
  wire [0:0] CLBLL_L_X2Y98_SLICE_X1Y98_DO6;
  wire [0:0] CLBLL_L_X2Y98_SLICE_X1Y98_D_CY;
  wire [0:0] CLBLL_L_X2Y98_SLICE_X1Y98_D_XOR;
  wire [0:0] CLBLL_L_X36Y113_SLICE_X54Y113_A;
  wire [0:0] CLBLL_L_X36Y113_SLICE_X54Y113_A1;
  wire [0:0] CLBLL_L_X36Y113_SLICE_X54Y113_A2;
  wire [0:0] CLBLL_L_X36Y113_SLICE_X54Y113_A3;
  wire [0:0] CLBLL_L_X36Y113_SLICE_X54Y113_A4;
  wire [0:0] CLBLL_L_X36Y113_SLICE_X54Y113_A5;
  wire [0:0] CLBLL_L_X36Y113_SLICE_X54Y113_A6;
  wire [0:0] CLBLL_L_X36Y113_SLICE_X54Y113_AO5;
  wire [0:0] CLBLL_L_X36Y113_SLICE_X54Y113_AO6;
  wire [0:0] CLBLL_L_X36Y113_SLICE_X54Y113_A_CY;
  wire [0:0] CLBLL_L_X36Y113_SLICE_X54Y113_A_XOR;
  wire [0:0] CLBLL_L_X36Y113_SLICE_X54Y113_B;
  wire [0:0] CLBLL_L_X36Y113_SLICE_X54Y113_B1;
  wire [0:0] CLBLL_L_X36Y113_SLICE_X54Y113_B2;
  wire [0:0] CLBLL_L_X36Y113_SLICE_X54Y113_B3;
  wire [0:0] CLBLL_L_X36Y113_SLICE_X54Y113_B4;
  wire [0:0] CLBLL_L_X36Y113_SLICE_X54Y113_B5;
  wire [0:0] CLBLL_L_X36Y113_SLICE_X54Y113_B6;
  wire [0:0] CLBLL_L_X36Y113_SLICE_X54Y113_BO5;
  wire [0:0] CLBLL_L_X36Y113_SLICE_X54Y113_BO6;
  wire [0:0] CLBLL_L_X36Y113_SLICE_X54Y113_B_CY;
  wire [0:0] CLBLL_L_X36Y113_SLICE_X54Y113_B_XOR;
  wire [0:0] CLBLL_L_X36Y113_SLICE_X54Y113_C;
  wire [0:0] CLBLL_L_X36Y113_SLICE_X54Y113_C1;
  wire [0:0] CLBLL_L_X36Y113_SLICE_X54Y113_C2;
  wire [0:0] CLBLL_L_X36Y113_SLICE_X54Y113_C3;
  wire [0:0] CLBLL_L_X36Y113_SLICE_X54Y113_C4;
  wire [0:0] CLBLL_L_X36Y113_SLICE_X54Y113_C5;
  wire [0:0] CLBLL_L_X36Y113_SLICE_X54Y113_C6;
  wire [0:0] CLBLL_L_X36Y113_SLICE_X54Y113_CO5;
  wire [0:0] CLBLL_L_X36Y113_SLICE_X54Y113_CO6;
  wire [0:0] CLBLL_L_X36Y113_SLICE_X54Y113_C_CY;
  wire [0:0] CLBLL_L_X36Y113_SLICE_X54Y113_C_XOR;
  wire [0:0] CLBLL_L_X36Y113_SLICE_X54Y113_D;
  wire [0:0] CLBLL_L_X36Y113_SLICE_X54Y113_D1;
  wire [0:0] CLBLL_L_X36Y113_SLICE_X54Y113_D2;
  wire [0:0] CLBLL_L_X36Y113_SLICE_X54Y113_D3;
  wire [0:0] CLBLL_L_X36Y113_SLICE_X54Y113_D4;
  wire [0:0] CLBLL_L_X36Y113_SLICE_X54Y113_D5;
  wire [0:0] CLBLL_L_X36Y113_SLICE_X54Y113_D6;
  wire [0:0] CLBLL_L_X36Y113_SLICE_X54Y113_DO5;
  wire [0:0] CLBLL_L_X36Y113_SLICE_X54Y113_DO6;
  wire [0:0] CLBLL_L_X36Y113_SLICE_X54Y113_D_CY;
  wire [0:0] CLBLL_L_X36Y113_SLICE_X54Y113_D_XOR;
  wire [0:0] CLBLL_L_X36Y113_SLICE_X55Y113_A;
  wire [0:0] CLBLL_L_X36Y113_SLICE_X55Y113_A1;
  wire [0:0] CLBLL_L_X36Y113_SLICE_X55Y113_A2;
  wire [0:0] CLBLL_L_X36Y113_SLICE_X55Y113_A3;
  wire [0:0] CLBLL_L_X36Y113_SLICE_X55Y113_A4;
  wire [0:0] CLBLL_L_X36Y113_SLICE_X55Y113_A5;
  wire [0:0] CLBLL_L_X36Y113_SLICE_X55Y113_A6;
  wire [0:0] CLBLL_L_X36Y113_SLICE_X55Y113_AO5;
  wire [0:0] CLBLL_L_X36Y113_SLICE_X55Y113_AO6;
  wire [0:0] CLBLL_L_X36Y113_SLICE_X55Y113_A_CY;
  wire [0:0] CLBLL_L_X36Y113_SLICE_X55Y113_A_XOR;
  wire [0:0] CLBLL_L_X36Y113_SLICE_X55Y113_B;
  wire [0:0] CLBLL_L_X36Y113_SLICE_X55Y113_B1;
  wire [0:0] CLBLL_L_X36Y113_SLICE_X55Y113_B2;
  wire [0:0] CLBLL_L_X36Y113_SLICE_X55Y113_B3;
  wire [0:0] CLBLL_L_X36Y113_SLICE_X55Y113_B4;
  wire [0:0] CLBLL_L_X36Y113_SLICE_X55Y113_B5;
  wire [0:0] CLBLL_L_X36Y113_SLICE_X55Y113_B6;
  wire [0:0] CLBLL_L_X36Y113_SLICE_X55Y113_BO5;
  wire [0:0] CLBLL_L_X36Y113_SLICE_X55Y113_BO6;
  wire [0:0] CLBLL_L_X36Y113_SLICE_X55Y113_B_CY;
  wire [0:0] CLBLL_L_X36Y113_SLICE_X55Y113_B_XOR;
  wire [0:0] CLBLL_L_X36Y113_SLICE_X55Y113_C;
  wire [0:0] CLBLL_L_X36Y113_SLICE_X55Y113_C1;
  wire [0:0] CLBLL_L_X36Y113_SLICE_X55Y113_C2;
  wire [0:0] CLBLL_L_X36Y113_SLICE_X55Y113_C3;
  wire [0:0] CLBLL_L_X36Y113_SLICE_X55Y113_C4;
  wire [0:0] CLBLL_L_X36Y113_SLICE_X55Y113_C5;
  wire [0:0] CLBLL_L_X36Y113_SLICE_X55Y113_C6;
  wire [0:0] CLBLL_L_X36Y113_SLICE_X55Y113_CO5;
  wire [0:0] CLBLL_L_X36Y113_SLICE_X55Y113_CO6;
  wire [0:0] CLBLL_L_X36Y113_SLICE_X55Y113_C_CY;
  wire [0:0] CLBLL_L_X36Y113_SLICE_X55Y113_C_XOR;
  wire [0:0] CLBLL_L_X36Y113_SLICE_X55Y113_D;
  wire [0:0] CLBLL_L_X36Y113_SLICE_X55Y113_D1;
  wire [0:0] CLBLL_L_X36Y113_SLICE_X55Y113_D2;
  wire [0:0] CLBLL_L_X36Y113_SLICE_X55Y113_D3;
  wire [0:0] CLBLL_L_X36Y113_SLICE_X55Y113_D4;
  wire [0:0] CLBLL_L_X36Y113_SLICE_X55Y113_D5;
  wire [0:0] CLBLL_L_X36Y113_SLICE_X55Y113_D6;
  wire [0:0] CLBLL_L_X36Y113_SLICE_X55Y113_DO5;
  wire [0:0] CLBLL_L_X36Y113_SLICE_X55Y113_DO6;
  wire [0:0] CLBLL_L_X36Y113_SLICE_X55Y113_D_CY;
  wire [0:0] CLBLL_L_X36Y113_SLICE_X55Y113_D_XOR;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X4Y107_A;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X4Y107_A1;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X4Y107_A2;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X4Y107_A3;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X4Y107_A4;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X4Y107_A5;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X4Y107_A6;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X4Y107_AO5;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X4Y107_AO6;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X4Y107_A_CY;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X4Y107_A_XOR;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X4Y107_B;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X4Y107_B1;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X4Y107_B2;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X4Y107_B3;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X4Y107_B4;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X4Y107_B5;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X4Y107_B6;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X4Y107_BO5;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X4Y107_BO6;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X4Y107_B_CY;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X4Y107_B_XOR;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X4Y107_C;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X4Y107_C1;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X4Y107_C2;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X4Y107_C3;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X4Y107_C4;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X4Y107_C5;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X4Y107_C6;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X4Y107_CO5;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X4Y107_CO6;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X4Y107_C_CY;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X4Y107_C_XOR;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X4Y107_D;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X4Y107_D1;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X4Y107_D2;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X4Y107_D3;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X4Y107_D4;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X4Y107_D5;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X4Y107_D6;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X4Y107_DO5;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X4Y107_DO6;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X4Y107_D_CY;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X4Y107_D_XOR;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X5Y107_A;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X5Y107_A1;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X5Y107_A2;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X5Y107_A3;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X5Y107_A4;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X5Y107_A5;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X5Y107_A6;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X5Y107_AO5;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X5Y107_AO6;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X5Y107_A_CY;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X5Y107_A_XOR;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X5Y107_B;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X5Y107_B1;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X5Y107_B2;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X5Y107_B3;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X5Y107_B4;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X5Y107_B5;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X5Y107_B6;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X5Y107_BO5;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X5Y107_BO6;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X5Y107_B_CY;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X5Y107_B_XOR;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X5Y107_C;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X5Y107_C1;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X5Y107_C2;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X5Y107_C3;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X5Y107_C4;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X5Y107_C5;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X5Y107_C6;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X5Y107_CO5;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X5Y107_CO6;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X5Y107_C_CY;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X5Y107_C_XOR;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X5Y107_D;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X5Y107_D1;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X5Y107_D2;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X5Y107_D3;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X5Y107_D4;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X5Y107_D5;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X5Y107_D6;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X5Y107_DO5;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X5Y107_DO6;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X5Y107_D_CY;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X5Y107_D_XOR;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X4Y109_A;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X4Y109_A1;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X4Y109_A2;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X4Y109_A3;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X4Y109_A4;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X4Y109_A5;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X4Y109_A6;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X4Y109_AMUX;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X4Y109_AO5;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X4Y109_AO6;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X4Y109_A_CY;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X4Y109_A_XOR;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X4Y109_B;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X4Y109_B1;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X4Y109_B2;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X4Y109_B3;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X4Y109_B4;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X4Y109_B5;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X4Y109_B6;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X4Y109_BMUX;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X4Y109_BO5;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X4Y109_BO6;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X4Y109_B_CY;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X4Y109_B_XOR;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X4Y109_C;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X4Y109_C1;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X4Y109_C2;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X4Y109_C3;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X4Y109_C4;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X4Y109_C5;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X4Y109_C6;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X4Y109_CO5;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X4Y109_CO6;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X4Y109_C_CY;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X4Y109_C_XOR;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X4Y109_D;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X4Y109_D1;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X4Y109_D2;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X4Y109_D3;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X4Y109_D4;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X4Y109_D5;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X4Y109_D6;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X4Y109_DO5;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X4Y109_DO6;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X4Y109_D_CY;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X4Y109_D_XOR;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X5Y109_A;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X5Y109_A1;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X5Y109_A2;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X5Y109_A3;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X5Y109_A4;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X5Y109_A5;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X5Y109_A6;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X5Y109_AO5;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X5Y109_AO6;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X5Y109_A_CY;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X5Y109_A_XOR;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X5Y109_B;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X5Y109_B1;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X5Y109_B2;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X5Y109_B3;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X5Y109_B4;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X5Y109_B5;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X5Y109_B6;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X5Y109_BO5;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X5Y109_BO6;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X5Y109_B_CY;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X5Y109_B_XOR;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X5Y109_C;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X5Y109_C1;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X5Y109_C2;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X5Y109_C3;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X5Y109_C4;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X5Y109_C5;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X5Y109_C6;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X5Y109_CO5;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X5Y109_CO6;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X5Y109_C_CY;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X5Y109_C_XOR;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X5Y109_D;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X5Y109_D1;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X5Y109_D2;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X5Y109_D3;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X5Y109_D4;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X5Y109_D5;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X5Y109_D6;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X5Y109_DO5;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X5Y109_DO6;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X5Y109_D_CY;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X5Y109_D_XOR;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X4Y110_A;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X4Y110_A1;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X4Y110_A2;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X4Y110_A3;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X4Y110_A4;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X4Y110_A5;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X4Y110_A6;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X4Y110_AMUX;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X4Y110_AO5;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X4Y110_AO6;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X4Y110_A_CY;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X4Y110_A_XOR;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X4Y110_B;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X4Y110_B1;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X4Y110_B2;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X4Y110_B3;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X4Y110_B4;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X4Y110_B5;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X4Y110_B6;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X4Y110_BMUX;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X4Y110_BO5;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X4Y110_BO6;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X4Y110_B_CY;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X4Y110_B_XOR;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X4Y110_C;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X4Y110_C1;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X4Y110_C2;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X4Y110_C3;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X4Y110_C4;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X4Y110_C5;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X4Y110_C6;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X4Y110_CMUX;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X4Y110_CO5;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X4Y110_CO6;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X4Y110_C_CY;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X4Y110_C_XOR;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X4Y110_D;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X4Y110_D1;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X4Y110_D2;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X4Y110_D3;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X4Y110_D4;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X4Y110_D5;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X4Y110_D6;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X4Y110_DO5;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X4Y110_DO6;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X4Y110_D_CY;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X4Y110_D_XOR;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X5Y110_A;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X5Y110_A1;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X5Y110_A2;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X5Y110_A3;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X5Y110_A4;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X5Y110_A5;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X5Y110_A6;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X5Y110_AO5;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X5Y110_AO6;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X5Y110_A_CY;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X5Y110_A_XOR;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X5Y110_B;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X5Y110_B1;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X5Y110_B2;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X5Y110_B3;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X5Y110_B4;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X5Y110_B5;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X5Y110_B6;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X5Y110_BO5;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X5Y110_BO6;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X5Y110_B_CY;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X5Y110_B_XOR;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X5Y110_C;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X5Y110_C1;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X5Y110_C2;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X5Y110_C3;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X5Y110_C4;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X5Y110_C5;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X5Y110_C6;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X5Y110_CO5;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X5Y110_CO6;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X5Y110_C_CY;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X5Y110_C_XOR;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X5Y110_D;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X5Y110_D1;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X5Y110_D2;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X5Y110_D3;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X5Y110_D4;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X5Y110_D5;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X5Y110_D6;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X5Y110_DO5;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X5Y110_DO6;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X5Y110_D_CY;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X5Y110_D_XOR;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X4Y111_A;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X4Y111_A1;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X4Y111_A2;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X4Y111_A3;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X4Y111_A4;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X4Y111_A5;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X4Y111_A6;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X4Y111_AMUX;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X4Y111_AO5;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X4Y111_AO6;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X4Y111_A_CY;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X4Y111_A_XOR;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X4Y111_B;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X4Y111_B1;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X4Y111_B2;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X4Y111_B3;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X4Y111_B4;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X4Y111_B5;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X4Y111_B6;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X4Y111_BMUX;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X4Y111_BO5;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X4Y111_BO6;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X4Y111_B_CY;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X4Y111_B_XOR;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X4Y111_C;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X4Y111_C1;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X4Y111_C2;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X4Y111_C3;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X4Y111_C4;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X4Y111_C5;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X4Y111_C6;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X4Y111_CO5;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X4Y111_CO6;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X4Y111_C_CY;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X4Y111_C_XOR;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X4Y111_D;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X4Y111_D1;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X4Y111_D2;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X4Y111_D3;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X4Y111_D4;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X4Y111_D5;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X4Y111_D6;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X4Y111_DO5;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X4Y111_DO6;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X4Y111_D_CY;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X4Y111_D_XOR;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X5Y111_A;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X5Y111_A1;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X5Y111_A2;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X5Y111_A3;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X5Y111_A4;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X5Y111_A5;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X5Y111_A6;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X5Y111_AMUX;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X5Y111_AO5;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X5Y111_AO6;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X5Y111_A_CY;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X5Y111_A_XOR;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X5Y111_B;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X5Y111_B1;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X5Y111_B2;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X5Y111_B3;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X5Y111_B4;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X5Y111_B5;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X5Y111_B6;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X5Y111_BMUX;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X5Y111_BO5;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X5Y111_BO6;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X5Y111_B_CY;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X5Y111_B_XOR;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X5Y111_C;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X5Y111_C1;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X5Y111_C2;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X5Y111_C3;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X5Y111_C4;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X5Y111_C5;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X5Y111_C6;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X5Y111_CO5;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X5Y111_CO6;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X5Y111_C_CY;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X5Y111_C_XOR;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X5Y111_D;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X5Y111_D1;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X5Y111_D2;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X5Y111_D3;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X5Y111_D4;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X5Y111_D5;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X5Y111_D6;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X5Y111_DO5;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X5Y111_DO6;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X5Y111_D_CY;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X5Y111_D_XOR;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X4Y112_A;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X4Y112_A1;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X4Y112_A2;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X4Y112_A3;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X4Y112_A4;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X4Y112_A5;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X4Y112_A6;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X4Y112_AMUX;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X4Y112_AO5;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X4Y112_AO6;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X4Y112_A_CY;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X4Y112_A_XOR;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X4Y112_B;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X4Y112_B1;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X4Y112_B2;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X4Y112_B3;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X4Y112_B4;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X4Y112_B5;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X4Y112_B6;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X4Y112_BO5;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X4Y112_BO6;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X4Y112_B_CY;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X4Y112_B_XOR;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X4Y112_C;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X4Y112_C1;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X4Y112_C2;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X4Y112_C3;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X4Y112_C4;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X4Y112_C5;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X4Y112_C6;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X4Y112_CO5;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X4Y112_CO6;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X4Y112_C_CY;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X4Y112_C_XOR;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X4Y112_D;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X4Y112_D1;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X4Y112_D2;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X4Y112_D3;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X4Y112_D4;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X4Y112_D5;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X4Y112_D6;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X4Y112_DO5;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X4Y112_DO6;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X4Y112_D_CY;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X4Y112_D_XOR;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X5Y112_A;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X5Y112_A1;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X5Y112_A2;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X5Y112_A3;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X5Y112_A4;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X5Y112_A5;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X5Y112_A6;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X5Y112_AMUX;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X5Y112_AO5;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X5Y112_AO6;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X5Y112_A_CY;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X5Y112_A_XOR;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X5Y112_B;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X5Y112_B1;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X5Y112_B2;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X5Y112_B3;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X5Y112_B4;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X5Y112_B5;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X5Y112_B6;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X5Y112_BMUX;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X5Y112_BO5;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X5Y112_BO6;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X5Y112_B_CY;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X5Y112_B_XOR;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X5Y112_C;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X5Y112_C1;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X5Y112_C2;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X5Y112_C3;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X5Y112_C4;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X5Y112_C5;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X5Y112_C6;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X5Y112_CO5;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X5Y112_CO6;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X5Y112_C_CY;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X5Y112_C_XOR;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X5Y112_D;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X5Y112_D1;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X5Y112_D2;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X5Y112_D3;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X5Y112_D4;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X5Y112_D5;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X5Y112_D6;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X5Y112_DO5;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X5Y112_DO6;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X5Y112_D_CY;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X5Y112_D_XOR;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_A;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_A1;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_A2;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_A3;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_A4;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_A5;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_A6;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_AO5;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_AO6;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_A_CY;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_A_XOR;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_B;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_B1;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_B2;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_B3;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_B4;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_B5;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_B6;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_BO5;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_BO6;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_B_CY;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_B_XOR;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_C;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_C1;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_C2;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_C3;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_C4;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_C5;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_C6;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_CO5;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_CO6;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_C_CY;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_C_XOR;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_D;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_D1;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_D2;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_D3;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_D4;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_D5;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_D6;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_DO5;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_DO6;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_D_CY;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_D_XOR;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_A;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_A1;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_A2;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_A3;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_A4;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_A5;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_A6;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_AO5;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_AO6;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_A_CY;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_A_XOR;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_B;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_B1;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_B2;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_B3;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_B4;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_B5;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_B6;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_BO5;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_BO6;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_B_CY;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_B_XOR;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_C;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_C1;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_C2;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_C3;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_C4;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_C5;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_C6;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_CO5;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_CO6;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_C_CY;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_C_XOR;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_D;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_D1;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_D2;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_D3;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_D4;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_D5;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_D6;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_DO5;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_DO6;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_D_CY;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_D_XOR;
  wire [0:0] CLBLL_L_X4Y141_SLICE_X4Y141_A;
  wire [0:0] CLBLL_L_X4Y141_SLICE_X4Y141_A1;
  wire [0:0] CLBLL_L_X4Y141_SLICE_X4Y141_A2;
  wire [0:0] CLBLL_L_X4Y141_SLICE_X4Y141_A3;
  wire [0:0] CLBLL_L_X4Y141_SLICE_X4Y141_A4;
  wire [0:0] CLBLL_L_X4Y141_SLICE_X4Y141_A5;
  wire [0:0] CLBLL_L_X4Y141_SLICE_X4Y141_A6;
  wire [0:0] CLBLL_L_X4Y141_SLICE_X4Y141_AO5;
  wire [0:0] CLBLL_L_X4Y141_SLICE_X4Y141_AO6;
  wire [0:0] CLBLL_L_X4Y141_SLICE_X4Y141_A_CY;
  wire [0:0] CLBLL_L_X4Y141_SLICE_X4Y141_A_XOR;
  wire [0:0] CLBLL_L_X4Y141_SLICE_X4Y141_B;
  wire [0:0] CLBLL_L_X4Y141_SLICE_X4Y141_B1;
  wire [0:0] CLBLL_L_X4Y141_SLICE_X4Y141_B2;
  wire [0:0] CLBLL_L_X4Y141_SLICE_X4Y141_B3;
  wire [0:0] CLBLL_L_X4Y141_SLICE_X4Y141_B4;
  wire [0:0] CLBLL_L_X4Y141_SLICE_X4Y141_B5;
  wire [0:0] CLBLL_L_X4Y141_SLICE_X4Y141_B6;
  wire [0:0] CLBLL_L_X4Y141_SLICE_X4Y141_BO5;
  wire [0:0] CLBLL_L_X4Y141_SLICE_X4Y141_BO6;
  wire [0:0] CLBLL_L_X4Y141_SLICE_X4Y141_B_CY;
  wire [0:0] CLBLL_L_X4Y141_SLICE_X4Y141_B_XOR;
  wire [0:0] CLBLL_L_X4Y141_SLICE_X4Y141_C;
  wire [0:0] CLBLL_L_X4Y141_SLICE_X4Y141_C1;
  wire [0:0] CLBLL_L_X4Y141_SLICE_X4Y141_C2;
  wire [0:0] CLBLL_L_X4Y141_SLICE_X4Y141_C3;
  wire [0:0] CLBLL_L_X4Y141_SLICE_X4Y141_C4;
  wire [0:0] CLBLL_L_X4Y141_SLICE_X4Y141_C5;
  wire [0:0] CLBLL_L_X4Y141_SLICE_X4Y141_C6;
  wire [0:0] CLBLL_L_X4Y141_SLICE_X4Y141_CO5;
  wire [0:0] CLBLL_L_X4Y141_SLICE_X4Y141_CO6;
  wire [0:0] CLBLL_L_X4Y141_SLICE_X4Y141_C_CY;
  wire [0:0] CLBLL_L_X4Y141_SLICE_X4Y141_C_XOR;
  wire [0:0] CLBLL_L_X4Y141_SLICE_X4Y141_D;
  wire [0:0] CLBLL_L_X4Y141_SLICE_X4Y141_D1;
  wire [0:0] CLBLL_L_X4Y141_SLICE_X4Y141_D2;
  wire [0:0] CLBLL_L_X4Y141_SLICE_X4Y141_D3;
  wire [0:0] CLBLL_L_X4Y141_SLICE_X4Y141_D4;
  wire [0:0] CLBLL_L_X4Y141_SLICE_X4Y141_D5;
  wire [0:0] CLBLL_L_X4Y141_SLICE_X4Y141_D6;
  wire [0:0] CLBLL_L_X4Y141_SLICE_X4Y141_DO5;
  wire [0:0] CLBLL_L_X4Y141_SLICE_X4Y141_DO6;
  wire [0:0] CLBLL_L_X4Y141_SLICE_X4Y141_D_CY;
  wire [0:0] CLBLL_L_X4Y141_SLICE_X4Y141_D_XOR;
  wire [0:0] CLBLL_L_X4Y141_SLICE_X5Y141_A;
  wire [0:0] CLBLL_L_X4Y141_SLICE_X5Y141_A1;
  wire [0:0] CLBLL_L_X4Y141_SLICE_X5Y141_A2;
  wire [0:0] CLBLL_L_X4Y141_SLICE_X5Y141_A3;
  wire [0:0] CLBLL_L_X4Y141_SLICE_X5Y141_A4;
  wire [0:0] CLBLL_L_X4Y141_SLICE_X5Y141_A5;
  wire [0:0] CLBLL_L_X4Y141_SLICE_X5Y141_A6;
  wire [0:0] CLBLL_L_X4Y141_SLICE_X5Y141_AO5;
  wire [0:0] CLBLL_L_X4Y141_SLICE_X5Y141_AO6;
  wire [0:0] CLBLL_L_X4Y141_SLICE_X5Y141_A_CY;
  wire [0:0] CLBLL_L_X4Y141_SLICE_X5Y141_A_XOR;
  wire [0:0] CLBLL_L_X4Y141_SLICE_X5Y141_B;
  wire [0:0] CLBLL_L_X4Y141_SLICE_X5Y141_B1;
  wire [0:0] CLBLL_L_X4Y141_SLICE_X5Y141_B2;
  wire [0:0] CLBLL_L_X4Y141_SLICE_X5Y141_B3;
  wire [0:0] CLBLL_L_X4Y141_SLICE_X5Y141_B4;
  wire [0:0] CLBLL_L_X4Y141_SLICE_X5Y141_B5;
  wire [0:0] CLBLL_L_X4Y141_SLICE_X5Y141_B6;
  wire [0:0] CLBLL_L_X4Y141_SLICE_X5Y141_BO5;
  wire [0:0] CLBLL_L_X4Y141_SLICE_X5Y141_BO6;
  wire [0:0] CLBLL_L_X4Y141_SLICE_X5Y141_B_CY;
  wire [0:0] CLBLL_L_X4Y141_SLICE_X5Y141_B_XOR;
  wire [0:0] CLBLL_L_X4Y141_SLICE_X5Y141_C;
  wire [0:0] CLBLL_L_X4Y141_SLICE_X5Y141_C1;
  wire [0:0] CLBLL_L_X4Y141_SLICE_X5Y141_C2;
  wire [0:0] CLBLL_L_X4Y141_SLICE_X5Y141_C3;
  wire [0:0] CLBLL_L_X4Y141_SLICE_X5Y141_C4;
  wire [0:0] CLBLL_L_X4Y141_SLICE_X5Y141_C5;
  wire [0:0] CLBLL_L_X4Y141_SLICE_X5Y141_C6;
  wire [0:0] CLBLL_L_X4Y141_SLICE_X5Y141_CO5;
  wire [0:0] CLBLL_L_X4Y141_SLICE_X5Y141_CO6;
  wire [0:0] CLBLL_L_X4Y141_SLICE_X5Y141_C_CY;
  wire [0:0] CLBLL_L_X4Y141_SLICE_X5Y141_C_XOR;
  wire [0:0] CLBLL_L_X4Y141_SLICE_X5Y141_D;
  wire [0:0] CLBLL_L_X4Y141_SLICE_X5Y141_D1;
  wire [0:0] CLBLL_L_X4Y141_SLICE_X5Y141_D2;
  wire [0:0] CLBLL_L_X4Y141_SLICE_X5Y141_D3;
  wire [0:0] CLBLL_L_X4Y141_SLICE_X5Y141_D4;
  wire [0:0] CLBLL_L_X4Y141_SLICE_X5Y141_D5;
  wire [0:0] CLBLL_L_X4Y141_SLICE_X5Y141_D6;
  wire [0:0] CLBLL_L_X4Y141_SLICE_X5Y141_DO5;
  wire [0:0] CLBLL_L_X4Y141_SLICE_X5Y141_DO6;
  wire [0:0] CLBLL_L_X4Y141_SLICE_X5Y141_D_CY;
  wire [0:0] CLBLL_L_X4Y141_SLICE_X5Y141_D_XOR;
  wire [0:0] CLBLL_R_X57Y113_SLICE_X86Y113_A;
  wire [0:0] CLBLL_R_X57Y113_SLICE_X86Y113_A1;
  wire [0:0] CLBLL_R_X57Y113_SLICE_X86Y113_A2;
  wire [0:0] CLBLL_R_X57Y113_SLICE_X86Y113_A3;
  wire [0:0] CLBLL_R_X57Y113_SLICE_X86Y113_A4;
  wire [0:0] CLBLL_R_X57Y113_SLICE_X86Y113_A5;
  wire [0:0] CLBLL_R_X57Y113_SLICE_X86Y113_A6;
  wire [0:0] CLBLL_R_X57Y113_SLICE_X86Y113_AO5;
  wire [0:0] CLBLL_R_X57Y113_SLICE_X86Y113_AO6;
  wire [0:0] CLBLL_R_X57Y113_SLICE_X86Y113_A_CY;
  wire [0:0] CLBLL_R_X57Y113_SLICE_X86Y113_A_XOR;
  wire [0:0] CLBLL_R_X57Y113_SLICE_X86Y113_B;
  wire [0:0] CLBLL_R_X57Y113_SLICE_X86Y113_B1;
  wire [0:0] CLBLL_R_X57Y113_SLICE_X86Y113_B2;
  wire [0:0] CLBLL_R_X57Y113_SLICE_X86Y113_B3;
  wire [0:0] CLBLL_R_X57Y113_SLICE_X86Y113_B4;
  wire [0:0] CLBLL_R_X57Y113_SLICE_X86Y113_B5;
  wire [0:0] CLBLL_R_X57Y113_SLICE_X86Y113_B6;
  wire [0:0] CLBLL_R_X57Y113_SLICE_X86Y113_BO5;
  wire [0:0] CLBLL_R_X57Y113_SLICE_X86Y113_BO6;
  wire [0:0] CLBLL_R_X57Y113_SLICE_X86Y113_B_CY;
  wire [0:0] CLBLL_R_X57Y113_SLICE_X86Y113_B_XOR;
  wire [0:0] CLBLL_R_X57Y113_SLICE_X86Y113_C;
  wire [0:0] CLBLL_R_X57Y113_SLICE_X86Y113_C1;
  wire [0:0] CLBLL_R_X57Y113_SLICE_X86Y113_C2;
  wire [0:0] CLBLL_R_X57Y113_SLICE_X86Y113_C3;
  wire [0:0] CLBLL_R_X57Y113_SLICE_X86Y113_C4;
  wire [0:0] CLBLL_R_X57Y113_SLICE_X86Y113_C5;
  wire [0:0] CLBLL_R_X57Y113_SLICE_X86Y113_C6;
  wire [0:0] CLBLL_R_X57Y113_SLICE_X86Y113_CO5;
  wire [0:0] CLBLL_R_X57Y113_SLICE_X86Y113_CO6;
  wire [0:0] CLBLL_R_X57Y113_SLICE_X86Y113_C_CY;
  wire [0:0] CLBLL_R_X57Y113_SLICE_X86Y113_C_XOR;
  wire [0:0] CLBLL_R_X57Y113_SLICE_X86Y113_D;
  wire [0:0] CLBLL_R_X57Y113_SLICE_X86Y113_D1;
  wire [0:0] CLBLL_R_X57Y113_SLICE_X86Y113_D2;
  wire [0:0] CLBLL_R_X57Y113_SLICE_X86Y113_D3;
  wire [0:0] CLBLL_R_X57Y113_SLICE_X86Y113_D4;
  wire [0:0] CLBLL_R_X57Y113_SLICE_X86Y113_D5;
  wire [0:0] CLBLL_R_X57Y113_SLICE_X86Y113_D6;
  wire [0:0] CLBLL_R_X57Y113_SLICE_X86Y113_DO5;
  wire [0:0] CLBLL_R_X57Y113_SLICE_X86Y113_DO6;
  wire [0:0] CLBLL_R_X57Y113_SLICE_X86Y113_D_CY;
  wire [0:0] CLBLL_R_X57Y113_SLICE_X86Y113_D_XOR;
  wire [0:0] CLBLL_R_X57Y113_SLICE_X87Y113_A;
  wire [0:0] CLBLL_R_X57Y113_SLICE_X87Y113_A1;
  wire [0:0] CLBLL_R_X57Y113_SLICE_X87Y113_A2;
  wire [0:0] CLBLL_R_X57Y113_SLICE_X87Y113_A3;
  wire [0:0] CLBLL_R_X57Y113_SLICE_X87Y113_A4;
  wire [0:0] CLBLL_R_X57Y113_SLICE_X87Y113_A5;
  wire [0:0] CLBLL_R_X57Y113_SLICE_X87Y113_A6;
  wire [0:0] CLBLL_R_X57Y113_SLICE_X87Y113_AO5;
  wire [0:0] CLBLL_R_X57Y113_SLICE_X87Y113_AO6;
  wire [0:0] CLBLL_R_X57Y113_SLICE_X87Y113_A_CY;
  wire [0:0] CLBLL_R_X57Y113_SLICE_X87Y113_A_XOR;
  wire [0:0] CLBLL_R_X57Y113_SLICE_X87Y113_B;
  wire [0:0] CLBLL_R_X57Y113_SLICE_X87Y113_B1;
  wire [0:0] CLBLL_R_X57Y113_SLICE_X87Y113_B2;
  wire [0:0] CLBLL_R_X57Y113_SLICE_X87Y113_B3;
  wire [0:0] CLBLL_R_X57Y113_SLICE_X87Y113_B4;
  wire [0:0] CLBLL_R_X57Y113_SLICE_X87Y113_B5;
  wire [0:0] CLBLL_R_X57Y113_SLICE_X87Y113_B6;
  wire [0:0] CLBLL_R_X57Y113_SLICE_X87Y113_BO5;
  wire [0:0] CLBLL_R_X57Y113_SLICE_X87Y113_BO6;
  wire [0:0] CLBLL_R_X57Y113_SLICE_X87Y113_B_CY;
  wire [0:0] CLBLL_R_X57Y113_SLICE_X87Y113_B_XOR;
  wire [0:0] CLBLL_R_X57Y113_SLICE_X87Y113_C;
  wire [0:0] CLBLL_R_X57Y113_SLICE_X87Y113_C1;
  wire [0:0] CLBLL_R_X57Y113_SLICE_X87Y113_C2;
  wire [0:0] CLBLL_R_X57Y113_SLICE_X87Y113_C3;
  wire [0:0] CLBLL_R_X57Y113_SLICE_X87Y113_C4;
  wire [0:0] CLBLL_R_X57Y113_SLICE_X87Y113_C5;
  wire [0:0] CLBLL_R_X57Y113_SLICE_X87Y113_C6;
  wire [0:0] CLBLL_R_X57Y113_SLICE_X87Y113_CO5;
  wire [0:0] CLBLL_R_X57Y113_SLICE_X87Y113_CO6;
  wire [0:0] CLBLL_R_X57Y113_SLICE_X87Y113_C_CY;
  wire [0:0] CLBLL_R_X57Y113_SLICE_X87Y113_C_XOR;
  wire [0:0] CLBLL_R_X57Y113_SLICE_X87Y113_D;
  wire [0:0] CLBLL_R_X57Y113_SLICE_X87Y113_D1;
  wire [0:0] CLBLL_R_X57Y113_SLICE_X87Y113_D2;
  wire [0:0] CLBLL_R_X57Y113_SLICE_X87Y113_D3;
  wire [0:0] CLBLL_R_X57Y113_SLICE_X87Y113_D4;
  wire [0:0] CLBLL_R_X57Y113_SLICE_X87Y113_D5;
  wire [0:0] CLBLL_R_X57Y113_SLICE_X87Y113_D6;
  wire [0:0] CLBLL_R_X57Y113_SLICE_X87Y113_DO5;
  wire [0:0] CLBLL_R_X57Y113_SLICE_X87Y113_DO6;
  wire [0:0] CLBLL_R_X57Y113_SLICE_X87Y113_D_CY;
  wire [0:0] CLBLL_R_X57Y113_SLICE_X87Y113_D_XOR;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X12Y113_A;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X12Y113_A1;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X12Y113_A2;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X12Y113_A3;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X12Y113_A4;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X12Y113_A5;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X12Y113_A6;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X12Y113_AO5;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X12Y113_AO6;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X12Y113_A_CY;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X12Y113_A_XOR;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X12Y113_B;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X12Y113_B1;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X12Y113_B2;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X12Y113_B3;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X12Y113_B4;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X12Y113_B5;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X12Y113_B6;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X12Y113_BO5;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X12Y113_BO6;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X12Y113_B_CY;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X12Y113_B_XOR;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X12Y113_C;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X12Y113_C1;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X12Y113_C2;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X12Y113_C3;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X12Y113_C4;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X12Y113_C5;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X12Y113_C6;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X12Y113_CO5;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X12Y113_CO6;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X12Y113_C_CY;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X12Y113_C_XOR;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X12Y113_D;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X12Y113_D1;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X12Y113_D2;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X12Y113_D3;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X12Y113_D4;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X12Y113_D5;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X12Y113_D6;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X12Y113_DO5;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X12Y113_DO6;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X12Y113_D_CY;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X12Y113_D_XOR;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X13Y113_A;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X13Y113_A1;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X13Y113_A2;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X13Y113_A3;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X13Y113_A4;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X13Y113_A5;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X13Y113_A6;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X13Y113_AO5;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X13Y113_AO6;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X13Y113_A_CY;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X13Y113_A_XOR;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X13Y113_B;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X13Y113_B1;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X13Y113_B2;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X13Y113_B3;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X13Y113_B4;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X13Y113_B5;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X13Y113_B6;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X13Y113_BO5;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X13Y113_BO6;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X13Y113_B_CY;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X13Y113_B_XOR;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X13Y113_C;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X13Y113_C1;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X13Y113_C2;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X13Y113_C3;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X13Y113_C4;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X13Y113_C5;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X13Y113_C6;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X13Y113_CO5;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X13Y113_CO6;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X13Y113_C_CY;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X13Y113_C_XOR;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X13Y113_D;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X13Y113_D1;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X13Y113_D2;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X13Y113_D3;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X13Y113_D4;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X13Y113_D5;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X13Y113_D6;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X13Y113_DO5;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X13Y113_DO6;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X13Y113_D_CY;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X13Y113_D_XOR;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X12Y114_A;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X12Y114_A1;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X12Y114_A2;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X12Y114_A3;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X12Y114_A4;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X12Y114_A5;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X12Y114_A6;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X12Y114_AO5;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X12Y114_AO6;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X12Y114_A_CY;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X12Y114_A_XOR;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X12Y114_B;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X12Y114_B1;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X12Y114_B2;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X12Y114_B3;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X12Y114_B4;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X12Y114_B5;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X12Y114_B6;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X12Y114_BO5;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X12Y114_BO6;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X12Y114_B_CY;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X12Y114_B_XOR;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X12Y114_C;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X12Y114_C1;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X12Y114_C2;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X12Y114_C3;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X12Y114_C4;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X12Y114_C5;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X12Y114_C6;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X12Y114_CO5;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X12Y114_CO6;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X12Y114_C_CY;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X12Y114_C_XOR;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X12Y114_D;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X12Y114_D1;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X12Y114_D2;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X12Y114_D3;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X12Y114_D4;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X12Y114_D5;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X12Y114_D6;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X12Y114_DO5;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X12Y114_DO6;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X12Y114_D_CY;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X12Y114_D_XOR;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X13Y114_A;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X13Y114_A1;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X13Y114_A2;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X13Y114_A3;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X13Y114_A4;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X13Y114_A5;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X13Y114_A6;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X13Y114_AO5;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X13Y114_AO6;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X13Y114_A_CY;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X13Y114_A_XOR;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X13Y114_B;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X13Y114_B1;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X13Y114_B2;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X13Y114_B3;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X13Y114_B4;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X13Y114_B5;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X13Y114_B6;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X13Y114_BO5;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X13Y114_BO6;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X13Y114_B_CY;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X13Y114_B_XOR;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X13Y114_C;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X13Y114_C1;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X13Y114_C2;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X13Y114_C3;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X13Y114_C4;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X13Y114_C5;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X13Y114_C6;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X13Y114_CO5;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X13Y114_CO6;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X13Y114_C_CY;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X13Y114_C_XOR;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X13Y114_D;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X13Y114_D1;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X13Y114_D2;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X13Y114_D3;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X13Y114_D4;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X13Y114_D5;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X13Y114_D6;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X13Y114_DO5;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X13Y114_DO6;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X13Y114_D_CY;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X13Y114_D_XOR;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X12Y123_A;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X12Y123_A1;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X12Y123_A2;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X12Y123_A3;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X12Y123_A4;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X12Y123_A5;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X12Y123_A6;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X12Y123_AO5;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X12Y123_AO6;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X12Y123_A_CY;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X12Y123_A_XOR;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X12Y123_B;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X12Y123_B1;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X12Y123_B2;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X12Y123_B3;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X12Y123_B4;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X12Y123_B5;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X12Y123_B6;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X12Y123_BO5;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X12Y123_BO6;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X12Y123_B_CY;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X12Y123_B_XOR;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X12Y123_C;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X12Y123_C1;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X12Y123_C2;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X12Y123_C3;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X12Y123_C4;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X12Y123_C5;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X12Y123_C6;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X12Y123_CO5;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X12Y123_CO6;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X12Y123_C_CY;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X12Y123_C_XOR;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X12Y123_D;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X12Y123_D1;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X12Y123_D2;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X12Y123_D3;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X12Y123_D4;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X12Y123_D5;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X12Y123_D6;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X12Y123_DO5;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X12Y123_DO6;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X12Y123_D_CY;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X12Y123_D_XOR;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X13Y123_A;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X13Y123_A1;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X13Y123_A2;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X13Y123_A3;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X13Y123_A4;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X13Y123_A5;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X13Y123_A6;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X13Y123_AO5;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X13Y123_AO6;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X13Y123_A_CY;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X13Y123_A_XOR;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X13Y123_B;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X13Y123_B1;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X13Y123_B2;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X13Y123_B3;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X13Y123_B4;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X13Y123_B5;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X13Y123_B6;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X13Y123_BO5;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X13Y123_BO6;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X13Y123_B_CY;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X13Y123_B_XOR;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X13Y123_C;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X13Y123_C1;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X13Y123_C2;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X13Y123_C3;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X13Y123_C4;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X13Y123_C5;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X13Y123_C6;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X13Y123_CO5;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X13Y123_CO6;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X13Y123_C_CY;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X13Y123_C_XOR;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X13Y123_D;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X13Y123_D1;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X13Y123_D2;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X13Y123_D3;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X13Y123_D4;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X13Y123_D5;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X13Y123_D6;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X13Y123_DO5;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X13Y123_DO6;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X13Y123_D_CY;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X13Y123_D_XOR;
  wire [0:0] CLBLM_L_X56Y119_SLICE_X84Y119_A;
  wire [0:0] CLBLM_L_X56Y119_SLICE_X84Y119_A1;
  wire [0:0] CLBLM_L_X56Y119_SLICE_X84Y119_A2;
  wire [0:0] CLBLM_L_X56Y119_SLICE_X84Y119_A3;
  wire [0:0] CLBLM_L_X56Y119_SLICE_X84Y119_A4;
  wire [0:0] CLBLM_L_X56Y119_SLICE_X84Y119_A5;
  wire [0:0] CLBLM_L_X56Y119_SLICE_X84Y119_A6;
  wire [0:0] CLBLM_L_X56Y119_SLICE_X84Y119_AMUX;
  wire [0:0] CLBLM_L_X56Y119_SLICE_X84Y119_AO5;
  wire [0:0] CLBLM_L_X56Y119_SLICE_X84Y119_AO6;
  wire [0:0] CLBLM_L_X56Y119_SLICE_X84Y119_A_CY;
  wire [0:0] CLBLM_L_X56Y119_SLICE_X84Y119_A_XOR;
  wire [0:0] CLBLM_L_X56Y119_SLICE_X84Y119_B;
  wire [0:0] CLBLM_L_X56Y119_SLICE_X84Y119_B1;
  wire [0:0] CLBLM_L_X56Y119_SLICE_X84Y119_B2;
  wire [0:0] CLBLM_L_X56Y119_SLICE_X84Y119_B3;
  wire [0:0] CLBLM_L_X56Y119_SLICE_X84Y119_B4;
  wire [0:0] CLBLM_L_X56Y119_SLICE_X84Y119_B5;
  wire [0:0] CLBLM_L_X56Y119_SLICE_X84Y119_B6;
  wire [0:0] CLBLM_L_X56Y119_SLICE_X84Y119_BO5;
  wire [0:0] CLBLM_L_X56Y119_SLICE_X84Y119_BO6;
  wire [0:0] CLBLM_L_X56Y119_SLICE_X84Y119_B_CY;
  wire [0:0] CLBLM_L_X56Y119_SLICE_X84Y119_B_XOR;
  wire [0:0] CLBLM_L_X56Y119_SLICE_X84Y119_C;
  wire [0:0] CLBLM_L_X56Y119_SLICE_X84Y119_C1;
  wire [0:0] CLBLM_L_X56Y119_SLICE_X84Y119_C2;
  wire [0:0] CLBLM_L_X56Y119_SLICE_X84Y119_C3;
  wire [0:0] CLBLM_L_X56Y119_SLICE_X84Y119_C4;
  wire [0:0] CLBLM_L_X56Y119_SLICE_X84Y119_C5;
  wire [0:0] CLBLM_L_X56Y119_SLICE_X84Y119_C6;
  wire [0:0] CLBLM_L_X56Y119_SLICE_X84Y119_CO5;
  wire [0:0] CLBLM_L_X56Y119_SLICE_X84Y119_CO6;
  wire [0:0] CLBLM_L_X56Y119_SLICE_X84Y119_C_CY;
  wire [0:0] CLBLM_L_X56Y119_SLICE_X84Y119_C_XOR;
  wire [0:0] CLBLM_L_X56Y119_SLICE_X84Y119_D;
  wire [0:0] CLBLM_L_X56Y119_SLICE_X84Y119_D1;
  wire [0:0] CLBLM_L_X56Y119_SLICE_X84Y119_D2;
  wire [0:0] CLBLM_L_X56Y119_SLICE_X84Y119_D3;
  wire [0:0] CLBLM_L_X56Y119_SLICE_X84Y119_D4;
  wire [0:0] CLBLM_L_X56Y119_SLICE_X84Y119_D5;
  wire [0:0] CLBLM_L_X56Y119_SLICE_X84Y119_D6;
  wire [0:0] CLBLM_L_X56Y119_SLICE_X84Y119_DO5;
  wire [0:0] CLBLM_L_X56Y119_SLICE_X84Y119_DO6;
  wire [0:0] CLBLM_L_X56Y119_SLICE_X84Y119_D_CY;
  wire [0:0] CLBLM_L_X56Y119_SLICE_X84Y119_D_XOR;
  wire [0:0] CLBLM_L_X56Y119_SLICE_X85Y119_A;
  wire [0:0] CLBLM_L_X56Y119_SLICE_X85Y119_A1;
  wire [0:0] CLBLM_L_X56Y119_SLICE_X85Y119_A2;
  wire [0:0] CLBLM_L_X56Y119_SLICE_X85Y119_A3;
  wire [0:0] CLBLM_L_X56Y119_SLICE_X85Y119_A4;
  wire [0:0] CLBLM_L_X56Y119_SLICE_X85Y119_A5;
  wire [0:0] CLBLM_L_X56Y119_SLICE_X85Y119_A6;
  wire [0:0] CLBLM_L_X56Y119_SLICE_X85Y119_AO5;
  wire [0:0] CLBLM_L_X56Y119_SLICE_X85Y119_AO6;
  wire [0:0] CLBLM_L_X56Y119_SLICE_X85Y119_A_CY;
  wire [0:0] CLBLM_L_X56Y119_SLICE_X85Y119_A_XOR;
  wire [0:0] CLBLM_L_X56Y119_SLICE_X85Y119_B;
  wire [0:0] CLBLM_L_X56Y119_SLICE_X85Y119_B1;
  wire [0:0] CLBLM_L_X56Y119_SLICE_X85Y119_B2;
  wire [0:0] CLBLM_L_X56Y119_SLICE_X85Y119_B3;
  wire [0:0] CLBLM_L_X56Y119_SLICE_X85Y119_B4;
  wire [0:0] CLBLM_L_X56Y119_SLICE_X85Y119_B5;
  wire [0:0] CLBLM_L_X56Y119_SLICE_X85Y119_B6;
  wire [0:0] CLBLM_L_X56Y119_SLICE_X85Y119_BO5;
  wire [0:0] CLBLM_L_X56Y119_SLICE_X85Y119_BO6;
  wire [0:0] CLBLM_L_X56Y119_SLICE_X85Y119_B_CY;
  wire [0:0] CLBLM_L_X56Y119_SLICE_X85Y119_B_XOR;
  wire [0:0] CLBLM_L_X56Y119_SLICE_X85Y119_C;
  wire [0:0] CLBLM_L_X56Y119_SLICE_X85Y119_C1;
  wire [0:0] CLBLM_L_X56Y119_SLICE_X85Y119_C2;
  wire [0:0] CLBLM_L_X56Y119_SLICE_X85Y119_C3;
  wire [0:0] CLBLM_L_X56Y119_SLICE_X85Y119_C4;
  wire [0:0] CLBLM_L_X56Y119_SLICE_X85Y119_C5;
  wire [0:0] CLBLM_L_X56Y119_SLICE_X85Y119_C6;
  wire [0:0] CLBLM_L_X56Y119_SLICE_X85Y119_CO5;
  wire [0:0] CLBLM_L_X56Y119_SLICE_X85Y119_CO6;
  wire [0:0] CLBLM_L_X56Y119_SLICE_X85Y119_C_CY;
  wire [0:0] CLBLM_L_X56Y119_SLICE_X85Y119_C_XOR;
  wire [0:0] CLBLM_L_X56Y119_SLICE_X85Y119_D;
  wire [0:0] CLBLM_L_X56Y119_SLICE_X85Y119_D1;
  wire [0:0] CLBLM_L_X56Y119_SLICE_X85Y119_D2;
  wire [0:0] CLBLM_L_X56Y119_SLICE_X85Y119_D3;
  wire [0:0] CLBLM_L_X56Y119_SLICE_X85Y119_D4;
  wire [0:0] CLBLM_L_X56Y119_SLICE_X85Y119_D5;
  wire [0:0] CLBLM_L_X56Y119_SLICE_X85Y119_D6;
  wire [0:0] CLBLM_L_X56Y119_SLICE_X85Y119_DO5;
  wire [0:0] CLBLM_L_X56Y119_SLICE_X85Y119_DO6;
  wire [0:0] CLBLM_L_X56Y119_SLICE_X85Y119_D_CY;
  wire [0:0] CLBLM_L_X56Y119_SLICE_X85Y119_D_XOR;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X10Y113_A;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X10Y113_A1;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X10Y113_A2;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X10Y113_A3;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X10Y113_A4;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X10Y113_A5;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X10Y113_A6;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X10Y113_AMUX;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X10Y113_AO5;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X10Y113_AO6;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X10Y113_A_CY;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X10Y113_A_XOR;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X10Y113_B;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X10Y113_B1;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X10Y113_B2;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X10Y113_B3;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X10Y113_B4;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X10Y113_B5;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X10Y113_B6;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X10Y113_BO5;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X10Y113_BO6;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X10Y113_B_CY;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X10Y113_B_XOR;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X10Y113_C;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X10Y113_C1;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X10Y113_C2;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X10Y113_C3;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X10Y113_C4;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X10Y113_C5;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X10Y113_C6;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X10Y113_CO5;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X10Y113_CO6;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X10Y113_C_CY;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X10Y113_C_XOR;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X10Y113_D;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X10Y113_D1;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X10Y113_D2;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X10Y113_D3;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X10Y113_D4;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X10Y113_D5;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X10Y113_D6;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X10Y113_DO5;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X10Y113_DO6;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X10Y113_D_CY;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X10Y113_D_XOR;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X11Y113_A;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X11Y113_A1;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X11Y113_A2;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X11Y113_A3;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X11Y113_A4;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X11Y113_A5;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X11Y113_A6;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X11Y113_AMUX;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X11Y113_AO5;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X11Y113_AO6;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X11Y113_A_CY;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X11Y113_A_XOR;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X11Y113_B;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X11Y113_B1;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X11Y113_B2;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X11Y113_B3;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X11Y113_B4;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X11Y113_B5;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X11Y113_B6;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X11Y113_BO5;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X11Y113_BO6;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X11Y113_B_CY;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X11Y113_B_XOR;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X11Y113_C;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X11Y113_C1;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X11Y113_C2;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X11Y113_C3;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X11Y113_C4;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X11Y113_C5;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X11Y113_C6;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X11Y113_CO5;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X11Y113_CO6;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X11Y113_C_CY;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X11Y113_C_XOR;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X11Y113_D;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X11Y113_D1;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X11Y113_D2;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X11Y113_D3;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X11Y113_D4;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X11Y113_D5;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X11Y113_D6;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X11Y113_DO5;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X11Y113_DO6;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X11Y113_D_CY;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X11Y113_D_XOR;
  wire [0:0] CLBLM_R_X101Y116_SLICE_X158Y116_A;
  wire [0:0] CLBLM_R_X101Y116_SLICE_X158Y116_A1;
  wire [0:0] CLBLM_R_X101Y116_SLICE_X158Y116_A2;
  wire [0:0] CLBLM_R_X101Y116_SLICE_X158Y116_A3;
  wire [0:0] CLBLM_R_X101Y116_SLICE_X158Y116_A4;
  wire [0:0] CLBLM_R_X101Y116_SLICE_X158Y116_A5;
  wire [0:0] CLBLM_R_X101Y116_SLICE_X158Y116_A6;
  wire [0:0] CLBLM_R_X101Y116_SLICE_X158Y116_AO5;
  wire [0:0] CLBLM_R_X101Y116_SLICE_X158Y116_AO6;
  wire [0:0] CLBLM_R_X101Y116_SLICE_X158Y116_A_CY;
  wire [0:0] CLBLM_R_X101Y116_SLICE_X158Y116_A_XOR;
  wire [0:0] CLBLM_R_X101Y116_SLICE_X158Y116_B;
  wire [0:0] CLBLM_R_X101Y116_SLICE_X158Y116_B1;
  wire [0:0] CLBLM_R_X101Y116_SLICE_X158Y116_B2;
  wire [0:0] CLBLM_R_X101Y116_SLICE_X158Y116_B3;
  wire [0:0] CLBLM_R_X101Y116_SLICE_X158Y116_B4;
  wire [0:0] CLBLM_R_X101Y116_SLICE_X158Y116_B5;
  wire [0:0] CLBLM_R_X101Y116_SLICE_X158Y116_B6;
  wire [0:0] CLBLM_R_X101Y116_SLICE_X158Y116_BO5;
  wire [0:0] CLBLM_R_X101Y116_SLICE_X158Y116_BO6;
  wire [0:0] CLBLM_R_X101Y116_SLICE_X158Y116_B_CY;
  wire [0:0] CLBLM_R_X101Y116_SLICE_X158Y116_B_XOR;
  wire [0:0] CLBLM_R_X101Y116_SLICE_X158Y116_C;
  wire [0:0] CLBLM_R_X101Y116_SLICE_X158Y116_C1;
  wire [0:0] CLBLM_R_X101Y116_SLICE_X158Y116_C2;
  wire [0:0] CLBLM_R_X101Y116_SLICE_X158Y116_C3;
  wire [0:0] CLBLM_R_X101Y116_SLICE_X158Y116_C4;
  wire [0:0] CLBLM_R_X101Y116_SLICE_X158Y116_C5;
  wire [0:0] CLBLM_R_X101Y116_SLICE_X158Y116_C6;
  wire [0:0] CLBLM_R_X101Y116_SLICE_X158Y116_CO5;
  wire [0:0] CLBLM_R_X101Y116_SLICE_X158Y116_CO6;
  wire [0:0] CLBLM_R_X101Y116_SLICE_X158Y116_C_CY;
  wire [0:0] CLBLM_R_X101Y116_SLICE_X158Y116_C_XOR;
  wire [0:0] CLBLM_R_X101Y116_SLICE_X158Y116_D;
  wire [0:0] CLBLM_R_X101Y116_SLICE_X158Y116_D1;
  wire [0:0] CLBLM_R_X101Y116_SLICE_X158Y116_D2;
  wire [0:0] CLBLM_R_X101Y116_SLICE_X158Y116_D3;
  wire [0:0] CLBLM_R_X101Y116_SLICE_X158Y116_D4;
  wire [0:0] CLBLM_R_X101Y116_SLICE_X158Y116_D5;
  wire [0:0] CLBLM_R_X101Y116_SLICE_X158Y116_D6;
  wire [0:0] CLBLM_R_X101Y116_SLICE_X158Y116_DO5;
  wire [0:0] CLBLM_R_X101Y116_SLICE_X158Y116_DO6;
  wire [0:0] CLBLM_R_X101Y116_SLICE_X158Y116_D_CY;
  wire [0:0] CLBLM_R_X101Y116_SLICE_X158Y116_D_XOR;
  wire [0:0] CLBLM_R_X101Y116_SLICE_X159Y116_A;
  wire [0:0] CLBLM_R_X101Y116_SLICE_X159Y116_A1;
  wire [0:0] CLBLM_R_X101Y116_SLICE_X159Y116_A2;
  wire [0:0] CLBLM_R_X101Y116_SLICE_X159Y116_A3;
  wire [0:0] CLBLM_R_X101Y116_SLICE_X159Y116_A4;
  wire [0:0] CLBLM_R_X101Y116_SLICE_X159Y116_A5;
  wire [0:0] CLBLM_R_X101Y116_SLICE_X159Y116_A6;
  wire [0:0] CLBLM_R_X101Y116_SLICE_X159Y116_AO5;
  wire [0:0] CLBLM_R_X101Y116_SLICE_X159Y116_AO6;
  wire [0:0] CLBLM_R_X101Y116_SLICE_X159Y116_A_CY;
  wire [0:0] CLBLM_R_X101Y116_SLICE_X159Y116_A_XOR;
  wire [0:0] CLBLM_R_X101Y116_SLICE_X159Y116_B;
  wire [0:0] CLBLM_R_X101Y116_SLICE_X159Y116_B1;
  wire [0:0] CLBLM_R_X101Y116_SLICE_X159Y116_B2;
  wire [0:0] CLBLM_R_X101Y116_SLICE_X159Y116_B3;
  wire [0:0] CLBLM_R_X101Y116_SLICE_X159Y116_B4;
  wire [0:0] CLBLM_R_X101Y116_SLICE_X159Y116_B5;
  wire [0:0] CLBLM_R_X101Y116_SLICE_X159Y116_B6;
  wire [0:0] CLBLM_R_X101Y116_SLICE_X159Y116_BO5;
  wire [0:0] CLBLM_R_X101Y116_SLICE_X159Y116_BO6;
  wire [0:0] CLBLM_R_X101Y116_SLICE_X159Y116_B_CY;
  wire [0:0] CLBLM_R_X101Y116_SLICE_X159Y116_B_XOR;
  wire [0:0] CLBLM_R_X101Y116_SLICE_X159Y116_C;
  wire [0:0] CLBLM_R_X101Y116_SLICE_X159Y116_C1;
  wire [0:0] CLBLM_R_X101Y116_SLICE_X159Y116_C2;
  wire [0:0] CLBLM_R_X101Y116_SLICE_X159Y116_C3;
  wire [0:0] CLBLM_R_X101Y116_SLICE_X159Y116_C4;
  wire [0:0] CLBLM_R_X101Y116_SLICE_X159Y116_C5;
  wire [0:0] CLBLM_R_X101Y116_SLICE_X159Y116_C6;
  wire [0:0] CLBLM_R_X101Y116_SLICE_X159Y116_CO5;
  wire [0:0] CLBLM_R_X101Y116_SLICE_X159Y116_CO6;
  wire [0:0] CLBLM_R_X101Y116_SLICE_X159Y116_C_CY;
  wire [0:0] CLBLM_R_X101Y116_SLICE_X159Y116_C_XOR;
  wire [0:0] CLBLM_R_X101Y116_SLICE_X159Y116_D;
  wire [0:0] CLBLM_R_X101Y116_SLICE_X159Y116_D1;
  wire [0:0] CLBLM_R_X101Y116_SLICE_X159Y116_D2;
  wire [0:0] CLBLM_R_X101Y116_SLICE_X159Y116_D3;
  wire [0:0] CLBLM_R_X101Y116_SLICE_X159Y116_D4;
  wire [0:0] CLBLM_R_X101Y116_SLICE_X159Y116_D5;
  wire [0:0] CLBLM_R_X101Y116_SLICE_X159Y116_D6;
  wire [0:0] CLBLM_R_X101Y116_SLICE_X159Y116_DO5;
  wire [0:0] CLBLM_R_X101Y116_SLICE_X159Y116_DO6;
  wire [0:0] CLBLM_R_X101Y116_SLICE_X159Y116_D_CY;
  wire [0:0] CLBLM_R_X101Y116_SLICE_X159Y116_D_XOR;
  wire [0:0] CLBLM_R_X101Y117_SLICE_X158Y117_A;
  wire [0:0] CLBLM_R_X101Y117_SLICE_X158Y117_A1;
  wire [0:0] CLBLM_R_X101Y117_SLICE_X158Y117_A2;
  wire [0:0] CLBLM_R_X101Y117_SLICE_X158Y117_A3;
  wire [0:0] CLBLM_R_X101Y117_SLICE_X158Y117_A4;
  wire [0:0] CLBLM_R_X101Y117_SLICE_X158Y117_A5;
  wire [0:0] CLBLM_R_X101Y117_SLICE_X158Y117_A6;
  wire [0:0] CLBLM_R_X101Y117_SLICE_X158Y117_AO5;
  wire [0:0] CLBLM_R_X101Y117_SLICE_X158Y117_AO6;
  wire [0:0] CLBLM_R_X101Y117_SLICE_X158Y117_A_CY;
  wire [0:0] CLBLM_R_X101Y117_SLICE_X158Y117_A_XOR;
  wire [0:0] CLBLM_R_X101Y117_SLICE_X158Y117_B;
  wire [0:0] CLBLM_R_X101Y117_SLICE_X158Y117_B1;
  wire [0:0] CLBLM_R_X101Y117_SLICE_X158Y117_B2;
  wire [0:0] CLBLM_R_X101Y117_SLICE_X158Y117_B3;
  wire [0:0] CLBLM_R_X101Y117_SLICE_X158Y117_B4;
  wire [0:0] CLBLM_R_X101Y117_SLICE_X158Y117_B5;
  wire [0:0] CLBLM_R_X101Y117_SLICE_X158Y117_B6;
  wire [0:0] CLBLM_R_X101Y117_SLICE_X158Y117_BO5;
  wire [0:0] CLBLM_R_X101Y117_SLICE_X158Y117_BO6;
  wire [0:0] CLBLM_R_X101Y117_SLICE_X158Y117_B_CY;
  wire [0:0] CLBLM_R_X101Y117_SLICE_X158Y117_B_XOR;
  wire [0:0] CLBLM_R_X101Y117_SLICE_X158Y117_C;
  wire [0:0] CLBLM_R_X101Y117_SLICE_X158Y117_C1;
  wire [0:0] CLBLM_R_X101Y117_SLICE_X158Y117_C2;
  wire [0:0] CLBLM_R_X101Y117_SLICE_X158Y117_C3;
  wire [0:0] CLBLM_R_X101Y117_SLICE_X158Y117_C4;
  wire [0:0] CLBLM_R_X101Y117_SLICE_X158Y117_C5;
  wire [0:0] CLBLM_R_X101Y117_SLICE_X158Y117_C6;
  wire [0:0] CLBLM_R_X101Y117_SLICE_X158Y117_CO5;
  wire [0:0] CLBLM_R_X101Y117_SLICE_X158Y117_CO6;
  wire [0:0] CLBLM_R_X101Y117_SLICE_X158Y117_C_CY;
  wire [0:0] CLBLM_R_X101Y117_SLICE_X158Y117_C_XOR;
  wire [0:0] CLBLM_R_X101Y117_SLICE_X158Y117_D;
  wire [0:0] CLBLM_R_X101Y117_SLICE_X158Y117_D1;
  wire [0:0] CLBLM_R_X101Y117_SLICE_X158Y117_D2;
  wire [0:0] CLBLM_R_X101Y117_SLICE_X158Y117_D3;
  wire [0:0] CLBLM_R_X101Y117_SLICE_X158Y117_D4;
  wire [0:0] CLBLM_R_X101Y117_SLICE_X158Y117_D5;
  wire [0:0] CLBLM_R_X101Y117_SLICE_X158Y117_D6;
  wire [0:0] CLBLM_R_X101Y117_SLICE_X158Y117_DO5;
  wire [0:0] CLBLM_R_X101Y117_SLICE_X158Y117_DO6;
  wire [0:0] CLBLM_R_X101Y117_SLICE_X158Y117_D_CY;
  wire [0:0] CLBLM_R_X101Y117_SLICE_X158Y117_D_XOR;
  wire [0:0] CLBLM_R_X101Y117_SLICE_X159Y117_A;
  wire [0:0] CLBLM_R_X101Y117_SLICE_X159Y117_A1;
  wire [0:0] CLBLM_R_X101Y117_SLICE_X159Y117_A2;
  wire [0:0] CLBLM_R_X101Y117_SLICE_X159Y117_A3;
  wire [0:0] CLBLM_R_X101Y117_SLICE_X159Y117_A4;
  wire [0:0] CLBLM_R_X101Y117_SLICE_X159Y117_A5;
  wire [0:0] CLBLM_R_X101Y117_SLICE_X159Y117_A6;
  wire [0:0] CLBLM_R_X101Y117_SLICE_X159Y117_AO5;
  wire [0:0] CLBLM_R_X101Y117_SLICE_X159Y117_AO6;
  wire [0:0] CLBLM_R_X101Y117_SLICE_X159Y117_A_CY;
  wire [0:0] CLBLM_R_X101Y117_SLICE_X159Y117_A_XOR;
  wire [0:0] CLBLM_R_X101Y117_SLICE_X159Y117_B;
  wire [0:0] CLBLM_R_X101Y117_SLICE_X159Y117_B1;
  wire [0:0] CLBLM_R_X101Y117_SLICE_X159Y117_B2;
  wire [0:0] CLBLM_R_X101Y117_SLICE_X159Y117_B3;
  wire [0:0] CLBLM_R_X101Y117_SLICE_X159Y117_B4;
  wire [0:0] CLBLM_R_X101Y117_SLICE_X159Y117_B5;
  wire [0:0] CLBLM_R_X101Y117_SLICE_X159Y117_B6;
  wire [0:0] CLBLM_R_X101Y117_SLICE_X159Y117_BO5;
  wire [0:0] CLBLM_R_X101Y117_SLICE_X159Y117_BO6;
  wire [0:0] CLBLM_R_X101Y117_SLICE_X159Y117_B_CY;
  wire [0:0] CLBLM_R_X101Y117_SLICE_X159Y117_B_XOR;
  wire [0:0] CLBLM_R_X101Y117_SLICE_X159Y117_C;
  wire [0:0] CLBLM_R_X101Y117_SLICE_X159Y117_C1;
  wire [0:0] CLBLM_R_X101Y117_SLICE_X159Y117_C2;
  wire [0:0] CLBLM_R_X101Y117_SLICE_X159Y117_C3;
  wire [0:0] CLBLM_R_X101Y117_SLICE_X159Y117_C4;
  wire [0:0] CLBLM_R_X101Y117_SLICE_X159Y117_C5;
  wire [0:0] CLBLM_R_X101Y117_SLICE_X159Y117_C6;
  wire [0:0] CLBLM_R_X101Y117_SLICE_X159Y117_CO5;
  wire [0:0] CLBLM_R_X101Y117_SLICE_X159Y117_CO6;
  wire [0:0] CLBLM_R_X101Y117_SLICE_X159Y117_C_CY;
  wire [0:0] CLBLM_R_X101Y117_SLICE_X159Y117_C_XOR;
  wire [0:0] CLBLM_R_X101Y117_SLICE_X159Y117_D;
  wire [0:0] CLBLM_R_X101Y117_SLICE_X159Y117_D1;
  wire [0:0] CLBLM_R_X101Y117_SLICE_X159Y117_D2;
  wire [0:0] CLBLM_R_X101Y117_SLICE_X159Y117_D3;
  wire [0:0] CLBLM_R_X101Y117_SLICE_X159Y117_D4;
  wire [0:0] CLBLM_R_X101Y117_SLICE_X159Y117_D5;
  wire [0:0] CLBLM_R_X101Y117_SLICE_X159Y117_D6;
  wire [0:0] CLBLM_R_X101Y117_SLICE_X159Y117_DO5;
  wire [0:0] CLBLM_R_X101Y117_SLICE_X159Y117_DO6;
  wire [0:0] CLBLM_R_X101Y117_SLICE_X159Y117_D_CY;
  wire [0:0] CLBLM_R_X101Y117_SLICE_X159Y117_D_XOR;
  wire [0:0] CLBLM_R_X101Y118_SLICE_X158Y118_A;
  wire [0:0] CLBLM_R_X101Y118_SLICE_X158Y118_A1;
  wire [0:0] CLBLM_R_X101Y118_SLICE_X158Y118_A2;
  wire [0:0] CLBLM_R_X101Y118_SLICE_X158Y118_A3;
  wire [0:0] CLBLM_R_X101Y118_SLICE_X158Y118_A4;
  wire [0:0] CLBLM_R_X101Y118_SLICE_X158Y118_A5;
  wire [0:0] CLBLM_R_X101Y118_SLICE_X158Y118_A6;
  wire [0:0] CLBLM_R_X101Y118_SLICE_X158Y118_AO5;
  wire [0:0] CLBLM_R_X101Y118_SLICE_X158Y118_AO6;
  wire [0:0] CLBLM_R_X101Y118_SLICE_X158Y118_A_CY;
  wire [0:0] CLBLM_R_X101Y118_SLICE_X158Y118_A_XOR;
  wire [0:0] CLBLM_R_X101Y118_SLICE_X158Y118_B;
  wire [0:0] CLBLM_R_X101Y118_SLICE_X158Y118_B1;
  wire [0:0] CLBLM_R_X101Y118_SLICE_X158Y118_B2;
  wire [0:0] CLBLM_R_X101Y118_SLICE_X158Y118_B3;
  wire [0:0] CLBLM_R_X101Y118_SLICE_X158Y118_B4;
  wire [0:0] CLBLM_R_X101Y118_SLICE_X158Y118_B5;
  wire [0:0] CLBLM_R_X101Y118_SLICE_X158Y118_B6;
  wire [0:0] CLBLM_R_X101Y118_SLICE_X158Y118_BO5;
  wire [0:0] CLBLM_R_X101Y118_SLICE_X158Y118_BO6;
  wire [0:0] CLBLM_R_X101Y118_SLICE_X158Y118_B_CY;
  wire [0:0] CLBLM_R_X101Y118_SLICE_X158Y118_B_XOR;
  wire [0:0] CLBLM_R_X101Y118_SLICE_X158Y118_C;
  wire [0:0] CLBLM_R_X101Y118_SLICE_X158Y118_C1;
  wire [0:0] CLBLM_R_X101Y118_SLICE_X158Y118_C2;
  wire [0:0] CLBLM_R_X101Y118_SLICE_X158Y118_C3;
  wire [0:0] CLBLM_R_X101Y118_SLICE_X158Y118_C4;
  wire [0:0] CLBLM_R_X101Y118_SLICE_X158Y118_C5;
  wire [0:0] CLBLM_R_X101Y118_SLICE_X158Y118_C6;
  wire [0:0] CLBLM_R_X101Y118_SLICE_X158Y118_CO5;
  wire [0:0] CLBLM_R_X101Y118_SLICE_X158Y118_CO6;
  wire [0:0] CLBLM_R_X101Y118_SLICE_X158Y118_C_CY;
  wire [0:0] CLBLM_R_X101Y118_SLICE_X158Y118_C_XOR;
  wire [0:0] CLBLM_R_X101Y118_SLICE_X158Y118_D;
  wire [0:0] CLBLM_R_X101Y118_SLICE_X158Y118_D1;
  wire [0:0] CLBLM_R_X101Y118_SLICE_X158Y118_D2;
  wire [0:0] CLBLM_R_X101Y118_SLICE_X158Y118_D3;
  wire [0:0] CLBLM_R_X101Y118_SLICE_X158Y118_D4;
  wire [0:0] CLBLM_R_X101Y118_SLICE_X158Y118_D5;
  wire [0:0] CLBLM_R_X101Y118_SLICE_X158Y118_D6;
  wire [0:0] CLBLM_R_X101Y118_SLICE_X158Y118_DO5;
  wire [0:0] CLBLM_R_X101Y118_SLICE_X158Y118_DO6;
  wire [0:0] CLBLM_R_X101Y118_SLICE_X158Y118_D_CY;
  wire [0:0] CLBLM_R_X101Y118_SLICE_X158Y118_D_XOR;
  wire [0:0] CLBLM_R_X101Y118_SLICE_X159Y118_A;
  wire [0:0] CLBLM_R_X101Y118_SLICE_X159Y118_A1;
  wire [0:0] CLBLM_R_X101Y118_SLICE_X159Y118_A2;
  wire [0:0] CLBLM_R_X101Y118_SLICE_X159Y118_A3;
  wire [0:0] CLBLM_R_X101Y118_SLICE_X159Y118_A4;
  wire [0:0] CLBLM_R_X101Y118_SLICE_X159Y118_A5;
  wire [0:0] CLBLM_R_X101Y118_SLICE_X159Y118_A6;
  wire [0:0] CLBLM_R_X101Y118_SLICE_X159Y118_AO5;
  wire [0:0] CLBLM_R_X101Y118_SLICE_X159Y118_AO6;
  wire [0:0] CLBLM_R_X101Y118_SLICE_X159Y118_A_CY;
  wire [0:0] CLBLM_R_X101Y118_SLICE_X159Y118_A_XOR;
  wire [0:0] CLBLM_R_X101Y118_SLICE_X159Y118_B;
  wire [0:0] CLBLM_R_X101Y118_SLICE_X159Y118_B1;
  wire [0:0] CLBLM_R_X101Y118_SLICE_X159Y118_B2;
  wire [0:0] CLBLM_R_X101Y118_SLICE_X159Y118_B3;
  wire [0:0] CLBLM_R_X101Y118_SLICE_X159Y118_B4;
  wire [0:0] CLBLM_R_X101Y118_SLICE_X159Y118_B5;
  wire [0:0] CLBLM_R_X101Y118_SLICE_X159Y118_B6;
  wire [0:0] CLBLM_R_X101Y118_SLICE_X159Y118_BO5;
  wire [0:0] CLBLM_R_X101Y118_SLICE_X159Y118_BO6;
  wire [0:0] CLBLM_R_X101Y118_SLICE_X159Y118_B_CY;
  wire [0:0] CLBLM_R_X101Y118_SLICE_X159Y118_B_XOR;
  wire [0:0] CLBLM_R_X101Y118_SLICE_X159Y118_C;
  wire [0:0] CLBLM_R_X101Y118_SLICE_X159Y118_C1;
  wire [0:0] CLBLM_R_X101Y118_SLICE_X159Y118_C2;
  wire [0:0] CLBLM_R_X101Y118_SLICE_X159Y118_C3;
  wire [0:0] CLBLM_R_X101Y118_SLICE_X159Y118_C4;
  wire [0:0] CLBLM_R_X101Y118_SLICE_X159Y118_C5;
  wire [0:0] CLBLM_R_X101Y118_SLICE_X159Y118_C6;
  wire [0:0] CLBLM_R_X101Y118_SLICE_X159Y118_CO5;
  wire [0:0] CLBLM_R_X101Y118_SLICE_X159Y118_CO6;
  wire [0:0] CLBLM_R_X101Y118_SLICE_X159Y118_C_CY;
  wire [0:0] CLBLM_R_X101Y118_SLICE_X159Y118_C_XOR;
  wire [0:0] CLBLM_R_X101Y118_SLICE_X159Y118_D;
  wire [0:0] CLBLM_R_X101Y118_SLICE_X159Y118_D1;
  wire [0:0] CLBLM_R_X101Y118_SLICE_X159Y118_D2;
  wire [0:0] CLBLM_R_X101Y118_SLICE_X159Y118_D3;
  wire [0:0] CLBLM_R_X101Y118_SLICE_X159Y118_D4;
  wire [0:0] CLBLM_R_X101Y118_SLICE_X159Y118_D5;
  wire [0:0] CLBLM_R_X101Y118_SLICE_X159Y118_D6;
  wire [0:0] CLBLM_R_X101Y118_SLICE_X159Y118_DO5;
  wire [0:0] CLBLM_R_X101Y118_SLICE_X159Y118_DO6;
  wire [0:0] CLBLM_R_X101Y118_SLICE_X159Y118_D_CY;
  wire [0:0] CLBLM_R_X101Y118_SLICE_X159Y118_D_XOR;
  wire [0:0] CLBLM_R_X101Y119_SLICE_X158Y119_A;
  wire [0:0] CLBLM_R_X101Y119_SLICE_X158Y119_A1;
  wire [0:0] CLBLM_R_X101Y119_SLICE_X158Y119_A2;
  wire [0:0] CLBLM_R_X101Y119_SLICE_X158Y119_A3;
  wire [0:0] CLBLM_R_X101Y119_SLICE_X158Y119_A4;
  wire [0:0] CLBLM_R_X101Y119_SLICE_X158Y119_A5;
  wire [0:0] CLBLM_R_X101Y119_SLICE_X158Y119_A6;
  wire [0:0] CLBLM_R_X101Y119_SLICE_X158Y119_AO5;
  wire [0:0] CLBLM_R_X101Y119_SLICE_X158Y119_AO6;
  wire [0:0] CLBLM_R_X101Y119_SLICE_X158Y119_A_CY;
  wire [0:0] CLBLM_R_X101Y119_SLICE_X158Y119_A_XOR;
  wire [0:0] CLBLM_R_X101Y119_SLICE_X158Y119_B;
  wire [0:0] CLBLM_R_X101Y119_SLICE_X158Y119_B1;
  wire [0:0] CLBLM_R_X101Y119_SLICE_X158Y119_B2;
  wire [0:0] CLBLM_R_X101Y119_SLICE_X158Y119_B3;
  wire [0:0] CLBLM_R_X101Y119_SLICE_X158Y119_B4;
  wire [0:0] CLBLM_R_X101Y119_SLICE_X158Y119_B5;
  wire [0:0] CLBLM_R_X101Y119_SLICE_X158Y119_B6;
  wire [0:0] CLBLM_R_X101Y119_SLICE_X158Y119_BO5;
  wire [0:0] CLBLM_R_X101Y119_SLICE_X158Y119_BO6;
  wire [0:0] CLBLM_R_X101Y119_SLICE_X158Y119_B_CY;
  wire [0:0] CLBLM_R_X101Y119_SLICE_X158Y119_B_XOR;
  wire [0:0] CLBLM_R_X101Y119_SLICE_X158Y119_C;
  wire [0:0] CLBLM_R_X101Y119_SLICE_X158Y119_C1;
  wire [0:0] CLBLM_R_X101Y119_SLICE_X158Y119_C2;
  wire [0:0] CLBLM_R_X101Y119_SLICE_X158Y119_C3;
  wire [0:0] CLBLM_R_X101Y119_SLICE_X158Y119_C4;
  wire [0:0] CLBLM_R_X101Y119_SLICE_X158Y119_C5;
  wire [0:0] CLBLM_R_X101Y119_SLICE_X158Y119_C6;
  wire [0:0] CLBLM_R_X101Y119_SLICE_X158Y119_CO5;
  wire [0:0] CLBLM_R_X101Y119_SLICE_X158Y119_CO6;
  wire [0:0] CLBLM_R_X101Y119_SLICE_X158Y119_C_CY;
  wire [0:0] CLBLM_R_X101Y119_SLICE_X158Y119_C_XOR;
  wire [0:0] CLBLM_R_X101Y119_SLICE_X158Y119_D;
  wire [0:0] CLBLM_R_X101Y119_SLICE_X158Y119_D1;
  wire [0:0] CLBLM_R_X101Y119_SLICE_X158Y119_D2;
  wire [0:0] CLBLM_R_X101Y119_SLICE_X158Y119_D3;
  wire [0:0] CLBLM_R_X101Y119_SLICE_X158Y119_D4;
  wire [0:0] CLBLM_R_X101Y119_SLICE_X158Y119_D5;
  wire [0:0] CLBLM_R_X101Y119_SLICE_X158Y119_D6;
  wire [0:0] CLBLM_R_X101Y119_SLICE_X158Y119_DO5;
  wire [0:0] CLBLM_R_X101Y119_SLICE_X158Y119_DO6;
  wire [0:0] CLBLM_R_X101Y119_SLICE_X158Y119_D_CY;
  wire [0:0] CLBLM_R_X101Y119_SLICE_X158Y119_D_XOR;
  wire [0:0] CLBLM_R_X101Y119_SLICE_X159Y119_A;
  wire [0:0] CLBLM_R_X101Y119_SLICE_X159Y119_A1;
  wire [0:0] CLBLM_R_X101Y119_SLICE_X159Y119_A2;
  wire [0:0] CLBLM_R_X101Y119_SLICE_X159Y119_A3;
  wire [0:0] CLBLM_R_X101Y119_SLICE_X159Y119_A4;
  wire [0:0] CLBLM_R_X101Y119_SLICE_X159Y119_A5;
  wire [0:0] CLBLM_R_X101Y119_SLICE_X159Y119_A6;
  wire [0:0] CLBLM_R_X101Y119_SLICE_X159Y119_AO5;
  wire [0:0] CLBLM_R_X101Y119_SLICE_X159Y119_AO6;
  wire [0:0] CLBLM_R_X101Y119_SLICE_X159Y119_A_CY;
  wire [0:0] CLBLM_R_X101Y119_SLICE_X159Y119_A_XOR;
  wire [0:0] CLBLM_R_X101Y119_SLICE_X159Y119_B;
  wire [0:0] CLBLM_R_X101Y119_SLICE_X159Y119_B1;
  wire [0:0] CLBLM_R_X101Y119_SLICE_X159Y119_B2;
  wire [0:0] CLBLM_R_X101Y119_SLICE_X159Y119_B3;
  wire [0:0] CLBLM_R_X101Y119_SLICE_X159Y119_B4;
  wire [0:0] CLBLM_R_X101Y119_SLICE_X159Y119_B5;
  wire [0:0] CLBLM_R_X101Y119_SLICE_X159Y119_B6;
  wire [0:0] CLBLM_R_X101Y119_SLICE_X159Y119_BO5;
  wire [0:0] CLBLM_R_X101Y119_SLICE_X159Y119_BO6;
  wire [0:0] CLBLM_R_X101Y119_SLICE_X159Y119_B_CY;
  wire [0:0] CLBLM_R_X101Y119_SLICE_X159Y119_B_XOR;
  wire [0:0] CLBLM_R_X101Y119_SLICE_X159Y119_C;
  wire [0:0] CLBLM_R_X101Y119_SLICE_X159Y119_C1;
  wire [0:0] CLBLM_R_X101Y119_SLICE_X159Y119_C2;
  wire [0:0] CLBLM_R_X101Y119_SLICE_X159Y119_C3;
  wire [0:0] CLBLM_R_X101Y119_SLICE_X159Y119_C4;
  wire [0:0] CLBLM_R_X101Y119_SLICE_X159Y119_C5;
  wire [0:0] CLBLM_R_X101Y119_SLICE_X159Y119_C6;
  wire [0:0] CLBLM_R_X101Y119_SLICE_X159Y119_CO5;
  wire [0:0] CLBLM_R_X101Y119_SLICE_X159Y119_CO6;
  wire [0:0] CLBLM_R_X101Y119_SLICE_X159Y119_C_CY;
  wire [0:0] CLBLM_R_X101Y119_SLICE_X159Y119_C_XOR;
  wire [0:0] CLBLM_R_X101Y119_SLICE_X159Y119_D;
  wire [0:0] CLBLM_R_X101Y119_SLICE_X159Y119_D1;
  wire [0:0] CLBLM_R_X101Y119_SLICE_X159Y119_D2;
  wire [0:0] CLBLM_R_X101Y119_SLICE_X159Y119_D3;
  wire [0:0] CLBLM_R_X101Y119_SLICE_X159Y119_D4;
  wire [0:0] CLBLM_R_X101Y119_SLICE_X159Y119_D5;
  wire [0:0] CLBLM_R_X101Y119_SLICE_X159Y119_D6;
  wire [0:0] CLBLM_R_X101Y119_SLICE_X159Y119_DO5;
  wire [0:0] CLBLM_R_X101Y119_SLICE_X159Y119_DO6;
  wire [0:0] CLBLM_R_X101Y119_SLICE_X159Y119_D_CY;
  wire [0:0] CLBLM_R_X101Y119_SLICE_X159Y119_D_XOR;
  wire [0:0] CLBLM_R_X101Y123_SLICE_X158Y123_A;
  wire [0:0] CLBLM_R_X101Y123_SLICE_X158Y123_A1;
  wire [0:0] CLBLM_R_X101Y123_SLICE_X158Y123_A2;
  wire [0:0] CLBLM_R_X101Y123_SLICE_X158Y123_A3;
  wire [0:0] CLBLM_R_X101Y123_SLICE_X158Y123_A4;
  wire [0:0] CLBLM_R_X101Y123_SLICE_X158Y123_A5;
  wire [0:0] CLBLM_R_X101Y123_SLICE_X158Y123_A6;
  wire [0:0] CLBLM_R_X101Y123_SLICE_X158Y123_AMUX;
  wire [0:0] CLBLM_R_X101Y123_SLICE_X158Y123_AO5;
  wire [0:0] CLBLM_R_X101Y123_SLICE_X158Y123_AO6;
  wire [0:0] CLBLM_R_X101Y123_SLICE_X158Y123_A_CY;
  wire [0:0] CLBLM_R_X101Y123_SLICE_X158Y123_A_XOR;
  wire [0:0] CLBLM_R_X101Y123_SLICE_X158Y123_B;
  wire [0:0] CLBLM_R_X101Y123_SLICE_X158Y123_B1;
  wire [0:0] CLBLM_R_X101Y123_SLICE_X158Y123_B2;
  wire [0:0] CLBLM_R_X101Y123_SLICE_X158Y123_B3;
  wire [0:0] CLBLM_R_X101Y123_SLICE_X158Y123_B4;
  wire [0:0] CLBLM_R_X101Y123_SLICE_X158Y123_B5;
  wire [0:0] CLBLM_R_X101Y123_SLICE_X158Y123_B6;
  wire [0:0] CLBLM_R_X101Y123_SLICE_X158Y123_BO5;
  wire [0:0] CLBLM_R_X101Y123_SLICE_X158Y123_BO6;
  wire [0:0] CLBLM_R_X101Y123_SLICE_X158Y123_B_CY;
  wire [0:0] CLBLM_R_X101Y123_SLICE_X158Y123_B_XOR;
  wire [0:0] CLBLM_R_X101Y123_SLICE_X158Y123_C;
  wire [0:0] CLBLM_R_X101Y123_SLICE_X158Y123_C1;
  wire [0:0] CLBLM_R_X101Y123_SLICE_X158Y123_C2;
  wire [0:0] CLBLM_R_X101Y123_SLICE_X158Y123_C3;
  wire [0:0] CLBLM_R_X101Y123_SLICE_X158Y123_C4;
  wire [0:0] CLBLM_R_X101Y123_SLICE_X158Y123_C5;
  wire [0:0] CLBLM_R_X101Y123_SLICE_X158Y123_C6;
  wire [0:0] CLBLM_R_X101Y123_SLICE_X158Y123_CO5;
  wire [0:0] CLBLM_R_X101Y123_SLICE_X158Y123_CO6;
  wire [0:0] CLBLM_R_X101Y123_SLICE_X158Y123_C_CY;
  wire [0:0] CLBLM_R_X101Y123_SLICE_X158Y123_C_XOR;
  wire [0:0] CLBLM_R_X101Y123_SLICE_X158Y123_D;
  wire [0:0] CLBLM_R_X101Y123_SLICE_X158Y123_D1;
  wire [0:0] CLBLM_R_X101Y123_SLICE_X158Y123_D2;
  wire [0:0] CLBLM_R_X101Y123_SLICE_X158Y123_D3;
  wire [0:0] CLBLM_R_X101Y123_SLICE_X158Y123_D4;
  wire [0:0] CLBLM_R_X101Y123_SLICE_X158Y123_D5;
  wire [0:0] CLBLM_R_X101Y123_SLICE_X158Y123_D6;
  wire [0:0] CLBLM_R_X101Y123_SLICE_X158Y123_DO5;
  wire [0:0] CLBLM_R_X101Y123_SLICE_X158Y123_DO6;
  wire [0:0] CLBLM_R_X101Y123_SLICE_X158Y123_D_CY;
  wire [0:0] CLBLM_R_X101Y123_SLICE_X158Y123_D_XOR;
  wire [0:0] CLBLM_R_X101Y123_SLICE_X159Y123_A;
  wire [0:0] CLBLM_R_X101Y123_SLICE_X159Y123_A1;
  wire [0:0] CLBLM_R_X101Y123_SLICE_X159Y123_A2;
  wire [0:0] CLBLM_R_X101Y123_SLICE_X159Y123_A3;
  wire [0:0] CLBLM_R_X101Y123_SLICE_X159Y123_A4;
  wire [0:0] CLBLM_R_X101Y123_SLICE_X159Y123_A5;
  wire [0:0] CLBLM_R_X101Y123_SLICE_X159Y123_A6;
  wire [0:0] CLBLM_R_X101Y123_SLICE_X159Y123_AO5;
  wire [0:0] CLBLM_R_X101Y123_SLICE_X159Y123_AO6;
  wire [0:0] CLBLM_R_X101Y123_SLICE_X159Y123_A_CY;
  wire [0:0] CLBLM_R_X101Y123_SLICE_X159Y123_A_XOR;
  wire [0:0] CLBLM_R_X101Y123_SLICE_X159Y123_B;
  wire [0:0] CLBLM_R_X101Y123_SLICE_X159Y123_B1;
  wire [0:0] CLBLM_R_X101Y123_SLICE_X159Y123_B2;
  wire [0:0] CLBLM_R_X101Y123_SLICE_X159Y123_B3;
  wire [0:0] CLBLM_R_X101Y123_SLICE_X159Y123_B4;
  wire [0:0] CLBLM_R_X101Y123_SLICE_X159Y123_B5;
  wire [0:0] CLBLM_R_X101Y123_SLICE_X159Y123_B6;
  wire [0:0] CLBLM_R_X101Y123_SLICE_X159Y123_BO5;
  wire [0:0] CLBLM_R_X101Y123_SLICE_X159Y123_BO6;
  wire [0:0] CLBLM_R_X101Y123_SLICE_X159Y123_B_CY;
  wire [0:0] CLBLM_R_X101Y123_SLICE_X159Y123_B_XOR;
  wire [0:0] CLBLM_R_X101Y123_SLICE_X159Y123_C;
  wire [0:0] CLBLM_R_X101Y123_SLICE_X159Y123_C1;
  wire [0:0] CLBLM_R_X101Y123_SLICE_X159Y123_C2;
  wire [0:0] CLBLM_R_X101Y123_SLICE_X159Y123_C3;
  wire [0:0] CLBLM_R_X101Y123_SLICE_X159Y123_C4;
  wire [0:0] CLBLM_R_X101Y123_SLICE_X159Y123_C5;
  wire [0:0] CLBLM_R_X101Y123_SLICE_X159Y123_C6;
  wire [0:0] CLBLM_R_X101Y123_SLICE_X159Y123_CO5;
  wire [0:0] CLBLM_R_X101Y123_SLICE_X159Y123_CO6;
  wire [0:0] CLBLM_R_X101Y123_SLICE_X159Y123_C_CY;
  wire [0:0] CLBLM_R_X101Y123_SLICE_X159Y123_C_XOR;
  wire [0:0] CLBLM_R_X101Y123_SLICE_X159Y123_D;
  wire [0:0] CLBLM_R_X101Y123_SLICE_X159Y123_D1;
  wire [0:0] CLBLM_R_X101Y123_SLICE_X159Y123_D2;
  wire [0:0] CLBLM_R_X101Y123_SLICE_X159Y123_D3;
  wire [0:0] CLBLM_R_X101Y123_SLICE_X159Y123_D4;
  wire [0:0] CLBLM_R_X101Y123_SLICE_X159Y123_D5;
  wire [0:0] CLBLM_R_X101Y123_SLICE_X159Y123_D6;
  wire [0:0] CLBLM_R_X101Y123_SLICE_X159Y123_DO5;
  wire [0:0] CLBLM_R_X101Y123_SLICE_X159Y123_DO6;
  wire [0:0] CLBLM_R_X101Y123_SLICE_X159Y123_D_CY;
  wire [0:0] CLBLM_R_X101Y123_SLICE_X159Y123_D_XOR;
  wire [0:0] CLBLM_R_X103Y102_SLICE_X162Y102_A;
  wire [0:0] CLBLM_R_X103Y102_SLICE_X162Y102_A1;
  wire [0:0] CLBLM_R_X103Y102_SLICE_X162Y102_A2;
  wire [0:0] CLBLM_R_X103Y102_SLICE_X162Y102_A3;
  wire [0:0] CLBLM_R_X103Y102_SLICE_X162Y102_A4;
  wire [0:0] CLBLM_R_X103Y102_SLICE_X162Y102_A5;
  wire [0:0] CLBLM_R_X103Y102_SLICE_X162Y102_A6;
  wire [0:0] CLBLM_R_X103Y102_SLICE_X162Y102_AO5;
  wire [0:0] CLBLM_R_X103Y102_SLICE_X162Y102_AO6;
  wire [0:0] CLBLM_R_X103Y102_SLICE_X162Y102_A_CY;
  wire [0:0] CLBLM_R_X103Y102_SLICE_X162Y102_A_XOR;
  wire [0:0] CLBLM_R_X103Y102_SLICE_X162Y102_B;
  wire [0:0] CLBLM_R_X103Y102_SLICE_X162Y102_B1;
  wire [0:0] CLBLM_R_X103Y102_SLICE_X162Y102_B2;
  wire [0:0] CLBLM_R_X103Y102_SLICE_X162Y102_B3;
  wire [0:0] CLBLM_R_X103Y102_SLICE_X162Y102_B4;
  wire [0:0] CLBLM_R_X103Y102_SLICE_X162Y102_B5;
  wire [0:0] CLBLM_R_X103Y102_SLICE_X162Y102_B6;
  wire [0:0] CLBLM_R_X103Y102_SLICE_X162Y102_BO5;
  wire [0:0] CLBLM_R_X103Y102_SLICE_X162Y102_BO6;
  wire [0:0] CLBLM_R_X103Y102_SLICE_X162Y102_B_CY;
  wire [0:0] CLBLM_R_X103Y102_SLICE_X162Y102_B_XOR;
  wire [0:0] CLBLM_R_X103Y102_SLICE_X162Y102_C;
  wire [0:0] CLBLM_R_X103Y102_SLICE_X162Y102_C1;
  wire [0:0] CLBLM_R_X103Y102_SLICE_X162Y102_C2;
  wire [0:0] CLBLM_R_X103Y102_SLICE_X162Y102_C3;
  wire [0:0] CLBLM_R_X103Y102_SLICE_X162Y102_C4;
  wire [0:0] CLBLM_R_X103Y102_SLICE_X162Y102_C5;
  wire [0:0] CLBLM_R_X103Y102_SLICE_X162Y102_C6;
  wire [0:0] CLBLM_R_X103Y102_SLICE_X162Y102_CO5;
  wire [0:0] CLBLM_R_X103Y102_SLICE_X162Y102_CO6;
  wire [0:0] CLBLM_R_X103Y102_SLICE_X162Y102_C_CY;
  wire [0:0] CLBLM_R_X103Y102_SLICE_X162Y102_C_XOR;
  wire [0:0] CLBLM_R_X103Y102_SLICE_X162Y102_D;
  wire [0:0] CLBLM_R_X103Y102_SLICE_X162Y102_D1;
  wire [0:0] CLBLM_R_X103Y102_SLICE_X162Y102_D2;
  wire [0:0] CLBLM_R_X103Y102_SLICE_X162Y102_D3;
  wire [0:0] CLBLM_R_X103Y102_SLICE_X162Y102_D4;
  wire [0:0] CLBLM_R_X103Y102_SLICE_X162Y102_D5;
  wire [0:0] CLBLM_R_X103Y102_SLICE_X162Y102_D6;
  wire [0:0] CLBLM_R_X103Y102_SLICE_X162Y102_DO5;
  wire [0:0] CLBLM_R_X103Y102_SLICE_X162Y102_DO6;
  wire [0:0] CLBLM_R_X103Y102_SLICE_X162Y102_D_CY;
  wire [0:0] CLBLM_R_X103Y102_SLICE_X162Y102_D_XOR;
  wire [0:0] CLBLM_R_X103Y102_SLICE_X163Y102_A;
  wire [0:0] CLBLM_R_X103Y102_SLICE_X163Y102_A1;
  wire [0:0] CLBLM_R_X103Y102_SLICE_X163Y102_A2;
  wire [0:0] CLBLM_R_X103Y102_SLICE_X163Y102_A3;
  wire [0:0] CLBLM_R_X103Y102_SLICE_X163Y102_A4;
  wire [0:0] CLBLM_R_X103Y102_SLICE_X163Y102_A5;
  wire [0:0] CLBLM_R_X103Y102_SLICE_X163Y102_A6;
  wire [0:0] CLBLM_R_X103Y102_SLICE_X163Y102_AO5;
  wire [0:0] CLBLM_R_X103Y102_SLICE_X163Y102_AO6;
  wire [0:0] CLBLM_R_X103Y102_SLICE_X163Y102_A_CY;
  wire [0:0] CLBLM_R_X103Y102_SLICE_X163Y102_A_XOR;
  wire [0:0] CLBLM_R_X103Y102_SLICE_X163Y102_B;
  wire [0:0] CLBLM_R_X103Y102_SLICE_X163Y102_B1;
  wire [0:0] CLBLM_R_X103Y102_SLICE_X163Y102_B2;
  wire [0:0] CLBLM_R_X103Y102_SLICE_X163Y102_B3;
  wire [0:0] CLBLM_R_X103Y102_SLICE_X163Y102_B4;
  wire [0:0] CLBLM_R_X103Y102_SLICE_X163Y102_B5;
  wire [0:0] CLBLM_R_X103Y102_SLICE_X163Y102_B6;
  wire [0:0] CLBLM_R_X103Y102_SLICE_X163Y102_BO5;
  wire [0:0] CLBLM_R_X103Y102_SLICE_X163Y102_BO6;
  wire [0:0] CLBLM_R_X103Y102_SLICE_X163Y102_B_CY;
  wire [0:0] CLBLM_R_X103Y102_SLICE_X163Y102_B_XOR;
  wire [0:0] CLBLM_R_X103Y102_SLICE_X163Y102_C;
  wire [0:0] CLBLM_R_X103Y102_SLICE_X163Y102_C1;
  wire [0:0] CLBLM_R_X103Y102_SLICE_X163Y102_C2;
  wire [0:0] CLBLM_R_X103Y102_SLICE_X163Y102_C3;
  wire [0:0] CLBLM_R_X103Y102_SLICE_X163Y102_C4;
  wire [0:0] CLBLM_R_X103Y102_SLICE_X163Y102_C5;
  wire [0:0] CLBLM_R_X103Y102_SLICE_X163Y102_C6;
  wire [0:0] CLBLM_R_X103Y102_SLICE_X163Y102_CO5;
  wire [0:0] CLBLM_R_X103Y102_SLICE_X163Y102_CO6;
  wire [0:0] CLBLM_R_X103Y102_SLICE_X163Y102_C_CY;
  wire [0:0] CLBLM_R_X103Y102_SLICE_X163Y102_C_XOR;
  wire [0:0] CLBLM_R_X103Y102_SLICE_X163Y102_D;
  wire [0:0] CLBLM_R_X103Y102_SLICE_X163Y102_D1;
  wire [0:0] CLBLM_R_X103Y102_SLICE_X163Y102_D2;
  wire [0:0] CLBLM_R_X103Y102_SLICE_X163Y102_D3;
  wire [0:0] CLBLM_R_X103Y102_SLICE_X163Y102_D4;
  wire [0:0] CLBLM_R_X103Y102_SLICE_X163Y102_D5;
  wire [0:0] CLBLM_R_X103Y102_SLICE_X163Y102_D6;
  wire [0:0] CLBLM_R_X103Y102_SLICE_X163Y102_DO5;
  wire [0:0] CLBLM_R_X103Y102_SLICE_X163Y102_DO6;
  wire [0:0] CLBLM_R_X103Y102_SLICE_X163Y102_D_CY;
  wire [0:0] CLBLM_R_X103Y102_SLICE_X163Y102_D_XOR;
  wire [0:0] CLBLM_R_X103Y107_SLICE_X162Y107_A;
  wire [0:0] CLBLM_R_X103Y107_SLICE_X162Y107_A1;
  wire [0:0] CLBLM_R_X103Y107_SLICE_X162Y107_A2;
  wire [0:0] CLBLM_R_X103Y107_SLICE_X162Y107_A3;
  wire [0:0] CLBLM_R_X103Y107_SLICE_X162Y107_A4;
  wire [0:0] CLBLM_R_X103Y107_SLICE_X162Y107_A5;
  wire [0:0] CLBLM_R_X103Y107_SLICE_X162Y107_A6;
  wire [0:0] CLBLM_R_X103Y107_SLICE_X162Y107_AO5;
  wire [0:0] CLBLM_R_X103Y107_SLICE_X162Y107_AO6;
  wire [0:0] CLBLM_R_X103Y107_SLICE_X162Y107_A_CY;
  wire [0:0] CLBLM_R_X103Y107_SLICE_X162Y107_A_XOR;
  wire [0:0] CLBLM_R_X103Y107_SLICE_X162Y107_B;
  wire [0:0] CLBLM_R_X103Y107_SLICE_X162Y107_B1;
  wire [0:0] CLBLM_R_X103Y107_SLICE_X162Y107_B2;
  wire [0:0] CLBLM_R_X103Y107_SLICE_X162Y107_B3;
  wire [0:0] CLBLM_R_X103Y107_SLICE_X162Y107_B4;
  wire [0:0] CLBLM_R_X103Y107_SLICE_X162Y107_B5;
  wire [0:0] CLBLM_R_X103Y107_SLICE_X162Y107_B6;
  wire [0:0] CLBLM_R_X103Y107_SLICE_X162Y107_BO5;
  wire [0:0] CLBLM_R_X103Y107_SLICE_X162Y107_BO6;
  wire [0:0] CLBLM_R_X103Y107_SLICE_X162Y107_B_CY;
  wire [0:0] CLBLM_R_X103Y107_SLICE_X162Y107_B_XOR;
  wire [0:0] CLBLM_R_X103Y107_SLICE_X162Y107_C;
  wire [0:0] CLBLM_R_X103Y107_SLICE_X162Y107_C1;
  wire [0:0] CLBLM_R_X103Y107_SLICE_X162Y107_C2;
  wire [0:0] CLBLM_R_X103Y107_SLICE_X162Y107_C3;
  wire [0:0] CLBLM_R_X103Y107_SLICE_X162Y107_C4;
  wire [0:0] CLBLM_R_X103Y107_SLICE_X162Y107_C5;
  wire [0:0] CLBLM_R_X103Y107_SLICE_X162Y107_C6;
  wire [0:0] CLBLM_R_X103Y107_SLICE_X162Y107_CO5;
  wire [0:0] CLBLM_R_X103Y107_SLICE_X162Y107_CO6;
  wire [0:0] CLBLM_R_X103Y107_SLICE_X162Y107_C_CY;
  wire [0:0] CLBLM_R_X103Y107_SLICE_X162Y107_C_XOR;
  wire [0:0] CLBLM_R_X103Y107_SLICE_X162Y107_D;
  wire [0:0] CLBLM_R_X103Y107_SLICE_X162Y107_D1;
  wire [0:0] CLBLM_R_X103Y107_SLICE_X162Y107_D2;
  wire [0:0] CLBLM_R_X103Y107_SLICE_X162Y107_D3;
  wire [0:0] CLBLM_R_X103Y107_SLICE_X162Y107_D4;
  wire [0:0] CLBLM_R_X103Y107_SLICE_X162Y107_D5;
  wire [0:0] CLBLM_R_X103Y107_SLICE_X162Y107_D6;
  wire [0:0] CLBLM_R_X103Y107_SLICE_X162Y107_DO5;
  wire [0:0] CLBLM_R_X103Y107_SLICE_X162Y107_DO6;
  wire [0:0] CLBLM_R_X103Y107_SLICE_X162Y107_D_CY;
  wire [0:0] CLBLM_R_X103Y107_SLICE_X162Y107_D_XOR;
  wire [0:0] CLBLM_R_X103Y107_SLICE_X163Y107_A;
  wire [0:0] CLBLM_R_X103Y107_SLICE_X163Y107_A1;
  wire [0:0] CLBLM_R_X103Y107_SLICE_X163Y107_A2;
  wire [0:0] CLBLM_R_X103Y107_SLICE_X163Y107_A3;
  wire [0:0] CLBLM_R_X103Y107_SLICE_X163Y107_A4;
  wire [0:0] CLBLM_R_X103Y107_SLICE_X163Y107_A5;
  wire [0:0] CLBLM_R_X103Y107_SLICE_X163Y107_A6;
  wire [0:0] CLBLM_R_X103Y107_SLICE_X163Y107_AMUX;
  wire [0:0] CLBLM_R_X103Y107_SLICE_X163Y107_AO5;
  wire [0:0] CLBLM_R_X103Y107_SLICE_X163Y107_AO6;
  wire [0:0] CLBLM_R_X103Y107_SLICE_X163Y107_A_CY;
  wire [0:0] CLBLM_R_X103Y107_SLICE_X163Y107_A_XOR;
  wire [0:0] CLBLM_R_X103Y107_SLICE_X163Y107_B;
  wire [0:0] CLBLM_R_X103Y107_SLICE_X163Y107_B1;
  wire [0:0] CLBLM_R_X103Y107_SLICE_X163Y107_B2;
  wire [0:0] CLBLM_R_X103Y107_SLICE_X163Y107_B3;
  wire [0:0] CLBLM_R_X103Y107_SLICE_X163Y107_B4;
  wire [0:0] CLBLM_R_X103Y107_SLICE_X163Y107_B5;
  wire [0:0] CLBLM_R_X103Y107_SLICE_X163Y107_B6;
  wire [0:0] CLBLM_R_X103Y107_SLICE_X163Y107_BO5;
  wire [0:0] CLBLM_R_X103Y107_SLICE_X163Y107_BO6;
  wire [0:0] CLBLM_R_X103Y107_SLICE_X163Y107_B_CY;
  wire [0:0] CLBLM_R_X103Y107_SLICE_X163Y107_B_XOR;
  wire [0:0] CLBLM_R_X103Y107_SLICE_X163Y107_C;
  wire [0:0] CLBLM_R_X103Y107_SLICE_X163Y107_C1;
  wire [0:0] CLBLM_R_X103Y107_SLICE_X163Y107_C2;
  wire [0:0] CLBLM_R_X103Y107_SLICE_X163Y107_C3;
  wire [0:0] CLBLM_R_X103Y107_SLICE_X163Y107_C4;
  wire [0:0] CLBLM_R_X103Y107_SLICE_X163Y107_C5;
  wire [0:0] CLBLM_R_X103Y107_SLICE_X163Y107_C6;
  wire [0:0] CLBLM_R_X103Y107_SLICE_X163Y107_CO5;
  wire [0:0] CLBLM_R_X103Y107_SLICE_X163Y107_CO6;
  wire [0:0] CLBLM_R_X103Y107_SLICE_X163Y107_C_CY;
  wire [0:0] CLBLM_R_X103Y107_SLICE_X163Y107_C_XOR;
  wire [0:0] CLBLM_R_X103Y107_SLICE_X163Y107_D;
  wire [0:0] CLBLM_R_X103Y107_SLICE_X163Y107_D1;
  wire [0:0] CLBLM_R_X103Y107_SLICE_X163Y107_D2;
  wire [0:0] CLBLM_R_X103Y107_SLICE_X163Y107_D3;
  wire [0:0] CLBLM_R_X103Y107_SLICE_X163Y107_D4;
  wire [0:0] CLBLM_R_X103Y107_SLICE_X163Y107_D5;
  wire [0:0] CLBLM_R_X103Y107_SLICE_X163Y107_D6;
  wire [0:0] CLBLM_R_X103Y107_SLICE_X163Y107_DO5;
  wire [0:0] CLBLM_R_X103Y107_SLICE_X163Y107_DO6;
  wire [0:0] CLBLM_R_X103Y107_SLICE_X163Y107_D_CY;
  wire [0:0] CLBLM_R_X103Y107_SLICE_X163Y107_D_XOR;
  wire [0:0] CLBLM_R_X103Y108_SLICE_X162Y108_A;
  wire [0:0] CLBLM_R_X103Y108_SLICE_X162Y108_A1;
  wire [0:0] CLBLM_R_X103Y108_SLICE_X162Y108_A2;
  wire [0:0] CLBLM_R_X103Y108_SLICE_X162Y108_A3;
  wire [0:0] CLBLM_R_X103Y108_SLICE_X162Y108_A4;
  wire [0:0] CLBLM_R_X103Y108_SLICE_X162Y108_A5;
  wire [0:0] CLBLM_R_X103Y108_SLICE_X162Y108_A6;
  wire [0:0] CLBLM_R_X103Y108_SLICE_X162Y108_AO5;
  wire [0:0] CLBLM_R_X103Y108_SLICE_X162Y108_AO6;
  wire [0:0] CLBLM_R_X103Y108_SLICE_X162Y108_A_CY;
  wire [0:0] CLBLM_R_X103Y108_SLICE_X162Y108_A_XOR;
  wire [0:0] CLBLM_R_X103Y108_SLICE_X162Y108_B;
  wire [0:0] CLBLM_R_X103Y108_SLICE_X162Y108_B1;
  wire [0:0] CLBLM_R_X103Y108_SLICE_X162Y108_B2;
  wire [0:0] CLBLM_R_X103Y108_SLICE_X162Y108_B3;
  wire [0:0] CLBLM_R_X103Y108_SLICE_X162Y108_B4;
  wire [0:0] CLBLM_R_X103Y108_SLICE_X162Y108_B5;
  wire [0:0] CLBLM_R_X103Y108_SLICE_X162Y108_B6;
  wire [0:0] CLBLM_R_X103Y108_SLICE_X162Y108_BO5;
  wire [0:0] CLBLM_R_X103Y108_SLICE_X162Y108_BO6;
  wire [0:0] CLBLM_R_X103Y108_SLICE_X162Y108_B_CY;
  wire [0:0] CLBLM_R_X103Y108_SLICE_X162Y108_B_XOR;
  wire [0:0] CLBLM_R_X103Y108_SLICE_X162Y108_C;
  wire [0:0] CLBLM_R_X103Y108_SLICE_X162Y108_C1;
  wire [0:0] CLBLM_R_X103Y108_SLICE_X162Y108_C2;
  wire [0:0] CLBLM_R_X103Y108_SLICE_X162Y108_C3;
  wire [0:0] CLBLM_R_X103Y108_SLICE_X162Y108_C4;
  wire [0:0] CLBLM_R_X103Y108_SLICE_X162Y108_C5;
  wire [0:0] CLBLM_R_X103Y108_SLICE_X162Y108_C6;
  wire [0:0] CLBLM_R_X103Y108_SLICE_X162Y108_CO5;
  wire [0:0] CLBLM_R_X103Y108_SLICE_X162Y108_CO6;
  wire [0:0] CLBLM_R_X103Y108_SLICE_X162Y108_C_CY;
  wire [0:0] CLBLM_R_X103Y108_SLICE_X162Y108_C_XOR;
  wire [0:0] CLBLM_R_X103Y108_SLICE_X162Y108_D;
  wire [0:0] CLBLM_R_X103Y108_SLICE_X162Y108_D1;
  wire [0:0] CLBLM_R_X103Y108_SLICE_X162Y108_D2;
  wire [0:0] CLBLM_R_X103Y108_SLICE_X162Y108_D3;
  wire [0:0] CLBLM_R_X103Y108_SLICE_X162Y108_D4;
  wire [0:0] CLBLM_R_X103Y108_SLICE_X162Y108_D5;
  wire [0:0] CLBLM_R_X103Y108_SLICE_X162Y108_D6;
  wire [0:0] CLBLM_R_X103Y108_SLICE_X162Y108_DO5;
  wire [0:0] CLBLM_R_X103Y108_SLICE_X162Y108_DO6;
  wire [0:0] CLBLM_R_X103Y108_SLICE_X162Y108_D_CY;
  wire [0:0] CLBLM_R_X103Y108_SLICE_X162Y108_D_XOR;
  wire [0:0] CLBLM_R_X103Y108_SLICE_X163Y108_A;
  wire [0:0] CLBLM_R_X103Y108_SLICE_X163Y108_A1;
  wire [0:0] CLBLM_R_X103Y108_SLICE_X163Y108_A2;
  wire [0:0] CLBLM_R_X103Y108_SLICE_X163Y108_A3;
  wire [0:0] CLBLM_R_X103Y108_SLICE_X163Y108_A4;
  wire [0:0] CLBLM_R_X103Y108_SLICE_X163Y108_A5;
  wire [0:0] CLBLM_R_X103Y108_SLICE_X163Y108_A6;
  wire [0:0] CLBLM_R_X103Y108_SLICE_X163Y108_AMUX;
  wire [0:0] CLBLM_R_X103Y108_SLICE_X163Y108_AO5;
  wire [0:0] CLBLM_R_X103Y108_SLICE_X163Y108_AO6;
  wire [0:0] CLBLM_R_X103Y108_SLICE_X163Y108_A_CY;
  wire [0:0] CLBLM_R_X103Y108_SLICE_X163Y108_A_XOR;
  wire [0:0] CLBLM_R_X103Y108_SLICE_X163Y108_B;
  wire [0:0] CLBLM_R_X103Y108_SLICE_X163Y108_B1;
  wire [0:0] CLBLM_R_X103Y108_SLICE_X163Y108_B2;
  wire [0:0] CLBLM_R_X103Y108_SLICE_X163Y108_B3;
  wire [0:0] CLBLM_R_X103Y108_SLICE_X163Y108_B4;
  wire [0:0] CLBLM_R_X103Y108_SLICE_X163Y108_B5;
  wire [0:0] CLBLM_R_X103Y108_SLICE_X163Y108_B6;
  wire [0:0] CLBLM_R_X103Y108_SLICE_X163Y108_BO5;
  wire [0:0] CLBLM_R_X103Y108_SLICE_X163Y108_BO6;
  wire [0:0] CLBLM_R_X103Y108_SLICE_X163Y108_B_CY;
  wire [0:0] CLBLM_R_X103Y108_SLICE_X163Y108_B_XOR;
  wire [0:0] CLBLM_R_X103Y108_SLICE_X163Y108_C;
  wire [0:0] CLBLM_R_X103Y108_SLICE_X163Y108_C1;
  wire [0:0] CLBLM_R_X103Y108_SLICE_X163Y108_C2;
  wire [0:0] CLBLM_R_X103Y108_SLICE_X163Y108_C3;
  wire [0:0] CLBLM_R_X103Y108_SLICE_X163Y108_C4;
  wire [0:0] CLBLM_R_X103Y108_SLICE_X163Y108_C5;
  wire [0:0] CLBLM_R_X103Y108_SLICE_X163Y108_C6;
  wire [0:0] CLBLM_R_X103Y108_SLICE_X163Y108_CO5;
  wire [0:0] CLBLM_R_X103Y108_SLICE_X163Y108_CO6;
  wire [0:0] CLBLM_R_X103Y108_SLICE_X163Y108_C_CY;
  wire [0:0] CLBLM_R_X103Y108_SLICE_X163Y108_C_XOR;
  wire [0:0] CLBLM_R_X103Y108_SLICE_X163Y108_D;
  wire [0:0] CLBLM_R_X103Y108_SLICE_X163Y108_D1;
  wire [0:0] CLBLM_R_X103Y108_SLICE_X163Y108_D2;
  wire [0:0] CLBLM_R_X103Y108_SLICE_X163Y108_D3;
  wire [0:0] CLBLM_R_X103Y108_SLICE_X163Y108_D4;
  wire [0:0] CLBLM_R_X103Y108_SLICE_X163Y108_D5;
  wire [0:0] CLBLM_R_X103Y108_SLICE_X163Y108_D6;
  wire [0:0] CLBLM_R_X103Y108_SLICE_X163Y108_DO5;
  wire [0:0] CLBLM_R_X103Y108_SLICE_X163Y108_DO6;
  wire [0:0] CLBLM_R_X103Y108_SLICE_X163Y108_D_CY;
  wire [0:0] CLBLM_R_X103Y108_SLICE_X163Y108_D_XOR;
  wire [0:0] CLBLM_R_X103Y115_SLICE_X162Y115_A;
  wire [0:0] CLBLM_R_X103Y115_SLICE_X162Y115_A1;
  wire [0:0] CLBLM_R_X103Y115_SLICE_X162Y115_A2;
  wire [0:0] CLBLM_R_X103Y115_SLICE_X162Y115_A3;
  wire [0:0] CLBLM_R_X103Y115_SLICE_X162Y115_A4;
  wire [0:0] CLBLM_R_X103Y115_SLICE_X162Y115_A5;
  wire [0:0] CLBLM_R_X103Y115_SLICE_X162Y115_A6;
  wire [0:0] CLBLM_R_X103Y115_SLICE_X162Y115_AO5;
  wire [0:0] CLBLM_R_X103Y115_SLICE_X162Y115_AO6;
  wire [0:0] CLBLM_R_X103Y115_SLICE_X162Y115_A_CY;
  wire [0:0] CLBLM_R_X103Y115_SLICE_X162Y115_A_XOR;
  wire [0:0] CLBLM_R_X103Y115_SLICE_X162Y115_B;
  wire [0:0] CLBLM_R_X103Y115_SLICE_X162Y115_B1;
  wire [0:0] CLBLM_R_X103Y115_SLICE_X162Y115_B2;
  wire [0:0] CLBLM_R_X103Y115_SLICE_X162Y115_B3;
  wire [0:0] CLBLM_R_X103Y115_SLICE_X162Y115_B4;
  wire [0:0] CLBLM_R_X103Y115_SLICE_X162Y115_B5;
  wire [0:0] CLBLM_R_X103Y115_SLICE_X162Y115_B6;
  wire [0:0] CLBLM_R_X103Y115_SLICE_X162Y115_BO5;
  wire [0:0] CLBLM_R_X103Y115_SLICE_X162Y115_BO6;
  wire [0:0] CLBLM_R_X103Y115_SLICE_X162Y115_B_CY;
  wire [0:0] CLBLM_R_X103Y115_SLICE_X162Y115_B_XOR;
  wire [0:0] CLBLM_R_X103Y115_SLICE_X162Y115_C;
  wire [0:0] CLBLM_R_X103Y115_SLICE_X162Y115_C1;
  wire [0:0] CLBLM_R_X103Y115_SLICE_X162Y115_C2;
  wire [0:0] CLBLM_R_X103Y115_SLICE_X162Y115_C3;
  wire [0:0] CLBLM_R_X103Y115_SLICE_X162Y115_C4;
  wire [0:0] CLBLM_R_X103Y115_SLICE_X162Y115_C5;
  wire [0:0] CLBLM_R_X103Y115_SLICE_X162Y115_C6;
  wire [0:0] CLBLM_R_X103Y115_SLICE_X162Y115_CO5;
  wire [0:0] CLBLM_R_X103Y115_SLICE_X162Y115_CO6;
  wire [0:0] CLBLM_R_X103Y115_SLICE_X162Y115_C_CY;
  wire [0:0] CLBLM_R_X103Y115_SLICE_X162Y115_C_XOR;
  wire [0:0] CLBLM_R_X103Y115_SLICE_X162Y115_D;
  wire [0:0] CLBLM_R_X103Y115_SLICE_X162Y115_D1;
  wire [0:0] CLBLM_R_X103Y115_SLICE_X162Y115_D2;
  wire [0:0] CLBLM_R_X103Y115_SLICE_X162Y115_D3;
  wire [0:0] CLBLM_R_X103Y115_SLICE_X162Y115_D4;
  wire [0:0] CLBLM_R_X103Y115_SLICE_X162Y115_D5;
  wire [0:0] CLBLM_R_X103Y115_SLICE_X162Y115_D6;
  wire [0:0] CLBLM_R_X103Y115_SLICE_X162Y115_DO5;
  wire [0:0] CLBLM_R_X103Y115_SLICE_X162Y115_DO6;
  wire [0:0] CLBLM_R_X103Y115_SLICE_X162Y115_D_CY;
  wire [0:0] CLBLM_R_X103Y115_SLICE_X162Y115_D_XOR;
  wire [0:0] CLBLM_R_X103Y115_SLICE_X163Y115_A;
  wire [0:0] CLBLM_R_X103Y115_SLICE_X163Y115_A1;
  wire [0:0] CLBLM_R_X103Y115_SLICE_X163Y115_A2;
  wire [0:0] CLBLM_R_X103Y115_SLICE_X163Y115_A3;
  wire [0:0] CLBLM_R_X103Y115_SLICE_X163Y115_A4;
  wire [0:0] CLBLM_R_X103Y115_SLICE_X163Y115_A5;
  wire [0:0] CLBLM_R_X103Y115_SLICE_X163Y115_A6;
  wire [0:0] CLBLM_R_X103Y115_SLICE_X163Y115_AO5;
  wire [0:0] CLBLM_R_X103Y115_SLICE_X163Y115_AO6;
  wire [0:0] CLBLM_R_X103Y115_SLICE_X163Y115_A_CY;
  wire [0:0] CLBLM_R_X103Y115_SLICE_X163Y115_A_XOR;
  wire [0:0] CLBLM_R_X103Y115_SLICE_X163Y115_B;
  wire [0:0] CLBLM_R_X103Y115_SLICE_X163Y115_B1;
  wire [0:0] CLBLM_R_X103Y115_SLICE_X163Y115_B2;
  wire [0:0] CLBLM_R_X103Y115_SLICE_X163Y115_B3;
  wire [0:0] CLBLM_R_X103Y115_SLICE_X163Y115_B4;
  wire [0:0] CLBLM_R_X103Y115_SLICE_X163Y115_B5;
  wire [0:0] CLBLM_R_X103Y115_SLICE_X163Y115_B6;
  wire [0:0] CLBLM_R_X103Y115_SLICE_X163Y115_BO5;
  wire [0:0] CLBLM_R_X103Y115_SLICE_X163Y115_BO6;
  wire [0:0] CLBLM_R_X103Y115_SLICE_X163Y115_B_CY;
  wire [0:0] CLBLM_R_X103Y115_SLICE_X163Y115_B_XOR;
  wire [0:0] CLBLM_R_X103Y115_SLICE_X163Y115_C;
  wire [0:0] CLBLM_R_X103Y115_SLICE_X163Y115_C1;
  wire [0:0] CLBLM_R_X103Y115_SLICE_X163Y115_C2;
  wire [0:0] CLBLM_R_X103Y115_SLICE_X163Y115_C3;
  wire [0:0] CLBLM_R_X103Y115_SLICE_X163Y115_C4;
  wire [0:0] CLBLM_R_X103Y115_SLICE_X163Y115_C5;
  wire [0:0] CLBLM_R_X103Y115_SLICE_X163Y115_C6;
  wire [0:0] CLBLM_R_X103Y115_SLICE_X163Y115_CO5;
  wire [0:0] CLBLM_R_X103Y115_SLICE_X163Y115_CO6;
  wire [0:0] CLBLM_R_X103Y115_SLICE_X163Y115_C_CY;
  wire [0:0] CLBLM_R_X103Y115_SLICE_X163Y115_C_XOR;
  wire [0:0] CLBLM_R_X103Y115_SLICE_X163Y115_D;
  wire [0:0] CLBLM_R_X103Y115_SLICE_X163Y115_D1;
  wire [0:0] CLBLM_R_X103Y115_SLICE_X163Y115_D2;
  wire [0:0] CLBLM_R_X103Y115_SLICE_X163Y115_D3;
  wire [0:0] CLBLM_R_X103Y115_SLICE_X163Y115_D4;
  wire [0:0] CLBLM_R_X103Y115_SLICE_X163Y115_D5;
  wire [0:0] CLBLM_R_X103Y115_SLICE_X163Y115_D6;
  wire [0:0] CLBLM_R_X103Y115_SLICE_X163Y115_DO5;
  wire [0:0] CLBLM_R_X103Y115_SLICE_X163Y115_DO6;
  wire [0:0] CLBLM_R_X103Y115_SLICE_X163Y115_D_CY;
  wire [0:0] CLBLM_R_X103Y115_SLICE_X163Y115_D_XOR;
  wire [0:0] CLBLM_R_X103Y122_SLICE_X162Y122_A;
  wire [0:0] CLBLM_R_X103Y122_SLICE_X162Y122_A1;
  wire [0:0] CLBLM_R_X103Y122_SLICE_X162Y122_A2;
  wire [0:0] CLBLM_R_X103Y122_SLICE_X162Y122_A3;
  wire [0:0] CLBLM_R_X103Y122_SLICE_X162Y122_A4;
  wire [0:0] CLBLM_R_X103Y122_SLICE_X162Y122_A5;
  wire [0:0] CLBLM_R_X103Y122_SLICE_X162Y122_A6;
  wire [0:0] CLBLM_R_X103Y122_SLICE_X162Y122_AO5;
  wire [0:0] CLBLM_R_X103Y122_SLICE_X162Y122_AO6;
  wire [0:0] CLBLM_R_X103Y122_SLICE_X162Y122_A_CY;
  wire [0:0] CLBLM_R_X103Y122_SLICE_X162Y122_A_XOR;
  wire [0:0] CLBLM_R_X103Y122_SLICE_X162Y122_B;
  wire [0:0] CLBLM_R_X103Y122_SLICE_X162Y122_B1;
  wire [0:0] CLBLM_R_X103Y122_SLICE_X162Y122_B2;
  wire [0:0] CLBLM_R_X103Y122_SLICE_X162Y122_B3;
  wire [0:0] CLBLM_R_X103Y122_SLICE_X162Y122_B4;
  wire [0:0] CLBLM_R_X103Y122_SLICE_X162Y122_B5;
  wire [0:0] CLBLM_R_X103Y122_SLICE_X162Y122_B6;
  wire [0:0] CLBLM_R_X103Y122_SLICE_X162Y122_BO5;
  wire [0:0] CLBLM_R_X103Y122_SLICE_X162Y122_BO6;
  wire [0:0] CLBLM_R_X103Y122_SLICE_X162Y122_B_CY;
  wire [0:0] CLBLM_R_X103Y122_SLICE_X162Y122_B_XOR;
  wire [0:0] CLBLM_R_X103Y122_SLICE_X162Y122_C;
  wire [0:0] CLBLM_R_X103Y122_SLICE_X162Y122_C1;
  wire [0:0] CLBLM_R_X103Y122_SLICE_X162Y122_C2;
  wire [0:0] CLBLM_R_X103Y122_SLICE_X162Y122_C3;
  wire [0:0] CLBLM_R_X103Y122_SLICE_X162Y122_C4;
  wire [0:0] CLBLM_R_X103Y122_SLICE_X162Y122_C5;
  wire [0:0] CLBLM_R_X103Y122_SLICE_X162Y122_C6;
  wire [0:0] CLBLM_R_X103Y122_SLICE_X162Y122_CO5;
  wire [0:0] CLBLM_R_X103Y122_SLICE_X162Y122_CO6;
  wire [0:0] CLBLM_R_X103Y122_SLICE_X162Y122_C_CY;
  wire [0:0] CLBLM_R_X103Y122_SLICE_X162Y122_C_XOR;
  wire [0:0] CLBLM_R_X103Y122_SLICE_X162Y122_D;
  wire [0:0] CLBLM_R_X103Y122_SLICE_X162Y122_D1;
  wire [0:0] CLBLM_R_X103Y122_SLICE_X162Y122_D2;
  wire [0:0] CLBLM_R_X103Y122_SLICE_X162Y122_D3;
  wire [0:0] CLBLM_R_X103Y122_SLICE_X162Y122_D4;
  wire [0:0] CLBLM_R_X103Y122_SLICE_X162Y122_D5;
  wire [0:0] CLBLM_R_X103Y122_SLICE_X162Y122_D6;
  wire [0:0] CLBLM_R_X103Y122_SLICE_X162Y122_DO5;
  wire [0:0] CLBLM_R_X103Y122_SLICE_X162Y122_DO6;
  wire [0:0] CLBLM_R_X103Y122_SLICE_X162Y122_D_CY;
  wire [0:0] CLBLM_R_X103Y122_SLICE_X162Y122_D_XOR;
  wire [0:0] CLBLM_R_X103Y122_SLICE_X163Y122_A;
  wire [0:0] CLBLM_R_X103Y122_SLICE_X163Y122_A1;
  wire [0:0] CLBLM_R_X103Y122_SLICE_X163Y122_A2;
  wire [0:0] CLBLM_R_X103Y122_SLICE_X163Y122_A3;
  wire [0:0] CLBLM_R_X103Y122_SLICE_X163Y122_A4;
  wire [0:0] CLBLM_R_X103Y122_SLICE_X163Y122_A5;
  wire [0:0] CLBLM_R_X103Y122_SLICE_X163Y122_A6;
  wire [0:0] CLBLM_R_X103Y122_SLICE_X163Y122_AMUX;
  wire [0:0] CLBLM_R_X103Y122_SLICE_X163Y122_AO5;
  wire [0:0] CLBLM_R_X103Y122_SLICE_X163Y122_AO6;
  wire [0:0] CLBLM_R_X103Y122_SLICE_X163Y122_A_CY;
  wire [0:0] CLBLM_R_X103Y122_SLICE_X163Y122_A_XOR;
  wire [0:0] CLBLM_R_X103Y122_SLICE_X163Y122_B;
  wire [0:0] CLBLM_R_X103Y122_SLICE_X163Y122_B1;
  wire [0:0] CLBLM_R_X103Y122_SLICE_X163Y122_B2;
  wire [0:0] CLBLM_R_X103Y122_SLICE_X163Y122_B3;
  wire [0:0] CLBLM_R_X103Y122_SLICE_X163Y122_B4;
  wire [0:0] CLBLM_R_X103Y122_SLICE_X163Y122_B5;
  wire [0:0] CLBLM_R_X103Y122_SLICE_X163Y122_B6;
  wire [0:0] CLBLM_R_X103Y122_SLICE_X163Y122_BMUX;
  wire [0:0] CLBLM_R_X103Y122_SLICE_X163Y122_BO5;
  wire [0:0] CLBLM_R_X103Y122_SLICE_X163Y122_BO6;
  wire [0:0] CLBLM_R_X103Y122_SLICE_X163Y122_B_CY;
  wire [0:0] CLBLM_R_X103Y122_SLICE_X163Y122_B_XOR;
  wire [0:0] CLBLM_R_X103Y122_SLICE_X163Y122_C;
  wire [0:0] CLBLM_R_X103Y122_SLICE_X163Y122_C1;
  wire [0:0] CLBLM_R_X103Y122_SLICE_X163Y122_C2;
  wire [0:0] CLBLM_R_X103Y122_SLICE_X163Y122_C3;
  wire [0:0] CLBLM_R_X103Y122_SLICE_X163Y122_C4;
  wire [0:0] CLBLM_R_X103Y122_SLICE_X163Y122_C5;
  wire [0:0] CLBLM_R_X103Y122_SLICE_X163Y122_C6;
  wire [0:0] CLBLM_R_X103Y122_SLICE_X163Y122_CMUX;
  wire [0:0] CLBLM_R_X103Y122_SLICE_X163Y122_CO5;
  wire [0:0] CLBLM_R_X103Y122_SLICE_X163Y122_CO6;
  wire [0:0] CLBLM_R_X103Y122_SLICE_X163Y122_C_CY;
  wire [0:0] CLBLM_R_X103Y122_SLICE_X163Y122_C_XOR;
  wire [0:0] CLBLM_R_X103Y122_SLICE_X163Y122_D;
  wire [0:0] CLBLM_R_X103Y122_SLICE_X163Y122_D1;
  wire [0:0] CLBLM_R_X103Y122_SLICE_X163Y122_D2;
  wire [0:0] CLBLM_R_X103Y122_SLICE_X163Y122_D3;
  wire [0:0] CLBLM_R_X103Y122_SLICE_X163Y122_D4;
  wire [0:0] CLBLM_R_X103Y122_SLICE_X163Y122_D5;
  wire [0:0] CLBLM_R_X103Y122_SLICE_X163Y122_D6;
  wire [0:0] CLBLM_R_X103Y122_SLICE_X163Y122_DMUX;
  wire [0:0] CLBLM_R_X103Y122_SLICE_X163Y122_DO5;
  wire [0:0] CLBLM_R_X103Y122_SLICE_X163Y122_DO6;
  wire [0:0] CLBLM_R_X103Y122_SLICE_X163Y122_D_CY;
  wire [0:0] CLBLM_R_X103Y122_SLICE_X163Y122_D_XOR;
  wire [0:0] CLBLM_R_X103Y123_SLICE_X162Y123_A;
  wire [0:0] CLBLM_R_X103Y123_SLICE_X162Y123_A1;
  wire [0:0] CLBLM_R_X103Y123_SLICE_X162Y123_A2;
  wire [0:0] CLBLM_R_X103Y123_SLICE_X162Y123_A3;
  wire [0:0] CLBLM_R_X103Y123_SLICE_X162Y123_A4;
  wire [0:0] CLBLM_R_X103Y123_SLICE_X162Y123_A5;
  wire [0:0] CLBLM_R_X103Y123_SLICE_X162Y123_A6;
  wire [0:0] CLBLM_R_X103Y123_SLICE_X162Y123_AO5;
  wire [0:0] CLBLM_R_X103Y123_SLICE_X162Y123_AO6;
  wire [0:0] CLBLM_R_X103Y123_SLICE_X162Y123_A_CY;
  wire [0:0] CLBLM_R_X103Y123_SLICE_X162Y123_A_XOR;
  wire [0:0] CLBLM_R_X103Y123_SLICE_X162Y123_B;
  wire [0:0] CLBLM_R_X103Y123_SLICE_X162Y123_B1;
  wire [0:0] CLBLM_R_X103Y123_SLICE_X162Y123_B2;
  wire [0:0] CLBLM_R_X103Y123_SLICE_X162Y123_B3;
  wire [0:0] CLBLM_R_X103Y123_SLICE_X162Y123_B4;
  wire [0:0] CLBLM_R_X103Y123_SLICE_X162Y123_B5;
  wire [0:0] CLBLM_R_X103Y123_SLICE_X162Y123_B6;
  wire [0:0] CLBLM_R_X103Y123_SLICE_X162Y123_BO5;
  wire [0:0] CLBLM_R_X103Y123_SLICE_X162Y123_BO6;
  wire [0:0] CLBLM_R_X103Y123_SLICE_X162Y123_B_CY;
  wire [0:0] CLBLM_R_X103Y123_SLICE_X162Y123_B_XOR;
  wire [0:0] CLBLM_R_X103Y123_SLICE_X162Y123_C;
  wire [0:0] CLBLM_R_X103Y123_SLICE_X162Y123_C1;
  wire [0:0] CLBLM_R_X103Y123_SLICE_X162Y123_C2;
  wire [0:0] CLBLM_R_X103Y123_SLICE_X162Y123_C3;
  wire [0:0] CLBLM_R_X103Y123_SLICE_X162Y123_C4;
  wire [0:0] CLBLM_R_X103Y123_SLICE_X162Y123_C5;
  wire [0:0] CLBLM_R_X103Y123_SLICE_X162Y123_C6;
  wire [0:0] CLBLM_R_X103Y123_SLICE_X162Y123_CO5;
  wire [0:0] CLBLM_R_X103Y123_SLICE_X162Y123_CO6;
  wire [0:0] CLBLM_R_X103Y123_SLICE_X162Y123_C_CY;
  wire [0:0] CLBLM_R_X103Y123_SLICE_X162Y123_C_XOR;
  wire [0:0] CLBLM_R_X103Y123_SLICE_X162Y123_D;
  wire [0:0] CLBLM_R_X103Y123_SLICE_X162Y123_D1;
  wire [0:0] CLBLM_R_X103Y123_SLICE_X162Y123_D2;
  wire [0:0] CLBLM_R_X103Y123_SLICE_X162Y123_D3;
  wire [0:0] CLBLM_R_X103Y123_SLICE_X162Y123_D4;
  wire [0:0] CLBLM_R_X103Y123_SLICE_X162Y123_D5;
  wire [0:0] CLBLM_R_X103Y123_SLICE_X162Y123_D6;
  wire [0:0] CLBLM_R_X103Y123_SLICE_X162Y123_DO5;
  wire [0:0] CLBLM_R_X103Y123_SLICE_X162Y123_DO6;
  wire [0:0] CLBLM_R_X103Y123_SLICE_X162Y123_D_CY;
  wire [0:0] CLBLM_R_X103Y123_SLICE_X162Y123_D_XOR;
  wire [0:0] CLBLM_R_X103Y123_SLICE_X163Y123_A;
  wire [0:0] CLBLM_R_X103Y123_SLICE_X163Y123_A1;
  wire [0:0] CLBLM_R_X103Y123_SLICE_X163Y123_A2;
  wire [0:0] CLBLM_R_X103Y123_SLICE_X163Y123_A3;
  wire [0:0] CLBLM_R_X103Y123_SLICE_X163Y123_A4;
  wire [0:0] CLBLM_R_X103Y123_SLICE_X163Y123_A5;
  wire [0:0] CLBLM_R_X103Y123_SLICE_X163Y123_A6;
  wire [0:0] CLBLM_R_X103Y123_SLICE_X163Y123_AMUX;
  wire [0:0] CLBLM_R_X103Y123_SLICE_X163Y123_AO5;
  wire [0:0] CLBLM_R_X103Y123_SLICE_X163Y123_AO6;
  wire [0:0] CLBLM_R_X103Y123_SLICE_X163Y123_A_CY;
  wire [0:0] CLBLM_R_X103Y123_SLICE_X163Y123_A_XOR;
  wire [0:0] CLBLM_R_X103Y123_SLICE_X163Y123_B;
  wire [0:0] CLBLM_R_X103Y123_SLICE_X163Y123_B1;
  wire [0:0] CLBLM_R_X103Y123_SLICE_X163Y123_B2;
  wire [0:0] CLBLM_R_X103Y123_SLICE_X163Y123_B3;
  wire [0:0] CLBLM_R_X103Y123_SLICE_X163Y123_B4;
  wire [0:0] CLBLM_R_X103Y123_SLICE_X163Y123_B5;
  wire [0:0] CLBLM_R_X103Y123_SLICE_X163Y123_B6;
  wire [0:0] CLBLM_R_X103Y123_SLICE_X163Y123_BO5;
  wire [0:0] CLBLM_R_X103Y123_SLICE_X163Y123_BO6;
  wire [0:0] CLBLM_R_X103Y123_SLICE_X163Y123_B_CY;
  wire [0:0] CLBLM_R_X103Y123_SLICE_X163Y123_B_XOR;
  wire [0:0] CLBLM_R_X103Y123_SLICE_X163Y123_C;
  wire [0:0] CLBLM_R_X103Y123_SLICE_X163Y123_C1;
  wire [0:0] CLBLM_R_X103Y123_SLICE_X163Y123_C2;
  wire [0:0] CLBLM_R_X103Y123_SLICE_X163Y123_C3;
  wire [0:0] CLBLM_R_X103Y123_SLICE_X163Y123_C4;
  wire [0:0] CLBLM_R_X103Y123_SLICE_X163Y123_C5;
  wire [0:0] CLBLM_R_X103Y123_SLICE_X163Y123_C6;
  wire [0:0] CLBLM_R_X103Y123_SLICE_X163Y123_CO5;
  wire [0:0] CLBLM_R_X103Y123_SLICE_X163Y123_CO6;
  wire [0:0] CLBLM_R_X103Y123_SLICE_X163Y123_C_CY;
  wire [0:0] CLBLM_R_X103Y123_SLICE_X163Y123_C_XOR;
  wire [0:0] CLBLM_R_X103Y123_SLICE_X163Y123_D;
  wire [0:0] CLBLM_R_X103Y123_SLICE_X163Y123_D1;
  wire [0:0] CLBLM_R_X103Y123_SLICE_X163Y123_D2;
  wire [0:0] CLBLM_R_X103Y123_SLICE_X163Y123_D3;
  wire [0:0] CLBLM_R_X103Y123_SLICE_X163Y123_D4;
  wire [0:0] CLBLM_R_X103Y123_SLICE_X163Y123_D5;
  wire [0:0] CLBLM_R_X103Y123_SLICE_X163Y123_D6;
  wire [0:0] CLBLM_R_X103Y123_SLICE_X163Y123_DO5;
  wire [0:0] CLBLM_R_X103Y123_SLICE_X163Y123_DO6;
  wire [0:0] CLBLM_R_X103Y123_SLICE_X163Y123_D_CY;
  wire [0:0] CLBLM_R_X103Y123_SLICE_X163Y123_D_XOR;
  wire [0:0] CLBLM_R_X103Y147_SLICE_X162Y147_A;
  wire [0:0] CLBLM_R_X103Y147_SLICE_X162Y147_A1;
  wire [0:0] CLBLM_R_X103Y147_SLICE_X162Y147_A2;
  wire [0:0] CLBLM_R_X103Y147_SLICE_X162Y147_A3;
  wire [0:0] CLBLM_R_X103Y147_SLICE_X162Y147_A4;
  wire [0:0] CLBLM_R_X103Y147_SLICE_X162Y147_A5;
  wire [0:0] CLBLM_R_X103Y147_SLICE_X162Y147_A6;
  wire [0:0] CLBLM_R_X103Y147_SLICE_X162Y147_AO5;
  wire [0:0] CLBLM_R_X103Y147_SLICE_X162Y147_AO6;
  wire [0:0] CLBLM_R_X103Y147_SLICE_X162Y147_A_CY;
  wire [0:0] CLBLM_R_X103Y147_SLICE_X162Y147_A_XOR;
  wire [0:0] CLBLM_R_X103Y147_SLICE_X162Y147_B;
  wire [0:0] CLBLM_R_X103Y147_SLICE_X162Y147_B1;
  wire [0:0] CLBLM_R_X103Y147_SLICE_X162Y147_B2;
  wire [0:0] CLBLM_R_X103Y147_SLICE_X162Y147_B3;
  wire [0:0] CLBLM_R_X103Y147_SLICE_X162Y147_B4;
  wire [0:0] CLBLM_R_X103Y147_SLICE_X162Y147_B5;
  wire [0:0] CLBLM_R_X103Y147_SLICE_X162Y147_B6;
  wire [0:0] CLBLM_R_X103Y147_SLICE_X162Y147_BO5;
  wire [0:0] CLBLM_R_X103Y147_SLICE_X162Y147_BO6;
  wire [0:0] CLBLM_R_X103Y147_SLICE_X162Y147_B_CY;
  wire [0:0] CLBLM_R_X103Y147_SLICE_X162Y147_B_XOR;
  wire [0:0] CLBLM_R_X103Y147_SLICE_X162Y147_C;
  wire [0:0] CLBLM_R_X103Y147_SLICE_X162Y147_C1;
  wire [0:0] CLBLM_R_X103Y147_SLICE_X162Y147_C2;
  wire [0:0] CLBLM_R_X103Y147_SLICE_X162Y147_C3;
  wire [0:0] CLBLM_R_X103Y147_SLICE_X162Y147_C4;
  wire [0:0] CLBLM_R_X103Y147_SLICE_X162Y147_C5;
  wire [0:0] CLBLM_R_X103Y147_SLICE_X162Y147_C6;
  wire [0:0] CLBLM_R_X103Y147_SLICE_X162Y147_CO5;
  wire [0:0] CLBLM_R_X103Y147_SLICE_X162Y147_CO6;
  wire [0:0] CLBLM_R_X103Y147_SLICE_X162Y147_C_CY;
  wire [0:0] CLBLM_R_X103Y147_SLICE_X162Y147_C_XOR;
  wire [0:0] CLBLM_R_X103Y147_SLICE_X162Y147_D;
  wire [0:0] CLBLM_R_X103Y147_SLICE_X162Y147_D1;
  wire [0:0] CLBLM_R_X103Y147_SLICE_X162Y147_D2;
  wire [0:0] CLBLM_R_X103Y147_SLICE_X162Y147_D3;
  wire [0:0] CLBLM_R_X103Y147_SLICE_X162Y147_D4;
  wire [0:0] CLBLM_R_X103Y147_SLICE_X162Y147_D5;
  wire [0:0] CLBLM_R_X103Y147_SLICE_X162Y147_D6;
  wire [0:0] CLBLM_R_X103Y147_SLICE_X162Y147_DO5;
  wire [0:0] CLBLM_R_X103Y147_SLICE_X162Y147_DO6;
  wire [0:0] CLBLM_R_X103Y147_SLICE_X162Y147_D_CY;
  wire [0:0] CLBLM_R_X103Y147_SLICE_X162Y147_D_XOR;
  wire [0:0] CLBLM_R_X103Y147_SLICE_X163Y147_A;
  wire [0:0] CLBLM_R_X103Y147_SLICE_X163Y147_A1;
  wire [0:0] CLBLM_R_X103Y147_SLICE_X163Y147_A2;
  wire [0:0] CLBLM_R_X103Y147_SLICE_X163Y147_A3;
  wire [0:0] CLBLM_R_X103Y147_SLICE_X163Y147_A4;
  wire [0:0] CLBLM_R_X103Y147_SLICE_X163Y147_A5;
  wire [0:0] CLBLM_R_X103Y147_SLICE_X163Y147_A6;
  wire [0:0] CLBLM_R_X103Y147_SLICE_X163Y147_AMUX;
  wire [0:0] CLBLM_R_X103Y147_SLICE_X163Y147_AO5;
  wire [0:0] CLBLM_R_X103Y147_SLICE_X163Y147_AO6;
  wire [0:0] CLBLM_R_X103Y147_SLICE_X163Y147_A_CY;
  wire [0:0] CLBLM_R_X103Y147_SLICE_X163Y147_A_XOR;
  wire [0:0] CLBLM_R_X103Y147_SLICE_X163Y147_B;
  wire [0:0] CLBLM_R_X103Y147_SLICE_X163Y147_B1;
  wire [0:0] CLBLM_R_X103Y147_SLICE_X163Y147_B2;
  wire [0:0] CLBLM_R_X103Y147_SLICE_X163Y147_B3;
  wire [0:0] CLBLM_R_X103Y147_SLICE_X163Y147_B4;
  wire [0:0] CLBLM_R_X103Y147_SLICE_X163Y147_B5;
  wire [0:0] CLBLM_R_X103Y147_SLICE_X163Y147_B6;
  wire [0:0] CLBLM_R_X103Y147_SLICE_X163Y147_BO5;
  wire [0:0] CLBLM_R_X103Y147_SLICE_X163Y147_BO6;
  wire [0:0] CLBLM_R_X103Y147_SLICE_X163Y147_B_CY;
  wire [0:0] CLBLM_R_X103Y147_SLICE_X163Y147_B_XOR;
  wire [0:0] CLBLM_R_X103Y147_SLICE_X163Y147_C;
  wire [0:0] CLBLM_R_X103Y147_SLICE_X163Y147_C1;
  wire [0:0] CLBLM_R_X103Y147_SLICE_X163Y147_C2;
  wire [0:0] CLBLM_R_X103Y147_SLICE_X163Y147_C3;
  wire [0:0] CLBLM_R_X103Y147_SLICE_X163Y147_C4;
  wire [0:0] CLBLM_R_X103Y147_SLICE_X163Y147_C5;
  wire [0:0] CLBLM_R_X103Y147_SLICE_X163Y147_C6;
  wire [0:0] CLBLM_R_X103Y147_SLICE_X163Y147_CO5;
  wire [0:0] CLBLM_R_X103Y147_SLICE_X163Y147_CO6;
  wire [0:0] CLBLM_R_X103Y147_SLICE_X163Y147_C_CY;
  wire [0:0] CLBLM_R_X103Y147_SLICE_X163Y147_C_XOR;
  wire [0:0] CLBLM_R_X103Y147_SLICE_X163Y147_D;
  wire [0:0] CLBLM_R_X103Y147_SLICE_X163Y147_D1;
  wire [0:0] CLBLM_R_X103Y147_SLICE_X163Y147_D2;
  wire [0:0] CLBLM_R_X103Y147_SLICE_X163Y147_D3;
  wire [0:0] CLBLM_R_X103Y147_SLICE_X163Y147_D4;
  wire [0:0] CLBLM_R_X103Y147_SLICE_X163Y147_D5;
  wire [0:0] CLBLM_R_X103Y147_SLICE_X163Y147_D6;
  wire [0:0] CLBLM_R_X103Y147_SLICE_X163Y147_DO5;
  wire [0:0] CLBLM_R_X103Y147_SLICE_X163Y147_DO6;
  wire [0:0] CLBLM_R_X103Y147_SLICE_X163Y147_D_CY;
  wire [0:0] CLBLM_R_X103Y147_SLICE_X163Y147_D_XOR;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X162Y177_A;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X162Y177_A1;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X162Y177_A2;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X162Y177_A3;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X162Y177_A4;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X162Y177_A5;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X162Y177_A6;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X162Y177_AO5;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X162Y177_AO6;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X162Y177_A_CY;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X162Y177_A_XOR;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X162Y177_B;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X162Y177_B1;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X162Y177_B2;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X162Y177_B3;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X162Y177_B4;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X162Y177_B5;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X162Y177_B6;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X162Y177_BO5;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X162Y177_BO6;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X162Y177_B_CY;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X162Y177_B_XOR;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X162Y177_C;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X162Y177_C1;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X162Y177_C2;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X162Y177_C3;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X162Y177_C4;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X162Y177_C5;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X162Y177_C6;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X162Y177_CO5;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X162Y177_CO6;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X162Y177_C_CY;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X162Y177_C_XOR;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X162Y177_D;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X162Y177_D1;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X162Y177_D2;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X162Y177_D3;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X162Y177_D4;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X162Y177_D5;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X162Y177_D6;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X162Y177_DO5;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X162Y177_DO6;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X162Y177_D_CY;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X162Y177_D_XOR;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X163Y177_A;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X163Y177_A1;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X163Y177_A2;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X163Y177_A3;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X163Y177_A4;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X163Y177_A5;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X163Y177_A6;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X163Y177_AMUX;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X163Y177_AO5;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X163Y177_AO6;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X163Y177_A_CY;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X163Y177_A_XOR;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X163Y177_B;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X163Y177_B1;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X163Y177_B2;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X163Y177_B3;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X163Y177_B4;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X163Y177_B5;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X163Y177_B6;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X163Y177_BO5;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X163Y177_BO6;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X163Y177_B_CY;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X163Y177_B_XOR;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X163Y177_C;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X163Y177_C1;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X163Y177_C2;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X163Y177_C3;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X163Y177_C4;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X163Y177_C5;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X163Y177_C6;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X163Y177_CO5;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X163Y177_CO6;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X163Y177_C_CY;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X163Y177_C_XOR;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X163Y177_D;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X163Y177_D1;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X163Y177_D2;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X163Y177_D3;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X163Y177_D4;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X163Y177_D5;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X163Y177_D6;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X163Y177_DO5;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X163Y177_DO6;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X163Y177_D_CY;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X163Y177_D_XOR;
  wire [0:0] CLBLM_R_X103Y185_SLICE_X162Y185_A;
  wire [0:0] CLBLM_R_X103Y185_SLICE_X162Y185_A1;
  wire [0:0] CLBLM_R_X103Y185_SLICE_X162Y185_A2;
  wire [0:0] CLBLM_R_X103Y185_SLICE_X162Y185_A3;
  wire [0:0] CLBLM_R_X103Y185_SLICE_X162Y185_A4;
  wire [0:0] CLBLM_R_X103Y185_SLICE_X162Y185_A5;
  wire [0:0] CLBLM_R_X103Y185_SLICE_X162Y185_A6;
  wire [0:0] CLBLM_R_X103Y185_SLICE_X162Y185_AO5;
  wire [0:0] CLBLM_R_X103Y185_SLICE_X162Y185_AO6;
  wire [0:0] CLBLM_R_X103Y185_SLICE_X162Y185_A_CY;
  wire [0:0] CLBLM_R_X103Y185_SLICE_X162Y185_A_XOR;
  wire [0:0] CLBLM_R_X103Y185_SLICE_X162Y185_B;
  wire [0:0] CLBLM_R_X103Y185_SLICE_X162Y185_B1;
  wire [0:0] CLBLM_R_X103Y185_SLICE_X162Y185_B2;
  wire [0:0] CLBLM_R_X103Y185_SLICE_X162Y185_B3;
  wire [0:0] CLBLM_R_X103Y185_SLICE_X162Y185_B4;
  wire [0:0] CLBLM_R_X103Y185_SLICE_X162Y185_B5;
  wire [0:0] CLBLM_R_X103Y185_SLICE_X162Y185_B6;
  wire [0:0] CLBLM_R_X103Y185_SLICE_X162Y185_BO5;
  wire [0:0] CLBLM_R_X103Y185_SLICE_X162Y185_BO6;
  wire [0:0] CLBLM_R_X103Y185_SLICE_X162Y185_B_CY;
  wire [0:0] CLBLM_R_X103Y185_SLICE_X162Y185_B_XOR;
  wire [0:0] CLBLM_R_X103Y185_SLICE_X162Y185_C;
  wire [0:0] CLBLM_R_X103Y185_SLICE_X162Y185_C1;
  wire [0:0] CLBLM_R_X103Y185_SLICE_X162Y185_C2;
  wire [0:0] CLBLM_R_X103Y185_SLICE_X162Y185_C3;
  wire [0:0] CLBLM_R_X103Y185_SLICE_X162Y185_C4;
  wire [0:0] CLBLM_R_X103Y185_SLICE_X162Y185_C5;
  wire [0:0] CLBLM_R_X103Y185_SLICE_X162Y185_C6;
  wire [0:0] CLBLM_R_X103Y185_SLICE_X162Y185_CO5;
  wire [0:0] CLBLM_R_X103Y185_SLICE_X162Y185_CO6;
  wire [0:0] CLBLM_R_X103Y185_SLICE_X162Y185_C_CY;
  wire [0:0] CLBLM_R_X103Y185_SLICE_X162Y185_C_XOR;
  wire [0:0] CLBLM_R_X103Y185_SLICE_X162Y185_D;
  wire [0:0] CLBLM_R_X103Y185_SLICE_X162Y185_D1;
  wire [0:0] CLBLM_R_X103Y185_SLICE_X162Y185_D2;
  wire [0:0] CLBLM_R_X103Y185_SLICE_X162Y185_D3;
  wire [0:0] CLBLM_R_X103Y185_SLICE_X162Y185_D4;
  wire [0:0] CLBLM_R_X103Y185_SLICE_X162Y185_D5;
  wire [0:0] CLBLM_R_X103Y185_SLICE_X162Y185_D6;
  wire [0:0] CLBLM_R_X103Y185_SLICE_X162Y185_DO5;
  wire [0:0] CLBLM_R_X103Y185_SLICE_X162Y185_DO6;
  wire [0:0] CLBLM_R_X103Y185_SLICE_X162Y185_D_CY;
  wire [0:0] CLBLM_R_X103Y185_SLICE_X162Y185_D_XOR;
  wire [0:0] CLBLM_R_X103Y185_SLICE_X163Y185_A;
  wire [0:0] CLBLM_R_X103Y185_SLICE_X163Y185_A1;
  wire [0:0] CLBLM_R_X103Y185_SLICE_X163Y185_A2;
  wire [0:0] CLBLM_R_X103Y185_SLICE_X163Y185_A3;
  wire [0:0] CLBLM_R_X103Y185_SLICE_X163Y185_A4;
  wire [0:0] CLBLM_R_X103Y185_SLICE_X163Y185_A5;
  wire [0:0] CLBLM_R_X103Y185_SLICE_X163Y185_A6;
  wire [0:0] CLBLM_R_X103Y185_SLICE_X163Y185_AO5;
  wire [0:0] CLBLM_R_X103Y185_SLICE_X163Y185_AO6;
  wire [0:0] CLBLM_R_X103Y185_SLICE_X163Y185_A_CY;
  wire [0:0] CLBLM_R_X103Y185_SLICE_X163Y185_A_XOR;
  wire [0:0] CLBLM_R_X103Y185_SLICE_X163Y185_B;
  wire [0:0] CLBLM_R_X103Y185_SLICE_X163Y185_B1;
  wire [0:0] CLBLM_R_X103Y185_SLICE_X163Y185_B2;
  wire [0:0] CLBLM_R_X103Y185_SLICE_X163Y185_B3;
  wire [0:0] CLBLM_R_X103Y185_SLICE_X163Y185_B4;
  wire [0:0] CLBLM_R_X103Y185_SLICE_X163Y185_B5;
  wire [0:0] CLBLM_R_X103Y185_SLICE_X163Y185_B6;
  wire [0:0] CLBLM_R_X103Y185_SLICE_X163Y185_BO5;
  wire [0:0] CLBLM_R_X103Y185_SLICE_X163Y185_BO6;
  wire [0:0] CLBLM_R_X103Y185_SLICE_X163Y185_B_CY;
  wire [0:0] CLBLM_R_X103Y185_SLICE_X163Y185_B_XOR;
  wire [0:0] CLBLM_R_X103Y185_SLICE_X163Y185_C;
  wire [0:0] CLBLM_R_X103Y185_SLICE_X163Y185_C1;
  wire [0:0] CLBLM_R_X103Y185_SLICE_X163Y185_C2;
  wire [0:0] CLBLM_R_X103Y185_SLICE_X163Y185_C3;
  wire [0:0] CLBLM_R_X103Y185_SLICE_X163Y185_C4;
  wire [0:0] CLBLM_R_X103Y185_SLICE_X163Y185_C5;
  wire [0:0] CLBLM_R_X103Y185_SLICE_X163Y185_C6;
  wire [0:0] CLBLM_R_X103Y185_SLICE_X163Y185_CO5;
  wire [0:0] CLBLM_R_X103Y185_SLICE_X163Y185_CO6;
  wire [0:0] CLBLM_R_X103Y185_SLICE_X163Y185_C_CY;
  wire [0:0] CLBLM_R_X103Y185_SLICE_X163Y185_C_XOR;
  wire [0:0] CLBLM_R_X103Y185_SLICE_X163Y185_D;
  wire [0:0] CLBLM_R_X103Y185_SLICE_X163Y185_D1;
  wire [0:0] CLBLM_R_X103Y185_SLICE_X163Y185_D2;
  wire [0:0] CLBLM_R_X103Y185_SLICE_X163Y185_D3;
  wire [0:0] CLBLM_R_X103Y185_SLICE_X163Y185_D4;
  wire [0:0] CLBLM_R_X103Y185_SLICE_X163Y185_D5;
  wire [0:0] CLBLM_R_X103Y185_SLICE_X163Y185_D6;
  wire [0:0] CLBLM_R_X103Y185_SLICE_X163Y185_DO5;
  wire [0:0] CLBLM_R_X103Y185_SLICE_X163Y185_DO6;
  wire [0:0] CLBLM_R_X103Y185_SLICE_X163Y185_D_CY;
  wire [0:0] CLBLM_R_X103Y185_SLICE_X163Y185_D_XOR;
  wire [0:0] CLBLM_R_X103Y193_SLICE_X162Y193_A;
  wire [0:0] CLBLM_R_X103Y193_SLICE_X162Y193_A1;
  wire [0:0] CLBLM_R_X103Y193_SLICE_X162Y193_A2;
  wire [0:0] CLBLM_R_X103Y193_SLICE_X162Y193_A3;
  wire [0:0] CLBLM_R_X103Y193_SLICE_X162Y193_A4;
  wire [0:0] CLBLM_R_X103Y193_SLICE_X162Y193_A5;
  wire [0:0] CLBLM_R_X103Y193_SLICE_X162Y193_A6;
  wire [0:0] CLBLM_R_X103Y193_SLICE_X162Y193_AO5;
  wire [0:0] CLBLM_R_X103Y193_SLICE_X162Y193_AO6;
  wire [0:0] CLBLM_R_X103Y193_SLICE_X162Y193_A_CY;
  wire [0:0] CLBLM_R_X103Y193_SLICE_X162Y193_A_XOR;
  wire [0:0] CLBLM_R_X103Y193_SLICE_X162Y193_B;
  wire [0:0] CLBLM_R_X103Y193_SLICE_X162Y193_B1;
  wire [0:0] CLBLM_R_X103Y193_SLICE_X162Y193_B2;
  wire [0:0] CLBLM_R_X103Y193_SLICE_X162Y193_B3;
  wire [0:0] CLBLM_R_X103Y193_SLICE_X162Y193_B4;
  wire [0:0] CLBLM_R_X103Y193_SLICE_X162Y193_B5;
  wire [0:0] CLBLM_R_X103Y193_SLICE_X162Y193_B6;
  wire [0:0] CLBLM_R_X103Y193_SLICE_X162Y193_BO5;
  wire [0:0] CLBLM_R_X103Y193_SLICE_X162Y193_BO6;
  wire [0:0] CLBLM_R_X103Y193_SLICE_X162Y193_B_CY;
  wire [0:0] CLBLM_R_X103Y193_SLICE_X162Y193_B_XOR;
  wire [0:0] CLBLM_R_X103Y193_SLICE_X162Y193_C;
  wire [0:0] CLBLM_R_X103Y193_SLICE_X162Y193_C1;
  wire [0:0] CLBLM_R_X103Y193_SLICE_X162Y193_C2;
  wire [0:0] CLBLM_R_X103Y193_SLICE_X162Y193_C3;
  wire [0:0] CLBLM_R_X103Y193_SLICE_X162Y193_C4;
  wire [0:0] CLBLM_R_X103Y193_SLICE_X162Y193_C5;
  wire [0:0] CLBLM_R_X103Y193_SLICE_X162Y193_C6;
  wire [0:0] CLBLM_R_X103Y193_SLICE_X162Y193_CO5;
  wire [0:0] CLBLM_R_X103Y193_SLICE_X162Y193_CO6;
  wire [0:0] CLBLM_R_X103Y193_SLICE_X162Y193_C_CY;
  wire [0:0] CLBLM_R_X103Y193_SLICE_X162Y193_C_XOR;
  wire [0:0] CLBLM_R_X103Y193_SLICE_X162Y193_D;
  wire [0:0] CLBLM_R_X103Y193_SLICE_X162Y193_D1;
  wire [0:0] CLBLM_R_X103Y193_SLICE_X162Y193_D2;
  wire [0:0] CLBLM_R_X103Y193_SLICE_X162Y193_D3;
  wire [0:0] CLBLM_R_X103Y193_SLICE_X162Y193_D4;
  wire [0:0] CLBLM_R_X103Y193_SLICE_X162Y193_D5;
  wire [0:0] CLBLM_R_X103Y193_SLICE_X162Y193_D6;
  wire [0:0] CLBLM_R_X103Y193_SLICE_X162Y193_DO5;
  wire [0:0] CLBLM_R_X103Y193_SLICE_X162Y193_DO6;
  wire [0:0] CLBLM_R_X103Y193_SLICE_X162Y193_D_CY;
  wire [0:0] CLBLM_R_X103Y193_SLICE_X162Y193_D_XOR;
  wire [0:0] CLBLM_R_X103Y193_SLICE_X163Y193_A;
  wire [0:0] CLBLM_R_X103Y193_SLICE_X163Y193_A1;
  wire [0:0] CLBLM_R_X103Y193_SLICE_X163Y193_A2;
  wire [0:0] CLBLM_R_X103Y193_SLICE_X163Y193_A3;
  wire [0:0] CLBLM_R_X103Y193_SLICE_X163Y193_A4;
  wire [0:0] CLBLM_R_X103Y193_SLICE_X163Y193_A5;
  wire [0:0] CLBLM_R_X103Y193_SLICE_X163Y193_A6;
  wire [0:0] CLBLM_R_X103Y193_SLICE_X163Y193_AO5;
  wire [0:0] CLBLM_R_X103Y193_SLICE_X163Y193_AO6;
  wire [0:0] CLBLM_R_X103Y193_SLICE_X163Y193_A_CY;
  wire [0:0] CLBLM_R_X103Y193_SLICE_X163Y193_A_XOR;
  wire [0:0] CLBLM_R_X103Y193_SLICE_X163Y193_B;
  wire [0:0] CLBLM_R_X103Y193_SLICE_X163Y193_B1;
  wire [0:0] CLBLM_R_X103Y193_SLICE_X163Y193_B2;
  wire [0:0] CLBLM_R_X103Y193_SLICE_X163Y193_B3;
  wire [0:0] CLBLM_R_X103Y193_SLICE_X163Y193_B4;
  wire [0:0] CLBLM_R_X103Y193_SLICE_X163Y193_B5;
  wire [0:0] CLBLM_R_X103Y193_SLICE_X163Y193_B6;
  wire [0:0] CLBLM_R_X103Y193_SLICE_X163Y193_BO5;
  wire [0:0] CLBLM_R_X103Y193_SLICE_X163Y193_BO6;
  wire [0:0] CLBLM_R_X103Y193_SLICE_X163Y193_B_CY;
  wire [0:0] CLBLM_R_X103Y193_SLICE_X163Y193_B_XOR;
  wire [0:0] CLBLM_R_X103Y193_SLICE_X163Y193_C;
  wire [0:0] CLBLM_R_X103Y193_SLICE_X163Y193_C1;
  wire [0:0] CLBLM_R_X103Y193_SLICE_X163Y193_C2;
  wire [0:0] CLBLM_R_X103Y193_SLICE_X163Y193_C3;
  wire [0:0] CLBLM_R_X103Y193_SLICE_X163Y193_C4;
  wire [0:0] CLBLM_R_X103Y193_SLICE_X163Y193_C5;
  wire [0:0] CLBLM_R_X103Y193_SLICE_X163Y193_C6;
  wire [0:0] CLBLM_R_X103Y193_SLICE_X163Y193_CO5;
  wire [0:0] CLBLM_R_X103Y193_SLICE_X163Y193_CO6;
  wire [0:0] CLBLM_R_X103Y193_SLICE_X163Y193_C_CY;
  wire [0:0] CLBLM_R_X103Y193_SLICE_X163Y193_C_XOR;
  wire [0:0] CLBLM_R_X103Y193_SLICE_X163Y193_D;
  wire [0:0] CLBLM_R_X103Y193_SLICE_X163Y193_D1;
  wire [0:0] CLBLM_R_X103Y193_SLICE_X163Y193_D2;
  wire [0:0] CLBLM_R_X103Y193_SLICE_X163Y193_D3;
  wire [0:0] CLBLM_R_X103Y193_SLICE_X163Y193_D4;
  wire [0:0] CLBLM_R_X103Y193_SLICE_X163Y193_D5;
  wire [0:0] CLBLM_R_X103Y193_SLICE_X163Y193_D6;
  wire [0:0] CLBLM_R_X103Y193_SLICE_X163Y193_DO5;
  wire [0:0] CLBLM_R_X103Y193_SLICE_X163Y193_DO6;
  wire [0:0] CLBLM_R_X103Y193_SLICE_X163Y193_D_CY;
  wire [0:0] CLBLM_R_X103Y193_SLICE_X163Y193_D_XOR;
  wire [0:0] CLBLM_R_X103Y97_SLICE_X162Y97_A;
  wire [0:0] CLBLM_R_X103Y97_SLICE_X162Y97_A1;
  wire [0:0] CLBLM_R_X103Y97_SLICE_X162Y97_A2;
  wire [0:0] CLBLM_R_X103Y97_SLICE_X162Y97_A3;
  wire [0:0] CLBLM_R_X103Y97_SLICE_X162Y97_A4;
  wire [0:0] CLBLM_R_X103Y97_SLICE_X162Y97_A5;
  wire [0:0] CLBLM_R_X103Y97_SLICE_X162Y97_A6;
  wire [0:0] CLBLM_R_X103Y97_SLICE_X162Y97_AO5;
  wire [0:0] CLBLM_R_X103Y97_SLICE_X162Y97_AO6;
  wire [0:0] CLBLM_R_X103Y97_SLICE_X162Y97_A_CY;
  wire [0:0] CLBLM_R_X103Y97_SLICE_X162Y97_A_XOR;
  wire [0:0] CLBLM_R_X103Y97_SLICE_X162Y97_B;
  wire [0:0] CLBLM_R_X103Y97_SLICE_X162Y97_B1;
  wire [0:0] CLBLM_R_X103Y97_SLICE_X162Y97_B2;
  wire [0:0] CLBLM_R_X103Y97_SLICE_X162Y97_B3;
  wire [0:0] CLBLM_R_X103Y97_SLICE_X162Y97_B4;
  wire [0:0] CLBLM_R_X103Y97_SLICE_X162Y97_B5;
  wire [0:0] CLBLM_R_X103Y97_SLICE_X162Y97_B6;
  wire [0:0] CLBLM_R_X103Y97_SLICE_X162Y97_BO5;
  wire [0:0] CLBLM_R_X103Y97_SLICE_X162Y97_BO6;
  wire [0:0] CLBLM_R_X103Y97_SLICE_X162Y97_B_CY;
  wire [0:0] CLBLM_R_X103Y97_SLICE_X162Y97_B_XOR;
  wire [0:0] CLBLM_R_X103Y97_SLICE_X162Y97_C;
  wire [0:0] CLBLM_R_X103Y97_SLICE_X162Y97_C1;
  wire [0:0] CLBLM_R_X103Y97_SLICE_X162Y97_C2;
  wire [0:0] CLBLM_R_X103Y97_SLICE_X162Y97_C3;
  wire [0:0] CLBLM_R_X103Y97_SLICE_X162Y97_C4;
  wire [0:0] CLBLM_R_X103Y97_SLICE_X162Y97_C5;
  wire [0:0] CLBLM_R_X103Y97_SLICE_X162Y97_C6;
  wire [0:0] CLBLM_R_X103Y97_SLICE_X162Y97_CO5;
  wire [0:0] CLBLM_R_X103Y97_SLICE_X162Y97_CO6;
  wire [0:0] CLBLM_R_X103Y97_SLICE_X162Y97_C_CY;
  wire [0:0] CLBLM_R_X103Y97_SLICE_X162Y97_C_XOR;
  wire [0:0] CLBLM_R_X103Y97_SLICE_X162Y97_D;
  wire [0:0] CLBLM_R_X103Y97_SLICE_X162Y97_D1;
  wire [0:0] CLBLM_R_X103Y97_SLICE_X162Y97_D2;
  wire [0:0] CLBLM_R_X103Y97_SLICE_X162Y97_D3;
  wire [0:0] CLBLM_R_X103Y97_SLICE_X162Y97_D4;
  wire [0:0] CLBLM_R_X103Y97_SLICE_X162Y97_D5;
  wire [0:0] CLBLM_R_X103Y97_SLICE_X162Y97_D6;
  wire [0:0] CLBLM_R_X103Y97_SLICE_X162Y97_DO5;
  wire [0:0] CLBLM_R_X103Y97_SLICE_X162Y97_DO6;
  wire [0:0] CLBLM_R_X103Y97_SLICE_X162Y97_D_CY;
  wire [0:0] CLBLM_R_X103Y97_SLICE_X162Y97_D_XOR;
  wire [0:0] CLBLM_R_X103Y97_SLICE_X163Y97_A;
  wire [0:0] CLBLM_R_X103Y97_SLICE_X163Y97_A1;
  wire [0:0] CLBLM_R_X103Y97_SLICE_X163Y97_A2;
  wire [0:0] CLBLM_R_X103Y97_SLICE_X163Y97_A3;
  wire [0:0] CLBLM_R_X103Y97_SLICE_X163Y97_A4;
  wire [0:0] CLBLM_R_X103Y97_SLICE_X163Y97_A5;
  wire [0:0] CLBLM_R_X103Y97_SLICE_X163Y97_A6;
  wire [0:0] CLBLM_R_X103Y97_SLICE_X163Y97_AO5;
  wire [0:0] CLBLM_R_X103Y97_SLICE_X163Y97_AO6;
  wire [0:0] CLBLM_R_X103Y97_SLICE_X163Y97_A_CY;
  wire [0:0] CLBLM_R_X103Y97_SLICE_X163Y97_A_XOR;
  wire [0:0] CLBLM_R_X103Y97_SLICE_X163Y97_B;
  wire [0:0] CLBLM_R_X103Y97_SLICE_X163Y97_B1;
  wire [0:0] CLBLM_R_X103Y97_SLICE_X163Y97_B2;
  wire [0:0] CLBLM_R_X103Y97_SLICE_X163Y97_B3;
  wire [0:0] CLBLM_R_X103Y97_SLICE_X163Y97_B4;
  wire [0:0] CLBLM_R_X103Y97_SLICE_X163Y97_B5;
  wire [0:0] CLBLM_R_X103Y97_SLICE_X163Y97_B6;
  wire [0:0] CLBLM_R_X103Y97_SLICE_X163Y97_BO5;
  wire [0:0] CLBLM_R_X103Y97_SLICE_X163Y97_BO6;
  wire [0:0] CLBLM_R_X103Y97_SLICE_X163Y97_B_CY;
  wire [0:0] CLBLM_R_X103Y97_SLICE_X163Y97_B_XOR;
  wire [0:0] CLBLM_R_X103Y97_SLICE_X163Y97_C;
  wire [0:0] CLBLM_R_X103Y97_SLICE_X163Y97_C1;
  wire [0:0] CLBLM_R_X103Y97_SLICE_X163Y97_C2;
  wire [0:0] CLBLM_R_X103Y97_SLICE_X163Y97_C3;
  wire [0:0] CLBLM_R_X103Y97_SLICE_X163Y97_C4;
  wire [0:0] CLBLM_R_X103Y97_SLICE_X163Y97_C5;
  wire [0:0] CLBLM_R_X103Y97_SLICE_X163Y97_C6;
  wire [0:0] CLBLM_R_X103Y97_SLICE_X163Y97_CO5;
  wire [0:0] CLBLM_R_X103Y97_SLICE_X163Y97_CO6;
  wire [0:0] CLBLM_R_X103Y97_SLICE_X163Y97_C_CY;
  wire [0:0] CLBLM_R_X103Y97_SLICE_X163Y97_C_XOR;
  wire [0:0] CLBLM_R_X103Y97_SLICE_X163Y97_D;
  wire [0:0] CLBLM_R_X103Y97_SLICE_X163Y97_D1;
  wire [0:0] CLBLM_R_X103Y97_SLICE_X163Y97_D2;
  wire [0:0] CLBLM_R_X103Y97_SLICE_X163Y97_D3;
  wire [0:0] CLBLM_R_X103Y97_SLICE_X163Y97_D4;
  wire [0:0] CLBLM_R_X103Y97_SLICE_X163Y97_D5;
  wire [0:0] CLBLM_R_X103Y97_SLICE_X163Y97_D6;
  wire [0:0] CLBLM_R_X103Y97_SLICE_X163Y97_DO5;
  wire [0:0] CLBLM_R_X103Y97_SLICE_X163Y97_DO6;
  wire [0:0] CLBLM_R_X103Y97_SLICE_X163Y97_D_CY;
  wire [0:0] CLBLM_R_X103Y97_SLICE_X163Y97_D_XOR;
  wire [0:0] CLBLM_R_X25Y115_SLICE_X36Y115_A;
  wire [0:0] CLBLM_R_X25Y115_SLICE_X36Y115_A1;
  wire [0:0] CLBLM_R_X25Y115_SLICE_X36Y115_A2;
  wire [0:0] CLBLM_R_X25Y115_SLICE_X36Y115_A3;
  wire [0:0] CLBLM_R_X25Y115_SLICE_X36Y115_A4;
  wire [0:0] CLBLM_R_X25Y115_SLICE_X36Y115_A5;
  wire [0:0] CLBLM_R_X25Y115_SLICE_X36Y115_A6;
  wire [0:0] CLBLM_R_X25Y115_SLICE_X36Y115_AMUX;
  wire [0:0] CLBLM_R_X25Y115_SLICE_X36Y115_AO5;
  wire [0:0] CLBLM_R_X25Y115_SLICE_X36Y115_AO6;
  wire [0:0] CLBLM_R_X25Y115_SLICE_X36Y115_A_CY;
  wire [0:0] CLBLM_R_X25Y115_SLICE_X36Y115_A_XOR;
  wire [0:0] CLBLM_R_X25Y115_SLICE_X36Y115_B;
  wire [0:0] CLBLM_R_X25Y115_SLICE_X36Y115_B1;
  wire [0:0] CLBLM_R_X25Y115_SLICE_X36Y115_B2;
  wire [0:0] CLBLM_R_X25Y115_SLICE_X36Y115_B3;
  wire [0:0] CLBLM_R_X25Y115_SLICE_X36Y115_B4;
  wire [0:0] CLBLM_R_X25Y115_SLICE_X36Y115_B5;
  wire [0:0] CLBLM_R_X25Y115_SLICE_X36Y115_B6;
  wire [0:0] CLBLM_R_X25Y115_SLICE_X36Y115_BO5;
  wire [0:0] CLBLM_R_X25Y115_SLICE_X36Y115_BO6;
  wire [0:0] CLBLM_R_X25Y115_SLICE_X36Y115_B_CY;
  wire [0:0] CLBLM_R_X25Y115_SLICE_X36Y115_B_XOR;
  wire [0:0] CLBLM_R_X25Y115_SLICE_X36Y115_C;
  wire [0:0] CLBLM_R_X25Y115_SLICE_X36Y115_C1;
  wire [0:0] CLBLM_R_X25Y115_SLICE_X36Y115_C2;
  wire [0:0] CLBLM_R_X25Y115_SLICE_X36Y115_C3;
  wire [0:0] CLBLM_R_X25Y115_SLICE_X36Y115_C4;
  wire [0:0] CLBLM_R_X25Y115_SLICE_X36Y115_C5;
  wire [0:0] CLBLM_R_X25Y115_SLICE_X36Y115_C6;
  wire [0:0] CLBLM_R_X25Y115_SLICE_X36Y115_CO5;
  wire [0:0] CLBLM_R_X25Y115_SLICE_X36Y115_CO6;
  wire [0:0] CLBLM_R_X25Y115_SLICE_X36Y115_C_CY;
  wire [0:0] CLBLM_R_X25Y115_SLICE_X36Y115_C_XOR;
  wire [0:0] CLBLM_R_X25Y115_SLICE_X36Y115_D;
  wire [0:0] CLBLM_R_X25Y115_SLICE_X36Y115_D1;
  wire [0:0] CLBLM_R_X25Y115_SLICE_X36Y115_D2;
  wire [0:0] CLBLM_R_X25Y115_SLICE_X36Y115_D3;
  wire [0:0] CLBLM_R_X25Y115_SLICE_X36Y115_D4;
  wire [0:0] CLBLM_R_X25Y115_SLICE_X36Y115_D5;
  wire [0:0] CLBLM_R_X25Y115_SLICE_X36Y115_D6;
  wire [0:0] CLBLM_R_X25Y115_SLICE_X36Y115_DO5;
  wire [0:0] CLBLM_R_X25Y115_SLICE_X36Y115_DO6;
  wire [0:0] CLBLM_R_X25Y115_SLICE_X36Y115_D_CY;
  wire [0:0] CLBLM_R_X25Y115_SLICE_X36Y115_D_XOR;
  wire [0:0] CLBLM_R_X25Y115_SLICE_X37Y115_A;
  wire [0:0] CLBLM_R_X25Y115_SLICE_X37Y115_A1;
  wire [0:0] CLBLM_R_X25Y115_SLICE_X37Y115_A2;
  wire [0:0] CLBLM_R_X25Y115_SLICE_X37Y115_A3;
  wire [0:0] CLBLM_R_X25Y115_SLICE_X37Y115_A4;
  wire [0:0] CLBLM_R_X25Y115_SLICE_X37Y115_A5;
  wire [0:0] CLBLM_R_X25Y115_SLICE_X37Y115_A6;
  wire [0:0] CLBLM_R_X25Y115_SLICE_X37Y115_AO5;
  wire [0:0] CLBLM_R_X25Y115_SLICE_X37Y115_AO6;
  wire [0:0] CLBLM_R_X25Y115_SLICE_X37Y115_A_CY;
  wire [0:0] CLBLM_R_X25Y115_SLICE_X37Y115_A_XOR;
  wire [0:0] CLBLM_R_X25Y115_SLICE_X37Y115_B;
  wire [0:0] CLBLM_R_X25Y115_SLICE_X37Y115_B1;
  wire [0:0] CLBLM_R_X25Y115_SLICE_X37Y115_B2;
  wire [0:0] CLBLM_R_X25Y115_SLICE_X37Y115_B3;
  wire [0:0] CLBLM_R_X25Y115_SLICE_X37Y115_B4;
  wire [0:0] CLBLM_R_X25Y115_SLICE_X37Y115_B5;
  wire [0:0] CLBLM_R_X25Y115_SLICE_X37Y115_B6;
  wire [0:0] CLBLM_R_X25Y115_SLICE_X37Y115_BO5;
  wire [0:0] CLBLM_R_X25Y115_SLICE_X37Y115_BO6;
  wire [0:0] CLBLM_R_X25Y115_SLICE_X37Y115_B_CY;
  wire [0:0] CLBLM_R_X25Y115_SLICE_X37Y115_B_XOR;
  wire [0:0] CLBLM_R_X25Y115_SLICE_X37Y115_C;
  wire [0:0] CLBLM_R_X25Y115_SLICE_X37Y115_C1;
  wire [0:0] CLBLM_R_X25Y115_SLICE_X37Y115_C2;
  wire [0:0] CLBLM_R_X25Y115_SLICE_X37Y115_C3;
  wire [0:0] CLBLM_R_X25Y115_SLICE_X37Y115_C4;
  wire [0:0] CLBLM_R_X25Y115_SLICE_X37Y115_C5;
  wire [0:0] CLBLM_R_X25Y115_SLICE_X37Y115_C6;
  wire [0:0] CLBLM_R_X25Y115_SLICE_X37Y115_CO5;
  wire [0:0] CLBLM_R_X25Y115_SLICE_X37Y115_CO6;
  wire [0:0] CLBLM_R_X25Y115_SLICE_X37Y115_C_CY;
  wire [0:0] CLBLM_R_X25Y115_SLICE_X37Y115_C_XOR;
  wire [0:0] CLBLM_R_X25Y115_SLICE_X37Y115_D;
  wire [0:0] CLBLM_R_X25Y115_SLICE_X37Y115_D1;
  wire [0:0] CLBLM_R_X25Y115_SLICE_X37Y115_D2;
  wire [0:0] CLBLM_R_X25Y115_SLICE_X37Y115_D3;
  wire [0:0] CLBLM_R_X25Y115_SLICE_X37Y115_D4;
  wire [0:0] CLBLM_R_X25Y115_SLICE_X37Y115_D5;
  wire [0:0] CLBLM_R_X25Y115_SLICE_X37Y115_D6;
  wire [0:0] CLBLM_R_X25Y115_SLICE_X37Y115_DO5;
  wire [0:0] CLBLM_R_X25Y115_SLICE_X37Y115_DO6;
  wire [0:0] CLBLM_R_X25Y115_SLICE_X37Y115_D_CY;
  wire [0:0] CLBLM_R_X25Y115_SLICE_X37Y115_D_XOR;
  wire [0:0] CLBLM_R_X25Y116_SLICE_X36Y116_A;
  wire [0:0] CLBLM_R_X25Y116_SLICE_X36Y116_A1;
  wire [0:0] CLBLM_R_X25Y116_SLICE_X36Y116_A2;
  wire [0:0] CLBLM_R_X25Y116_SLICE_X36Y116_A3;
  wire [0:0] CLBLM_R_X25Y116_SLICE_X36Y116_A4;
  wire [0:0] CLBLM_R_X25Y116_SLICE_X36Y116_A5;
  wire [0:0] CLBLM_R_X25Y116_SLICE_X36Y116_A6;
  wire [0:0] CLBLM_R_X25Y116_SLICE_X36Y116_AMUX;
  wire [0:0] CLBLM_R_X25Y116_SLICE_X36Y116_AO5;
  wire [0:0] CLBLM_R_X25Y116_SLICE_X36Y116_AO6;
  wire [0:0] CLBLM_R_X25Y116_SLICE_X36Y116_A_CY;
  wire [0:0] CLBLM_R_X25Y116_SLICE_X36Y116_A_XOR;
  wire [0:0] CLBLM_R_X25Y116_SLICE_X36Y116_B;
  wire [0:0] CLBLM_R_X25Y116_SLICE_X36Y116_B1;
  wire [0:0] CLBLM_R_X25Y116_SLICE_X36Y116_B2;
  wire [0:0] CLBLM_R_X25Y116_SLICE_X36Y116_B3;
  wire [0:0] CLBLM_R_X25Y116_SLICE_X36Y116_B4;
  wire [0:0] CLBLM_R_X25Y116_SLICE_X36Y116_B5;
  wire [0:0] CLBLM_R_X25Y116_SLICE_X36Y116_B6;
  wire [0:0] CLBLM_R_X25Y116_SLICE_X36Y116_BO5;
  wire [0:0] CLBLM_R_X25Y116_SLICE_X36Y116_BO6;
  wire [0:0] CLBLM_R_X25Y116_SLICE_X36Y116_B_CY;
  wire [0:0] CLBLM_R_X25Y116_SLICE_X36Y116_B_XOR;
  wire [0:0] CLBLM_R_X25Y116_SLICE_X36Y116_C;
  wire [0:0] CLBLM_R_X25Y116_SLICE_X36Y116_C1;
  wire [0:0] CLBLM_R_X25Y116_SLICE_X36Y116_C2;
  wire [0:0] CLBLM_R_X25Y116_SLICE_X36Y116_C3;
  wire [0:0] CLBLM_R_X25Y116_SLICE_X36Y116_C4;
  wire [0:0] CLBLM_R_X25Y116_SLICE_X36Y116_C5;
  wire [0:0] CLBLM_R_X25Y116_SLICE_X36Y116_C6;
  wire [0:0] CLBLM_R_X25Y116_SLICE_X36Y116_CO5;
  wire [0:0] CLBLM_R_X25Y116_SLICE_X36Y116_CO6;
  wire [0:0] CLBLM_R_X25Y116_SLICE_X36Y116_C_CY;
  wire [0:0] CLBLM_R_X25Y116_SLICE_X36Y116_C_XOR;
  wire [0:0] CLBLM_R_X25Y116_SLICE_X36Y116_D;
  wire [0:0] CLBLM_R_X25Y116_SLICE_X36Y116_D1;
  wire [0:0] CLBLM_R_X25Y116_SLICE_X36Y116_D2;
  wire [0:0] CLBLM_R_X25Y116_SLICE_X36Y116_D3;
  wire [0:0] CLBLM_R_X25Y116_SLICE_X36Y116_D4;
  wire [0:0] CLBLM_R_X25Y116_SLICE_X36Y116_D5;
  wire [0:0] CLBLM_R_X25Y116_SLICE_X36Y116_D6;
  wire [0:0] CLBLM_R_X25Y116_SLICE_X36Y116_DO5;
  wire [0:0] CLBLM_R_X25Y116_SLICE_X36Y116_DO6;
  wire [0:0] CLBLM_R_X25Y116_SLICE_X36Y116_D_CY;
  wire [0:0] CLBLM_R_X25Y116_SLICE_X36Y116_D_XOR;
  wire [0:0] CLBLM_R_X25Y116_SLICE_X37Y116_A;
  wire [0:0] CLBLM_R_X25Y116_SLICE_X37Y116_A1;
  wire [0:0] CLBLM_R_X25Y116_SLICE_X37Y116_A2;
  wire [0:0] CLBLM_R_X25Y116_SLICE_X37Y116_A3;
  wire [0:0] CLBLM_R_X25Y116_SLICE_X37Y116_A4;
  wire [0:0] CLBLM_R_X25Y116_SLICE_X37Y116_A5;
  wire [0:0] CLBLM_R_X25Y116_SLICE_X37Y116_A6;
  wire [0:0] CLBLM_R_X25Y116_SLICE_X37Y116_AO5;
  wire [0:0] CLBLM_R_X25Y116_SLICE_X37Y116_AO6;
  wire [0:0] CLBLM_R_X25Y116_SLICE_X37Y116_A_CY;
  wire [0:0] CLBLM_R_X25Y116_SLICE_X37Y116_A_XOR;
  wire [0:0] CLBLM_R_X25Y116_SLICE_X37Y116_B;
  wire [0:0] CLBLM_R_X25Y116_SLICE_X37Y116_B1;
  wire [0:0] CLBLM_R_X25Y116_SLICE_X37Y116_B2;
  wire [0:0] CLBLM_R_X25Y116_SLICE_X37Y116_B3;
  wire [0:0] CLBLM_R_X25Y116_SLICE_X37Y116_B4;
  wire [0:0] CLBLM_R_X25Y116_SLICE_X37Y116_B5;
  wire [0:0] CLBLM_R_X25Y116_SLICE_X37Y116_B6;
  wire [0:0] CLBLM_R_X25Y116_SLICE_X37Y116_BO5;
  wire [0:0] CLBLM_R_X25Y116_SLICE_X37Y116_BO6;
  wire [0:0] CLBLM_R_X25Y116_SLICE_X37Y116_B_CY;
  wire [0:0] CLBLM_R_X25Y116_SLICE_X37Y116_B_XOR;
  wire [0:0] CLBLM_R_X25Y116_SLICE_X37Y116_C;
  wire [0:0] CLBLM_R_X25Y116_SLICE_X37Y116_C1;
  wire [0:0] CLBLM_R_X25Y116_SLICE_X37Y116_C2;
  wire [0:0] CLBLM_R_X25Y116_SLICE_X37Y116_C3;
  wire [0:0] CLBLM_R_X25Y116_SLICE_X37Y116_C4;
  wire [0:0] CLBLM_R_X25Y116_SLICE_X37Y116_C5;
  wire [0:0] CLBLM_R_X25Y116_SLICE_X37Y116_C6;
  wire [0:0] CLBLM_R_X25Y116_SLICE_X37Y116_CO5;
  wire [0:0] CLBLM_R_X25Y116_SLICE_X37Y116_CO6;
  wire [0:0] CLBLM_R_X25Y116_SLICE_X37Y116_C_CY;
  wire [0:0] CLBLM_R_X25Y116_SLICE_X37Y116_C_XOR;
  wire [0:0] CLBLM_R_X25Y116_SLICE_X37Y116_D;
  wire [0:0] CLBLM_R_X25Y116_SLICE_X37Y116_D1;
  wire [0:0] CLBLM_R_X25Y116_SLICE_X37Y116_D2;
  wire [0:0] CLBLM_R_X25Y116_SLICE_X37Y116_D3;
  wire [0:0] CLBLM_R_X25Y116_SLICE_X37Y116_D4;
  wire [0:0] CLBLM_R_X25Y116_SLICE_X37Y116_D5;
  wire [0:0] CLBLM_R_X25Y116_SLICE_X37Y116_D6;
  wire [0:0] CLBLM_R_X25Y116_SLICE_X37Y116_DO5;
  wire [0:0] CLBLM_R_X25Y116_SLICE_X37Y116_DO6;
  wire [0:0] CLBLM_R_X25Y116_SLICE_X37Y116_D_CY;
  wire [0:0] CLBLM_R_X25Y116_SLICE_X37Y116_D_XOR;
  wire [0:0] CLBLM_R_X29Y115_SLICE_X42Y115_A;
  wire [0:0] CLBLM_R_X29Y115_SLICE_X42Y115_A1;
  wire [0:0] CLBLM_R_X29Y115_SLICE_X42Y115_A2;
  wire [0:0] CLBLM_R_X29Y115_SLICE_X42Y115_A3;
  wire [0:0] CLBLM_R_X29Y115_SLICE_X42Y115_A4;
  wire [0:0] CLBLM_R_X29Y115_SLICE_X42Y115_A5;
  wire [0:0] CLBLM_R_X29Y115_SLICE_X42Y115_A6;
  wire [0:0] CLBLM_R_X29Y115_SLICE_X42Y115_AO5;
  wire [0:0] CLBLM_R_X29Y115_SLICE_X42Y115_AO6;
  wire [0:0] CLBLM_R_X29Y115_SLICE_X42Y115_A_CY;
  wire [0:0] CLBLM_R_X29Y115_SLICE_X42Y115_A_XOR;
  wire [0:0] CLBLM_R_X29Y115_SLICE_X42Y115_B;
  wire [0:0] CLBLM_R_X29Y115_SLICE_X42Y115_B1;
  wire [0:0] CLBLM_R_X29Y115_SLICE_X42Y115_B2;
  wire [0:0] CLBLM_R_X29Y115_SLICE_X42Y115_B3;
  wire [0:0] CLBLM_R_X29Y115_SLICE_X42Y115_B4;
  wire [0:0] CLBLM_R_X29Y115_SLICE_X42Y115_B5;
  wire [0:0] CLBLM_R_X29Y115_SLICE_X42Y115_B6;
  wire [0:0] CLBLM_R_X29Y115_SLICE_X42Y115_BO5;
  wire [0:0] CLBLM_R_X29Y115_SLICE_X42Y115_BO6;
  wire [0:0] CLBLM_R_X29Y115_SLICE_X42Y115_B_CY;
  wire [0:0] CLBLM_R_X29Y115_SLICE_X42Y115_B_XOR;
  wire [0:0] CLBLM_R_X29Y115_SLICE_X42Y115_C;
  wire [0:0] CLBLM_R_X29Y115_SLICE_X42Y115_C1;
  wire [0:0] CLBLM_R_X29Y115_SLICE_X42Y115_C2;
  wire [0:0] CLBLM_R_X29Y115_SLICE_X42Y115_C3;
  wire [0:0] CLBLM_R_X29Y115_SLICE_X42Y115_C4;
  wire [0:0] CLBLM_R_X29Y115_SLICE_X42Y115_C5;
  wire [0:0] CLBLM_R_X29Y115_SLICE_X42Y115_C6;
  wire [0:0] CLBLM_R_X29Y115_SLICE_X42Y115_CO5;
  wire [0:0] CLBLM_R_X29Y115_SLICE_X42Y115_CO6;
  wire [0:0] CLBLM_R_X29Y115_SLICE_X42Y115_C_CY;
  wire [0:0] CLBLM_R_X29Y115_SLICE_X42Y115_C_XOR;
  wire [0:0] CLBLM_R_X29Y115_SLICE_X42Y115_D;
  wire [0:0] CLBLM_R_X29Y115_SLICE_X42Y115_D1;
  wire [0:0] CLBLM_R_X29Y115_SLICE_X42Y115_D2;
  wire [0:0] CLBLM_R_X29Y115_SLICE_X42Y115_D3;
  wire [0:0] CLBLM_R_X29Y115_SLICE_X42Y115_D4;
  wire [0:0] CLBLM_R_X29Y115_SLICE_X42Y115_D5;
  wire [0:0] CLBLM_R_X29Y115_SLICE_X42Y115_D6;
  wire [0:0] CLBLM_R_X29Y115_SLICE_X42Y115_DO5;
  wire [0:0] CLBLM_R_X29Y115_SLICE_X42Y115_DO6;
  wire [0:0] CLBLM_R_X29Y115_SLICE_X42Y115_D_CY;
  wire [0:0] CLBLM_R_X29Y115_SLICE_X42Y115_D_XOR;
  wire [0:0] CLBLM_R_X29Y115_SLICE_X43Y115_A;
  wire [0:0] CLBLM_R_X29Y115_SLICE_X43Y115_A1;
  wire [0:0] CLBLM_R_X29Y115_SLICE_X43Y115_A2;
  wire [0:0] CLBLM_R_X29Y115_SLICE_X43Y115_A3;
  wire [0:0] CLBLM_R_X29Y115_SLICE_X43Y115_A4;
  wire [0:0] CLBLM_R_X29Y115_SLICE_X43Y115_A5;
  wire [0:0] CLBLM_R_X29Y115_SLICE_X43Y115_A6;
  wire [0:0] CLBLM_R_X29Y115_SLICE_X43Y115_AO5;
  wire [0:0] CLBLM_R_X29Y115_SLICE_X43Y115_AO6;
  wire [0:0] CLBLM_R_X29Y115_SLICE_X43Y115_A_CY;
  wire [0:0] CLBLM_R_X29Y115_SLICE_X43Y115_A_XOR;
  wire [0:0] CLBLM_R_X29Y115_SLICE_X43Y115_B;
  wire [0:0] CLBLM_R_X29Y115_SLICE_X43Y115_B1;
  wire [0:0] CLBLM_R_X29Y115_SLICE_X43Y115_B2;
  wire [0:0] CLBLM_R_X29Y115_SLICE_X43Y115_B3;
  wire [0:0] CLBLM_R_X29Y115_SLICE_X43Y115_B4;
  wire [0:0] CLBLM_R_X29Y115_SLICE_X43Y115_B5;
  wire [0:0] CLBLM_R_X29Y115_SLICE_X43Y115_B6;
  wire [0:0] CLBLM_R_X29Y115_SLICE_X43Y115_BO5;
  wire [0:0] CLBLM_R_X29Y115_SLICE_X43Y115_BO6;
  wire [0:0] CLBLM_R_X29Y115_SLICE_X43Y115_B_CY;
  wire [0:0] CLBLM_R_X29Y115_SLICE_X43Y115_B_XOR;
  wire [0:0] CLBLM_R_X29Y115_SLICE_X43Y115_C;
  wire [0:0] CLBLM_R_X29Y115_SLICE_X43Y115_C1;
  wire [0:0] CLBLM_R_X29Y115_SLICE_X43Y115_C2;
  wire [0:0] CLBLM_R_X29Y115_SLICE_X43Y115_C3;
  wire [0:0] CLBLM_R_X29Y115_SLICE_X43Y115_C4;
  wire [0:0] CLBLM_R_X29Y115_SLICE_X43Y115_C5;
  wire [0:0] CLBLM_R_X29Y115_SLICE_X43Y115_C6;
  wire [0:0] CLBLM_R_X29Y115_SLICE_X43Y115_CO5;
  wire [0:0] CLBLM_R_X29Y115_SLICE_X43Y115_CO6;
  wire [0:0] CLBLM_R_X29Y115_SLICE_X43Y115_C_CY;
  wire [0:0] CLBLM_R_X29Y115_SLICE_X43Y115_C_XOR;
  wire [0:0] CLBLM_R_X29Y115_SLICE_X43Y115_D;
  wire [0:0] CLBLM_R_X29Y115_SLICE_X43Y115_D1;
  wire [0:0] CLBLM_R_X29Y115_SLICE_X43Y115_D2;
  wire [0:0] CLBLM_R_X29Y115_SLICE_X43Y115_D3;
  wire [0:0] CLBLM_R_X29Y115_SLICE_X43Y115_D4;
  wire [0:0] CLBLM_R_X29Y115_SLICE_X43Y115_D5;
  wire [0:0] CLBLM_R_X29Y115_SLICE_X43Y115_D6;
  wire [0:0] CLBLM_R_X29Y115_SLICE_X43Y115_DO5;
  wire [0:0] CLBLM_R_X29Y115_SLICE_X43Y115_DO6;
  wire [0:0] CLBLM_R_X29Y115_SLICE_X43Y115_D_CY;
  wire [0:0] CLBLM_R_X29Y115_SLICE_X43Y115_D_XOR;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X2Y110_A;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X2Y110_A1;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X2Y110_A2;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X2Y110_A3;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X2Y110_A4;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X2Y110_A5;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X2Y110_A6;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X2Y110_AO5;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X2Y110_AO6;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X2Y110_A_CY;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X2Y110_A_XOR;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X2Y110_B;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X2Y110_B1;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X2Y110_B2;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X2Y110_B3;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X2Y110_B4;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X2Y110_B5;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X2Y110_B6;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X2Y110_BO5;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X2Y110_BO6;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X2Y110_B_CY;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X2Y110_B_XOR;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X2Y110_C;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X2Y110_C1;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X2Y110_C2;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X2Y110_C3;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X2Y110_C4;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X2Y110_C5;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X2Y110_C6;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X2Y110_CO5;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X2Y110_CO6;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X2Y110_C_CY;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X2Y110_C_XOR;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X2Y110_D;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X2Y110_D1;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X2Y110_D2;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X2Y110_D3;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X2Y110_D4;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X2Y110_D5;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X2Y110_D6;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X2Y110_DO5;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X2Y110_DO6;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X2Y110_D_CY;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X2Y110_D_XOR;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X3Y110_A;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X3Y110_A1;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X3Y110_A2;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X3Y110_A3;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X3Y110_A4;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X3Y110_A5;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X3Y110_A6;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X3Y110_AMUX;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X3Y110_AO5;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X3Y110_AO6;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X3Y110_A_CY;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X3Y110_A_XOR;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X3Y110_B;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X3Y110_B1;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X3Y110_B2;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X3Y110_B3;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X3Y110_B4;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X3Y110_B5;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X3Y110_B6;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X3Y110_BO5;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X3Y110_BO6;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X3Y110_B_CY;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X3Y110_B_XOR;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X3Y110_C;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X3Y110_C1;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X3Y110_C2;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X3Y110_C3;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X3Y110_C4;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X3Y110_C5;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X3Y110_C6;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X3Y110_CO5;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X3Y110_CO6;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X3Y110_C_CY;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X3Y110_C_XOR;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X3Y110_D;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X3Y110_D1;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X3Y110_D2;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X3Y110_D3;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X3Y110_D4;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X3Y110_D5;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X3Y110_D6;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X3Y110_DO5;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X3Y110_DO6;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X3Y110_D_CY;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X3Y110_D_XOR;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X2Y111_A;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X2Y111_A1;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X2Y111_A2;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X2Y111_A3;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X2Y111_A4;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X2Y111_A5;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X2Y111_A6;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X2Y111_AMUX;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X2Y111_AO5;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X2Y111_AO6;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X2Y111_A_CY;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X2Y111_A_XOR;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X2Y111_B;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X2Y111_B1;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X2Y111_B2;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X2Y111_B3;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X2Y111_B4;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X2Y111_B5;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X2Y111_B6;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X2Y111_BO5;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X2Y111_BO6;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X2Y111_B_CY;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X2Y111_B_XOR;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X2Y111_C;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X2Y111_C1;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X2Y111_C2;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X2Y111_C3;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X2Y111_C4;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X2Y111_C5;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X2Y111_C6;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X2Y111_CO5;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X2Y111_CO6;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X2Y111_C_CY;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X2Y111_C_XOR;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X2Y111_D;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X2Y111_D1;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X2Y111_D2;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X2Y111_D3;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X2Y111_D4;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X2Y111_D5;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X2Y111_D6;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X2Y111_DO5;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X2Y111_DO6;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X2Y111_D_CY;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X2Y111_D_XOR;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X3Y111_A;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X3Y111_A1;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X3Y111_A2;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X3Y111_A3;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X3Y111_A4;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X3Y111_A5;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X3Y111_A6;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X3Y111_AMUX;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X3Y111_AO5;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X3Y111_AO6;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X3Y111_A_CY;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X3Y111_A_XOR;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X3Y111_B;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X3Y111_B1;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X3Y111_B2;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X3Y111_B3;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X3Y111_B4;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X3Y111_B5;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X3Y111_B6;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X3Y111_BMUX;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X3Y111_BO5;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X3Y111_BO6;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X3Y111_B_CY;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X3Y111_B_XOR;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X3Y111_C;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X3Y111_C1;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X3Y111_C2;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X3Y111_C3;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X3Y111_C4;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X3Y111_C5;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X3Y111_C6;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X3Y111_CMUX;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X3Y111_CO5;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X3Y111_CO6;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X3Y111_C_CY;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X3Y111_C_XOR;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X3Y111_D;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X3Y111_D1;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X3Y111_D2;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X3Y111_D3;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X3Y111_D4;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X3Y111_D5;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X3Y111_D6;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X3Y111_DMUX;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X3Y111_DO5;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X3Y111_DO6;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X3Y111_D_CY;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X3Y111_D_XOR;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X2Y112_A;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X2Y112_A1;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X2Y112_A2;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X2Y112_A3;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X2Y112_A4;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X2Y112_A5;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X2Y112_A6;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X2Y112_AO5;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X2Y112_AO6;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X2Y112_A_CY;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X2Y112_A_XOR;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X2Y112_B;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X2Y112_B1;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X2Y112_B2;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X2Y112_B3;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X2Y112_B4;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X2Y112_B5;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X2Y112_B6;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X2Y112_BO5;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X2Y112_BO6;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X2Y112_B_CY;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X2Y112_B_XOR;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X2Y112_C;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X2Y112_C1;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X2Y112_C2;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X2Y112_C3;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X2Y112_C4;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X2Y112_C5;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X2Y112_C6;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X2Y112_CO5;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X2Y112_CO6;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X2Y112_C_CY;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X2Y112_C_XOR;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X2Y112_D;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X2Y112_D1;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X2Y112_D2;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X2Y112_D3;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X2Y112_D4;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X2Y112_D5;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X2Y112_D6;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X2Y112_DO5;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X2Y112_DO6;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X2Y112_D_CY;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X2Y112_D_XOR;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X3Y112_A;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X3Y112_A1;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X3Y112_A2;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X3Y112_A3;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X3Y112_A4;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X3Y112_A5;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X3Y112_A6;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X3Y112_AMUX;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X3Y112_AO5;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X3Y112_AO6;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X3Y112_A_CY;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X3Y112_A_XOR;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X3Y112_B;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X3Y112_B1;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X3Y112_B2;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X3Y112_B3;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X3Y112_B4;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X3Y112_B5;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X3Y112_B6;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X3Y112_BO5;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X3Y112_BO6;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X3Y112_B_CY;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X3Y112_B_XOR;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X3Y112_C;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X3Y112_C1;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X3Y112_C2;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X3Y112_C3;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X3Y112_C4;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X3Y112_C5;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X3Y112_C6;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X3Y112_CO5;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X3Y112_CO6;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X3Y112_C_CY;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X3Y112_C_XOR;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X3Y112_D;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X3Y112_D1;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X3Y112_D2;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X3Y112_D3;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X3Y112_D4;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X3Y112_D5;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X3Y112_D6;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X3Y112_DO5;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X3Y112_DO6;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X3Y112_D_CY;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X3Y112_D_XOR;
  wire [0:0] CLBLM_R_X49Y101_SLICE_X74Y101_A;
  wire [0:0] CLBLM_R_X49Y101_SLICE_X74Y101_A1;
  wire [0:0] CLBLM_R_X49Y101_SLICE_X74Y101_A2;
  wire [0:0] CLBLM_R_X49Y101_SLICE_X74Y101_A3;
  wire [0:0] CLBLM_R_X49Y101_SLICE_X74Y101_A4;
  wire [0:0] CLBLM_R_X49Y101_SLICE_X74Y101_A5;
  wire [0:0] CLBLM_R_X49Y101_SLICE_X74Y101_A6;
  wire [0:0] CLBLM_R_X49Y101_SLICE_X74Y101_AMUX;
  wire [0:0] CLBLM_R_X49Y101_SLICE_X74Y101_AO5;
  wire [0:0] CLBLM_R_X49Y101_SLICE_X74Y101_AO6;
  wire [0:0] CLBLM_R_X49Y101_SLICE_X74Y101_A_CY;
  wire [0:0] CLBLM_R_X49Y101_SLICE_X74Y101_A_XOR;
  wire [0:0] CLBLM_R_X49Y101_SLICE_X74Y101_B;
  wire [0:0] CLBLM_R_X49Y101_SLICE_X74Y101_B1;
  wire [0:0] CLBLM_R_X49Y101_SLICE_X74Y101_B2;
  wire [0:0] CLBLM_R_X49Y101_SLICE_X74Y101_B3;
  wire [0:0] CLBLM_R_X49Y101_SLICE_X74Y101_B4;
  wire [0:0] CLBLM_R_X49Y101_SLICE_X74Y101_B5;
  wire [0:0] CLBLM_R_X49Y101_SLICE_X74Y101_B6;
  wire [0:0] CLBLM_R_X49Y101_SLICE_X74Y101_BO5;
  wire [0:0] CLBLM_R_X49Y101_SLICE_X74Y101_BO6;
  wire [0:0] CLBLM_R_X49Y101_SLICE_X74Y101_B_CY;
  wire [0:0] CLBLM_R_X49Y101_SLICE_X74Y101_B_XOR;
  wire [0:0] CLBLM_R_X49Y101_SLICE_X74Y101_C;
  wire [0:0] CLBLM_R_X49Y101_SLICE_X74Y101_C1;
  wire [0:0] CLBLM_R_X49Y101_SLICE_X74Y101_C2;
  wire [0:0] CLBLM_R_X49Y101_SLICE_X74Y101_C3;
  wire [0:0] CLBLM_R_X49Y101_SLICE_X74Y101_C4;
  wire [0:0] CLBLM_R_X49Y101_SLICE_X74Y101_C5;
  wire [0:0] CLBLM_R_X49Y101_SLICE_X74Y101_C6;
  wire [0:0] CLBLM_R_X49Y101_SLICE_X74Y101_CO5;
  wire [0:0] CLBLM_R_X49Y101_SLICE_X74Y101_CO6;
  wire [0:0] CLBLM_R_X49Y101_SLICE_X74Y101_C_CY;
  wire [0:0] CLBLM_R_X49Y101_SLICE_X74Y101_C_XOR;
  wire [0:0] CLBLM_R_X49Y101_SLICE_X74Y101_D;
  wire [0:0] CLBLM_R_X49Y101_SLICE_X74Y101_D1;
  wire [0:0] CLBLM_R_X49Y101_SLICE_X74Y101_D2;
  wire [0:0] CLBLM_R_X49Y101_SLICE_X74Y101_D3;
  wire [0:0] CLBLM_R_X49Y101_SLICE_X74Y101_D4;
  wire [0:0] CLBLM_R_X49Y101_SLICE_X74Y101_D5;
  wire [0:0] CLBLM_R_X49Y101_SLICE_X74Y101_D6;
  wire [0:0] CLBLM_R_X49Y101_SLICE_X74Y101_DO5;
  wire [0:0] CLBLM_R_X49Y101_SLICE_X74Y101_DO6;
  wire [0:0] CLBLM_R_X49Y101_SLICE_X74Y101_D_CY;
  wire [0:0] CLBLM_R_X49Y101_SLICE_X74Y101_D_XOR;
  wire [0:0] CLBLM_R_X49Y101_SLICE_X75Y101_A;
  wire [0:0] CLBLM_R_X49Y101_SLICE_X75Y101_A1;
  wire [0:0] CLBLM_R_X49Y101_SLICE_X75Y101_A2;
  wire [0:0] CLBLM_R_X49Y101_SLICE_X75Y101_A3;
  wire [0:0] CLBLM_R_X49Y101_SLICE_X75Y101_A4;
  wire [0:0] CLBLM_R_X49Y101_SLICE_X75Y101_A5;
  wire [0:0] CLBLM_R_X49Y101_SLICE_X75Y101_A6;
  wire [0:0] CLBLM_R_X49Y101_SLICE_X75Y101_AO5;
  wire [0:0] CLBLM_R_X49Y101_SLICE_X75Y101_AO6;
  wire [0:0] CLBLM_R_X49Y101_SLICE_X75Y101_A_CY;
  wire [0:0] CLBLM_R_X49Y101_SLICE_X75Y101_A_XOR;
  wire [0:0] CLBLM_R_X49Y101_SLICE_X75Y101_B;
  wire [0:0] CLBLM_R_X49Y101_SLICE_X75Y101_B1;
  wire [0:0] CLBLM_R_X49Y101_SLICE_X75Y101_B2;
  wire [0:0] CLBLM_R_X49Y101_SLICE_X75Y101_B3;
  wire [0:0] CLBLM_R_X49Y101_SLICE_X75Y101_B4;
  wire [0:0] CLBLM_R_X49Y101_SLICE_X75Y101_B5;
  wire [0:0] CLBLM_R_X49Y101_SLICE_X75Y101_B6;
  wire [0:0] CLBLM_R_X49Y101_SLICE_X75Y101_BO5;
  wire [0:0] CLBLM_R_X49Y101_SLICE_X75Y101_BO6;
  wire [0:0] CLBLM_R_X49Y101_SLICE_X75Y101_B_CY;
  wire [0:0] CLBLM_R_X49Y101_SLICE_X75Y101_B_XOR;
  wire [0:0] CLBLM_R_X49Y101_SLICE_X75Y101_C;
  wire [0:0] CLBLM_R_X49Y101_SLICE_X75Y101_C1;
  wire [0:0] CLBLM_R_X49Y101_SLICE_X75Y101_C2;
  wire [0:0] CLBLM_R_X49Y101_SLICE_X75Y101_C3;
  wire [0:0] CLBLM_R_X49Y101_SLICE_X75Y101_C4;
  wire [0:0] CLBLM_R_X49Y101_SLICE_X75Y101_C5;
  wire [0:0] CLBLM_R_X49Y101_SLICE_X75Y101_C6;
  wire [0:0] CLBLM_R_X49Y101_SLICE_X75Y101_CO5;
  wire [0:0] CLBLM_R_X49Y101_SLICE_X75Y101_CO6;
  wire [0:0] CLBLM_R_X49Y101_SLICE_X75Y101_C_CY;
  wire [0:0] CLBLM_R_X49Y101_SLICE_X75Y101_C_XOR;
  wire [0:0] CLBLM_R_X49Y101_SLICE_X75Y101_D;
  wire [0:0] CLBLM_R_X49Y101_SLICE_X75Y101_D1;
  wire [0:0] CLBLM_R_X49Y101_SLICE_X75Y101_D2;
  wire [0:0] CLBLM_R_X49Y101_SLICE_X75Y101_D3;
  wire [0:0] CLBLM_R_X49Y101_SLICE_X75Y101_D4;
  wire [0:0] CLBLM_R_X49Y101_SLICE_X75Y101_D5;
  wire [0:0] CLBLM_R_X49Y101_SLICE_X75Y101_D6;
  wire [0:0] CLBLM_R_X49Y101_SLICE_X75Y101_DO5;
  wire [0:0] CLBLM_R_X49Y101_SLICE_X75Y101_DO6;
  wire [0:0] CLBLM_R_X49Y101_SLICE_X75Y101_D_CY;
  wire [0:0] CLBLM_R_X49Y101_SLICE_X75Y101_D_XOR;
  wire [0:0] CLBLM_R_X49Y95_SLICE_X74Y95_A;
  wire [0:0] CLBLM_R_X49Y95_SLICE_X74Y95_A1;
  wire [0:0] CLBLM_R_X49Y95_SLICE_X74Y95_A2;
  wire [0:0] CLBLM_R_X49Y95_SLICE_X74Y95_A3;
  wire [0:0] CLBLM_R_X49Y95_SLICE_X74Y95_A4;
  wire [0:0] CLBLM_R_X49Y95_SLICE_X74Y95_A5;
  wire [0:0] CLBLM_R_X49Y95_SLICE_X74Y95_A6;
  wire [0:0] CLBLM_R_X49Y95_SLICE_X74Y95_AMUX;
  wire [0:0] CLBLM_R_X49Y95_SLICE_X74Y95_AO5;
  wire [0:0] CLBLM_R_X49Y95_SLICE_X74Y95_AO6;
  wire [0:0] CLBLM_R_X49Y95_SLICE_X74Y95_A_CY;
  wire [0:0] CLBLM_R_X49Y95_SLICE_X74Y95_A_XOR;
  wire [0:0] CLBLM_R_X49Y95_SLICE_X74Y95_B;
  wire [0:0] CLBLM_R_X49Y95_SLICE_X74Y95_B1;
  wire [0:0] CLBLM_R_X49Y95_SLICE_X74Y95_B2;
  wire [0:0] CLBLM_R_X49Y95_SLICE_X74Y95_B3;
  wire [0:0] CLBLM_R_X49Y95_SLICE_X74Y95_B4;
  wire [0:0] CLBLM_R_X49Y95_SLICE_X74Y95_B5;
  wire [0:0] CLBLM_R_X49Y95_SLICE_X74Y95_B6;
  wire [0:0] CLBLM_R_X49Y95_SLICE_X74Y95_BO5;
  wire [0:0] CLBLM_R_X49Y95_SLICE_X74Y95_BO6;
  wire [0:0] CLBLM_R_X49Y95_SLICE_X74Y95_B_CY;
  wire [0:0] CLBLM_R_X49Y95_SLICE_X74Y95_B_XOR;
  wire [0:0] CLBLM_R_X49Y95_SLICE_X74Y95_C;
  wire [0:0] CLBLM_R_X49Y95_SLICE_X74Y95_C1;
  wire [0:0] CLBLM_R_X49Y95_SLICE_X74Y95_C2;
  wire [0:0] CLBLM_R_X49Y95_SLICE_X74Y95_C3;
  wire [0:0] CLBLM_R_X49Y95_SLICE_X74Y95_C4;
  wire [0:0] CLBLM_R_X49Y95_SLICE_X74Y95_C5;
  wire [0:0] CLBLM_R_X49Y95_SLICE_X74Y95_C6;
  wire [0:0] CLBLM_R_X49Y95_SLICE_X74Y95_CO5;
  wire [0:0] CLBLM_R_X49Y95_SLICE_X74Y95_CO6;
  wire [0:0] CLBLM_R_X49Y95_SLICE_X74Y95_C_CY;
  wire [0:0] CLBLM_R_X49Y95_SLICE_X74Y95_C_XOR;
  wire [0:0] CLBLM_R_X49Y95_SLICE_X74Y95_D;
  wire [0:0] CLBLM_R_X49Y95_SLICE_X74Y95_D1;
  wire [0:0] CLBLM_R_X49Y95_SLICE_X74Y95_D2;
  wire [0:0] CLBLM_R_X49Y95_SLICE_X74Y95_D3;
  wire [0:0] CLBLM_R_X49Y95_SLICE_X74Y95_D4;
  wire [0:0] CLBLM_R_X49Y95_SLICE_X74Y95_D5;
  wire [0:0] CLBLM_R_X49Y95_SLICE_X74Y95_D6;
  wire [0:0] CLBLM_R_X49Y95_SLICE_X74Y95_DO5;
  wire [0:0] CLBLM_R_X49Y95_SLICE_X74Y95_DO6;
  wire [0:0] CLBLM_R_X49Y95_SLICE_X74Y95_D_CY;
  wire [0:0] CLBLM_R_X49Y95_SLICE_X74Y95_D_XOR;
  wire [0:0] CLBLM_R_X49Y95_SLICE_X75Y95_A;
  wire [0:0] CLBLM_R_X49Y95_SLICE_X75Y95_A1;
  wire [0:0] CLBLM_R_X49Y95_SLICE_X75Y95_A2;
  wire [0:0] CLBLM_R_X49Y95_SLICE_X75Y95_A3;
  wire [0:0] CLBLM_R_X49Y95_SLICE_X75Y95_A4;
  wire [0:0] CLBLM_R_X49Y95_SLICE_X75Y95_A5;
  wire [0:0] CLBLM_R_X49Y95_SLICE_X75Y95_A6;
  wire [0:0] CLBLM_R_X49Y95_SLICE_X75Y95_AO5;
  wire [0:0] CLBLM_R_X49Y95_SLICE_X75Y95_AO6;
  wire [0:0] CLBLM_R_X49Y95_SLICE_X75Y95_A_CY;
  wire [0:0] CLBLM_R_X49Y95_SLICE_X75Y95_A_XOR;
  wire [0:0] CLBLM_R_X49Y95_SLICE_X75Y95_B;
  wire [0:0] CLBLM_R_X49Y95_SLICE_X75Y95_B1;
  wire [0:0] CLBLM_R_X49Y95_SLICE_X75Y95_B2;
  wire [0:0] CLBLM_R_X49Y95_SLICE_X75Y95_B3;
  wire [0:0] CLBLM_R_X49Y95_SLICE_X75Y95_B4;
  wire [0:0] CLBLM_R_X49Y95_SLICE_X75Y95_B5;
  wire [0:0] CLBLM_R_X49Y95_SLICE_X75Y95_B6;
  wire [0:0] CLBLM_R_X49Y95_SLICE_X75Y95_BO5;
  wire [0:0] CLBLM_R_X49Y95_SLICE_X75Y95_BO6;
  wire [0:0] CLBLM_R_X49Y95_SLICE_X75Y95_B_CY;
  wire [0:0] CLBLM_R_X49Y95_SLICE_X75Y95_B_XOR;
  wire [0:0] CLBLM_R_X49Y95_SLICE_X75Y95_C;
  wire [0:0] CLBLM_R_X49Y95_SLICE_X75Y95_C1;
  wire [0:0] CLBLM_R_X49Y95_SLICE_X75Y95_C2;
  wire [0:0] CLBLM_R_X49Y95_SLICE_X75Y95_C3;
  wire [0:0] CLBLM_R_X49Y95_SLICE_X75Y95_C4;
  wire [0:0] CLBLM_R_X49Y95_SLICE_X75Y95_C5;
  wire [0:0] CLBLM_R_X49Y95_SLICE_X75Y95_C6;
  wire [0:0] CLBLM_R_X49Y95_SLICE_X75Y95_CO5;
  wire [0:0] CLBLM_R_X49Y95_SLICE_X75Y95_CO6;
  wire [0:0] CLBLM_R_X49Y95_SLICE_X75Y95_C_CY;
  wire [0:0] CLBLM_R_X49Y95_SLICE_X75Y95_C_XOR;
  wire [0:0] CLBLM_R_X49Y95_SLICE_X75Y95_D;
  wire [0:0] CLBLM_R_X49Y95_SLICE_X75Y95_D1;
  wire [0:0] CLBLM_R_X49Y95_SLICE_X75Y95_D2;
  wire [0:0] CLBLM_R_X49Y95_SLICE_X75Y95_D3;
  wire [0:0] CLBLM_R_X49Y95_SLICE_X75Y95_D4;
  wire [0:0] CLBLM_R_X49Y95_SLICE_X75Y95_D5;
  wire [0:0] CLBLM_R_X49Y95_SLICE_X75Y95_D6;
  wire [0:0] CLBLM_R_X49Y95_SLICE_X75Y95_DO5;
  wire [0:0] CLBLM_R_X49Y95_SLICE_X75Y95_DO6;
  wire [0:0] CLBLM_R_X49Y95_SLICE_X75Y95_D_CY;
  wire [0:0] CLBLM_R_X49Y95_SLICE_X75Y95_D_XOR;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X6Y109_A;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X6Y109_A1;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X6Y109_A2;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X6Y109_A3;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X6Y109_A4;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X6Y109_A5;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X6Y109_A6;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X6Y109_AO5;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X6Y109_AO6;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X6Y109_A_CY;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X6Y109_A_XOR;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X6Y109_B;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X6Y109_B1;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X6Y109_B2;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X6Y109_B3;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X6Y109_B4;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X6Y109_B5;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X6Y109_B6;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X6Y109_BO5;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X6Y109_BO6;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X6Y109_B_CY;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X6Y109_B_XOR;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X6Y109_C;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X6Y109_C1;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X6Y109_C2;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X6Y109_C3;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X6Y109_C4;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X6Y109_C5;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X6Y109_C6;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X6Y109_CO5;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X6Y109_CO6;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X6Y109_C_CY;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X6Y109_C_XOR;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X6Y109_D;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X6Y109_D1;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X6Y109_D2;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X6Y109_D3;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X6Y109_D4;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X6Y109_D5;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X6Y109_D6;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X6Y109_DO5;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X6Y109_DO6;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X6Y109_D_CY;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X6Y109_D_XOR;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X7Y109_A;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X7Y109_A1;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X7Y109_A2;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X7Y109_A3;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X7Y109_A4;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X7Y109_A5;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X7Y109_A6;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X7Y109_AO5;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X7Y109_AO6;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X7Y109_A_CY;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X7Y109_A_XOR;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X7Y109_B;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X7Y109_B1;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X7Y109_B2;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X7Y109_B3;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X7Y109_B4;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X7Y109_B5;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X7Y109_B6;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X7Y109_BO5;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X7Y109_BO6;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X7Y109_B_CY;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X7Y109_B_XOR;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X7Y109_C;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X7Y109_C1;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X7Y109_C2;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X7Y109_C3;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X7Y109_C4;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X7Y109_C5;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X7Y109_C6;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X7Y109_CO5;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X7Y109_CO6;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X7Y109_C_CY;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X7Y109_C_XOR;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X7Y109_D;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X7Y109_D1;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X7Y109_D2;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X7Y109_D3;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X7Y109_D4;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X7Y109_D5;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X7Y109_D6;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X7Y109_DO5;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X7Y109_DO6;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X7Y109_D_CY;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X7Y109_D_XOR;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X6Y110_A;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X6Y110_A1;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X6Y110_A2;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X6Y110_A3;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X6Y110_A4;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X6Y110_A5;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X6Y110_A6;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X6Y110_AMUX;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X6Y110_AO5;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X6Y110_AO6;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X6Y110_A_CY;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X6Y110_A_XOR;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X6Y110_B;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X6Y110_B1;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X6Y110_B2;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X6Y110_B3;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X6Y110_B4;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X6Y110_B5;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X6Y110_B6;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X6Y110_BO5;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X6Y110_BO6;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X6Y110_B_CY;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X6Y110_B_XOR;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X6Y110_C;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X6Y110_C1;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X6Y110_C2;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X6Y110_C3;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X6Y110_C4;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X6Y110_C5;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X6Y110_C6;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X6Y110_CO5;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X6Y110_CO6;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X6Y110_C_CY;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X6Y110_C_XOR;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X6Y110_D;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X6Y110_D1;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X6Y110_D2;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X6Y110_D3;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X6Y110_D4;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X6Y110_D5;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X6Y110_D6;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X6Y110_DO5;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X6Y110_DO6;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X6Y110_D_CY;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X6Y110_D_XOR;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X7Y110_A;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X7Y110_A1;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X7Y110_A2;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X7Y110_A3;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X7Y110_A4;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X7Y110_A5;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X7Y110_A6;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X7Y110_AO5;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X7Y110_AO6;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X7Y110_A_CY;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X7Y110_A_XOR;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X7Y110_B;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X7Y110_B1;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X7Y110_B2;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X7Y110_B3;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X7Y110_B4;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X7Y110_B5;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X7Y110_B6;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X7Y110_BO5;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X7Y110_BO6;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X7Y110_B_CY;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X7Y110_B_XOR;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X7Y110_C;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X7Y110_C1;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X7Y110_C2;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X7Y110_C3;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X7Y110_C4;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X7Y110_C5;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X7Y110_C6;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X7Y110_CO5;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X7Y110_CO6;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X7Y110_C_CY;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X7Y110_C_XOR;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X7Y110_D;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X7Y110_D1;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X7Y110_D2;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X7Y110_D3;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X7Y110_D4;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X7Y110_D5;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X7Y110_D6;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X7Y110_DO5;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X7Y110_DO6;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X7Y110_D_CY;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X7Y110_D_XOR;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X6Y111_A;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X6Y111_A1;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X6Y111_A2;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X6Y111_A3;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X6Y111_A4;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X6Y111_A5;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X6Y111_A6;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X6Y111_AMUX;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X6Y111_AO5;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X6Y111_AO6;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X6Y111_A_CY;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X6Y111_A_XOR;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X6Y111_B;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X6Y111_B1;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X6Y111_B2;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X6Y111_B3;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X6Y111_B4;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X6Y111_B5;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X6Y111_B6;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X6Y111_BO5;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X6Y111_BO6;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X6Y111_B_CY;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X6Y111_B_XOR;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X6Y111_C;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X6Y111_C1;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X6Y111_C2;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X6Y111_C3;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X6Y111_C4;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X6Y111_C5;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X6Y111_C6;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X6Y111_CO5;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X6Y111_CO6;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X6Y111_C_CY;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X6Y111_C_XOR;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X6Y111_D;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X6Y111_D1;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X6Y111_D2;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X6Y111_D3;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X6Y111_D4;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X6Y111_D5;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X6Y111_D6;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X6Y111_DO5;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X6Y111_DO6;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X6Y111_D_CY;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X6Y111_D_XOR;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X7Y111_A;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X7Y111_A1;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X7Y111_A2;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X7Y111_A3;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X7Y111_A4;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X7Y111_A5;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X7Y111_A6;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X7Y111_AMUX;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X7Y111_AO5;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X7Y111_AO6;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X7Y111_A_CY;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X7Y111_A_XOR;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X7Y111_B;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X7Y111_B1;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X7Y111_B2;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X7Y111_B3;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X7Y111_B4;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X7Y111_B5;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X7Y111_B6;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X7Y111_BO5;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X7Y111_BO6;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X7Y111_B_CY;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X7Y111_B_XOR;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X7Y111_C;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X7Y111_C1;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X7Y111_C2;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X7Y111_C3;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X7Y111_C4;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X7Y111_C5;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X7Y111_C6;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X7Y111_CO5;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X7Y111_CO6;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X7Y111_C_CY;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X7Y111_C_XOR;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X7Y111_D;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X7Y111_D1;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X7Y111_D2;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X7Y111_D3;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X7Y111_D4;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X7Y111_D5;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X7Y111_D6;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X7Y111_DO5;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X7Y111_DO6;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X7Y111_D_CY;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X7Y111_D_XOR;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X6Y112_A;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X6Y112_A1;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X6Y112_A2;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X6Y112_A3;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X6Y112_A4;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X6Y112_A5;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X6Y112_A6;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X6Y112_AO5;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X6Y112_AO6;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X6Y112_A_CY;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X6Y112_A_XOR;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X6Y112_B;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X6Y112_B1;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X6Y112_B2;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X6Y112_B3;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X6Y112_B4;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X6Y112_B5;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X6Y112_B6;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X6Y112_BO5;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X6Y112_BO6;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X6Y112_B_CY;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X6Y112_B_XOR;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X6Y112_C;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X6Y112_C1;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X6Y112_C2;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X6Y112_C3;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X6Y112_C4;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X6Y112_C5;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X6Y112_C6;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X6Y112_CO5;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X6Y112_CO6;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X6Y112_C_CY;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X6Y112_C_XOR;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X6Y112_D;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X6Y112_D1;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X6Y112_D2;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X6Y112_D3;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X6Y112_D4;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X6Y112_D5;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X6Y112_D6;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X6Y112_DO5;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X6Y112_DO6;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X6Y112_D_CY;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X6Y112_D_XOR;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X7Y112_A;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X7Y112_A1;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X7Y112_A2;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X7Y112_A3;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X7Y112_A4;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X7Y112_A5;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X7Y112_A6;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X7Y112_AMUX;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X7Y112_AO5;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X7Y112_AO6;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X7Y112_A_CY;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X7Y112_A_XOR;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X7Y112_B;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X7Y112_B1;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X7Y112_B2;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X7Y112_B3;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X7Y112_B4;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X7Y112_B5;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X7Y112_B6;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X7Y112_BO5;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X7Y112_BO6;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X7Y112_B_CY;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X7Y112_B_XOR;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X7Y112_C;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X7Y112_C1;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X7Y112_C2;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X7Y112_C3;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X7Y112_C4;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X7Y112_C5;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X7Y112_C6;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X7Y112_CO5;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X7Y112_CO6;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X7Y112_C_CY;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X7Y112_C_XOR;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X7Y112_D;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X7Y112_D1;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X7Y112_D2;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X7Y112_D3;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X7Y112_D4;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X7Y112_D5;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X7Y112_D6;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X7Y112_DO5;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X7Y112_DO6;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X7Y112_D_CY;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X7Y112_D_XOR;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X6Y113_A;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X6Y113_A1;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X6Y113_A2;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X6Y113_A3;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X6Y113_A4;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X6Y113_A5;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X6Y113_A6;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X6Y113_AMUX;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X6Y113_AO5;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X6Y113_AO6;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X6Y113_A_CY;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X6Y113_A_XOR;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X6Y113_B;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X6Y113_B1;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X6Y113_B2;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X6Y113_B3;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X6Y113_B4;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X6Y113_B5;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X6Y113_B6;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X6Y113_BO5;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X6Y113_BO6;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X6Y113_B_CY;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X6Y113_B_XOR;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X6Y113_C;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X6Y113_C1;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X6Y113_C2;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X6Y113_C3;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X6Y113_C4;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X6Y113_C5;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X6Y113_C6;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X6Y113_CO5;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X6Y113_CO6;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X6Y113_C_CY;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X6Y113_C_XOR;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X6Y113_D;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X6Y113_D1;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X6Y113_D2;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X6Y113_D3;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X6Y113_D4;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X6Y113_D5;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X6Y113_D6;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X6Y113_DO5;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X6Y113_DO6;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X6Y113_D_CY;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X6Y113_D_XOR;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X7Y113_A;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X7Y113_A1;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X7Y113_A2;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X7Y113_A3;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X7Y113_A4;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X7Y113_A5;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X7Y113_A6;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X7Y113_AO5;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X7Y113_AO6;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X7Y113_A_CY;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X7Y113_A_XOR;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X7Y113_B;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X7Y113_B1;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X7Y113_B2;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X7Y113_B3;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X7Y113_B4;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X7Y113_B5;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X7Y113_B6;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X7Y113_BO5;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X7Y113_BO6;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X7Y113_B_CY;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X7Y113_B_XOR;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X7Y113_C;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X7Y113_C1;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X7Y113_C2;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X7Y113_C3;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X7Y113_C4;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X7Y113_C5;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X7Y113_C6;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X7Y113_CO5;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X7Y113_CO6;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X7Y113_C_CY;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X7Y113_C_XOR;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X7Y113_D;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X7Y113_D1;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X7Y113_D2;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X7Y113_D3;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X7Y113_D4;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X7Y113_D5;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X7Y113_D6;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X7Y113_DO5;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X7Y113_DO6;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X7Y113_D_CY;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X7Y113_D_XOR;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X6Y114_A;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X6Y114_A1;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X6Y114_A2;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X6Y114_A3;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X6Y114_A4;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X6Y114_A5;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X6Y114_A6;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X6Y114_AO5;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X6Y114_AO6;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X6Y114_A_CY;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X6Y114_A_XOR;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X6Y114_B;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X6Y114_B1;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X6Y114_B2;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X6Y114_B3;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X6Y114_B4;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X6Y114_B5;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X6Y114_B6;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X6Y114_BO5;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X6Y114_BO6;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X6Y114_B_CY;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X6Y114_B_XOR;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X6Y114_C;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X6Y114_C1;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X6Y114_C2;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X6Y114_C3;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X6Y114_C4;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X6Y114_C5;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X6Y114_C6;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X6Y114_CO5;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X6Y114_CO6;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X6Y114_C_CY;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X6Y114_C_XOR;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X6Y114_D;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X6Y114_D1;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X6Y114_D2;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X6Y114_D3;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X6Y114_D4;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X6Y114_D5;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X6Y114_D6;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X6Y114_DO5;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X6Y114_DO6;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X6Y114_D_CY;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X6Y114_D_XOR;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X7Y114_A;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X7Y114_A1;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X7Y114_A2;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X7Y114_A3;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X7Y114_A4;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X7Y114_A5;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X7Y114_A6;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X7Y114_AMUX;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X7Y114_AO5;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X7Y114_AO6;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X7Y114_A_CY;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X7Y114_A_XOR;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X7Y114_B;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X7Y114_B1;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X7Y114_B2;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X7Y114_B3;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X7Y114_B4;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X7Y114_B5;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X7Y114_B6;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X7Y114_BO5;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X7Y114_BO6;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X7Y114_B_CY;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X7Y114_B_XOR;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X7Y114_C;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X7Y114_C1;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X7Y114_C2;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X7Y114_C3;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X7Y114_C4;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X7Y114_C5;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X7Y114_C6;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X7Y114_CO5;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X7Y114_CO6;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X7Y114_C_CY;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X7Y114_C_XOR;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X7Y114_D;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X7Y114_D1;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X7Y114_D2;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X7Y114_D3;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X7Y114_D4;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X7Y114_D5;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X7Y114_D6;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X7Y114_DO5;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X7Y114_DO6;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X7Y114_D_CY;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X7Y114_D_XOR;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X6Y115_A;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X6Y115_A1;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X6Y115_A2;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X6Y115_A3;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X6Y115_A4;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X6Y115_A5;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X6Y115_A6;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X6Y115_AMUX;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X6Y115_AO5;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X6Y115_AO6;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X6Y115_A_CY;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X6Y115_A_XOR;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X6Y115_B;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X6Y115_B1;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X6Y115_B2;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X6Y115_B3;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X6Y115_B4;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X6Y115_B5;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X6Y115_B6;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X6Y115_BMUX;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X6Y115_BO5;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X6Y115_BO6;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X6Y115_B_CY;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X6Y115_B_XOR;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X6Y115_C;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X6Y115_C1;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X6Y115_C2;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X6Y115_C3;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X6Y115_C4;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X6Y115_C5;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X6Y115_C6;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X6Y115_CO5;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X6Y115_CO6;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X6Y115_C_CY;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X6Y115_C_XOR;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X6Y115_D;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X6Y115_D1;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X6Y115_D2;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X6Y115_D3;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X6Y115_D4;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X6Y115_D5;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X6Y115_D6;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X6Y115_DO5;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X6Y115_DO6;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X6Y115_D_CY;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X6Y115_D_XOR;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X7Y115_A;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X7Y115_A1;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X7Y115_A2;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X7Y115_A3;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X7Y115_A4;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X7Y115_A5;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X7Y115_A6;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X7Y115_AO5;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X7Y115_AO6;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X7Y115_A_CY;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X7Y115_A_XOR;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X7Y115_B;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X7Y115_B1;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X7Y115_B2;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X7Y115_B3;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X7Y115_B4;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X7Y115_B5;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X7Y115_B6;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X7Y115_BO5;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X7Y115_BO6;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X7Y115_B_CY;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X7Y115_B_XOR;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X7Y115_C;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X7Y115_C1;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X7Y115_C2;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X7Y115_C3;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X7Y115_C4;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X7Y115_C5;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X7Y115_C6;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X7Y115_CO5;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X7Y115_CO6;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X7Y115_C_CY;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X7Y115_C_XOR;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X7Y115_D;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X7Y115_D1;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X7Y115_D2;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X7Y115_D3;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X7Y115_D4;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X7Y115_D5;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X7Y115_D6;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X7Y115_DO5;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X7Y115_DO6;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X7Y115_D_CY;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X7Y115_D_XOR;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X8Y113_A;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X8Y113_A1;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X8Y113_A2;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X8Y113_A3;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X8Y113_A4;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X8Y113_A5;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X8Y113_A6;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X8Y113_AMUX;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X8Y113_AO5;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X8Y113_AO6;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X8Y113_A_CY;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X8Y113_A_XOR;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X8Y113_B;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X8Y113_B1;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X8Y113_B2;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X8Y113_B3;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X8Y113_B4;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X8Y113_B5;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X8Y113_B6;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X8Y113_BMUX;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X8Y113_BO5;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X8Y113_BO6;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X8Y113_B_CY;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X8Y113_B_XOR;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X8Y113_C;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X8Y113_C1;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X8Y113_C2;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X8Y113_C3;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X8Y113_C4;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X8Y113_C5;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X8Y113_C6;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X8Y113_CO5;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X8Y113_CO6;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X8Y113_C_CY;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X8Y113_C_XOR;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X8Y113_D;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X8Y113_D1;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X8Y113_D2;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X8Y113_D3;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X8Y113_D4;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X8Y113_D5;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X8Y113_D6;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X8Y113_DO5;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X8Y113_DO6;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X8Y113_D_CY;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X8Y113_D_XOR;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X9Y113_A;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X9Y113_A1;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X9Y113_A2;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X9Y113_A3;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X9Y113_A4;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X9Y113_A5;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X9Y113_A6;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X9Y113_AO5;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X9Y113_AO6;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X9Y113_A_CY;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X9Y113_A_XOR;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X9Y113_B;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X9Y113_B1;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X9Y113_B2;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X9Y113_B3;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X9Y113_B4;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X9Y113_B5;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X9Y113_B6;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X9Y113_BO5;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X9Y113_BO6;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X9Y113_B_CY;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X9Y113_B_XOR;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X9Y113_C;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X9Y113_C1;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X9Y113_C2;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X9Y113_C3;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X9Y113_C4;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X9Y113_C5;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X9Y113_C6;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X9Y113_CO5;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X9Y113_CO6;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X9Y113_C_CY;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X9Y113_C_XOR;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X9Y113_D;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X9Y113_D1;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X9Y113_D2;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X9Y113_D3;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X9Y113_D4;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X9Y113_D5;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X9Y113_D6;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X9Y113_DO5;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X9Y113_DO6;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X9Y113_D_CY;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X9Y113_D_XOR;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X8Y114_A;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X8Y114_A1;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X8Y114_A2;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X8Y114_A3;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X8Y114_A4;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X8Y114_A5;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X8Y114_A6;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X8Y114_AMUX;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X8Y114_AO5;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X8Y114_AO6;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X8Y114_A_CY;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X8Y114_A_XOR;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X8Y114_B;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X8Y114_B1;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X8Y114_B2;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X8Y114_B3;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X8Y114_B4;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X8Y114_B5;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X8Y114_B6;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X8Y114_BMUX;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X8Y114_BO5;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X8Y114_BO6;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X8Y114_B_CY;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X8Y114_B_XOR;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X8Y114_C;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X8Y114_C1;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X8Y114_C2;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X8Y114_C3;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X8Y114_C4;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X8Y114_C5;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X8Y114_C6;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X8Y114_CO5;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X8Y114_CO6;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X8Y114_C_CY;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X8Y114_C_XOR;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X8Y114_D;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X8Y114_D1;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X8Y114_D2;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X8Y114_D3;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X8Y114_D4;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X8Y114_D5;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X8Y114_D6;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X8Y114_DO5;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X8Y114_DO6;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X8Y114_D_CY;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X8Y114_D_XOR;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X9Y114_A;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X9Y114_A1;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X9Y114_A2;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X9Y114_A3;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X9Y114_A4;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X9Y114_A5;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X9Y114_A6;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X9Y114_AO5;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X9Y114_AO6;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X9Y114_A_CY;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X9Y114_A_XOR;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X9Y114_B;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X9Y114_B1;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X9Y114_B2;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X9Y114_B3;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X9Y114_B4;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X9Y114_B5;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X9Y114_B6;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X9Y114_BO5;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X9Y114_BO6;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X9Y114_B_CY;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X9Y114_B_XOR;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X9Y114_C;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X9Y114_C1;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X9Y114_C2;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X9Y114_C3;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X9Y114_C4;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X9Y114_C5;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X9Y114_C6;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X9Y114_CO5;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X9Y114_CO6;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X9Y114_C_CY;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X9Y114_C_XOR;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X9Y114_D;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X9Y114_D1;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X9Y114_D2;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X9Y114_D3;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X9Y114_D4;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X9Y114_D5;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X9Y114_D6;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X9Y114_DO5;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X9Y114_DO6;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X9Y114_D_CY;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X9Y114_D_XOR;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X8Y121_A;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X8Y121_A1;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X8Y121_A2;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X8Y121_A3;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X8Y121_A4;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X8Y121_A5;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X8Y121_A6;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X8Y121_AO5;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X8Y121_AO6;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X8Y121_A_CY;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X8Y121_A_XOR;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X8Y121_B;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X8Y121_B1;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X8Y121_B2;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X8Y121_B3;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X8Y121_B4;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X8Y121_B5;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X8Y121_B6;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X8Y121_BO5;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X8Y121_BO6;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X8Y121_B_CY;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X8Y121_B_XOR;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X8Y121_C;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X8Y121_C1;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X8Y121_C2;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X8Y121_C3;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X8Y121_C4;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X8Y121_C5;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X8Y121_C6;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X8Y121_CO5;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X8Y121_CO6;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X8Y121_C_CY;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X8Y121_C_XOR;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X8Y121_D;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X8Y121_D1;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X8Y121_D2;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X8Y121_D3;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X8Y121_D4;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X8Y121_D5;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X8Y121_D6;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X8Y121_DO5;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X8Y121_DO6;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X8Y121_D_CY;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X8Y121_D_XOR;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X9Y121_A;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X9Y121_A1;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X9Y121_A2;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X9Y121_A3;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X9Y121_A4;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X9Y121_A5;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X9Y121_A6;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X9Y121_AMUX;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X9Y121_AO5;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X9Y121_AO6;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X9Y121_A_CY;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X9Y121_A_XOR;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X9Y121_B;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X9Y121_B1;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X9Y121_B2;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X9Y121_B3;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X9Y121_B4;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X9Y121_B5;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X9Y121_B6;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X9Y121_BO5;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X9Y121_BO6;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X9Y121_B_CY;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X9Y121_B_XOR;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X9Y121_C;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X9Y121_C1;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X9Y121_C2;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X9Y121_C3;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X9Y121_C4;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X9Y121_C5;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X9Y121_C6;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X9Y121_CO5;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X9Y121_CO6;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X9Y121_C_CY;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X9Y121_C_XOR;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X9Y121_D;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X9Y121_D1;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X9Y121_D2;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X9Y121_D3;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X9Y121_D4;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X9Y121_D5;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X9Y121_D6;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X9Y121_DO5;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X9Y121_DO6;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X9Y121_D_CY;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X9Y121_D_XOR;
  wire [0:0] LIOB33_SING_X0Y100_IOB_X0Y100_I;
  wire [0:0] LIOB33_SING_X0Y149_IOB_X0Y149_I;
  wire [0:0] LIOB33_SING_X0Y150_IOB_X0Y150_I;
  wire [0:0] LIOB33_SING_X0Y199_IOB_X0Y199_O;
  wire [0:0] LIOB33_SING_X0Y200_IOB_X0Y200_O;
  wire [0:0] LIOB33_SING_X0Y50_IOB_X0Y50_I;
  wire [0:0] LIOB33_SING_X0Y99_IOB_X0Y99_I;
  wire [0:0] LIOB33_X0Y101_IOB_X0Y101_I;
  wire [0:0] LIOB33_X0Y101_IOB_X0Y102_I;
  wire [0:0] LIOB33_X0Y103_IOB_X0Y103_I;
  wire [0:0] LIOB33_X0Y103_IOB_X0Y104_I;
  wire [0:0] LIOB33_X0Y105_IOB_X0Y105_I;
  wire [0:0] LIOB33_X0Y105_IOB_X0Y106_I;
  wire [0:0] LIOB33_X0Y107_IOB_X0Y107_I;
  wire [0:0] LIOB33_X0Y107_IOB_X0Y108_I;
  wire [0:0] LIOB33_X0Y109_IOB_X0Y109_I;
  wire [0:0] LIOB33_X0Y109_IOB_X0Y110_I;
  wire [0:0] LIOB33_X0Y111_IOB_X0Y111_I;
  wire [0:0] LIOB33_X0Y111_IOB_X0Y112_I;
  wire [0:0] LIOB33_X0Y113_IOB_X0Y113_I;
  wire [0:0] LIOB33_X0Y113_IOB_X0Y114_I;
  wire [0:0] LIOB33_X0Y115_IOB_X0Y115_I;
  wire [0:0] LIOB33_X0Y115_IOB_X0Y116_I;
  wire [0:0] LIOB33_X0Y117_IOB_X0Y117_I;
  wire [0:0] LIOB33_X0Y117_IOB_X0Y118_I;
  wire [0:0] LIOB33_X0Y119_IOB_X0Y119_I;
  wire [0:0] LIOB33_X0Y119_IOB_X0Y120_I;
  wire [0:0] LIOB33_X0Y121_IOB_X0Y121_I;
  wire [0:0] LIOB33_X0Y121_IOB_X0Y122_I;
  wire [0:0] LIOB33_X0Y123_IOB_X0Y123_I;
  wire [0:0] LIOB33_X0Y123_IOB_X0Y124_I;
  wire [0:0] LIOB33_X0Y125_IOB_X0Y125_I;
  wire [0:0] LIOB33_X0Y125_IOB_X0Y126_I;
  wire [0:0] LIOB33_X0Y127_IOB_X0Y127_I;
  wire [0:0] LIOB33_X0Y127_IOB_X0Y128_I;
  wire [0:0] LIOB33_X0Y129_IOB_X0Y129_I;
  wire [0:0] LIOB33_X0Y129_IOB_X0Y130_I;
  wire [0:0] LIOB33_X0Y131_IOB_X0Y131_I;
  wire [0:0] LIOB33_X0Y131_IOB_X0Y132_I;
  wire [0:0] LIOB33_X0Y133_IOB_X0Y133_I;
  wire [0:0] LIOB33_X0Y133_IOB_X0Y134_I;
  wire [0:0] LIOB33_X0Y135_IOB_X0Y135_I;
  wire [0:0] LIOB33_X0Y135_IOB_X0Y136_I;
  wire [0:0] LIOB33_X0Y137_IOB_X0Y137_I;
  wire [0:0] LIOB33_X0Y137_IOB_X0Y138_I;
  wire [0:0] LIOB33_X0Y139_IOB_X0Y139_I;
  wire [0:0] LIOB33_X0Y139_IOB_X0Y140_I;
  wire [0:0] LIOB33_X0Y141_IOB_X0Y141_I;
  wire [0:0] LIOB33_X0Y141_IOB_X0Y142_I;
  wire [0:0] LIOB33_X0Y143_IOB_X0Y143_I;
  wire [0:0] LIOB33_X0Y145_IOB_X0Y145_I;
  wire [0:0] LIOB33_X0Y145_IOB_X0Y146_I;
  wire [0:0] LIOB33_X0Y147_IOB_X0Y147_I;
  wire [0:0] LIOB33_X0Y147_IOB_X0Y148_I;
  wire [0:0] LIOB33_X0Y151_IOB_X0Y151_I;
  wire [0:0] LIOB33_X0Y151_IOB_X0Y152_I;
  wire [0:0] LIOB33_X0Y153_IOB_X0Y153_I;
  wire [0:0] LIOB33_X0Y153_IOB_X0Y154_I;
  wire [0:0] LIOB33_X0Y155_IOB_X0Y155_I;
  wire [0:0] LIOB33_X0Y155_IOB_X0Y156_I;
  wire [0:0] LIOB33_X0Y157_IOB_X0Y157_I;
  wire [0:0] LIOB33_X0Y157_IOB_X0Y158_I;
  wire [0:0] LIOB33_X0Y159_IOB_X0Y159_I;
  wire [0:0] LIOB33_X0Y159_IOB_X0Y160_I;
  wire [0:0] LIOB33_X0Y161_IOB_X0Y161_I;
  wire [0:0] LIOB33_X0Y161_IOB_X0Y162_I;
  wire [0:0] LIOB33_X0Y163_IOB_X0Y163_I;
  wire [0:0] LIOB33_X0Y163_IOB_X0Y164_I;
  wire [0:0] LIOB33_X0Y165_IOB_X0Y165_I;
  wire [0:0] LIOB33_X0Y165_IOB_X0Y166_I;
  wire [0:0] LIOB33_X0Y167_IOB_X0Y167_I;
  wire [0:0] LIOB33_X0Y167_IOB_X0Y168_I;
  wire [0:0] LIOB33_X0Y169_IOB_X0Y169_I;
  wire [0:0] LIOB33_X0Y169_IOB_X0Y170_I;
  wire [0:0] LIOB33_X0Y171_IOB_X0Y171_I;
  wire [0:0] LIOB33_X0Y171_IOB_X0Y172_I;
  wire [0:0] LIOB33_X0Y173_IOB_X0Y173_I;
  wire [0:0] LIOB33_X0Y173_IOB_X0Y174_I;
  wire [0:0] LIOB33_X0Y175_IOB_X0Y175_I;
  wire [0:0] LIOB33_X0Y175_IOB_X0Y176_I;
  wire [0:0] LIOB33_X0Y177_IOB_X0Y177_I;
  wire [0:0] LIOB33_X0Y177_IOB_X0Y178_O;
  wire [0:0] LIOB33_X0Y179_IOB_X0Y179_O;
  wire [0:0] LIOB33_X0Y179_IOB_X0Y180_O;
  wire [0:0] LIOB33_X0Y181_IOB_X0Y181_O;
  wire [0:0] LIOB33_X0Y181_IOB_X0Y182_O;
  wire [0:0] LIOB33_X0Y183_IOB_X0Y183_O;
  wire [0:0] LIOB33_X0Y183_IOB_X0Y184_O;
  wire [0:0] LIOB33_X0Y185_IOB_X0Y185_O;
  wire [0:0] LIOB33_X0Y185_IOB_X0Y186_O;
  wire [0:0] LIOB33_X0Y187_IOB_X0Y187_O;
  wire [0:0] LIOB33_X0Y187_IOB_X0Y188_O;
  wire [0:0] LIOB33_X0Y189_IOB_X0Y189_O;
  wire [0:0] LIOB33_X0Y189_IOB_X0Y190_O;
  wire [0:0] LIOB33_X0Y191_IOB_X0Y191_O;
  wire [0:0] LIOB33_X0Y191_IOB_X0Y192_O;
  wire [0:0] LIOB33_X0Y193_IOB_X0Y193_O;
  wire [0:0] LIOB33_X0Y193_IOB_X0Y194_O;
  wire [0:0] LIOB33_X0Y195_IOB_X0Y195_O;
  wire [0:0] LIOB33_X0Y195_IOB_X0Y196_O;
  wire [0:0] LIOB33_X0Y197_IOB_X0Y197_O;
  wire [0:0] LIOB33_X0Y197_IOB_X0Y198_O;
  wire [0:0] LIOB33_X0Y51_IOB_X0Y51_I;
  wire [0:0] LIOB33_X0Y51_IOB_X0Y52_I;
  wire [0:0] LIOB33_X0Y53_IOB_X0Y53_I;
  wire [0:0] LIOB33_X0Y53_IOB_X0Y54_I;
  wire [0:0] LIOB33_X0Y55_IOB_X0Y55_I;
  wire [0:0] LIOB33_X0Y55_IOB_X0Y56_I;
  wire [0:0] LIOB33_X0Y57_IOB_X0Y57_I;
  wire [0:0] LIOB33_X0Y57_IOB_X0Y58_I;
  wire [0:0] LIOB33_X0Y59_IOB_X0Y59_I;
  wire [0:0] LIOB33_X0Y59_IOB_X0Y60_I;
  wire [0:0] LIOB33_X0Y61_IOB_X0Y61_I;
  wire [0:0] LIOB33_X0Y61_IOB_X0Y62_I;
  wire [0:0] LIOB33_X0Y63_IOB_X0Y63_I;
  wire [0:0] LIOB33_X0Y63_IOB_X0Y64_I;
  wire [0:0] LIOB33_X0Y65_IOB_X0Y65_I;
  wire [0:0] LIOB33_X0Y65_IOB_X0Y66_I;
  wire [0:0] LIOB33_X0Y67_IOB_X0Y67_I;
  wire [0:0] LIOB33_X0Y67_IOB_X0Y68_I;
  wire [0:0] LIOB33_X0Y69_IOB_X0Y69_I;
  wire [0:0] LIOB33_X0Y69_IOB_X0Y70_I;
  wire [0:0] LIOB33_X0Y71_IOB_X0Y71_I;
  wire [0:0] LIOB33_X0Y71_IOB_X0Y72_I;
  wire [0:0] LIOB33_X0Y73_IOB_X0Y73_I;
  wire [0:0] LIOB33_X0Y73_IOB_X0Y74_I;
  wire [0:0] LIOB33_X0Y75_IOB_X0Y75_I;
  wire [0:0] LIOB33_X0Y75_IOB_X0Y76_I;
  wire [0:0] LIOB33_X0Y77_IOB_X0Y77_I;
  wire [0:0] LIOB33_X0Y77_IOB_X0Y78_I;
  wire [0:0] LIOB33_X0Y79_IOB_X0Y79_I;
  wire [0:0] LIOB33_X0Y79_IOB_X0Y80_I;
  wire [0:0] LIOB33_X0Y81_IOB_X0Y81_I;
  wire [0:0] LIOB33_X0Y81_IOB_X0Y82_I;
  wire [0:0] LIOB33_X0Y83_IOB_X0Y83_I;
  wire [0:0] LIOB33_X0Y83_IOB_X0Y84_I;
  wire [0:0] LIOB33_X0Y85_IOB_X0Y85_I;
  wire [0:0] LIOB33_X0Y85_IOB_X0Y86_I;
  wire [0:0] LIOB33_X0Y87_IOB_X0Y87_I;
  wire [0:0] LIOB33_X0Y87_IOB_X0Y88_I;
  wire [0:0] LIOB33_X0Y89_IOB_X0Y89_I;
  wire [0:0] LIOB33_X0Y89_IOB_X0Y90_I;
  wire [0:0] LIOB33_X0Y91_IOB_X0Y91_I;
  wire [0:0] LIOB33_X0Y91_IOB_X0Y92_I;
  wire [0:0] LIOB33_X0Y93_IOB_X0Y93_I;
  wire [0:0] LIOB33_X0Y93_IOB_X0Y94_I;
  wire [0:0] LIOB33_X0Y95_IOB_X0Y95_I;
  wire [0:0] LIOB33_X0Y95_IOB_X0Y96_I;
  wire [0:0] LIOB33_X0Y97_IOB_X0Y97_I;
  wire [0:0] LIOB33_X0Y97_IOB_X0Y98_I;
  wire [0:0] LIOI3_SING_X0Y100_ILOGIC_X0Y100_D;
  wire [0:0] LIOI3_SING_X0Y100_ILOGIC_X0Y100_O;
  wire [0:0] LIOI3_SING_X0Y150_ILOGIC_X0Y150_D;
  wire [0:0] LIOI3_SING_X0Y150_ILOGIC_X0Y150_O;
  wire [0:0] LIOI3_SING_X0Y199_OLOGIC_X0Y199_D1;
  wire [0:0] LIOI3_SING_X0Y199_OLOGIC_X0Y199_OQ;
  wire [0:0] LIOI3_SING_X0Y199_OLOGIC_X0Y199_T1;
  wire [0:0] LIOI3_SING_X0Y199_OLOGIC_X0Y199_TQ;
  wire [0:0] LIOI3_SING_X0Y200_OLOGIC_X0Y200_D1;
  wire [0:0] LIOI3_SING_X0Y200_OLOGIC_X0Y200_OQ;
  wire [0:0] LIOI3_SING_X0Y200_OLOGIC_X0Y200_T1;
  wire [0:0] LIOI3_SING_X0Y200_OLOGIC_X0Y200_TQ;
  wire [0:0] LIOI3_SING_X0Y50_ILOGIC_X0Y50_D;
  wire [0:0] LIOI3_SING_X0Y50_ILOGIC_X0Y50_O;
  wire [0:0] LIOI3_SING_X0Y99_ILOGIC_X0Y99_D;
  wire [0:0] LIOI3_SING_X0Y99_ILOGIC_X0Y99_O;
  wire [0:0] LIOI3_TBYTESRC_X0Y107_ILOGIC_X0Y107_D;
  wire [0:0] LIOI3_TBYTESRC_X0Y107_ILOGIC_X0Y107_O;
  wire [0:0] LIOI3_TBYTESRC_X0Y107_ILOGIC_X0Y108_D;
  wire [0:0] LIOI3_TBYTESRC_X0Y107_ILOGIC_X0Y108_O;
  wire [0:0] LIOI3_TBYTESRC_X0Y119_ILOGIC_X0Y119_D;
  wire [0:0] LIOI3_TBYTESRC_X0Y119_ILOGIC_X0Y119_O;
  wire [0:0] LIOI3_TBYTESRC_X0Y119_ILOGIC_X0Y120_D;
  wire [0:0] LIOI3_TBYTESRC_X0Y119_ILOGIC_X0Y120_O;
  wire [0:0] LIOI3_TBYTESRC_X0Y131_ILOGIC_X0Y131_D;
  wire [0:0] LIOI3_TBYTESRC_X0Y131_ILOGIC_X0Y131_O;
  wire [0:0] LIOI3_TBYTESRC_X0Y131_ILOGIC_X0Y132_D;
  wire [0:0] LIOI3_TBYTESRC_X0Y131_ILOGIC_X0Y132_O;
  wire [0:0] LIOI3_TBYTESRC_X0Y143_ILOGIC_X0Y143_D;
  wire [0:0] LIOI3_TBYTESRC_X0Y143_ILOGIC_X0Y143_O;
  wire [0:0] LIOI3_TBYTESRC_X0Y157_ILOGIC_X0Y157_D;
  wire [0:0] LIOI3_TBYTESRC_X0Y157_ILOGIC_X0Y157_O;
  wire [0:0] LIOI3_TBYTESRC_X0Y157_ILOGIC_X0Y158_D;
  wire [0:0] LIOI3_TBYTESRC_X0Y157_ILOGIC_X0Y158_O;
  wire [0:0] LIOI3_TBYTESRC_X0Y181_OLOGIC_X0Y181_D1;
  wire [0:0] LIOI3_TBYTESRC_X0Y181_OLOGIC_X0Y181_OQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y181_OLOGIC_X0Y181_T1;
  wire [0:0] LIOI3_TBYTESRC_X0Y181_OLOGIC_X0Y181_TQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y181_OLOGIC_X0Y182_D1;
  wire [0:0] LIOI3_TBYTESRC_X0Y181_OLOGIC_X0Y182_OQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y181_OLOGIC_X0Y182_T1;
  wire [0:0] LIOI3_TBYTESRC_X0Y181_OLOGIC_X0Y182_TQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y193_OLOGIC_X0Y193_D1;
  wire [0:0] LIOI3_TBYTESRC_X0Y193_OLOGIC_X0Y193_OQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y193_OLOGIC_X0Y193_T1;
  wire [0:0] LIOI3_TBYTESRC_X0Y193_OLOGIC_X0Y193_TQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y193_OLOGIC_X0Y194_D1;
  wire [0:0] LIOI3_TBYTESRC_X0Y193_OLOGIC_X0Y194_OQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y193_OLOGIC_X0Y194_T1;
  wire [0:0] LIOI3_TBYTESRC_X0Y193_OLOGIC_X0Y194_TQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y57_ILOGIC_X0Y57_D;
  wire [0:0] LIOI3_TBYTESRC_X0Y57_ILOGIC_X0Y57_O;
  wire [0:0] LIOI3_TBYTESRC_X0Y57_ILOGIC_X0Y58_D;
  wire [0:0] LIOI3_TBYTESRC_X0Y57_ILOGIC_X0Y58_O;
  wire [0:0] LIOI3_TBYTESRC_X0Y69_ILOGIC_X0Y70_D;
  wire [0:0] LIOI3_TBYTESRC_X0Y69_ILOGIC_X0Y70_O;
  wire [0:0] LIOI3_TBYTESRC_X0Y81_ILOGIC_X0Y81_D;
  wire [0:0] LIOI3_TBYTESRC_X0Y81_ILOGIC_X0Y81_O;
  wire [0:0] LIOI3_TBYTESRC_X0Y81_ILOGIC_X0Y82_D;
  wire [0:0] LIOI3_TBYTESRC_X0Y81_ILOGIC_X0Y82_O;
  wire [0:0] LIOI3_TBYTESRC_X0Y93_ILOGIC_X0Y93_D;
  wire [0:0] LIOI3_TBYTESRC_X0Y93_ILOGIC_X0Y93_O;
  wire [0:0] LIOI3_TBYTESRC_X0Y93_ILOGIC_X0Y94_D;
  wire [0:0] LIOI3_TBYTESRC_X0Y93_ILOGIC_X0Y94_O;
  wire [0:0] LIOI3_TBYTETERM_X0Y113_ILOGIC_X0Y113_D;
  wire [0:0] LIOI3_TBYTETERM_X0Y113_ILOGIC_X0Y113_O;
  wire [0:0] LIOI3_TBYTETERM_X0Y113_ILOGIC_X0Y114_D;
  wire [0:0] LIOI3_TBYTETERM_X0Y113_ILOGIC_X0Y114_O;
  wire [0:0] LIOI3_TBYTETERM_X0Y137_ILOGIC_X0Y137_D;
  wire [0:0] LIOI3_TBYTETERM_X0Y137_ILOGIC_X0Y137_O;
  wire [0:0] LIOI3_TBYTETERM_X0Y137_ILOGIC_X0Y138_D;
  wire [0:0] LIOI3_TBYTETERM_X0Y137_ILOGIC_X0Y138_O;
  wire [0:0] LIOI3_TBYTETERM_X0Y163_ILOGIC_X0Y163_D;
  wire [0:0] LIOI3_TBYTETERM_X0Y163_ILOGIC_X0Y163_O;
  wire [0:0] LIOI3_TBYTETERM_X0Y163_ILOGIC_X0Y164_D;
  wire [0:0] LIOI3_TBYTETERM_X0Y163_ILOGIC_X0Y164_O;
  wire [0:0] LIOI3_TBYTETERM_X0Y187_OLOGIC_X0Y187_D1;
  wire [0:0] LIOI3_TBYTETERM_X0Y187_OLOGIC_X0Y187_OQ;
  wire [0:0] LIOI3_TBYTETERM_X0Y187_OLOGIC_X0Y187_T1;
  wire [0:0] LIOI3_TBYTETERM_X0Y187_OLOGIC_X0Y187_TQ;
  wire [0:0] LIOI3_TBYTETERM_X0Y187_OLOGIC_X0Y188_D1;
  wire [0:0] LIOI3_TBYTETERM_X0Y187_OLOGIC_X0Y188_OQ;
  wire [0:0] LIOI3_TBYTETERM_X0Y187_OLOGIC_X0Y188_T1;
  wire [0:0] LIOI3_TBYTETERM_X0Y187_OLOGIC_X0Y188_TQ;
  wire [0:0] LIOI3_TBYTETERM_X0Y63_ILOGIC_X0Y63_D;
  wire [0:0] LIOI3_TBYTETERM_X0Y63_ILOGIC_X0Y63_O;
  wire [0:0] LIOI3_TBYTETERM_X0Y87_ILOGIC_X0Y87_D;
  wire [0:0] LIOI3_TBYTETERM_X0Y87_ILOGIC_X0Y87_O;
  wire [0:0] LIOI3_TBYTETERM_X0Y87_ILOGIC_X0Y88_D;
  wire [0:0] LIOI3_TBYTETERM_X0Y87_ILOGIC_X0Y88_O;
  wire [0:0] LIOI3_X0Y101_ILOGIC_X0Y101_D;
  wire [0:0] LIOI3_X0Y101_ILOGIC_X0Y101_O;
  wire [0:0] LIOI3_X0Y101_ILOGIC_X0Y102_D;
  wire [0:0] LIOI3_X0Y101_ILOGIC_X0Y102_O;
  wire [0:0] LIOI3_X0Y103_ILOGIC_X0Y103_D;
  wire [0:0] LIOI3_X0Y103_ILOGIC_X0Y103_O;
  wire [0:0] LIOI3_X0Y103_ILOGIC_X0Y104_D;
  wire [0:0] LIOI3_X0Y103_ILOGIC_X0Y104_O;
  wire [0:0] LIOI3_X0Y105_ILOGIC_X0Y105_D;
  wire [0:0] LIOI3_X0Y105_ILOGIC_X0Y105_O;
  wire [0:0] LIOI3_X0Y105_ILOGIC_X0Y106_D;
  wire [0:0] LIOI3_X0Y105_ILOGIC_X0Y106_O;
  wire [0:0] LIOI3_X0Y109_ILOGIC_X0Y109_D;
  wire [0:0] LIOI3_X0Y109_ILOGIC_X0Y109_O;
  wire [0:0] LIOI3_X0Y109_ILOGIC_X0Y110_D;
  wire [0:0] LIOI3_X0Y109_ILOGIC_X0Y110_O;
  wire [0:0] LIOI3_X0Y111_ILOGIC_X0Y111_D;
  wire [0:0] LIOI3_X0Y111_ILOGIC_X0Y111_O;
  wire [0:0] LIOI3_X0Y111_ILOGIC_X0Y112_D;
  wire [0:0] LIOI3_X0Y111_ILOGIC_X0Y112_O;
  wire [0:0] LIOI3_X0Y115_ILOGIC_X0Y115_D;
  wire [0:0] LIOI3_X0Y115_ILOGIC_X0Y115_O;
  wire [0:0] LIOI3_X0Y115_ILOGIC_X0Y116_D;
  wire [0:0] LIOI3_X0Y115_ILOGIC_X0Y116_O;
  wire [0:0] LIOI3_X0Y117_ILOGIC_X0Y117_D;
  wire [0:0] LIOI3_X0Y117_ILOGIC_X0Y117_O;
  wire [0:0] LIOI3_X0Y117_ILOGIC_X0Y118_D;
  wire [0:0] LIOI3_X0Y117_ILOGIC_X0Y118_O;
  wire [0:0] LIOI3_X0Y121_ILOGIC_X0Y121_D;
  wire [0:0] LIOI3_X0Y121_ILOGIC_X0Y121_O;
  wire [0:0] LIOI3_X0Y121_ILOGIC_X0Y122_D;
  wire [0:0] LIOI3_X0Y121_ILOGIC_X0Y122_O;
  wire [0:0] LIOI3_X0Y123_ILOGIC_X0Y123_D;
  wire [0:0] LIOI3_X0Y123_ILOGIC_X0Y123_O;
  wire [0:0] LIOI3_X0Y123_ILOGIC_X0Y124_D;
  wire [0:0] LIOI3_X0Y123_ILOGIC_X0Y124_O;
  wire [0:0] LIOI3_X0Y125_ILOGIC_X0Y125_D;
  wire [0:0] LIOI3_X0Y125_ILOGIC_X0Y125_O;
  wire [0:0] LIOI3_X0Y125_ILOGIC_X0Y126_D;
  wire [0:0] LIOI3_X0Y125_ILOGIC_X0Y126_O;
  wire [0:0] LIOI3_X0Y127_ILOGIC_X0Y127_D;
  wire [0:0] LIOI3_X0Y127_ILOGIC_X0Y127_O;
  wire [0:0] LIOI3_X0Y127_ILOGIC_X0Y128_D;
  wire [0:0] LIOI3_X0Y127_ILOGIC_X0Y128_O;
  wire [0:0] LIOI3_X0Y129_ILOGIC_X0Y129_D;
  wire [0:0] LIOI3_X0Y129_ILOGIC_X0Y129_O;
  wire [0:0] LIOI3_X0Y129_ILOGIC_X0Y130_D;
  wire [0:0] LIOI3_X0Y129_ILOGIC_X0Y130_O;
  wire [0:0] LIOI3_X0Y133_ILOGIC_X0Y133_D;
  wire [0:0] LIOI3_X0Y133_ILOGIC_X0Y133_O;
  wire [0:0] LIOI3_X0Y133_ILOGIC_X0Y134_D;
  wire [0:0] LIOI3_X0Y133_ILOGIC_X0Y134_O;
  wire [0:0] LIOI3_X0Y135_ILOGIC_X0Y135_D;
  wire [0:0] LIOI3_X0Y135_ILOGIC_X0Y135_O;
  wire [0:0] LIOI3_X0Y135_ILOGIC_X0Y136_D;
  wire [0:0] LIOI3_X0Y135_ILOGIC_X0Y136_O;
  wire [0:0] LIOI3_X0Y139_ILOGIC_X0Y139_D;
  wire [0:0] LIOI3_X0Y139_ILOGIC_X0Y139_O;
  wire [0:0] LIOI3_X0Y139_ILOGIC_X0Y140_D;
  wire [0:0] LIOI3_X0Y139_ILOGIC_X0Y140_O;
  wire [0:0] LIOI3_X0Y141_ILOGIC_X0Y141_D;
  wire [0:0] LIOI3_X0Y141_ILOGIC_X0Y141_O;
  wire [0:0] LIOI3_X0Y141_ILOGIC_X0Y142_D;
  wire [0:0] LIOI3_X0Y141_ILOGIC_X0Y142_O;
  wire [0:0] LIOI3_X0Y145_ILOGIC_X0Y145_D;
  wire [0:0] LIOI3_X0Y145_ILOGIC_X0Y145_O;
  wire [0:0] LIOI3_X0Y145_ILOGIC_X0Y146_D;
  wire [0:0] LIOI3_X0Y145_ILOGIC_X0Y146_O;
  wire [0:0] LIOI3_X0Y147_ILOGIC_X0Y147_D;
  wire [0:0] LIOI3_X0Y147_ILOGIC_X0Y147_O;
  wire [0:0] LIOI3_X0Y151_ILOGIC_X0Y151_D;
  wire [0:0] LIOI3_X0Y151_ILOGIC_X0Y151_O;
  wire [0:0] LIOI3_X0Y151_ILOGIC_X0Y152_D;
  wire [0:0] LIOI3_X0Y151_ILOGIC_X0Y152_O;
  wire [0:0] LIOI3_X0Y153_ILOGIC_X0Y153_D;
  wire [0:0] LIOI3_X0Y153_ILOGIC_X0Y153_O;
  wire [0:0] LIOI3_X0Y153_ILOGIC_X0Y154_D;
  wire [0:0] LIOI3_X0Y153_ILOGIC_X0Y154_O;
  wire [0:0] LIOI3_X0Y155_ILOGIC_X0Y155_D;
  wire [0:0] LIOI3_X0Y155_ILOGIC_X0Y155_O;
  wire [0:0] LIOI3_X0Y155_ILOGIC_X0Y156_D;
  wire [0:0] LIOI3_X0Y155_ILOGIC_X0Y156_O;
  wire [0:0] LIOI3_X0Y159_ILOGIC_X0Y159_D;
  wire [0:0] LIOI3_X0Y159_ILOGIC_X0Y159_O;
  wire [0:0] LIOI3_X0Y159_ILOGIC_X0Y160_D;
  wire [0:0] LIOI3_X0Y159_ILOGIC_X0Y160_O;
  wire [0:0] LIOI3_X0Y161_ILOGIC_X0Y161_D;
  wire [0:0] LIOI3_X0Y161_ILOGIC_X0Y161_O;
  wire [0:0] LIOI3_X0Y161_ILOGIC_X0Y162_D;
  wire [0:0] LIOI3_X0Y161_ILOGIC_X0Y162_O;
  wire [0:0] LIOI3_X0Y165_ILOGIC_X0Y165_D;
  wire [0:0] LIOI3_X0Y165_ILOGIC_X0Y165_O;
  wire [0:0] LIOI3_X0Y165_ILOGIC_X0Y166_D;
  wire [0:0] LIOI3_X0Y165_ILOGIC_X0Y166_O;
  wire [0:0] LIOI3_X0Y171_ILOGIC_X0Y171_D;
  wire [0:0] LIOI3_X0Y171_ILOGIC_X0Y171_O;
  wire [0:0] LIOI3_X0Y171_ILOGIC_X0Y172_D;
  wire [0:0] LIOI3_X0Y171_ILOGIC_X0Y172_O;
  wire [0:0] LIOI3_X0Y173_ILOGIC_X0Y173_D;
  wire [0:0] LIOI3_X0Y173_ILOGIC_X0Y173_O;
  wire [0:0] LIOI3_X0Y173_ILOGIC_X0Y174_D;
  wire [0:0] LIOI3_X0Y173_ILOGIC_X0Y174_O;
  wire [0:0] LIOI3_X0Y175_ILOGIC_X0Y175_D;
  wire [0:0] LIOI3_X0Y175_ILOGIC_X0Y175_O;
  wire [0:0] LIOI3_X0Y175_ILOGIC_X0Y176_D;
  wire [0:0] LIOI3_X0Y175_ILOGIC_X0Y176_O;
  wire [0:0] LIOI3_X0Y177_ILOGIC_X0Y177_D;
  wire [0:0] LIOI3_X0Y177_ILOGIC_X0Y177_O;
  wire [0:0] LIOI3_X0Y177_OLOGIC_X0Y178_D1;
  wire [0:0] LIOI3_X0Y177_OLOGIC_X0Y178_OQ;
  wire [0:0] LIOI3_X0Y177_OLOGIC_X0Y178_T1;
  wire [0:0] LIOI3_X0Y177_OLOGIC_X0Y178_TQ;
  wire [0:0] LIOI3_X0Y179_OLOGIC_X0Y179_D1;
  wire [0:0] LIOI3_X0Y179_OLOGIC_X0Y179_OQ;
  wire [0:0] LIOI3_X0Y179_OLOGIC_X0Y179_T1;
  wire [0:0] LIOI3_X0Y179_OLOGIC_X0Y179_TQ;
  wire [0:0] LIOI3_X0Y179_OLOGIC_X0Y180_D1;
  wire [0:0] LIOI3_X0Y179_OLOGIC_X0Y180_OQ;
  wire [0:0] LIOI3_X0Y179_OLOGIC_X0Y180_T1;
  wire [0:0] LIOI3_X0Y179_OLOGIC_X0Y180_TQ;
  wire [0:0] LIOI3_X0Y183_OLOGIC_X0Y183_D1;
  wire [0:0] LIOI3_X0Y183_OLOGIC_X0Y183_OQ;
  wire [0:0] LIOI3_X0Y183_OLOGIC_X0Y183_T1;
  wire [0:0] LIOI3_X0Y183_OLOGIC_X0Y183_TQ;
  wire [0:0] LIOI3_X0Y183_OLOGIC_X0Y184_D1;
  wire [0:0] LIOI3_X0Y183_OLOGIC_X0Y184_OQ;
  wire [0:0] LIOI3_X0Y183_OLOGIC_X0Y184_T1;
  wire [0:0] LIOI3_X0Y183_OLOGIC_X0Y184_TQ;
  wire [0:0] LIOI3_X0Y185_OLOGIC_X0Y185_D1;
  wire [0:0] LIOI3_X0Y185_OLOGIC_X0Y185_OQ;
  wire [0:0] LIOI3_X0Y185_OLOGIC_X0Y185_T1;
  wire [0:0] LIOI3_X0Y185_OLOGIC_X0Y185_TQ;
  wire [0:0] LIOI3_X0Y185_OLOGIC_X0Y186_D1;
  wire [0:0] LIOI3_X0Y185_OLOGIC_X0Y186_OQ;
  wire [0:0] LIOI3_X0Y185_OLOGIC_X0Y186_T1;
  wire [0:0] LIOI3_X0Y185_OLOGIC_X0Y186_TQ;
  wire [0:0] LIOI3_X0Y189_OLOGIC_X0Y189_D1;
  wire [0:0] LIOI3_X0Y189_OLOGIC_X0Y189_OQ;
  wire [0:0] LIOI3_X0Y189_OLOGIC_X0Y189_T1;
  wire [0:0] LIOI3_X0Y189_OLOGIC_X0Y189_TQ;
  wire [0:0] LIOI3_X0Y189_OLOGIC_X0Y190_D1;
  wire [0:0] LIOI3_X0Y189_OLOGIC_X0Y190_OQ;
  wire [0:0] LIOI3_X0Y189_OLOGIC_X0Y190_T1;
  wire [0:0] LIOI3_X0Y189_OLOGIC_X0Y190_TQ;
  wire [0:0] LIOI3_X0Y191_OLOGIC_X0Y191_D1;
  wire [0:0] LIOI3_X0Y191_OLOGIC_X0Y191_OQ;
  wire [0:0] LIOI3_X0Y191_OLOGIC_X0Y191_T1;
  wire [0:0] LIOI3_X0Y191_OLOGIC_X0Y191_TQ;
  wire [0:0] LIOI3_X0Y191_OLOGIC_X0Y192_D1;
  wire [0:0] LIOI3_X0Y191_OLOGIC_X0Y192_OQ;
  wire [0:0] LIOI3_X0Y191_OLOGIC_X0Y192_T1;
  wire [0:0] LIOI3_X0Y191_OLOGIC_X0Y192_TQ;
  wire [0:0] LIOI3_X0Y195_OLOGIC_X0Y195_D1;
  wire [0:0] LIOI3_X0Y195_OLOGIC_X0Y195_OQ;
  wire [0:0] LIOI3_X0Y195_OLOGIC_X0Y195_T1;
  wire [0:0] LIOI3_X0Y195_OLOGIC_X0Y195_TQ;
  wire [0:0] LIOI3_X0Y195_OLOGIC_X0Y196_D1;
  wire [0:0] LIOI3_X0Y195_OLOGIC_X0Y196_OQ;
  wire [0:0] LIOI3_X0Y195_OLOGIC_X0Y196_T1;
  wire [0:0] LIOI3_X0Y195_OLOGIC_X0Y196_TQ;
  wire [0:0] LIOI3_X0Y197_OLOGIC_X0Y197_D1;
  wire [0:0] LIOI3_X0Y197_OLOGIC_X0Y197_OQ;
  wire [0:0] LIOI3_X0Y197_OLOGIC_X0Y197_T1;
  wire [0:0] LIOI3_X0Y197_OLOGIC_X0Y197_TQ;
  wire [0:0] LIOI3_X0Y197_OLOGIC_X0Y198_D1;
  wire [0:0] LIOI3_X0Y197_OLOGIC_X0Y198_OQ;
  wire [0:0] LIOI3_X0Y197_OLOGIC_X0Y198_T1;
  wire [0:0] LIOI3_X0Y197_OLOGIC_X0Y198_TQ;
  wire [0:0] LIOI3_X0Y51_ILOGIC_X0Y51_D;
  wire [0:0] LIOI3_X0Y51_ILOGIC_X0Y51_O;
  wire [0:0] LIOI3_X0Y51_ILOGIC_X0Y52_D;
  wire [0:0] LIOI3_X0Y51_ILOGIC_X0Y52_O;
  wire [0:0] LIOI3_X0Y53_ILOGIC_X0Y53_D;
  wire [0:0] LIOI3_X0Y53_ILOGIC_X0Y53_O;
  wire [0:0] LIOI3_X0Y53_ILOGIC_X0Y54_D;
  wire [0:0] LIOI3_X0Y53_ILOGIC_X0Y54_O;
  wire [0:0] LIOI3_X0Y55_ILOGIC_X0Y55_D;
  wire [0:0] LIOI3_X0Y55_ILOGIC_X0Y55_O;
  wire [0:0] LIOI3_X0Y55_ILOGIC_X0Y56_D;
  wire [0:0] LIOI3_X0Y55_ILOGIC_X0Y56_O;
  wire [0:0] LIOI3_X0Y59_ILOGIC_X0Y59_D;
  wire [0:0] LIOI3_X0Y59_ILOGIC_X0Y59_O;
  wire [0:0] LIOI3_X0Y59_ILOGIC_X0Y60_D;
  wire [0:0] LIOI3_X0Y59_ILOGIC_X0Y60_O;
  wire [0:0] LIOI3_X0Y61_ILOGIC_X0Y62_D;
  wire [0:0] LIOI3_X0Y61_ILOGIC_X0Y62_O;
  wire [0:0] LIOI3_X0Y65_ILOGIC_X0Y65_D;
  wire [0:0] LIOI3_X0Y65_ILOGIC_X0Y65_O;
  wire [0:0] LIOI3_X0Y65_ILOGIC_X0Y66_D;
  wire [0:0] LIOI3_X0Y65_ILOGIC_X0Y66_O;
  wire [0:0] LIOI3_X0Y67_ILOGIC_X0Y67_D;
  wire [0:0] LIOI3_X0Y67_ILOGIC_X0Y67_O;
  wire [0:0] LIOI3_X0Y67_ILOGIC_X0Y68_D;
  wire [0:0] LIOI3_X0Y67_ILOGIC_X0Y68_O;
  wire [0:0] LIOI3_X0Y71_ILOGIC_X0Y71_D;
  wire [0:0] LIOI3_X0Y71_ILOGIC_X0Y71_O;
  wire [0:0] LIOI3_X0Y71_ILOGIC_X0Y72_D;
  wire [0:0] LIOI3_X0Y71_ILOGIC_X0Y72_O;
  wire [0:0] LIOI3_X0Y73_ILOGIC_X0Y74_D;
  wire [0:0] LIOI3_X0Y73_ILOGIC_X0Y74_O;
  wire [0:0] LIOI3_X0Y75_ILOGIC_X0Y75_D;
  wire [0:0] LIOI3_X0Y75_ILOGIC_X0Y75_O;
  wire [0:0] LIOI3_X0Y75_ILOGIC_X0Y76_D;
  wire [0:0] LIOI3_X0Y75_ILOGIC_X0Y76_O;
  wire [0:0] LIOI3_X0Y77_ILOGIC_X0Y77_D;
  wire [0:0] LIOI3_X0Y77_ILOGIC_X0Y77_O;
  wire [0:0] LIOI3_X0Y77_ILOGIC_X0Y78_D;
  wire [0:0] LIOI3_X0Y77_ILOGIC_X0Y78_O;
  wire [0:0] LIOI3_X0Y79_ILOGIC_X0Y79_D;
  wire [0:0] LIOI3_X0Y79_ILOGIC_X0Y79_O;
  wire [0:0] LIOI3_X0Y79_ILOGIC_X0Y80_D;
  wire [0:0] LIOI3_X0Y79_ILOGIC_X0Y80_O;
  wire [0:0] LIOI3_X0Y83_ILOGIC_X0Y83_D;
  wire [0:0] LIOI3_X0Y83_ILOGIC_X0Y83_O;
  wire [0:0] LIOI3_X0Y83_ILOGIC_X0Y84_D;
  wire [0:0] LIOI3_X0Y83_ILOGIC_X0Y84_O;
  wire [0:0] LIOI3_X0Y85_ILOGIC_X0Y85_D;
  wire [0:0] LIOI3_X0Y85_ILOGIC_X0Y85_O;
  wire [0:0] LIOI3_X0Y85_ILOGIC_X0Y86_D;
  wire [0:0] LIOI3_X0Y85_ILOGIC_X0Y86_O;
  wire [0:0] LIOI3_X0Y89_ILOGIC_X0Y89_D;
  wire [0:0] LIOI3_X0Y89_ILOGIC_X0Y89_O;
  wire [0:0] LIOI3_X0Y89_ILOGIC_X0Y90_D;
  wire [0:0] LIOI3_X0Y89_ILOGIC_X0Y90_O;
  wire [0:0] LIOI3_X0Y91_ILOGIC_X0Y91_D;
  wire [0:0] LIOI3_X0Y91_ILOGIC_X0Y91_O;
  wire [0:0] LIOI3_X0Y91_ILOGIC_X0Y92_D;
  wire [0:0] LIOI3_X0Y91_ILOGIC_X0Y92_O;
  wire [0:0] LIOI3_X0Y95_ILOGIC_X0Y95_D;
  wire [0:0] LIOI3_X0Y95_ILOGIC_X0Y95_O;
  wire [0:0] LIOI3_X0Y95_ILOGIC_X0Y96_D;
  wire [0:0] LIOI3_X0Y95_ILOGIC_X0Y96_O;
  wire [0:0] LIOI3_X0Y97_ILOGIC_X0Y97_D;
  wire [0:0] LIOI3_X0Y97_ILOGIC_X0Y97_O;
  wire [0:0] LIOI3_X0Y97_ILOGIC_X0Y98_D;
  wire [0:0] LIOI3_X0Y97_ILOGIC_X0Y98_O;
  wire [0:0] RIOB33_SING_X105Y100_IOB_X1Y100_I;
  wire [0:0] RIOB33_SING_X105Y149_IOB_X1Y149_O;
  wire [0:0] RIOB33_SING_X105Y150_IOB_X1Y150_I;
  wire [0:0] RIOB33_SING_X105Y199_IOB_X1Y199_O;
  wire [0:0] RIOB33_SING_X105Y50_IOB_X1Y50_O;
  wire [0:0] RIOB33_SING_X105Y99_IOB_X1Y99_O;
  wire [0:0] RIOB33_X105Y101_IOB_X1Y101_I;
  wire [0:0] RIOB33_X105Y101_IOB_X1Y102_I;
  wire [0:0] RIOB33_X105Y103_IOB_X1Y103_I;
  wire [0:0] RIOB33_X105Y103_IOB_X1Y104_I;
  wire [0:0] RIOB33_X105Y105_IOB_X1Y105_I;
  wire [0:0] RIOB33_X105Y105_IOB_X1Y106_I;
  wire [0:0] RIOB33_X105Y107_IOB_X1Y107_I;
  wire [0:0] RIOB33_X105Y107_IOB_X1Y108_I;
  wire [0:0] RIOB33_X105Y109_IOB_X1Y109_I;
  wire [0:0] RIOB33_X105Y109_IOB_X1Y110_I;
  wire [0:0] RIOB33_X105Y111_IOB_X1Y111_I;
  wire [0:0] RIOB33_X105Y111_IOB_X1Y112_I;
  wire [0:0] RIOB33_X105Y113_IOB_X1Y113_I;
  wire [0:0] RIOB33_X105Y113_IOB_X1Y114_I;
  wire [0:0] RIOB33_X105Y115_IOB_X1Y115_I;
  wire [0:0] RIOB33_X105Y115_IOB_X1Y116_I;
  wire [0:0] RIOB33_X105Y117_IOB_X1Y117_I;
  wire [0:0] RIOB33_X105Y117_IOB_X1Y118_I;
  wire [0:0] RIOB33_X105Y119_IOB_X1Y119_I;
  wire [0:0] RIOB33_X105Y119_IOB_X1Y120_I;
  wire [0:0] RIOB33_X105Y121_IOB_X1Y121_I;
  wire [0:0] RIOB33_X105Y121_IOB_X1Y122_I;
  wire [0:0] RIOB33_X105Y123_IOB_X1Y123_I;
  wire [0:0] RIOB33_X105Y123_IOB_X1Y124_I;
  wire [0:0] RIOB33_X105Y125_IOB_X1Y125_I;
  wire [0:0] RIOB33_X105Y125_IOB_X1Y126_I;
  wire [0:0] RIOB33_X105Y127_IOB_X1Y127_O;
  wire [0:0] RIOB33_X105Y127_IOB_X1Y128_O;
  wire [0:0] RIOB33_X105Y129_IOB_X1Y129_O;
  wire [0:0] RIOB33_X105Y129_IOB_X1Y130_O;
  wire [0:0] RIOB33_X105Y131_IOB_X1Y131_O;
  wire [0:0] RIOB33_X105Y131_IOB_X1Y132_O;
  wire [0:0] RIOB33_X105Y133_IOB_X1Y133_O;
  wire [0:0] RIOB33_X105Y133_IOB_X1Y134_O;
  wire [0:0] RIOB33_X105Y135_IOB_X1Y135_O;
  wire [0:0] RIOB33_X105Y135_IOB_X1Y136_O;
  wire [0:0] RIOB33_X105Y137_IOB_X1Y137_O;
  wire [0:0] RIOB33_X105Y137_IOB_X1Y138_O;
  wire [0:0] RIOB33_X105Y139_IOB_X1Y139_O;
  wire [0:0] RIOB33_X105Y139_IOB_X1Y140_O;
  wire [0:0] RIOB33_X105Y141_IOB_X1Y141_O;
  wire [0:0] RIOB33_X105Y141_IOB_X1Y142_O;
  wire [0:0] RIOB33_X105Y143_IOB_X1Y143_O;
  wire [0:0] RIOB33_X105Y143_IOB_X1Y144_O;
  wire [0:0] RIOB33_X105Y145_IOB_X1Y145_O;
  wire [0:0] RIOB33_X105Y145_IOB_X1Y146_O;
  wire [0:0] RIOB33_X105Y147_IOB_X1Y147_O;
  wire [0:0] RIOB33_X105Y147_IOB_X1Y148_O;
  wire [0:0] RIOB33_X105Y151_IOB_X1Y151_I;
  wire [0:0] RIOB33_X105Y151_IOB_X1Y152_I;
  wire [0:0] RIOB33_X105Y153_IOB_X1Y153_I;
  wire [0:0] RIOB33_X105Y153_IOB_X1Y154_I;
  wire [0:0] RIOB33_X105Y155_IOB_X1Y155_I;
  wire [0:0] RIOB33_X105Y155_IOB_X1Y156_I;
  wire [0:0] RIOB33_X105Y157_IOB_X1Y157_I;
  wire [0:0] RIOB33_X105Y157_IOB_X1Y158_I;
  wire [0:0] RIOB33_X105Y159_IOB_X1Y159_I;
  wire [0:0] RIOB33_X105Y159_IOB_X1Y160_I;
  wire [0:0] RIOB33_X105Y161_IOB_X1Y161_I;
  wire [0:0] RIOB33_X105Y161_IOB_X1Y162_I;
  wire [0:0] RIOB33_X105Y163_IOB_X1Y163_I;
  wire [0:0] RIOB33_X105Y163_IOB_X1Y164_I;
  wire [0:0] RIOB33_X105Y165_IOB_X1Y165_I;
  wire [0:0] RIOB33_X105Y165_IOB_X1Y166_I;
  wire [0:0] RIOB33_X105Y167_IOB_X1Y167_I;
  wire [0:0] RIOB33_X105Y167_IOB_X1Y168_I;
  wire [0:0] RIOB33_X105Y169_IOB_X1Y169_I;
  wire [0:0] RIOB33_X105Y169_IOB_X1Y170_I;
  wire [0:0] RIOB33_X105Y171_IOB_X1Y171_I;
  wire [0:0] RIOB33_X105Y171_IOB_X1Y172_I;
  wire [0:0] RIOB33_X105Y173_IOB_X1Y173_O;
  wire [0:0] RIOB33_X105Y173_IOB_X1Y174_O;
  wire [0:0] RIOB33_X105Y175_IOB_X1Y175_O;
  wire [0:0] RIOB33_X105Y175_IOB_X1Y176_O;
  wire [0:0] RIOB33_X105Y177_IOB_X1Y177_O;
  wire [0:0] RIOB33_X105Y177_IOB_X1Y178_O;
  wire [0:0] RIOB33_X105Y179_IOB_X1Y179_O;
  wire [0:0] RIOB33_X105Y179_IOB_X1Y180_O;
  wire [0:0] RIOB33_X105Y181_IOB_X1Y181_O;
  wire [0:0] RIOB33_X105Y181_IOB_X1Y182_O;
  wire [0:0] RIOB33_X105Y183_IOB_X1Y183_O;
  wire [0:0] RIOB33_X105Y183_IOB_X1Y184_O;
  wire [0:0] RIOB33_X105Y185_IOB_X1Y185_O;
  wire [0:0] RIOB33_X105Y185_IOB_X1Y186_O;
  wire [0:0] RIOB33_X105Y187_IOB_X1Y187_O;
  wire [0:0] RIOB33_X105Y187_IOB_X1Y188_O;
  wire [0:0] RIOB33_X105Y189_IOB_X1Y189_O;
  wire [0:0] RIOB33_X105Y189_IOB_X1Y190_O;
  wire [0:0] RIOB33_X105Y191_IOB_X1Y191_O;
  wire [0:0] RIOB33_X105Y191_IOB_X1Y192_O;
  wire [0:0] RIOB33_X105Y193_IOB_X1Y193_O;
  wire [0:0] RIOB33_X105Y193_IOB_X1Y194_O;
  wire [0:0] RIOB33_X105Y195_IOB_X1Y195_O;
  wire [0:0] RIOB33_X105Y195_IOB_X1Y196_O;
  wire [0:0] RIOB33_X105Y197_IOB_X1Y197_O;
  wire [0:0] RIOB33_X105Y197_IOB_X1Y198_O;
  wire [0:0] RIOB33_X105Y51_IOB_X1Y51_O;
  wire [0:0] RIOB33_X105Y51_IOB_X1Y52_O;
  wire [0:0] RIOB33_X105Y53_IOB_X1Y53_O;
  wire [0:0] RIOB33_X105Y53_IOB_X1Y54_O;
  wire [0:0] RIOB33_X105Y55_IOB_X1Y55_O;
  wire [0:0] RIOB33_X105Y55_IOB_X1Y56_O;
  wire [0:0] RIOB33_X105Y57_IOB_X1Y57_O;
  wire [0:0] RIOB33_X105Y57_IOB_X1Y58_O;
  wire [0:0] RIOB33_X105Y59_IOB_X1Y59_O;
  wire [0:0] RIOB33_X105Y59_IOB_X1Y60_O;
  wire [0:0] RIOB33_X105Y61_IOB_X1Y61_O;
  wire [0:0] RIOB33_X105Y61_IOB_X1Y62_O;
  wire [0:0] RIOB33_X105Y63_IOB_X1Y63_O;
  wire [0:0] RIOB33_X105Y63_IOB_X1Y64_O;
  wire [0:0] RIOB33_X105Y65_IOB_X1Y65_O;
  wire [0:0] RIOB33_X105Y65_IOB_X1Y66_O;
  wire [0:0] RIOB33_X105Y67_IOB_X1Y67_O;
  wire [0:0] RIOB33_X105Y67_IOB_X1Y68_O;
  wire [0:0] RIOB33_X105Y69_IOB_X1Y69_O;
  wire [0:0] RIOB33_X105Y69_IOB_X1Y70_O;
  wire [0:0] RIOB33_X105Y71_IOB_X1Y71_O;
  wire [0:0] RIOB33_X105Y71_IOB_X1Y72_O;
  wire [0:0] RIOB33_X105Y73_IOB_X1Y73_O;
  wire [0:0] RIOB33_X105Y73_IOB_X1Y74_O;
  wire [0:0] RIOB33_X105Y75_IOB_X1Y75_O;
  wire [0:0] RIOB33_X105Y75_IOB_X1Y76_O;
  wire [0:0] RIOB33_X105Y77_IOB_X1Y77_O;
  wire [0:0] RIOB33_X105Y77_IOB_X1Y78_O;
  wire [0:0] RIOB33_X105Y79_IOB_X1Y79_O;
  wire [0:0] RIOB33_X105Y79_IOB_X1Y80_O;
  wire [0:0] RIOB33_X105Y81_IOB_X1Y81_O;
  wire [0:0] RIOB33_X105Y81_IOB_X1Y82_O;
  wire [0:0] RIOB33_X105Y83_IOB_X1Y83_O;
  wire [0:0] RIOB33_X105Y83_IOB_X1Y84_O;
  wire [0:0] RIOB33_X105Y85_IOB_X1Y85_O;
  wire [0:0] RIOB33_X105Y85_IOB_X1Y86_O;
  wire [0:0] RIOB33_X105Y87_IOB_X1Y87_O;
  wire [0:0] RIOB33_X105Y87_IOB_X1Y88_O;
  wire [0:0] RIOB33_X105Y89_IOB_X1Y89_O;
  wire [0:0] RIOB33_X105Y89_IOB_X1Y90_O;
  wire [0:0] RIOB33_X105Y91_IOB_X1Y91_O;
  wire [0:0] RIOB33_X105Y91_IOB_X1Y92_O;
  wire [0:0] RIOB33_X105Y93_IOB_X1Y93_O;
  wire [0:0] RIOB33_X105Y93_IOB_X1Y94_O;
  wire [0:0] RIOB33_X105Y95_IOB_X1Y95_O;
  wire [0:0] RIOB33_X105Y95_IOB_X1Y96_O;
  wire [0:0] RIOB33_X105Y97_IOB_X1Y97_O;
  wire [0:0] RIOB33_X105Y97_IOB_X1Y98_O;
  wire [0:0] RIOI3_SING_X105Y100_ILOGIC_X1Y100_D;
  wire [0:0] RIOI3_SING_X105Y100_ILOGIC_X1Y100_O;
  wire [0:0] RIOI3_SING_X105Y149_OLOGIC_X1Y149_D1;
  wire [0:0] RIOI3_SING_X105Y149_OLOGIC_X1Y149_OQ;
  wire [0:0] RIOI3_SING_X105Y149_OLOGIC_X1Y149_T1;
  wire [0:0] RIOI3_SING_X105Y149_OLOGIC_X1Y149_TQ;
  wire [0:0] RIOI3_SING_X105Y150_ILOGIC_X1Y150_D;
  wire [0:0] RIOI3_SING_X105Y150_ILOGIC_X1Y150_O;
  wire [0:0] RIOI3_SING_X105Y199_OLOGIC_X1Y199_D1;
  wire [0:0] RIOI3_SING_X105Y199_OLOGIC_X1Y199_OQ;
  wire [0:0] RIOI3_SING_X105Y199_OLOGIC_X1Y199_T1;
  wire [0:0] RIOI3_SING_X105Y199_OLOGIC_X1Y199_TQ;
  wire [0:0] RIOI3_SING_X105Y50_OLOGIC_X1Y50_D1;
  wire [0:0] RIOI3_SING_X105Y50_OLOGIC_X1Y50_OQ;
  wire [0:0] RIOI3_SING_X105Y50_OLOGIC_X1Y50_T1;
  wire [0:0] RIOI3_SING_X105Y50_OLOGIC_X1Y50_TQ;
  wire [0:0] RIOI3_SING_X105Y99_OLOGIC_X1Y99_D1;
  wire [0:0] RIOI3_SING_X105Y99_OLOGIC_X1Y99_OQ;
  wire [0:0] RIOI3_SING_X105Y99_OLOGIC_X1Y99_T1;
  wire [0:0] RIOI3_SING_X105Y99_OLOGIC_X1Y99_TQ;
  wire [0:0] RIOI3_TBYTESRC_X105Y107_ILOGIC_X1Y107_D;
  wire [0:0] RIOI3_TBYTESRC_X105Y107_ILOGIC_X1Y107_O;
  wire [0:0] RIOI3_TBYTESRC_X105Y107_ILOGIC_X1Y108_D;
  wire [0:0] RIOI3_TBYTESRC_X105Y107_ILOGIC_X1Y108_O;
  wire [0:0] RIOI3_TBYTESRC_X105Y119_ILOGIC_X1Y119_D;
  wire [0:0] RIOI3_TBYTESRC_X105Y119_ILOGIC_X1Y119_O;
  wire [0:0] RIOI3_TBYTESRC_X105Y119_ILOGIC_X1Y120_D;
  wire [0:0] RIOI3_TBYTESRC_X105Y119_ILOGIC_X1Y120_O;
  wire [0:0] RIOI3_TBYTESRC_X105Y131_OLOGIC_X1Y131_D1;
  wire [0:0] RIOI3_TBYTESRC_X105Y131_OLOGIC_X1Y131_OQ;
  wire [0:0] RIOI3_TBYTESRC_X105Y131_OLOGIC_X1Y131_T1;
  wire [0:0] RIOI3_TBYTESRC_X105Y131_OLOGIC_X1Y131_TQ;
  wire [0:0] RIOI3_TBYTESRC_X105Y131_OLOGIC_X1Y132_D1;
  wire [0:0] RIOI3_TBYTESRC_X105Y131_OLOGIC_X1Y132_OQ;
  wire [0:0] RIOI3_TBYTESRC_X105Y131_OLOGIC_X1Y132_T1;
  wire [0:0] RIOI3_TBYTESRC_X105Y131_OLOGIC_X1Y132_TQ;
  wire [0:0] RIOI3_TBYTESRC_X105Y143_OLOGIC_X1Y143_D1;
  wire [0:0] RIOI3_TBYTESRC_X105Y143_OLOGIC_X1Y143_OQ;
  wire [0:0] RIOI3_TBYTESRC_X105Y143_OLOGIC_X1Y143_T1;
  wire [0:0] RIOI3_TBYTESRC_X105Y143_OLOGIC_X1Y143_TQ;
  wire [0:0] RIOI3_TBYTESRC_X105Y143_OLOGIC_X1Y144_D1;
  wire [0:0] RIOI3_TBYTESRC_X105Y143_OLOGIC_X1Y144_OQ;
  wire [0:0] RIOI3_TBYTESRC_X105Y143_OLOGIC_X1Y144_T1;
  wire [0:0] RIOI3_TBYTESRC_X105Y143_OLOGIC_X1Y144_TQ;
  wire [0:0] RIOI3_TBYTESRC_X105Y157_ILOGIC_X1Y157_D;
  wire [0:0] RIOI3_TBYTESRC_X105Y157_ILOGIC_X1Y157_O;
  wire [0:0] RIOI3_TBYTESRC_X105Y157_ILOGIC_X1Y158_D;
  wire [0:0] RIOI3_TBYTESRC_X105Y157_ILOGIC_X1Y158_O;
  wire [0:0] RIOI3_TBYTESRC_X105Y169_ILOGIC_X1Y169_D;
  wire [0:0] RIOI3_TBYTESRC_X105Y169_ILOGIC_X1Y169_O;
  wire [0:0] RIOI3_TBYTESRC_X105Y169_ILOGIC_X1Y170_D;
  wire [0:0] RIOI3_TBYTESRC_X105Y169_ILOGIC_X1Y170_O;
  wire [0:0] RIOI3_TBYTESRC_X105Y181_OLOGIC_X1Y181_D1;
  wire [0:0] RIOI3_TBYTESRC_X105Y181_OLOGIC_X1Y181_OQ;
  wire [0:0] RIOI3_TBYTESRC_X105Y181_OLOGIC_X1Y181_T1;
  wire [0:0] RIOI3_TBYTESRC_X105Y181_OLOGIC_X1Y181_TQ;
  wire [0:0] RIOI3_TBYTESRC_X105Y181_OLOGIC_X1Y182_D1;
  wire [0:0] RIOI3_TBYTESRC_X105Y181_OLOGIC_X1Y182_OQ;
  wire [0:0] RIOI3_TBYTESRC_X105Y181_OLOGIC_X1Y182_T1;
  wire [0:0] RIOI3_TBYTESRC_X105Y181_OLOGIC_X1Y182_TQ;
  wire [0:0] RIOI3_TBYTESRC_X105Y193_OLOGIC_X1Y193_D1;
  wire [0:0] RIOI3_TBYTESRC_X105Y193_OLOGIC_X1Y193_OQ;
  wire [0:0] RIOI3_TBYTESRC_X105Y193_OLOGIC_X1Y193_T1;
  wire [0:0] RIOI3_TBYTESRC_X105Y193_OLOGIC_X1Y193_TQ;
  wire [0:0] RIOI3_TBYTESRC_X105Y193_OLOGIC_X1Y194_D1;
  wire [0:0] RIOI3_TBYTESRC_X105Y193_OLOGIC_X1Y194_OQ;
  wire [0:0] RIOI3_TBYTESRC_X105Y193_OLOGIC_X1Y194_T1;
  wire [0:0] RIOI3_TBYTESRC_X105Y193_OLOGIC_X1Y194_TQ;
  wire [0:0] RIOI3_TBYTESRC_X105Y57_OLOGIC_X1Y57_D1;
  wire [0:0] RIOI3_TBYTESRC_X105Y57_OLOGIC_X1Y57_OQ;
  wire [0:0] RIOI3_TBYTESRC_X105Y57_OLOGIC_X1Y57_T1;
  wire [0:0] RIOI3_TBYTESRC_X105Y57_OLOGIC_X1Y57_TQ;
  wire [0:0] RIOI3_TBYTESRC_X105Y57_OLOGIC_X1Y58_D1;
  wire [0:0] RIOI3_TBYTESRC_X105Y57_OLOGIC_X1Y58_OQ;
  wire [0:0] RIOI3_TBYTESRC_X105Y57_OLOGIC_X1Y58_T1;
  wire [0:0] RIOI3_TBYTESRC_X105Y57_OLOGIC_X1Y58_TQ;
  wire [0:0] RIOI3_TBYTESRC_X105Y69_OLOGIC_X1Y69_D1;
  wire [0:0] RIOI3_TBYTESRC_X105Y69_OLOGIC_X1Y69_OQ;
  wire [0:0] RIOI3_TBYTESRC_X105Y69_OLOGIC_X1Y69_T1;
  wire [0:0] RIOI3_TBYTESRC_X105Y69_OLOGIC_X1Y69_TQ;
  wire [0:0] RIOI3_TBYTESRC_X105Y69_OLOGIC_X1Y70_D1;
  wire [0:0] RIOI3_TBYTESRC_X105Y69_OLOGIC_X1Y70_OQ;
  wire [0:0] RIOI3_TBYTESRC_X105Y69_OLOGIC_X1Y70_T1;
  wire [0:0] RIOI3_TBYTESRC_X105Y69_OLOGIC_X1Y70_TQ;
  wire [0:0] RIOI3_TBYTESRC_X105Y81_OLOGIC_X1Y81_D1;
  wire [0:0] RIOI3_TBYTESRC_X105Y81_OLOGIC_X1Y81_OQ;
  wire [0:0] RIOI3_TBYTESRC_X105Y81_OLOGIC_X1Y81_T1;
  wire [0:0] RIOI3_TBYTESRC_X105Y81_OLOGIC_X1Y81_TQ;
  wire [0:0] RIOI3_TBYTESRC_X105Y81_OLOGIC_X1Y82_D1;
  wire [0:0] RIOI3_TBYTESRC_X105Y81_OLOGIC_X1Y82_OQ;
  wire [0:0] RIOI3_TBYTESRC_X105Y81_OLOGIC_X1Y82_T1;
  wire [0:0] RIOI3_TBYTESRC_X105Y81_OLOGIC_X1Y82_TQ;
  wire [0:0] RIOI3_TBYTESRC_X105Y93_OLOGIC_X1Y93_D1;
  wire [0:0] RIOI3_TBYTESRC_X105Y93_OLOGIC_X1Y93_OQ;
  wire [0:0] RIOI3_TBYTESRC_X105Y93_OLOGIC_X1Y93_T1;
  wire [0:0] RIOI3_TBYTESRC_X105Y93_OLOGIC_X1Y93_TQ;
  wire [0:0] RIOI3_TBYTESRC_X105Y93_OLOGIC_X1Y94_D1;
  wire [0:0] RIOI3_TBYTESRC_X105Y93_OLOGIC_X1Y94_OQ;
  wire [0:0] RIOI3_TBYTESRC_X105Y93_OLOGIC_X1Y94_T1;
  wire [0:0] RIOI3_TBYTESRC_X105Y93_OLOGIC_X1Y94_TQ;
  wire [0:0] RIOI3_TBYTETERM_X105Y113_ILOGIC_X1Y113_D;
  wire [0:0] RIOI3_TBYTETERM_X105Y113_ILOGIC_X1Y113_O;
  wire [0:0] RIOI3_TBYTETERM_X105Y113_ILOGIC_X1Y114_D;
  wire [0:0] RIOI3_TBYTETERM_X105Y113_ILOGIC_X1Y114_O;
  wire [0:0] RIOI3_TBYTETERM_X105Y137_OLOGIC_X1Y137_D1;
  wire [0:0] RIOI3_TBYTETERM_X105Y137_OLOGIC_X1Y137_OQ;
  wire [0:0] RIOI3_TBYTETERM_X105Y137_OLOGIC_X1Y137_T1;
  wire [0:0] RIOI3_TBYTETERM_X105Y137_OLOGIC_X1Y137_TQ;
  wire [0:0] RIOI3_TBYTETERM_X105Y137_OLOGIC_X1Y138_D1;
  wire [0:0] RIOI3_TBYTETERM_X105Y137_OLOGIC_X1Y138_OQ;
  wire [0:0] RIOI3_TBYTETERM_X105Y137_OLOGIC_X1Y138_T1;
  wire [0:0] RIOI3_TBYTETERM_X105Y137_OLOGIC_X1Y138_TQ;
  wire [0:0] RIOI3_TBYTETERM_X105Y163_ILOGIC_X1Y163_D;
  wire [0:0] RIOI3_TBYTETERM_X105Y163_ILOGIC_X1Y163_O;
  wire [0:0] RIOI3_TBYTETERM_X105Y187_OLOGIC_X1Y187_D1;
  wire [0:0] RIOI3_TBYTETERM_X105Y187_OLOGIC_X1Y187_OQ;
  wire [0:0] RIOI3_TBYTETERM_X105Y187_OLOGIC_X1Y187_T1;
  wire [0:0] RIOI3_TBYTETERM_X105Y187_OLOGIC_X1Y187_TQ;
  wire [0:0] RIOI3_TBYTETERM_X105Y187_OLOGIC_X1Y188_D1;
  wire [0:0] RIOI3_TBYTETERM_X105Y187_OLOGIC_X1Y188_OQ;
  wire [0:0] RIOI3_TBYTETERM_X105Y187_OLOGIC_X1Y188_T1;
  wire [0:0] RIOI3_TBYTETERM_X105Y187_OLOGIC_X1Y188_TQ;
  wire [0:0] RIOI3_TBYTETERM_X105Y63_OLOGIC_X1Y63_D1;
  wire [0:0] RIOI3_TBYTETERM_X105Y63_OLOGIC_X1Y63_OQ;
  wire [0:0] RIOI3_TBYTETERM_X105Y63_OLOGIC_X1Y63_T1;
  wire [0:0] RIOI3_TBYTETERM_X105Y63_OLOGIC_X1Y63_TQ;
  wire [0:0] RIOI3_TBYTETERM_X105Y63_OLOGIC_X1Y64_D1;
  wire [0:0] RIOI3_TBYTETERM_X105Y63_OLOGIC_X1Y64_OQ;
  wire [0:0] RIOI3_TBYTETERM_X105Y63_OLOGIC_X1Y64_T1;
  wire [0:0] RIOI3_TBYTETERM_X105Y63_OLOGIC_X1Y64_TQ;
  wire [0:0] RIOI3_TBYTETERM_X105Y87_OLOGIC_X1Y87_D1;
  wire [0:0] RIOI3_TBYTETERM_X105Y87_OLOGIC_X1Y87_OQ;
  wire [0:0] RIOI3_TBYTETERM_X105Y87_OLOGIC_X1Y87_T1;
  wire [0:0] RIOI3_TBYTETERM_X105Y87_OLOGIC_X1Y87_TQ;
  wire [0:0] RIOI3_TBYTETERM_X105Y87_OLOGIC_X1Y88_D1;
  wire [0:0] RIOI3_TBYTETERM_X105Y87_OLOGIC_X1Y88_OQ;
  wire [0:0] RIOI3_TBYTETERM_X105Y87_OLOGIC_X1Y88_T1;
  wire [0:0] RIOI3_TBYTETERM_X105Y87_OLOGIC_X1Y88_TQ;
  wire [0:0] RIOI3_X105Y101_ILOGIC_X1Y101_D;
  wire [0:0] RIOI3_X105Y101_ILOGIC_X1Y101_O;
  wire [0:0] RIOI3_X105Y101_ILOGIC_X1Y102_D;
  wire [0:0] RIOI3_X105Y101_ILOGIC_X1Y102_O;
  wire [0:0] RIOI3_X105Y103_ILOGIC_X1Y103_D;
  wire [0:0] RIOI3_X105Y103_ILOGIC_X1Y103_O;
  wire [0:0] RIOI3_X105Y103_ILOGIC_X1Y104_D;
  wire [0:0] RIOI3_X105Y103_ILOGIC_X1Y104_O;
  wire [0:0] RIOI3_X105Y105_ILOGIC_X1Y105_D;
  wire [0:0] RIOI3_X105Y105_ILOGIC_X1Y105_O;
  wire [0:0] RIOI3_X105Y105_ILOGIC_X1Y106_D;
  wire [0:0] RIOI3_X105Y105_ILOGIC_X1Y106_O;
  wire [0:0] RIOI3_X105Y109_ILOGIC_X1Y109_D;
  wire [0:0] RIOI3_X105Y109_ILOGIC_X1Y109_O;
  wire [0:0] RIOI3_X105Y109_ILOGIC_X1Y110_D;
  wire [0:0] RIOI3_X105Y109_ILOGIC_X1Y110_O;
  wire [0:0] RIOI3_X105Y111_ILOGIC_X1Y111_D;
  wire [0:0] RIOI3_X105Y111_ILOGIC_X1Y111_O;
  wire [0:0] RIOI3_X105Y111_ILOGIC_X1Y112_D;
  wire [0:0] RIOI3_X105Y111_ILOGIC_X1Y112_O;
  wire [0:0] RIOI3_X105Y115_ILOGIC_X1Y115_D;
  wire [0:0] RIOI3_X105Y115_ILOGIC_X1Y115_O;
  wire [0:0] RIOI3_X105Y115_ILOGIC_X1Y116_D;
  wire [0:0] RIOI3_X105Y115_ILOGIC_X1Y116_O;
  wire [0:0] RIOI3_X105Y117_ILOGIC_X1Y117_D;
  wire [0:0] RIOI3_X105Y117_ILOGIC_X1Y117_O;
  wire [0:0] RIOI3_X105Y117_ILOGIC_X1Y118_D;
  wire [0:0] RIOI3_X105Y117_ILOGIC_X1Y118_O;
  wire [0:0] RIOI3_X105Y121_ILOGIC_X1Y121_D;
  wire [0:0] RIOI3_X105Y121_ILOGIC_X1Y121_O;
  wire [0:0] RIOI3_X105Y121_ILOGIC_X1Y122_D;
  wire [0:0] RIOI3_X105Y121_ILOGIC_X1Y122_O;
  wire [0:0] RIOI3_X105Y123_ILOGIC_X1Y123_D;
  wire [0:0] RIOI3_X105Y123_ILOGIC_X1Y123_O;
  wire [0:0] RIOI3_X105Y123_ILOGIC_X1Y124_D;
  wire [0:0] RIOI3_X105Y123_ILOGIC_X1Y124_O;
  wire [0:0] RIOI3_X105Y125_ILOGIC_X1Y125_D;
  wire [0:0] RIOI3_X105Y125_ILOGIC_X1Y125_O;
  wire [0:0] RIOI3_X105Y125_ILOGIC_X1Y126_D;
  wire [0:0] RIOI3_X105Y125_ILOGIC_X1Y126_O;
  wire [0:0] RIOI3_X105Y127_OLOGIC_X1Y127_D1;
  wire [0:0] RIOI3_X105Y127_OLOGIC_X1Y127_OQ;
  wire [0:0] RIOI3_X105Y127_OLOGIC_X1Y127_T1;
  wire [0:0] RIOI3_X105Y127_OLOGIC_X1Y127_TQ;
  wire [0:0] RIOI3_X105Y127_OLOGIC_X1Y128_D1;
  wire [0:0] RIOI3_X105Y127_OLOGIC_X1Y128_OQ;
  wire [0:0] RIOI3_X105Y127_OLOGIC_X1Y128_T1;
  wire [0:0] RIOI3_X105Y127_OLOGIC_X1Y128_TQ;
  wire [0:0] RIOI3_X105Y129_OLOGIC_X1Y129_D1;
  wire [0:0] RIOI3_X105Y129_OLOGIC_X1Y129_OQ;
  wire [0:0] RIOI3_X105Y129_OLOGIC_X1Y129_T1;
  wire [0:0] RIOI3_X105Y129_OLOGIC_X1Y129_TQ;
  wire [0:0] RIOI3_X105Y129_OLOGIC_X1Y130_D1;
  wire [0:0] RIOI3_X105Y129_OLOGIC_X1Y130_OQ;
  wire [0:0] RIOI3_X105Y129_OLOGIC_X1Y130_T1;
  wire [0:0] RIOI3_X105Y129_OLOGIC_X1Y130_TQ;
  wire [0:0] RIOI3_X105Y133_OLOGIC_X1Y133_D1;
  wire [0:0] RIOI3_X105Y133_OLOGIC_X1Y133_OQ;
  wire [0:0] RIOI3_X105Y133_OLOGIC_X1Y133_T1;
  wire [0:0] RIOI3_X105Y133_OLOGIC_X1Y133_TQ;
  wire [0:0] RIOI3_X105Y133_OLOGIC_X1Y134_D1;
  wire [0:0] RIOI3_X105Y133_OLOGIC_X1Y134_OQ;
  wire [0:0] RIOI3_X105Y133_OLOGIC_X1Y134_T1;
  wire [0:0] RIOI3_X105Y133_OLOGIC_X1Y134_TQ;
  wire [0:0] RIOI3_X105Y135_OLOGIC_X1Y135_D1;
  wire [0:0] RIOI3_X105Y135_OLOGIC_X1Y135_OQ;
  wire [0:0] RIOI3_X105Y135_OLOGIC_X1Y135_T1;
  wire [0:0] RIOI3_X105Y135_OLOGIC_X1Y135_TQ;
  wire [0:0] RIOI3_X105Y135_OLOGIC_X1Y136_D1;
  wire [0:0] RIOI3_X105Y135_OLOGIC_X1Y136_OQ;
  wire [0:0] RIOI3_X105Y135_OLOGIC_X1Y136_T1;
  wire [0:0] RIOI3_X105Y135_OLOGIC_X1Y136_TQ;
  wire [0:0] RIOI3_X105Y139_OLOGIC_X1Y139_D1;
  wire [0:0] RIOI3_X105Y139_OLOGIC_X1Y139_OQ;
  wire [0:0] RIOI3_X105Y139_OLOGIC_X1Y139_T1;
  wire [0:0] RIOI3_X105Y139_OLOGIC_X1Y139_TQ;
  wire [0:0] RIOI3_X105Y139_OLOGIC_X1Y140_D1;
  wire [0:0] RIOI3_X105Y139_OLOGIC_X1Y140_OQ;
  wire [0:0] RIOI3_X105Y139_OLOGIC_X1Y140_T1;
  wire [0:0] RIOI3_X105Y139_OLOGIC_X1Y140_TQ;
  wire [0:0] RIOI3_X105Y141_OLOGIC_X1Y141_D1;
  wire [0:0] RIOI3_X105Y141_OLOGIC_X1Y141_OQ;
  wire [0:0] RIOI3_X105Y141_OLOGIC_X1Y141_T1;
  wire [0:0] RIOI3_X105Y141_OLOGIC_X1Y141_TQ;
  wire [0:0] RIOI3_X105Y141_OLOGIC_X1Y142_D1;
  wire [0:0] RIOI3_X105Y141_OLOGIC_X1Y142_OQ;
  wire [0:0] RIOI3_X105Y141_OLOGIC_X1Y142_T1;
  wire [0:0] RIOI3_X105Y141_OLOGIC_X1Y142_TQ;
  wire [0:0] RIOI3_X105Y145_OLOGIC_X1Y145_D1;
  wire [0:0] RIOI3_X105Y145_OLOGIC_X1Y145_OQ;
  wire [0:0] RIOI3_X105Y145_OLOGIC_X1Y145_T1;
  wire [0:0] RIOI3_X105Y145_OLOGIC_X1Y145_TQ;
  wire [0:0] RIOI3_X105Y145_OLOGIC_X1Y146_D1;
  wire [0:0] RIOI3_X105Y145_OLOGIC_X1Y146_OQ;
  wire [0:0] RIOI3_X105Y145_OLOGIC_X1Y146_T1;
  wire [0:0] RIOI3_X105Y145_OLOGIC_X1Y146_TQ;
  wire [0:0] RIOI3_X105Y147_OLOGIC_X1Y147_D1;
  wire [0:0] RIOI3_X105Y147_OLOGIC_X1Y147_OQ;
  wire [0:0] RIOI3_X105Y147_OLOGIC_X1Y147_T1;
  wire [0:0] RIOI3_X105Y147_OLOGIC_X1Y147_TQ;
  wire [0:0] RIOI3_X105Y147_OLOGIC_X1Y148_D1;
  wire [0:0] RIOI3_X105Y147_OLOGIC_X1Y148_OQ;
  wire [0:0] RIOI3_X105Y147_OLOGIC_X1Y148_T1;
  wire [0:0] RIOI3_X105Y147_OLOGIC_X1Y148_TQ;
  wire [0:0] RIOI3_X105Y151_ILOGIC_X1Y151_D;
  wire [0:0] RIOI3_X105Y151_ILOGIC_X1Y151_O;
  wire [0:0] RIOI3_X105Y151_ILOGIC_X1Y152_D;
  wire [0:0] RIOI3_X105Y151_ILOGIC_X1Y152_O;
  wire [0:0] RIOI3_X105Y153_ILOGIC_X1Y153_D;
  wire [0:0] RIOI3_X105Y153_ILOGIC_X1Y153_O;
  wire [0:0] RIOI3_X105Y153_ILOGIC_X1Y154_D;
  wire [0:0] RIOI3_X105Y153_ILOGIC_X1Y154_O;
  wire [0:0] RIOI3_X105Y155_ILOGIC_X1Y155_D;
  wire [0:0] RIOI3_X105Y155_ILOGIC_X1Y155_O;
  wire [0:0] RIOI3_X105Y155_ILOGIC_X1Y156_D;
  wire [0:0] RIOI3_X105Y155_ILOGIC_X1Y156_O;
  wire [0:0] RIOI3_X105Y159_ILOGIC_X1Y159_D;
  wire [0:0] RIOI3_X105Y159_ILOGIC_X1Y159_O;
  wire [0:0] RIOI3_X105Y159_ILOGIC_X1Y160_D;
  wire [0:0] RIOI3_X105Y159_ILOGIC_X1Y160_O;
  wire [0:0] RIOI3_X105Y161_ILOGIC_X1Y161_D;
  wire [0:0] RIOI3_X105Y161_ILOGIC_X1Y161_O;
  wire [0:0] RIOI3_X105Y165_ILOGIC_X1Y165_D;
  wire [0:0] RIOI3_X105Y165_ILOGIC_X1Y165_O;
  wire [0:0] RIOI3_X105Y165_ILOGIC_X1Y166_D;
  wire [0:0] RIOI3_X105Y165_ILOGIC_X1Y166_O;
  wire [0:0] RIOI3_X105Y167_ILOGIC_X1Y167_D;
  wire [0:0] RIOI3_X105Y167_ILOGIC_X1Y167_O;
  wire [0:0] RIOI3_X105Y167_ILOGIC_X1Y168_D;
  wire [0:0] RIOI3_X105Y167_ILOGIC_X1Y168_O;
  wire [0:0] RIOI3_X105Y171_ILOGIC_X1Y171_D;
  wire [0:0] RIOI3_X105Y171_ILOGIC_X1Y171_O;
  wire [0:0] RIOI3_X105Y171_ILOGIC_X1Y172_D;
  wire [0:0] RIOI3_X105Y171_ILOGIC_X1Y172_O;
  wire [0:0] RIOI3_X105Y173_OLOGIC_X1Y173_D1;
  wire [0:0] RIOI3_X105Y173_OLOGIC_X1Y173_OQ;
  wire [0:0] RIOI3_X105Y173_OLOGIC_X1Y173_T1;
  wire [0:0] RIOI3_X105Y173_OLOGIC_X1Y173_TQ;
  wire [0:0] RIOI3_X105Y173_OLOGIC_X1Y174_D1;
  wire [0:0] RIOI3_X105Y173_OLOGIC_X1Y174_OQ;
  wire [0:0] RIOI3_X105Y173_OLOGIC_X1Y174_T1;
  wire [0:0] RIOI3_X105Y173_OLOGIC_X1Y174_TQ;
  wire [0:0] RIOI3_X105Y175_OLOGIC_X1Y175_D1;
  wire [0:0] RIOI3_X105Y175_OLOGIC_X1Y175_OQ;
  wire [0:0] RIOI3_X105Y175_OLOGIC_X1Y175_T1;
  wire [0:0] RIOI3_X105Y175_OLOGIC_X1Y175_TQ;
  wire [0:0] RIOI3_X105Y175_OLOGIC_X1Y176_D1;
  wire [0:0] RIOI3_X105Y175_OLOGIC_X1Y176_OQ;
  wire [0:0] RIOI3_X105Y175_OLOGIC_X1Y176_T1;
  wire [0:0] RIOI3_X105Y175_OLOGIC_X1Y176_TQ;
  wire [0:0] RIOI3_X105Y177_OLOGIC_X1Y177_D1;
  wire [0:0] RIOI3_X105Y177_OLOGIC_X1Y177_OQ;
  wire [0:0] RIOI3_X105Y177_OLOGIC_X1Y177_T1;
  wire [0:0] RIOI3_X105Y177_OLOGIC_X1Y177_TQ;
  wire [0:0] RIOI3_X105Y177_OLOGIC_X1Y178_D1;
  wire [0:0] RIOI3_X105Y177_OLOGIC_X1Y178_OQ;
  wire [0:0] RIOI3_X105Y177_OLOGIC_X1Y178_T1;
  wire [0:0] RIOI3_X105Y177_OLOGIC_X1Y178_TQ;
  wire [0:0] RIOI3_X105Y179_OLOGIC_X1Y179_D1;
  wire [0:0] RIOI3_X105Y179_OLOGIC_X1Y179_OQ;
  wire [0:0] RIOI3_X105Y179_OLOGIC_X1Y179_T1;
  wire [0:0] RIOI3_X105Y179_OLOGIC_X1Y179_TQ;
  wire [0:0] RIOI3_X105Y179_OLOGIC_X1Y180_D1;
  wire [0:0] RIOI3_X105Y179_OLOGIC_X1Y180_OQ;
  wire [0:0] RIOI3_X105Y179_OLOGIC_X1Y180_T1;
  wire [0:0] RIOI3_X105Y179_OLOGIC_X1Y180_TQ;
  wire [0:0] RIOI3_X105Y183_OLOGIC_X1Y183_D1;
  wire [0:0] RIOI3_X105Y183_OLOGIC_X1Y183_OQ;
  wire [0:0] RIOI3_X105Y183_OLOGIC_X1Y183_T1;
  wire [0:0] RIOI3_X105Y183_OLOGIC_X1Y183_TQ;
  wire [0:0] RIOI3_X105Y183_OLOGIC_X1Y184_D1;
  wire [0:0] RIOI3_X105Y183_OLOGIC_X1Y184_OQ;
  wire [0:0] RIOI3_X105Y183_OLOGIC_X1Y184_T1;
  wire [0:0] RIOI3_X105Y183_OLOGIC_X1Y184_TQ;
  wire [0:0] RIOI3_X105Y185_OLOGIC_X1Y185_D1;
  wire [0:0] RIOI3_X105Y185_OLOGIC_X1Y185_OQ;
  wire [0:0] RIOI3_X105Y185_OLOGIC_X1Y185_T1;
  wire [0:0] RIOI3_X105Y185_OLOGIC_X1Y185_TQ;
  wire [0:0] RIOI3_X105Y185_OLOGIC_X1Y186_D1;
  wire [0:0] RIOI3_X105Y185_OLOGIC_X1Y186_OQ;
  wire [0:0] RIOI3_X105Y185_OLOGIC_X1Y186_T1;
  wire [0:0] RIOI3_X105Y185_OLOGIC_X1Y186_TQ;
  wire [0:0] RIOI3_X105Y189_OLOGIC_X1Y189_D1;
  wire [0:0] RIOI3_X105Y189_OLOGIC_X1Y189_OQ;
  wire [0:0] RIOI3_X105Y189_OLOGIC_X1Y189_T1;
  wire [0:0] RIOI3_X105Y189_OLOGIC_X1Y189_TQ;
  wire [0:0] RIOI3_X105Y189_OLOGIC_X1Y190_D1;
  wire [0:0] RIOI3_X105Y189_OLOGIC_X1Y190_OQ;
  wire [0:0] RIOI3_X105Y189_OLOGIC_X1Y190_T1;
  wire [0:0] RIOI3_X105Y189_OLOGIC_X1Y190_TQ;
  wire [0:0] RIOI3_X105Y191_OLOGIC_X1Y191_D1;
  wire [0:0] RIOI3_X105Y191_OLOGIC_X1Y191_OQ;
  wire [0:0] RIOI3_X105Y191_OLOGIC_X1Y191_T1;
  wire [0:0] RIOI3_X105Y191_OLOGIC_X1Y191_TQ;
  wire [0:0] RIOI3_X105Y191_OLOGIC_X1Y192_D1;
  wire [0:0] RIOI3_X105Y191_OLOGIC_X1Y192_OQ;
  wire [0:0] RIOI3_X105Y191_OLOGIC_X1Y192_T1;
  wire [0:0] RIOI3_X105Y191_OLOGIC_X1Y192_TQ;
  wire [0:0] RIOI3_X105Y195_OLOGIC_X1Y195_D1;
  wire [0:0] RIOI3_X105Y195_OLOGIC_X1Y195_OQ;
  wire [0:0] RIOI3_X105Y195_OLOGIC_X1Y195_T1;
  wire [0:0] RIOI3_X105Y195_OLOGIC_X1Y195_TQ;
  wire [0:0] RIOI3_X105Y195_OLOGIC_X1Y196_D1;
  wire [0:0] RIOI3_X105Y195_OLOGIC_X1Y196_OQ;
  wire [0:0] RIOI3_X105Y195_OLOGIC_X1Y196_T1;
  wire [0:0] RIOI3_X105Y195_OLOGIC_X1Y196_TQ;
  wire [0:0] RIOI3_X105Y197_OLOGIC_X1Y197_D1;
  wire [0:0] RIOI3_X105Y197_OLOGIC_X1Y197_OQ;
  wire [0:0] RIOI3_X105Y197_OLOGIC_X1Y197_T1;
  wire [0:0] RIOI3_X105Y197_OLOGIC_X1Y197_TQ;
  wire [0:0] RIOI3_X105Y197_OLOGIC_X1Y198_D1;
  wire [0:0] RIOI3_X105Y197_OLOGIC_X1Y198_OQ;
  wire [0:0] RIOI3_X105Y197_OLOGIC_X1Y198_T1;
  wire [0:0] RIOI3_X105Y197_OLOGIC_X1Y198_TQ;
  wire [0:0] RIOI3_X105Y51_OLOGIC_X1Y51_D1;
  wire [0:0] RIOI3_X105Y51_OLOGIC_X1Y51_OQ;
  wire [0:0] RIOI3_X105Y51_OLOGIC_X1Y51_T1;
  wire [0:0] RIOI3_X105Y51_OLOGIC_X1Y51_TQ;
  wire [0:0] RIOI3_X105Y51_OLOGIC_X1Y52_D1;
  wire [0:0] RIOI3_X105Y51_OLOGIC_X1Y52_OQ;
  wire [0:0] RIOI3_X105Y51_OLOGIC_X1Y52_T1;
  wire [0:0] RIOI3_X105Y51_OLOGIC_X1Y52_TQ;
  wire [0:0] RIOI3_X105Y53_OLOGIC_X1Y53_D1;
  wire [0:0] RIOI3_X105Y53_OLOGIC_X1Y53_OQ;
  wire [0:0] RIOI3_X105Y53_OLOGIC_X1Y53_T1;
  wire [0:0] RIOI3_X105Y53_OLOGIC_X1Y53_TQ;
  wire [0:0] RIOI3_X105Y53_OLOGIC_X1Y54_D1;
  wire [0:0] RIOI3_X105Y53_OLOGIC_X1Y54_OQ;
  wire [0:0] RIOI3_X105Y53_OLOGIC_X1Y54_T1;
  wire [0:0] RIOI3_X105Y53_OLOGIC_X1Y54_TQ;
  wire [0:0] RIOI3_X105Y55_OLOGIC_X1Y55_D1;
  wire [0:0] RIOI3_X105Y55_OLOGIC_X1Y55_OQ;
  wire [0:0] RIOI3_X105Y55_OLOGIC_X1Y55_T1;
  wire [0:0] RIOI3_X105Y55_OLOGIC_X1Y55_TQ;
  wire [0:0] RIOI3_X105Y55_OLOGIC_X1Y56_D1;
  wire [0:0] RIOI3_X105Y55_OLOGIC_X1Y56_OQ;
  wire [0:0] RIOI3_X105Y55_OLOGIC_X1Y56_T1;
  wire [0:0] RIOI3_X105Y55_OLOGIC_X1Y56_TQ;
  wire [0:0] RIOI3_X105Y59_OLOGIC_X1Y59_D1;
  wire [0:0] RIOI3_X105Y59_OLOGIC_X1Y59_OQ;
  wire [0:0] RIOI3_X105Y59_OLOGIC_X1Y59_T1;
  wire [0:0] RIOI3_X105Y59_OLOGIC_X1Y59_TQ;
  wire [0:0] RIOI3_X105Y59_OLOGIC_X1Y60_D1;
  wire [0:0] RIOI3_X105Y59_OLOGIC_X1Y60_OQ;
  wire [0:0] RIOI3_X105Y59_OLOGIC_X1Y60_T1;
  wire [0:0] RIOI3_X105Y59_OLOGIC_X1Y60_TQ;
  wire [0:0] RIOI3_X105Y61_OLOGIC_X1Y61_D1;
  wire [0:0] RIOI3_X105Y61_OLOGIC_X1Y61_OQ;
  wire [0:0] RIOI3_X105Y61_OLOGIC_X1Y61_T1;
  wire [0:0] RIOI3_X105Y61_OLOGIC_X1Y61_TQ;
  wire [0:0] RIOI3_X105Y61_OLOGIC_X1Y62_D1;
  wire [0:0] RIOI3_X105Y61_OLOGIC_X1Y62_OQ;
  wire [0:0] RIOI3_X105Y61_OLOGIC_X1Y62_T1;
  wire [0:0] RIOI3_X105Y61_OLOGIC_X1Y62_TQ;
  wire [0:0] RIOI3_X105Y65_OLOGIC_X1Y65_D1;
  wire [0:0] RIOI3_X105Y65_OLOGIC_X1Y65_OQ;
  wire [0:0] RIOI3_X105Y65_OLOGIC_X1Y65_T1;
  wire [0:0] RIOI3_X105Y65_OLOGIC_X1Y65_TQ;
  wire [0:0] RIOI3_X105Y65_OLOGIC_X1Y66_D1;
  wire [0:0] RIOI3_X105Y65_OLOGIC_X1Y66_OQ;
  wire [0:0] RIOI3_X105Y65_OLOGIC_X1Y66_T1;
  wire [0:0] RIOI3_X105Y65_OLOGIC_X1Y66_TQ;
  wire [0:0] RIOI3_X105Y67_OLOGIC_X1Y67_D1;
  wire [0:0] RIOI3_X105Y67_OLOGIC_X1Y67_OQ;
  wire [0:0] RIOI3_X105Y67_OLOGIC_X1Y67_T1;
  wire [0:0] RIOI3_X105Y67_OLOGIC_X1Y67_TQ;
  wire [0:0] RIOI3_X105Y67_OLOGIC_X1Y68_D1;
  wire [0:0] RIOI3_X105Y67_OLOGIC_X1Y68_OQ;
  wire [0:0] RIOI3_X105Y67_OLOGIC_X1Y68_T1;
  wire [0:0] RIOI3_X105Y67_OLOGIC_X1Y68_TQ;
  wire [0:0] RIOI3_X105Y71_OLOGIC_X1Y71_D1;
  wire [0:0] RIOI3_X105Y71_OLOGIC_X1Y71_OQ;
  wire [0:0] RIOI3_X105Y71_OLOGIC_X1Y71_T1;
  wire [0:0] RIOI3_X105Y71_OLOGIC_X1Y71_TQ;
  wire [0:0] RIOI3_X105Y71_OLOGIC_X1Y72_D1;
  wire [0:0] RIOI3_X105Y71_OLOGIC_X1Y72_OQ;
  wire [0:0] RIOI3_X105Y71_OLOGIC_X1Y72_T1;
  wire [0:0] RIOI3_X105Y71_OLOGIC_X1Y72_TQ;
  wire [0:0] RIOI3_X105Y73_OLOGIC_X1Y73_D1;
  wire [0:0] RIOI3_X105Y73_OLOGIC_X1Y73_OQ;
  wire [0:0] RIOI3_X105Y73_OLOGIC_X1Y73_T1;
  wire [0:0] RIOI3_X105Y73_OLOGIC_X1Y73_TQ;
  wire [0:0] RIOI3_X105Y73_OLOGIC_X1Y74_D1;
  wire [0:0] RIOI3_X105Y73_OLOGIC_X1Y74_OQ;
  wire [0:0] RIOI3_X105Y73_OLOGIC_X1Y74_T1;
  wire [0:0] RIOI3_X105Y73_OLOGIC_X1Y74_TQ;
  wire [0:0] RIOI3_X105Y75_OLOGIC_X1Y75_D1;
  wire [0:0] RIOI3_X105Y75_OLOGIC_X1Y75_OQ;
  wire [0:0] RIOI3_X105Y75_OLOGIC_X1Y75_T1;
  wire [0:0] RIOI3_X105Y75_OLOGIC_X1Y75_TQ;
  wire [0:0] RIOI3_X105Y75_OLOGIC_X1Y76_D1;
  wire [0:0] RIOI3_X105Y75_OLOGIC_X1Y76_OQ;
  wire [0:0] RIOI3_X105Y75_OLOGIC_X1Y76_T1;
  wire [0:0] RIOI3_X105Y75_OLOGIC_X1Y76_TQ;
  wire [0:0] RIOI3_X105Y77_OLOGIC_X1Y77_D1;
  wire [0:0] RIOI3_X105Y77_OLOGIC_X1Y77_OQ;
  wire [0:0] RIOI3_X105Y77_OLOGIC_X1Y77_T1;
  wire [0:0] RIOI3_X105Y77_OLOGIC_X1Y77_TQ;
  wire [0:0] RIOI3_X105Y77_OLOGIC_X1Y78_D1;
  wire [0:0] RIOI3_X105Y77_OLOGIC_X1Y78_OQ;
  wire [0:0] RIOI3_X105Y77_OLOGIC_X1Y78_T1;
  wire [0:0] RIOI3_X105Y77_OLOGIC_X1Y78_TQ;
  wire [0:0] RIOI3_X105Y79_OLOGIC_X1Y79_D1;
  wire [0:0] RIOI3_X105Y79_OLOGIC_X1Y79_OQ;
  wire [0:0] RIOI3_X105Y79_OLOGIC_X1Y79_T1;
  wire [0:0] RIOI3_X105Y79_OLOGIC_X1Y79_TQ;
  wire [0:0] RIOI3_X105Y79_OLOGIC_X1Y80_D1;
  wire [0:0] RIOI3_X105Y79_OLOGIC_X1Y80_OQ;
  wire [0:0] RIOI3_X105Y79_OLOGIC_X1Y80_T1;
  wire [0:0] RIOI3_X105Y79_OLOGIC_X1Y80_TQ;
  wire [0:0] RIOI3_X105Y83_OLOGIC_X1Y83_D1;
  wire [0:0] RIOI3_X105Y83_OLOGIC_X1Y83_OQ;
  wire [0:0] RIOI3_X105Y83_OLOGIC_X1Y83_T1;
  wire [0:0] RIOI3_X105Y83_OLOGIC_X1Y83_TQ;
  wire [0:0] RIOI3_X105Y83_OLOGIC_X1Y84_D1;
  wire [0:0] RIOI3_X105Y83_OLOGIC_X1Y84_OQ;
  wire [0:0] RIOI3_X105Y83_OLOGIC_X1Y84_T1;
  wire [0:0] RIOI3_X105Y83_OLOGIC_X1Y84_TQ;
  wire [0:0] RIOI3_X105Y85_OLOGIC_X1Y85_D1;
  wire [0:0] RIOI3_X105Y85_OLOGIC_X1Y85_OQ;
  wire [0:0] RIOI3_X105Y85_OLOGIC_X1Y85_T1;
  wire [0:0] RIOI3_X105Y85_OLOGIC_X1Y85_TQ;
  wire [0:0] RIOI3_X105Y85_OLOGIC_X1Y86_D1;
  wire [0:0] RIOI3_X105Y85_OLOGIC_X1Y86_OQ;
  wire [0:0] RIOI3_X105Y85_OLOGIC_X1Y86_T1;
  wire [0:0] RIOI3_X105Y85_OLOGIC_X1Y86_TQ;
  wire [0:0] RIOI3_X105Y89_OLOGIC_X1Y89_D1;
  wire [0:0] RIOI3_X105Y89_OLOGIC_X1Y89_OQ;
  wire [0:0] RIOI3_X105Y89_OLOGIC_X1Y89_T1;
  wire [0:0] RIOI3_X105Y89_OLOGIC_X1Y89_TQ;
  wire [0:0] RIOI3_X105Y89_OLOGIC_X1Y90_D1;
  wire [0:0] RIOI3_X105Y89_OLOGIC_X1Y90_OQ;
  wire [0:0] RIOI3_X105Y89_OLOGIC_X1Y90_T1;
  wire [0:0] RIOI3_X105Y89_OLOGIC_X1Y90_TQ;
  wire [0:0] RIOI3_X105Y91_OLOGIC_X1Y91_D1;
  wire [0:0] RIOI3_X105Y91_OLOGIC_X1Y91_OQ;
  wire [0:0] RIOI3_X105Y91_OLOGIC_X1Y91_T1;
  wire [0:0] RIOI3_X105Y91_OLOGIC_X1Y91_TQ;
  wire [0:0] RIOI3_X105Y91_OLOGIC_X1Y92_D1;
  wire [0:0] RIOI3_X105Y91_OLOGIC_X1Y92_OQ;
  wire [0:0] RIOI3_X105Y91_OLOGIC_X1Y92_T1;
  wire [0:0] RIOI3_X105Y91_OLOGIC_X1Y92_TQ;
  wire [0:0] RIOI3_X105Y95_OLOGIC_X1Y95_D1;
  wire [0:0] RIOI3_X105Y95_OLOGIC_X1Y95_OQ;
  wire [0:0] RIOI3_X105Y95_OLOGIC_X1Y95_T1;
  wire [0:0] RIOI3_X105Y95_OLOGIC_X1Y95_TQ;
  wire [0:0] RIOI3_X105Y95_OLOGIC_X1Y96_D1;
  wire [0:0] RIOI3_X105Y95_OLOGIC_X1Y96_OQ;
  wire [0:0] RIOI3_X105Y95_OLOGIC_X1Y96_T1;
  wire [0:0] RIOI3_X105Y95_OLOGIC_X1Y96_TQ;
  wire [0:0] RIOI3_X105Y97_OLOGIC_X1Y97_D1;
  wire [0:0] RIOI3_X105Y97_OLOGIC_X1Y97_OQ;
  wire [0:0] RIOI3_X105Y97_OLOGIC_X1Y97_T1;
  wire [0:0] RIOI3_X105Y97_OLOGIC_X1Y97_TQ;
  wire [0:0] RIOI3_X105Y97_OLOGIC_X1Y98_D1;
  wire [0:0] RIOI3_X105Y97_OLOGIC_X1Y98_OQ;
  wire [0:0] RIOI3_X105Y97_OLOGIC_X1Y98_T1;
  wire [0:0] RIOI3_X105Y97_OLOGIC_X1Y98_TQ;


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y98_SLICE_X0Y98_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y98_SLICE_X0Y98_DO5),
.O6(CLBLL_L_X2Y98_SLICE_X0Y98_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y98_SLICE_X0Y98_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y98_SLICE_X0Y98_CO5),
.O6(CLBLL_L_X2Y98_SLICE_X0Y98_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y98_SLICE_X0Y98_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y98_SLICE_X0Y98_BO5),
.O6(CLBLL_L_X2Y98_SLICE_X0Y98_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000005050500)
  ) CLBLL_L_X2Y98_SLICE_X0Y98_ALUT (
.I0(LIOB33_X0Y53_IOB_X0Y54_I),
.I1(1'b1),
.I2(LIOB33_X0Y95_IOB_X0Y96_I),
.I3(LIOB33_X0Y81_IOB_X0Y82_I),
.I4(LIOB33_X0Y83_IOB_X0Y83_I),
.I5(LIOB33_X0Y55_IOB_X0Y55_I),
.O5(CLBLL_L_X2Y98_SLICE_X0Y98_AO5),
.O6(CLBLL_L_X2Y98_SLICE_X0Y98_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y98_SLICE_X1Y98_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y98_SLICE_X1Y98_DO5),
.O6(CLBLL_L_X2Y98_SLICE_X1Y98_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y98_SLICE_X1Y98_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y98_SLICE_X1Y98_CO5),
.O6(CLBLL_L_X2Y98_SLICE_X1Y98_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y98_SLICE_X1Y98_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y98_SLICE_X1Y98_BO5),
.O6(CLBLL_L_X2Y98_SLICE_X1Y98_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y98_SLICE_X1Y98_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y98_SLICE_X1Y98_AO5),
.O6(CLBLL_L_X2Y98_SLICE_X1Y98_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y102_SLICE_X0Y102_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y102_SLICE_X0Y102_DO5),
.O6(CLBLL_L_X2Y102_SLICE_X0Y102_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y102_SLICE_X0Y102_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y102_SLICE_X0Y102_CO5),
.O6(CLBLL_L_X2Y102_SLICE_X0Y102_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffffffffffffc)
  ) CLBLL_L_X2Y102_SLICE_X0Y102_BLUT (
.I0(1'b1),
.I1(LIOB33_X0Y81_IOB_X0Y82_I),
.I2(LIOB33_X0Y77_IOB_X0Y78_I),
.I3(LIOB33_X0Y55_IOB_X0Y56_I),
.I4(CLBLL_L_X2Y102_SLICE_X0Y102_AO6),
.I5(LIOB33_X0Y59_IOB_X0Y60_I),
.O5(CLBLL_L_X2Y102_SLICE_X0Y102_BO5),
.O6(CLBLL_L_X2Y102_SLICE_X0Y102_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffffffff1ffff)
  ) CLBLL_L_X2Y102_SLICE_X0Y102_ALUT (
.I0(LIOB33_X0Y63_IOB_X0Y63_I),
.I1(LIOB33_X0Y71_IOB_X0Y72_I),
.I2(LIOB33_X0Y75_IOB_X0Y75_I),
.I3(LIOB33_X0Y57_IOB_X0Y58_I),
.I4(LIOB33_X0Y53_IOB_X0Y54_I),
.I5(LIOB33_X0Y79_IOB_X0Y80_I),
.O5(CLBLL_L_X2Y102_SLICE_X0Y102_AO5),
.O6(CLBLL_L_X2Y102_SLICE_X0Y102_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y102_SLICE_X1Y102_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y102_SLICE_X1Y102_DO5),
.O6(CLBLL_L_X2Y102_SLICE_X1Y102_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y102_SLICE_X1Y102_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y102_SLICE_X1Y102_CO5),
.O6(CLBLL_L_X2Y102_SLICE_X1Y102_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y102_SLICE_X1Y102_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y102_SLICE_X1Y102_BO5),
.O6(CLBLL_L_X2Y102_SLICE_X1Y102_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y102_SLICE_X1Y102_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y102_SLICE_X1Y102_AO5),
.O6(CLBLL_L_X2Y102_SLICE_X1Y102_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y136_SLICE_X0Y136_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y136_SLICE_X0Y136_DO5),
.O6(CLBLL_L_X2Y136_SLICE_X0Y136_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y136_SLICE_X0Y136_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y136_SLICE_X0Y136_CO5),
.O6(CLBLL_L_X2Y136_SLICE_X0Y136_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f00000f0f00000)
  ) CLBLL_L_X2Y136_SLICE_X0Y136_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(LIOB33_X0Y109_IOB_X0Y110_I),
.I3(1'b1),
.I4(LIOB33_X0Y135_IOB_X0Y136_I),
.I5(1'b1),
.O5(CLBLL_L_X2Y136_SLICE_X0Y136_BO5),
.O6(CLBLL_L_X2Y136_SLICE_X0Y136_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h7fffffffffffffff)
  ) CLBLL_L_X2Y136_SLICE_X0Y136_ALUT (
.I0(LIOB33_X0Y137_IOB_X0Y138_I),
.I1(LIOB33_X0Y109_IOB_X0Y110_I),
.I2(LIOB33_X0Y135_IOB_X0Y136_I),
.I3(LIOB33_X0Y135_IOB_X0Y135_I),
.I4(LIOB33_X0Y67_IOB_X0Y67_I),
.I5(LIOB33_X0Y137_IOB_X0Y137_I),
.O5(CLBLL_L_X2Y136_SLICE_X0Y136_AO5),
.O6(CLBLL_L_X2Y136_SLICE_X0Y136_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y136_SLICE_X1Y136_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y136_SLICE_X1Y136_DO5),
.O6(CLBLL_L_X2Y136_SLICE_X1Y136_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y136_SLICE_X1Y136_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y136_SLICE_X1Y136_CO5),
.O6(CLBLL_L_X2Y136_SLICE_X1Y136_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y136_SLICE_X1Y136_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y136_SLICE_X1Y136_BO5),
.O6(CLBLL_L_X2Y136_SLICE_X1Y136_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y136_SLICE_X1Y136_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y136_SLICE_X1Y136_AO5),
.O6(CLBLL_L_X2Y136_SLICE_X1Y136_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y146_SLICE_X0Y146_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y146_SLICE_X0Y146_DO5),
.O6(CLBLL_L_X2Y146_SLICE_X0Y146_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y146_SLICE_X0Y146_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y146_SLICE_X0Y146_CO5),
.O6(CLBLL_L_X2Y146_SLICE_X0Y146_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y146_SLICE_X0Y146_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y146_SLICE_X0Y146_BO5),
.O6(CLBLL_L_X2Y146_SLICE_X0Y146_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y146_SLICE_X0Y146_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y146_SLICE_X0Y146_AO5),
.O6(CLBLL_L_X2Y146_SLICE_X0Y146_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y146_SLICE_X1Y146_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y146_SLICE_X1Y146_DO5),
.O6(CLBLL_L_X2Y146_SLICE_X1Y146_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y146_SLICE_X1Y146_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y146_SLICE_X1Y146_CO5),
.O6(CLBLL_L_X2Y146_SLICE_X1Y146_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y146_SLICE_X1Y146_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y146_SLICE_X1Y146_BO5),
.O6(CLBLL_L_X2Y146_SLICE_X1Y146_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h5fff5fffaaaa0000)
  ) CLBLL_L_X2Y146_SLICE_X1Y146_ALUT (
.I0(LIOB33_X0Y75_IOB_X0Y76_I),
.I1(1'b1),
.I2(LIOB33_X0Y89_IOB_X0Y89_I),
.I3(RIOB33_X105Y105_IOB_X1Y106_I),
.I4(LIOB33_X0Y145_IOB_X0Y146_I),
.I5(1'b1),
.O5(CLBLL_L_X2Y146_SLICE_X1Y146_AO5),
.O6(CLBLL_L_X2Y146_SLICE_X1Y146_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y173_SLICE_X0Y173_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y173_SLICE_X0Y173_DO5),
.O6(CLBLL_L_X2Y173_SLICE_X0Y173_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y173_SLICE_X0Y173_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y173_SLICE_X0Y173_CO5),
.O6(CLBLL_L_X2Y173_SLICE_X0Y173_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y173_SLICE_X0Y173_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y173_SLICE_X0Y173_BO5),
.O6(CLBLL_L_X2Y173_SLICE_X0Y173_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'haa00a00000000000)
  ) CLBLL_L_X2Y173_SLICE_X0Y173_ALUT (
.I0(LIOB33_X0Y145_IOB_X0Y145_I),
.I1(1'b1),
.I2(LIOB33_X0Y171_IOB_X0Y172_I),
.I3(LIOB33_X0Y75_IOB_X0Y76_I),
.I4(LIOB33_X0Y173_IOB_X0Y173_I),
.I5(LIOB33_X0Y89_IOB_X0Y89_I),
.O5(CLBLL_L_X2Y173_SLICE_X0Y173_AO5),
.O6(CLBLL_L_X2Y173_SLICE_X0Y173_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y173_SLICE_X1Y173_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y173_SLICE_X1Y173_DO5),
.O6(CLBLL_L_X2Y173_SLICE_X1Y173_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y173_SLICE_X1Y173_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y173_SLICE_X1Y173_CO5),
.O6(CLBLL_L_X2Y173_SLICE_X1Y173_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h4000400088000000)
  ) CLBLL_L_X2Y173_SLICE_X1Y173_BLUT (
.I0(LIOB33_X0Y145_IOB_X0Y145_I),
.I1(LIOB33_X0Y75_IOB_X0Y76_I),
.I2(RIOB33_X105Y107_IOB_X1Y107_I),
.I3(LIOB33_X0Y89_IOB_X0Y89_I),
.I4(LIOB33_X0Y171_IOB_X0Y171_I),
.I5(1'b1),
.O5(CLBLL_L_X2Y173_SLICE_X1Y173_BO5),
.O6(CLBLL_L_X2Y173_SLICE_X1Y173_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h88008000cc00cc00)
  ) CLBLL_L_X2Y173_SLICE_X1Y173_ALUT (
.I0(LIOB33_X0Y145_IOB_X0Y145_I),
.I1(LIOB33_X0Y75_IOB_X0Y76_I),
.I2(LIOB33_X0Y173_IOB_X0Y174_I),
.I3(LIOB33_X0Y89_IOB_X0Y89_I),
.I4(LIOB33_X0Y97_IOB_X0Y98_I),
.I5(1'b1),
.O5(CLBLL_L_X2Y173_SLICE_X1Y173_AO5),
.O6(CLBLL_L_X2Y173_SLICE_X1Y173_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y175_SLICE_X0Y175_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y175_SLICE_X0Y175_DO5),
.O6(CLBLL_L_X2Y175_SLICE_X0Y175_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y175_SLICE_X0Y175_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y175_SLICE_X0Y175_CO5),
.O6(CLBLL_L_X2Y175_SLICE_X0Y175_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y175_SLICE_X0Y175_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y175_SLICE_X0Y175_BO5),
.O6(CLBLL_L_X2Y175_SLICE_X0Y175_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f00000f0f00000)
  ) CLBLL_L_X2Y175_SLICE_X0Y175_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(LIOB33_X0Y137_IOB_X0Y138_I),
.I3(1'b1),
.I4(LIOB33_X0Y135_IOB_X0Y135_I),
.I5(1'b1),
.O5(CLBLL_L_X2Y175_SLICE_X0Y175_AO5),
.O6(CLBLL_L_X2Y175_SLICE_X0Y175_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y175_SLICE_X1Y175_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y175_SLICE_X1Y175_DO5),
.O6(CLBLL_L_X2Y175_SLICE_X1Y175_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y175_SLICE_X1Y175_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y175_SLICE_X1Y175_CO5),
.O6(CLBLL_L_X2Y175_SLICE_X1Y175_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y175_SLICE_X1Y175_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y175_SLICE_X1Y175_BO5),
.O6(CLBLL_L_X2Y175_SLICE_X1Y175_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y175_SLICE_X1Y175_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y175_SLICE_X1Y175_AO5),
.O6(CLBLL_L_X2Y175_SLICE_X1Y175_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X4Y107_SLICE_X4Y107_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y107_SLICE_X4Y107_DO5),
.O6(CLBLL_L_X4Y107_SLICE_X4Y107_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X4Y107_SLICE_X4Y107_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y107_SLICE_X4Y107_CO5),
.O6(CLBLL_L_X4Y107_SLICE_X4Y107_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h000f000f000f000f)
  ) CLBLL_L_X4Y107_SLICE_X4Y107_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(LIOB33_X0Y103_IOB_X0Y103_I),
.I3(LIOB33_X0Y103_IOB_X0Y104_I),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y107_SLICE_X4Y107_BO5),
.O6(CLBLL_L_X4Y107_SLICE_X4Y107_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffafffffffbff)
  ) CLBLL_L_X4Y107_SLICE_X4Y107_ALUT (
.I0(LIOB33_X0Y83_IOB_X0Y84_I),
.I1(LIOB33_X0Y105_IOB_X0Y105_I),
.I2(LIOB33_X0Y95_IOB_X0Y95_I),
.I3(CLBLL_L_X4Y107_SLICE_X4Y107_BO6),
.I4(LIOB33_X0Y85_IOB_X0Y85_I),
.I5(LIOB33_X0Y107_IOB_X0Y107_I),
.O5(CLBLL_L_X4Y107_SLICE_X4Y107_AO5),
.O6(CLBLL_L_X4Y107_SLICE_X4Y107_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X4Y107_SLICE_X5Y107_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y107_SLICE_X5Y107_DO5),
.O6(CLBLL_L_X4Y107_SLICE_X5Y107_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X4Y107_SLICE_X5Y107_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y107_SLICE_X5Y107_CO5),
.O6(CLBLL_L_X4Y107_SLICE_X5Y107_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X4Y107_SLICE_X5Y107_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y107_SLICE_X5Y107_BO5),
.O6(CLBLL_L_X4Y107_SLICE_X5Y107_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X4Y107_SLICE_X5Y107_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y107_SLICE_X5Y107_AO5),
.O6(CLBLL_L_X4Y107_SLICE_X5Y107_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffffffffffefe)
  ) CLBLL_L_X4Y109_SLICE_X4Y109_DLUT (
.I0(LIOB33_X0Y103_IOB_X0Y103_I),
.I1(LIOB33_X0Y93_IOB_X0Y93_I),
.I2(LIOB33_SING_X0Y99_IOB_X0Y99_I),
.I3(1'b1),
.I4(LIOB33_X0Y101_IOB_X0Y101_I),
.I5(LIOB33_X0Y105_IOB_X0Y105_I),
.O5(CLBLL_L_X4Y109_SLICE_X4Y109_DO5),
.O6(CLBLL_L_X4Y109_SLICE_X4Y109_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000003301)
  ) CLBLL_L_X4Y109_SLICE_X4Y109_CLUT (
.I0(LIOB33_X0Y75_IOB_X0Y75_I),
.I1(CLBLL_L_X4Y110_SLICE_X4Y110_AO5),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(LIOB33_X0Y95_IOB_X0Y96_I),
.I4(CLBLL_L_X4Y109_SLICE_X4Y109_BO5),
.I5(CLBLL_L_X4Y109_SLICE_X4Y109_BO6),
.O5(CLBLL_L_X4Y109_SLICE_X4Y109_CO5),
.O6(CLBLL_L_X4Y109_SLICE_X4Y109_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h00ee00ee00ff00f0)
  ) CLBLL_L_X4Y109_SLICE_X4Y109_BLUT (
.I0(LIOB33_X0Y81_IOB_X0Y81_I),
.I1(LIOB33_X0Y79_IOB_X0Y80_I),
.I2(LIOB33_X0Y77_IOB_X0Y78_I),
.I3(LIOB33_X0Y95_IOB_X0Y96_I),
.I4(LIOB33_X0Y79_IOB_X0Y79_I),
.I5(1'b1),
.O5(CLBLL_L_X4Y109_SLICE_X4Y109_BO5),
.O6(CLBLL_L_X4Y109_SLICE_X4Y109_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h5555555500000002)
  ) CLBLL_L_X4Y109_SLICE_X4Y109_ALUT (
.I0(CLBLL_L_X4Y110_SLICE_X4Y110_DO6),
.I1(CLBLM_R_X5Y109_SLICE_X6Y109_AO6),
.I2(CLBLL_L_X2Y136_SLICE_X0Y136_AO6),
.I3(CLBLL_L_X4Y110_SLICE_X4Y110_CO5),
.I4(CLBLL_L_X2Y102_SLICE_X0Y102_BO6),
.I5(1'b1),
.O5(CLBLL_L_X4Y109_SLICE_X4Y109_AO5),
.O6(CLBLL_L_X4Y109_SLICE_X4Y109_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X4Y109_SLICE_X5Y109_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y109_SLICE_X5Y109_DO5),
.O6(CLBLL_L_X4Y109_SLICE_X5Y109_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X4Y109_SLICE_X5Y109_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y109_SLICE_X5Y109_CO5),
.O6(CLBLL_L_X4Y109_SLICE_X5Y109_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X4Y109_SLICE_X5Y109_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y109_SLICE_X5Y109_BO5),
.O6(CLBLL_L_X4Y109_SLICE_X5Y109_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X4Y109_SLICE_X5Y109_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y109_SLICE_X5Y109_AO5),
.O6(CLBLL_L_X4Y109_SLICE_X5Y109_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000100)
  ) CLBLL_L_X4Y110_SLICE_X4Y110_DLUT (
.I0(CLBLM_R_X3Y111_SLICE_X2Y111_AO6),
.I1(CLBLL_L_X2Y98_SLICE_X0Y98_AO6),
.I2(CLBLM_R_X3Y111_SLICE_X3Y111_BO6),
.I3(CLBLL_L_X4Y109_SLICE_X4Y109_CO6),
.I4(CLBLM_R_X3Y110_SLICE_X3Y110_AO5),
.I5(CLBLM_R_X3Y110_SLICE_X3Y110_AO6),
.O5(CLBLL_L_X4Y110_SLICE_X4Y110_DO5),
.O6(CLBLL_L_X4Y110_SLICE_X4Y110_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h33333333fffffffe)
  ) CLBLL_L_X4Y110_SLICE_X4Y110_CLUT (
.I0(LIOB33_X0Y91_IOB_X0Y91_I),
.I1(LIOB33_X0Y83_IOB_X0Y84_I),
.I2(LIOB33_X0Y87_IOB_X0Y88_I),
.I3(CLBLL_L_X4Y109_SLICE_X4Y109_DO6),
.I4(LIOB33_X0Y85_IOB_X0Y86_I),
.I5(1'b1),
.O5(CLBLL_L_X4Y110_SLICE_X4Y110_CO5),
.O6(CLBLL_L_X4Y110_SLICE_X4Y110_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf01eff1fffff0f01)
  ) CLBLL_L_X4Y110_SLICE_X4Y110_BLUT (
.I0(LIOB33_X0Y81_IOB_X0Y81_I),
.I1(LIOB33_X0Y79_IOB_X0Y80_I),
.I2(LIOB33_X0Y109_IOB_X0Y109_I),
.I3(LIOB33_X0Y95_IOB_X0Y96_I),
.I4(LIOB33_X0Y111_IOB_X0Y112_I),
.I5(1'b1),
.O5(CLBLL_L_X4Y110_SLICE_X4Y110_BO5),
.O6(CLBLL_L_X4Y110_SLICE_X4Y110_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f0f0ff0e0e0e0e)
  ) CLBLL_L_X4Y110_SLICE_X4Y110_ALUT (
.I0(LIOB33_X0Y73_IOB_X0Y74_I),
.I1(LIOB33_X0Y71_IOB_X0Y72_I),
.I2(LIOB33_X0Y95_IOB_X0Y96_I),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(LIOB33_X0Y75_IOB_X0Y75_I),
.I5(1'b1),
.O5(CLBLL_L_X4Y110_SLICE_X4Y110_AO5),
.O6(CLBLL_L_X4Y110_SLICE_X4Y110_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X4Y110_SLICE_X5Y110_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y110_SLICE_X5Y110_DO5),
.O6(CLBLL_L_X4Y110_SLICE_X5Y110_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X4Y110_SLICE_X5Y110_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y110_SLICE_X5Y110_CO5),
.O6(CLBLL_L_X4Y110_SLICE_X5Y110_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X4Y110_SLICE_X5Y110_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y110_SLICE_X5Y110_BO5),
.O6(CLBLL_L_X4Y110_SLICE_X5Y110_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X4Y110_SLICE_X5Y110_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y110_SLICE_X5Y110_AO5),
.O6(CLBLL_L_X4Y110_SLICE_X5Y110_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffff8fffff8f8)
  ) CLBLL_L_X4Y111_SLICE_X4Y111_DLUT (
.I0(LIOB33_X0Y111_IOB_X0Y111_I),
.I1(CLBLL_L_X4Y110_SLICE_X4Y110_AO5),
.I2(CLBLL_L_X4Y111_SLICE_X4Y111_AO5),
.I3(LIOB33_X0Y115_IOB_X0Y116_I),
.I4(CLBLM_R_X3Y111_SLICE_X3Y111_AO5),
.I5(CLBLM_R_X3Y110_SLICE_X3Y110_AO6),
.O5(CLBLL_L_X4Y111_SLICE_X4Y111_DO5),
.O6(CLBLL_L_X4Y111_SLICE_X4Y111_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffffffaa03fe)
  ) CLBLL_L_X4Y111_SLICE_X4Y111_CLUT (
.I0(CLBLL_L_X4Y110_SLICE_X4Y110_BO6),
.I1(LIOB33_X0Y77_IOB_X0Y78_I),
.I2(LIOB33_X0Y79_IOB_X0Y79_I),
.I3(LIOB33_X0Y115_IOB_X0Y115_I),
.I4(LIOB33_X0Y95_IOB_X0Y96_I),
.I5(CLBLM_R_X3Y111_SLICE_X3Y111_AO6),
.O5(CLBLL_L_X4Y111_SLICE_X4Y111_CO5),
.O6(CLBLL_L_X4Y111_SLICE_X4Y111_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h00000000f1000000)
  ) CLBLL_L_X4Y111_SLICE_X4Y111_BLUT (
.I0(LIOB33_X0Y61_IOB_X0Y62_I),
.I1(LIOB33_X0Y59_IOB_X0Y60_I),
.I2(LIOB33_X0Y95_IOB_X0Y96_I),
.I3(CLBLL_L_X4Y111_SLICE_X5Y111_AO5),
.I4(CLBLL_L_X4Y111_SLICE_X4Y111_AO6),
.I5(LIOB33_X0Y115_IOB_X0Y116_I),
.O5(CLBLL_L_X4Y111_SLICE_X4Y111_BO5),
.O6(CLBLL_L_X4Y111_SLICE_X4Y111_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0f0001000f0f0101)
  ) CLBLL_L_X4Y111_SLICE_X4Y111_ALUT (
.I0(LIOB33_X0Y59_IOB_X0Y59_I),
.I1(LIOB33_X0Y57_IOB_X0Y58_I),
.I2(LIOB33_X0Y121_IOB_X0Y122_I),
.I3(CLBLM_R_X3Y111_SLICE_X2Y111_AO5),
.I4(LIOB33_X0Y95_IOB_X0Y96_I),
.I5(1'b1),
.O5(CLBLL_L_X4Y111_SLICE_X4Y111_AO5),
.O6(CLBLL_L_X4Y111_SLICE_X4Y111_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0e0e00000e0e0000)
  ) CLBLL_L_X4Y111_SLICE_X5Y111_DLUT (
.I0(LIOB33_X0Y55_IOB_X0Y55_I),
.I1(LIOB33_X0Y53_IOB_X0Y54_I),
.I2(LIOB33_X0Y95_IOB_X0Y96_I),
.I3(1'b1),
.I4(LIOB33_X0Y119_IOB_X0Y119_I),
.I5(1'b1),
.O5(CLBLL_L_X4Y111_SLICE_X5Y111_DO5),
.O6(CLBLL_L_X4Y111_SLICE_X5Y111_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffeaeaffffaaba)
  ) CLBLL_L_X4Y111_SLICE_X5Y111_CLUT (
.I0(CLBLL_L_X4Y111_SLICE_X5Y111_AO6),
.I1(CLBLM_R_X3Y111_SLICE_X3Y111_BO6),
.I2(CLBLL_L_X4Y111_SLICE_X4Y111_BO6),
.I3(CLBLL_L_X4Y112_SLICE_X4Y112_BO6),
.I4(CLBLL_L_X4Y111_SLICE_X5Y111_DO6),
.I5(LIOB33_X0Y117_IOB_X0Y118_I),
.O5(CLBLL_L_X4Y111_SLICE_X5Y111_CO5),
.O6(CLBLL_L_X4Y111_SLICE_X5Y111_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hffccfffeff00fffa)
  ) CLBLL_L_X4Y111_SLICE_X5Y111_BLUT (
.I0(LIOB33_X0Y73_IOB_X0Y74_I),
.I1(CLBLL_L_X4Y112_SLICE_X5Y112_BO6),
.I2(LIOB33_X0Y71_IOB_X0Y72_I),
.I3(LIOB33_X0Y111_IOB_X0Y111_I),
.I4(LIOB33_X0Y95_IOB_X0Y96_I),
.I5(1'b1),
.O5(CLBLL_L_X4Y111_SLICE_X5Y111_BO5),
.O6(CLBLL_L_X4Y111_SLICE_X5Y111_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h3030001033330011)
  ) CLBLL_L_X4Y111_SLICE_X5Y111_ALUT (
.I0(LIOB33_X0Y53_IOB_X0Y54_I),
.I1(LIOB33_X0Y119_IOB_X0Y119_I),
.I2(CLBLM_R_X3Y111_SLICE_X3Y111_DO6),
.I3(LIOB33_X0Y55_IOB_X0Y55_I),
.I4(LIOB33_X0Y95_IOB_X0Y96_I),
.I5(1'b1),
.O5(CLBLL_L_X4Y111_SLICE_X5Y111_AO5),
.O6(CLBLL_L_X4Y111_SLICE_X5Y111_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0011001100000000)
  ) CLBLL_L_X4Y112_SLICE_X4Y112_DLUT (
.I0(CLBLL_L_X4Y112_SLICE_X4Y112_AO6),
.I1(CLBLL_L_X4Y112_SLICE_X5Y112_AO5),
.I2(1'b1),
.I3(CLBLL_L_X4Y111_SLICE_X5Y111_BO5),
.I4(1'b1),
.I5(CLBLM_R_X3Y111_SLICE_X3Y111_AO6),
.O5(CLBLL_L_X4Y112_SLICE_X4Y112_DO5),
.O6(CLBLL_L_X4Y112_SLICE_X4Y112_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h90b099bbffffffff)
  ) CLBLL_L_X4Y112_SLICE_X4Y112_CLUT (
.I0(CLBLL_L_X4Y110_SLICE_X4Y110_AO6),
.I1(LIOB33_X0Y113_IOB_X0Y114_I),
.I2(CLBLL_L_X4Y112_SLICE_X5Y112_BO6),
.I3(CLBLL_L_X4Y112_SLICE_X4Y112_AO5),
.I4(LIOB33_X0Y111_IOB_X0Y112_I),
.I5(CLBLL_L_X4Y111_SLICE_X5Y111_BO5),
.O5(CLBLL_L_X4Y112_SLICE_X4Y112_CO5),
.O6(CLBLL_L_X4Y112_SLICE_X4Y112_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000555555555141)
  ) CLBLL_L_X4Y112_SLICE_X4Y112_BLUT (
.I0(CLBLL_L_X4Y112_SLICE_X4Y112_DO6),
.I1(LIOB33_X0Y113_IOB_X0Y114_I),
.I2(CLBLL_L_X4Y110_SLICE_X4Y110_AO6),
.I3(CLBLM_R_X3Y112_SLICE_X3Y112_AO6),
.I4(LIOB33_X0Y111_IOB_X0Y111_I),
.I5(CLBLL_L_X4Y110_SLICE_X4Y110_AO5),
.O5(CLBLL_L_X4Y112_SLICE_X4Y112_BO5),
.O6(CLBLL_L_X4Y112_SLICE_X4Y112_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hff00fffc0055fc01)
  ) CLBLL_L_X4Y112_SLICE_X4Y112_ALUT (
.I0(CLBLL_L_X4Y112_SLICE_X5Y112_AO5),
.I1(LIOB33_X0Y77_IOB_X0Y78_I),
.I2(LIOB33_X0Y79_IOB_X0Y79_I),
.I3(LIOB33_X0Y115_IOB_X0Y115_I),
.I4(LIOB33_X0Y95_IOB_X0Y96_I),
.I5(1'b1),
.O5(CLBLL_L_X4Y112_SLICE_X4Y112_AO5),
.O6(CLBLL_L_X4Y112_SLICE_X4Y112_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hafafafafefefefff)
  ) CLBLL_L_X4Y112_SLICE_X5Y112_DLUT (
.I0(CLBLM_R_X3Y111_SLICE_X3Y111_BO5),
.I1(LIOB33_X0Y95_IOB_X0Y96_I),
.I2(CLBLL_L_X4Y112_SLICE_X5Y112_AO5),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(LIOB33_X0Y75_IOB_X0Y75_I),
.I5(LIOB33_X0Y113_IOB_X0Y114_I),
.O5(CLBLL_L_X4Y112_SLICE_X5Y112_DO5),
.O6(CLBLL_L_X4Y112_SLICE_X5Y112_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000004)
  ) CLBLL_L_X4Y112_SLICE_X5Y112_CLUT (
.I0(CLBLM_R_X3Y111_SLICE_X3Y111_DO6),
.I1(CLBLL_L_X4Y112_SLICE_X4Y112_AO5),
.I2(CLBLL_L_X4Y111_SLICE_X4Y111_DO6),
.I3(CLBLL_L_X4Y113_SLICE_X5Y113_BO6),
.I4(CLBLL_L_X4Y112_SLICE_X5Y112_DO6),
.I5(CLBLM_R_X5Y112_SLICE_X6Y112_CO6),
.O5(CLBLL_L_X4Y112_SLICE_X5Y112_CO5),
.O6(CLBLL_L_X4Y112_SLICE_X5Y112_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffff0fffffffe)
  ) CLBLL_L_X4Y112_SLICE_X5Y112_BLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(LIOB33_X0Y75_IOB_X0Y75_I),
.I2(CLBLL_L_X4Y112_SLICE_X4Y112_AO6),
.I3(LIOB33_X0Y113_IOB_X0Y114_I),
.I4(CLBLL_L_X4Y112_SLICE_X5Y112_AO6),
.I5(LIOB33_X0Y95_IOB_X0Y96_I),
.O5(CLBLL_L_X4Y112_SLICE_X5Y112_BO5),
.O6(CLBLL_L_X4Y112_SLICE_X5Y112_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f0fffaffff0f5f)
  ) CLBLL_L_X4Y112_SLICE_X5Y112_ALUT (
.I0(LIOB33_X0Y81_IOB_X0Y81_I),
.I1(1'b1),
.I2(LIOB33_X0Y109_IOB_X0Y109_I),
.I3(LIOB33_X0Y79_IOB_X0Y80_I),
.I4(LIOB33_X0Y95_IOB_X0Y96_I),
.I5(1'b1),
.O5(CLBLL_L_X4Y112_SLICE_X5Y112_AO5),
.O6(CLBLL_L_X4Y112_SLICE_X5Y112_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X4Y113_SLICE_X4Y113_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y113_SLICE_X4Y113_DO5),
.O6(CLBLL_L_X4Y113_SLICE_X4Y113_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X4Y113_SLICE_X4Y113_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y113_SLICE_X4Y113_CO5),
.O6(CLBLL_L_X4Y113_SLICE_X4Y113_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X4Y113_SLICE_X4Y113_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y113_SLICE_X4Y113_BO5),
.O6(CLBLL_L_X4Y113_SLICE_X4Y113_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X4Y113_SLICE_X4Y113_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y113_SLICE_X4Y113_AO5),
.O6(CLBLL_L_X4Y113_SLICE_X4Y113_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X4Y113_SLICE_X5Y113_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y113_SLICE_X5Y113_DO5),
.O6(CLBLL_L_X4Y113_SLICE_X5Y113_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X4Y113_SLICE_X5Y113_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y113_SLICE_X5Y113_CO5),
.O6(CLBLL_L_X4Y113_SLICE_X5Y113_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hcfffffffdfffffff)
  ) CLBLL_L_X4Y113_SLICE_X5Y113_BLUT (
.I0(LIOB33_X0Y111_IOB_X0Y111_I),
.I1(CLBLM_R_X3Y111_SLICE_X2Y111_AO5),
.I2(CLBLM_R_X3Y110_SLICE_X3Y110_AO5),
.I3(CLBLL_L_X4Y112_SLICE_X5Y112_AO6),
.I4(LIOB33_X0Y121_IOB_X0Y122_I),
.I5(CLBLL_L_X4Y110_SLICE_X4Y110_AO5),
.O5(CLBLL_L_X4Y113_SLICE_X5Y113_BO5),
.O6(CLBLL_L_X4Y113_SLICE_X5Y113_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffffffffdfff)
  ) CLBLL_L_X4Y113_SLICE_X5Y113_ALUT (
.I0(LIOB33_X0Y119_IOB_X0Y120_I),
.I1(LIOB33_X0Y59_IOB_X0Y60_I),
.I2(LIOB33_X0Y115_IOB_X0Y116_I),
.I3(LIOB33_X0Y115_IOB_X0Y115_I),
.I4(LIOB33_X0Y77_IOB_X0Y78_I),
.I5(LIOB33_X0Y55_IOB_X0Y56_I),
.O5(CLBLL_L_X4Y113_SLICE_X5Y113_AO5),
.O6(CLBLL_L_X4Y113_SLICE_X5Y113_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X4Y141_SLICE_X4Y141_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y141_SLICE_X4Y141_DO5),
.O6(CLBLL_L_X4Y141_SLICE_X4Y141_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X4Y141_SLICE_X4Y141_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y141_SLICE_X4Y141_CO5),
.O6(CLBLL_L_X4Y141_SLICE_X4Y141_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X4Y141_SLICE_X4Y141_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y141_SLICE_X4Y141_BO5),
.O6(CLBLL_L_X4Y141_SLICE_X4Y141_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0f000f000f000f00)
  ) CLBLL_L_X4Y141_SLICE_X4Y141_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(LIOB33_X0Y159_IOB_X0Y160_I),
.I3(LIOB33_X0Y175_IOB_X0Y176_I),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y141_SLICE_X4Y141_AO5),
.O6(CLBLL_L_X4Y141_SLICE_X4Y141_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X4Y141_SLICE_X5Y141_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y141_SLICE_X5Y141_DO5),
.O6(CLBLL_L_X4Y141_SLICE_X5Y141_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X4Y141_SLICE_X5Y141_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y141_SLICE_X5Y141_CO5),
.O6(CLBLL_L_X4Y141_SLICE_X5Y141_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X4Y141_SLICE_X5Y141_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y141_SLICE_X5Y141_BO5),
.O6(CLBLL_L_X4Y141_SLICE_X5Y141_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X4Y141_SLICE_X5Y141_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y141_SLICE_X5Y141_AO5),
.O6(CLBLL_L_X4Y141_SLICE_X5Y141_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X36Y113_SLICE_X54Y113_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X36Y113_SLICE_X54Y113_DO5),
.O6(CLBLL_L_X36Y113_SLICE_X54Y113_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X36Y113_SLICE_X54Y113_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X36Y113_SLICE_X54Y113_CO5),
.O6(CLBLL_L_X36Y113_SLICE_X54Y113_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000555500005554)
  ) CLBLL_L_X36Y113_SLICE_X54Y113_BLUT (
.I0(LIOB33_X0Y157_IOB_X0Y157_I),
.I1(CLBLM_L_X10Y113_SLICE_X12Y113_BO6),
.I2(CLBLM_R_X5Y113_SLICE_X6Y113_CO6),
.I3(LIOB33_X0Y51_IOB_X0Y51_I),
.I4(LIOB33_X0Y157_IOB_X0Y158_I),
.I5(LIOB33_X0Y165_IOB_X0Y166_I),
.O5(CLBLL_L_X36Y113_SLICE_X54Y113_BO5),
.O6(CLBLL_L_X36Y113_SLICE_X54Y113_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h000000000000fffe)
  ) CLBLL_L_X36Y113_SLICE_X54Y113_ALUT (
.I0(LIOB33_X0Y165_IOB_X0Y166_I),
.I1(CLBLM_R_X5Y113_SLICE_X6Y113_CO6),
.I2(LIOB33_X0Y51_IOB_X0Y51_I),
.I3(CLBLM_L_X10Y113_SLICE_X12Y113_BO6),
.I4(LIOB33_X0Y153_IOB_X0Y154_I),
.I5(LIOB33_X0Y155_IOB_X0Y156_I),
.O5(CLBLL_L_X36Y113_SLICE_X54Y113_AO5),
.O6(CLBLL_L_X36Y113_SLICE_X54Y113_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X36Y113_SLICE_X55Y113_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X36Y113_SLICE_X55Y113_DO5),
.O6(CLBLL_L_X36Y113_SLICE_X55Y113_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X36Y113_SLICE_X55Y113_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X36Y113_SLICE_X55Y113_CO5),
.O6(CLBLL_L_X36Y113_SLICE_X55Y113_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X36Y113_SLICE_X55Y113_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X36Y113_SLICE_X55Y113_BO5),
.O6(CLBLL_L_X36Y113_SLICE_X55Y113_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X36Y113_SLICE_X55Y113_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X36Y113_SLICE_X55Y113_AO5),
.O6(CLBLL_L_X36Y113_SLICE_X55Y113_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X100Y113_SLICE_X156Y113_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X100Y113_SLICE_X156Y113_DO5),
.O6(CLBLL_L_X100Y113_SLICE_X156Y113_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X100Y113_SLICE_X156Y113_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X100Y113_SLICE_X156Y113_CO5),
.O6(CLBLL_L_X100Y113_SLICE_X156Y113_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000555500005551)
  ) CLBLL_L_X100Y113_SLICE_X156Y113_BLUT (
.I0(LIOB33_X0Y157_IOB_X0Y157_I),
.I1(CLBLM_R_X5Y111_SLICE_X7Y111_CO6),
.I2(LIOB33_X0Y165_IOB_X0Y165_I),
.I3(CLBLM_L_X8Y113_SLICE_X11Y113_BO6),
.I4(LIOB33_X0Y157_IOB_X0Y158_I),
.I5(RIOB33_X105Y117_IOB_X1Y117_I),
.O5(CLBLL_L_X100Y113_SLICE_X156Y113_BO5),
.O6(CLBLL_L_X100Y113_SLICE_X156Y113_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000555500005551)
  ) CLBLL_L_X100Y113_SLICE_X156Y113_ALUT (
.I0(LIOB33_X0Y153_IOB_X0Y154_I),
.I1(CLBLM_R_X5Y111_SLICE_X7Y111_CO6),
.I2(LIOB33_X0Y165_IOB_X0Y165_I),
.I3(CLBLM_L_X8Y113_SLICE_X11Y113_BO6),
.I4(LIOB33_X0Y155_IOB_X0Y156_I),
.I5(RIOB33_X105Y117_IOB_X1Y117_I),
.O5(CLBLL_L_X100Y113_SLICE_X156Y113_AO5),
.O6(CLBLL_L_X100Y113_SLICE_X156Y113_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X100Y113_SLICE_X157Y113_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X100Y113_SLICE_X157Y113_DO5),
.O6(CLBLL_L_X100Y113_SLICE_X157Y113_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X100Y113_SLICE_X157Y113_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X100Y113_SLICE_X157Y113_CO5),
.O6(CLBLL_L_X100Y113_SLICE_X157Y113_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X100Y113_SLICE_X157Y113_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X100Y113_SLICE_X157Y113_BO5),
.O6(CLBLL_L_X100Y113_SLICE_X157Y113_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X100Y113_SLICE_X157Y113_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X100Y113_SLICE_X157Y113_AO5),
.O6(CLBLL_L_X100Y113_SLICE_X157Y113_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X100Y121_SLICE_X156Y121_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X100Y121_SLICE_X156Y121_DO5),
.O6(CLBLL_L_X100Y121_SLICE_X156Y121_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X100Y121_SLICE_X156Y121_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X100Y121_SLICE_X156Y121_CO5),
.O6(CLBLL_L_X100Y121_SLICE_X156Y121_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0505050505050504)
  ) CLBLL_L_X100Y121_SLICE_X156Y121_BLUT (
.I0(LIOB33_X0Y157_IOB_X0Y157_I),
.I1(CLBLM_R_X5Y111_SLICE_X7Y111_BO6),
.I2(LIOB33_X0Y157_IOB_X0Y158_I),
.I3(CLBLM_L_X10Y113_SLICE_X12Y113_AO6),
.I4(LIOB33_X0Y155_IOB_X0Y155_I),
.I5(RIOB33_X105Y155_IOB_X1Y155_I),
.O5(CLBLL_L_X100Y121_SLICE_X156Y121_BO5),
.O6(CLBLL_L_X100Y121_SLICE_X156Y121_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000055555554)
  ) CLBLL_L_X100Y121_SLICE_X156Y121_ALUT (
.I0(LIOB33_X0Y153_IOB_X0Y154_I),
.I1(CLBLM_R_X5Y111_SLICE_X7Y111_BO6),
.I2(CLBLM_L_X10Y113_SLICE_X12Y113_AO6),
.I3(RIOB33_X105Y155_IOB_X1Y155_I),
.I4(LIOB33_X0Y155_IOB_X0Y155_I),
.I5(LIOB33_X0Y155_IOB_X0Y156_I),
.O5(CLBLL_L_X100Y121_SLICE_X156Y121_AO5),
.O6(CLBLL_L_X100Y121_SLICE_X156Y121_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X100Y121_SLICE_X157Y121_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X100Y121_SLICE_X157Y121_DO5),
.O6(CLBLL_L_X100Y121_SLICE_X157Y121_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X100Y121_SLICE_X157Y121_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X100Y121_SLICE_X157Y121_CO5),
.O6(CLBLL_L_X100Y121_SLICE_X157Y121_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X100Y121_SLICE_X157Y121_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X100Y121_SLICE_X157Y121_BO5),
.O6(CLBLL_L_X100Y121_SLICE_X157Y121_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X100Y121_SLICE_X157Y121_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X100Y121_SLICE_X157Y121_AO5),
.O6(CLBLL_L_X100Y121_SLICE_X157Y121_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X100Y123_SLICE_X156Y123_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X100Y123_SLICE_X156Y123_DO5),
.O6(CLBLL_L_X100Y123_SLICE_X156Y123_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X100Y123_SLICE_X156Y123_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X100Y123_SLICE_X156Y123_CO5),
.O6(CLBLL_L_X100Y123_SLICE_X156Y123_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000555500001111)
  ) CLBLL_L_X100Y123_SLICE_X156Y123_BLUT (
.I0(LIOB33_X0Y153_IOB_X0Y154_I),
.I1(CLBLM_R_X7Y121_SLICE_X8Y121_AO6),
.I2(1'b1),
.I3(1'b1),
.I4(LIOB33_X0Y155_IOB_X0Y156_I),
.I5(1'b1),
.O5(CLBLL_L_X100Y123_SLICE_X156Y123_BO5),
.O6(CLBLL_L_X100Y123_SLICE_X156Y123_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000333300000033)
  ) CLBLL_L_X100Y123_SLICE_X156Y123_ALUT (
.I0(1'b1),
.I1(LIOB33_X0Y157_IOB_X0Y157_I),
.I2(1'b1),
.I3(CLBLM_R_X7Y121_SLICE_X8Y121_AO6),
.I4(LIOB33_X0Y157_IOB_X0Y158_I),
.I5(1'b1),
.O5(CLBLL_L_X100Y123_SLICE_X156Y123_AO5),
.O6(CLBLL_L_X100Y123_SLICE_X156Y123_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X100Y123_SLICE_X157Y123_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X100Y123_SLICE_X157Y123_DO5),
.O6(CLBLL_L_X100Y123_SLICE_X157Y123_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X100Y123_SLICE_X157Y123_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X100Y123_SLICE_X157Y123_CO5),
.O6(CLBLL_L_X100Y123_SLICE_X157Y123_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X100Y123_SLICE_X157Y123_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X100Y123_SLICE_X157Y123_BO5),
.O6(CLBLL_L_X100Y123_SLICE_X157Y123_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X100Y123_SLICE_X157Y123_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X100Y123_SLICE_X157Y123_AO5),
.O6(CLBLL_L_X100Y123_SLICE_X157Y123_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_R_X57Y113_SLICE_X86Y113_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X57Y113_SLICE_X86Y113_DO5),
.O6(CLBLL_R_X57Y113_SLICE_X86Y113_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_R_X57Y113_SLICE_X86Y113_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X57Y113_SLICE_X86Y113_CO5),
.O6(CLBLL_R_X57Y113_SLICE_X86Y113_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000555500005554)
  ) CLBLL_R_X57Y113_SLICE_X86Y113_BLUT (
.I0(LIOB33_X0Y157_IOB_X0Y158_I),
.I1(CLBLM_R_X5Y111_SLICE_X6Y111_BO6),
.I2(LIOB33_X0Y105_IOB_X0Y106_I),
.I3(CLBLM_R_X5Y113_SLICE_X6Y113_BO6),
.I4(LIOB33_X0Y157_IOB_X0Y157_I),
.I5(LIOB33_X0Y117_IOB_X0Y117_I),
.O5(CLBLL_R_X57Y113_SLICE_X86Y113_BO5),
.O6(CLBLL_R_X57Y113_SLICE_X86Y113_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h1111111111111110)
  ) CLBLL_R_X57Y113_SLICE_X86Y113_ALUT (
.I0(LIOB33_X0Y153_IOB_X0Y154_I),
.I1(LIOB33_X0Y155_IOB_X0Y156_I),
.I2(LIOB33_X0Y105_IOB_X0Y106_I),
.I3(CLBLM_R_X5Y111_SLICE_X6Y111_BO6),
.I4(CLBLM_R_X5Y113_SLICE_X6Y113_BO6),
.I5(LIOB33_X0Y117_IOB_X0Y117_I),
.O5(CLBLL_R_X57Y113_SLICE_X86Y113_AO5),
.O6(CLBLL_R_X57Y113_SLICE_X86Y113_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_R_X57Y113_SLICE_X87Y113_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X57Y113_SLICE_X87Y113_DO5),
.O6(CLBLL_R_X57Y113_SLICE_X87Y113_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_R_X57Y113_SLICE_X87Y113_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X57Y113_SLICE_X87Y113_CO5),
.O6(CLBLL_R_X57Y113_SLICE_X87Y113_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_R_X57Y113_SLICE_X87Y113_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X57Y113_SLICE_X87Y113_BO5),
.O6(CLBLL_R_X57Y113_SLICE_X87Y113_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_R_X57Y113_SLICE_X87Y113_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X57Y113_SLICE_X87Y113_AO5),
.O6(CLBLL_R_X57Y113_SLICE_X87Y113_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000ff00f4)
  ) CLBLM_L_X8Y113_SLICE_X10Y113_DLUT (
.I0(CLBLM_R_X5Y113_SLICE_X6Y113_AO6),
.I1(CLBLM_L_X8Y113_SLICE_X11Y113_AO5),
.I2(CLBLM_R_X7Y113_SLICE_X9Y113_CO6),
.I3(LIOB33_X0Y159_IOB_X0Y159_I),
.I4(RIOB33_X105Y167_IOB_X1Y167_I),
.I5(LIOB33_X0Y159_IOB_X0Y160_I),
.O5(CLBLM_L_X8Y113_SLICE_X10Y113_DO5),
.O6(CLBLM_L_X8Y113_SLICE_X10Y113_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000055500000111)
  ) CLBLM_L_X8Y113_SLICE_X10Y113_CLUT (
.I0(LIOB33_X0Y83_IOB_X0Y84_I),
.I1(CLBLM_L_X8Y113_SLICE_X11Y113_AO5),
.I2(LIOB33_X0Y65_IOB_X0Y66_I),
.I3(LIOB33_X0Y71_IOB_X0Y71_I),
.I4(RIOB33_X105Y167_IOB_X1Y167_I),
.I5(CLBLM_R_X5Y113_SLICE_X6Y113_AO6),
.O5(CLBLM_L_X8Y113_SLICE_X10Y113_CO5),
.O6(CLBLM_L_X8Y113_SLICE_X10Y113_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0800000088000000)
  ) CLBLM_L_X8Y113_SLICE_X10Y113_BLUT (
.I0(LIOB33_X0Y153_IOB_X0Y153_I),
.I1(RIOB33_X105Y101_IOB_X1Y102_I),
.I2(CLBLM_R_X49Y101_SLICE_X74Y101_AO6),
.I3(LIOB33_X0Y151_IOB_X0Y152_I),
.I4(LIOB33_X0Y161_IOB_X0Y161_I),
.I5(CLBLM_L_X8Y113_SLICE_X10Y113_CO6),
.O5(CLBLM_L_X8Y113_SLICE_X10Y113_BO5),
.O6(CLBLM_L_X8Y113_SLICE_X10Y113_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hccffccfc00ff00f0)
  ) CLBLM_L_X8Y113_SLICE_X10Y113_ALUT (
.I0(1'b1),
.I1(CLBLM_R_X5Y113_SLICE_X6Y113_AO6),
.I2(LIOB33_X0Y87_IOB_X0Y87_I),
.I3(LIOB33_X0Y95_IOB_X0Y95_I),
.I4(LIOB33_X0Y85_IOB_X0Y86_I),
.I5(1'b1),
.O5(CLBLM_L_X8Y113_SLICE_X10Y113_AO5),
.O6(CLBLM_L_X8Y113_SLICE_X10Y113_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffffffffffeff)
  ) CLBLM_L_X8Y113_SLICE_X11Y113_DLUT (
.I0(CLBLM_L_X8Y113_SLICE_X11Y113_AO6),
.I1(LIOB33_X0Y125_IOB_X0Y125_I),
.I2(CLBLM_R_X7Y114_SLICE_X8Y114_BO5),
.I3(CLBLM_L_X8Y113_SLICE_X11Y113_AO5),
.I4(CLBLM_R_X5Y110_SLICE_X6Y110_AO6),
.I5(LIOB33_X0Y131_IOB_X0Y132_I),
.O5(CLBLM_L_X8Y113_SLICE_X11Y113_DO5),
.O6(CLBLM_L_X8Y113_SLICE_X11Y113_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000001)
  ) CLBLM_L_X8Y113_SLICE_X11Y113_CLUT (
.I0(CLBLM_R_X7Y113_SLICE_X8Y113_AO5),
.I1(CLBLM_R_X7Y113_SLICE_X8Y113_DO6),
.I2(CLBLM_R_X7Y113_SLICE_X8Y113_CO6),
.I3(CLBLM_L_X8Y113_SLICE_X10Y113_AO6),
.I4(CLBLM_L_X8Y113_SLICE_X11Y113_DO6),
.I5(CLBLM_R_X5Y113_SLICE_X6Y113_AO5),
.O5(CLBLM_L_X8Y113_SLICE_X11Y113_CO5),
.O6(CLBLM_L_X8Y113_SLICE_X11Y113_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff000010ff0000)
  ) CLBLM_L_X8Y113_SLICE_X11Y113_BLUT (
.I0(LIOB33_SING_X0Y99_IOB_X0Y99_I),
.I1(CLBLM_R_X5Y115_SLICE_X6Y115_AO6),
.I2(LIOB33_X0Y129_IOB_X0Y129_I),
.I3(CLBLM_R_X7Y113_SLICE_X8Y113_AO5),
.I4(CLBLM_L_X10Y123_SLICE_X12Y123_AO6),
.I5(RIOB33_X105Y163_IOB_X1Y163_I),
.O5(CLBLM_L_X8Y113_SLICE_X11Y113_BO5),
.O6(CLBLM_L_X8Y113_SLICE_X11Y113_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h33223322cccccfcf)
  ) CLBLM_L_X8Y113_SLICE_X11Y113_ALUT (
.I0(LIOB33_X0Y103_IOB_X0Y103_I),
.I1(LIOB33_X0Y95_IOB_X0Y95_I),
.I2(LIOB33_X0Y85_IOB_X0Y85_I),
.I3(LIOB33_X0Y103_IOB_X0Y104_I),
.I4(LIOB33_X0Y83_IOB_X0Y84_I),
.I5(1'b1),
.O5(CLBLM_L_X8Y113_SLICE_X11Y113_AO5),
.O6(CLBLM_L_X8Y113_SLICE_X11Y113_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X10Y113_SLICE_X12Y113_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X10Y113_SLICE_X12Y113_DO5),
.O6(CLBLM_L_X10Y113_SLICE_X12Y113_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'haa00aa0aaa22aa2a)
  ) CLBLM_L_X10Y113_SLICE_X12Y113_CLUT (
.I0(CLBLM_L_X10Y123_SLICE_X12Y123_AO6),
.I1(CLBLM_L_X8Y113_SLICE_X10Y113_AO5),
.I2(CLBLM_R_X7Y114_SLICE_X8Y114_AO6),
.I3(RIOB33_X105Y165_IOB_X1Y165_I),
.I4(LIOB33_X0Y85_IOB_X0Y86_I),
.I5(CLBLM_R_X5Y113_SLICE_X6Y113_AO6),
.O5(CLBLM_L_X10Y113_SLICE_X12Y113_CO5),
.O6(CLBLM_L_X10Y113_SLICE_X12Y113_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000033313131)
  ) CLBLM_L_X10Y113_SLICE_X12Y113_BLUT (
.I0(CLBLM_R_X7Y113_SLICE_X8Y113_CO6),
.I1(LIOB33_X0Y159_IOB_X0Y160_I),
.I2(RIOB33_X105Y171_IOB_X1Y172_I),
.I3(LIOB33_X0Y151_IOB_X0Y151_I),
.I4(LIOB33_X0Y127_IOB_X0Y127_I),
.I5(LIOB33_X0Y159_IOB_X0Y159_I),
.O5(CLBLM_L_X10Y113_SLICE_X12Y113_BO5),
.O6(CLBLM_L_X10Y113_SLICE_X12Y113_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f50000f3f70000)
  ) CLBLM_L_X10Y113_SLICE_X12Y113_ALUT (
.I0(CLBLM_R_X7Y114_SLICE_X8Y114_AO6),
.I1(CLBLM_L_X8Y113_SLICE_X11Y113_AO6),
.I2(RIOB33_SING_X105Y100_IOB_X1Y100_I),
.I3(LIOB33_X0Y103_IOB_X0Y103_I),
.I4(CLBLM_L_X10Y123_SLICE_X12Y123_AO6),
.I5(LIOB33_X0Y131_IOB_X0Y132_I),
.O5(CLBLM_L_X10Y113_SLICE_X12Y113_AO5),
.O6(CLBLM_L_X10Y113_SLICE_X12Y113_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X10Y113_SLICE_X13Y113_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X10Y113_SLICE_X13Y113_DO5),
.O6(CLBLM_L_X10Y113_SLICE_X13Y113_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X10Y113_SLICE_X13Y113_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X10Y113_SLICE_X13Y113_CO5),
.O6(CLBLM_L_X10Y113_SLICE_X13Y113_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f0f0f0f000f010)
  ) CLBLM_L_X10Y113_SLICE_X13Y113_BLUT (
.I0(CLBLM_R_X5Y110_SLICE_X6Y110_AO6),
.I1(CLBLM_R_X5Y113_SLICE_X6Y113_AO6),
.I2(CLBLM_L_X10Y123_SLICE_X12Y123_AO6),
.I3(RIOB33_X105Y155_IOB_X1Y156_I),
.I4(LIOB33_X0Y125_IOB_X0Y125_I),
.I5(CLBLM_R_X5Y112_SLICE_X7Y112_AO6),
.O5(CLBLM_L_X10Y113_SLICE_X13Y113_BO5),
.O6(CLBLM_L_X10Y113_SLICE_X13Y113_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hcccccc00cccccc4c)
  ) CLBLM_L_X10Y113_SLICE_X13Y113_ALUT (
.I0(CLBLM_R_X5Y110_SLICE_X6Y110_AO6),
.I1(CLBLM_L_X10Y123_SLICE_X12Y123_AO6),
.I2(LIOB33_X0Y125_IOB_X0Y125_I),
.I3(RIOB33_X105Y159_IOB_X1Y160_I),
.I4(CLBLM_R_X7Y113_SLICE_X8Y113_BO6),
.I5(CLBLM_R_X7Y113_SLICE_X8Y113_DO6),
.O5(CLBLM_L_X10Y113_SLICE_X13Y113_AO5),
.O6(CLBLM_L_X10Y113_SLICE_X13Y113_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X10Y114_SLICE_X12Y114_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X10Y114_SLICE_X12Y114_DO5),
.O6(CLBLM_L_X10Y114_SLICE_X12Y114_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X10Y114_SLICE_X12Y114_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X10Y114_SLICE_X12Y114_CO5),
.O6(CLBLM_L_X10Y114_SLICE_X12Y114_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000fc00fd)
  ) CLBLM_L_X10Y114_SLICE_X12Y114_BLUT (
.I0(CLBLL_L_X4Y111_SLICE_X5Y111_AO5),
.I1(CLBLM_R_X5Y114_SLICE_X7Y114_AO5),
.I2(RIOB33_X105Y159_IOB_X1Y159_I),
.I3(LIOB33_X0Y159_IOB_X0Y160_I),
.I4(CLBLM_R_X5Y111_SLICE_X6Y111_AO6),
.I5(LIOB33_X0Y159_IOB_X0Y159_I),
.O5(CLBLM_L_X10Y114_SLICE_X12Y114_BO5),
.O6(CLBLM_L_X10Y114_SLICE_X12Y114_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0a0f0a0f0e0f0f0)
  ) CLBLM_L_X10Y114_SLICE_X12Y114_ALUT (
.I0(RIOB33_X105Y171_IOB_X1Y171_I),
.I1(LIOB33_X0Y131_IOB_X0Y132_I),
.I2(CLBLM_L_X10Y123_SLICE_X12Y123_AO6),
.I3(CLBLM_R_X7Y114_SLICE_X9Y114_AO6),
.I4(CLBLM_L_X8Y113_SLICE_X11Y113_AO6),
.I5(CLBLM_R_X7Y114_SLICE_X8Y114_BO5),
.O5(CLBLM_L_X10Y114_SLICE_X12Y114_AO5),
.O6(CLBLM_L_X10Y114_SLICE_X12Y114_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X10Y114_SLICE_X13Y114_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X10Y114_SLICE_X13Y114_DO5),
.O6(CLBLM_L_X10Y114_SLICE_X13Y114_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X10Y114_SLICE_X13Y114_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X10Y114_SLICE_X13Y114_CO5),
.O6(CLBLM_L_X10Y114_SLICE_X13Y114_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X10Y114_SLICE_X13Y114_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X10Y114_SLICE_X13Y114_BO5),
.O6(CLBLM_L_X10Y114_SLICE_X13Y114_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X10Y114_SLICE_X13Y114_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X10Y114_SLICE_X13Y114_AO5),
.O6(CLBLM_L_X10Y114_SLICE_X13Y114_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X10Y123_SLICE_X12Y123_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X10Y123_SLICE_X12Y123_DO5),
.O6(CLBLM_L_X10Y123_SLICE_X12Y123_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X10Y123_SLICE_X12Y123_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X10Y123_SLICE_X12Y123_CO5),
.O6(CLBLM_L_X10Y123_SLICE_X12Y123_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X10Y123_SLICE_X12Y123_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X10Y123_SLICE_X12Y123_BO5),
.O6(CLBLM_L_X10Y123_SLICE_X12Y123_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h00000f0f00000f0f)
  ) CLBLM_L_X10Y123_SLICE_X12Y123_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(LIOB33_X0Y159_IOB_X0Y160_I),
.I3(1'b1),
.I4(LIOB33_X0Y159_IOB_X0Y159_I),
.I5(1'b1),
.O5(CLBLM_L_X10Y123_SLICE_X12Y123_AO5),
.O6(CLBLM_L_X10Y123_SLICE_X12Y123_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X10Y123_SLICE_X13Y123_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X10Y123_SLICE_X13Y123_DO5),
.O6(CLBLM_L_X10Y123_SLICE_X13Y123_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X10Y123_SLICE_X13Y123_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X10Y123_SLICE_X13Y123_CO5),
.O6(CLBLM_L_X10Y123_SLICE_X13Y123_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X10Y123_SLICE_X13Y123_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X10Y123_SLICE_X13Y123_BO5),
.O6(CLBLM_L_X10Y123_SLICE_X13Y123_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X10Y123_SLICE_X13Y123_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X10Y123_SLICE_X13Y123_AO5),
.O6(CLBLM_L_X10Y123_SLICE_X13Y123_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X56Y119_SLICE_X84Y119_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X56Y119_SLICE_X84Y119_DO5),
.O6(CLBLM_L_X56Y119_SLICE_X84Y119_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X56Y119_SLICE_X84Y119_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X56Y119_SLICE_X84Y119_CO5),
.O6(CLBLM_L_X56Y119_SLICE_X84Y119_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X56Y119_SLICE_X84Y119_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X56Y119_SLICE_X84Y119_BO5),
.O6(CLBLM_L_X56Y119_SLICE_X84Y119_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffafffaffffffcc)
  ) CLBLM_L_X56Y119_SLICE_X84Y119_ALUT (
.I0(LIOB33_X0Y175_IOB_X0Y175_I),
.I1(RIOB33_X105Y119_IOB_X1Y119_I),
.I2(LIOB33_X0Y113_IOB_X0Y113_I),
.I3(CLBLM_L_X10Y113_SLICE_X13Y113_BO6),
.I4(LIOB33_X0Y53_IOB_X0Y53_I),
.I5(1'b1),
.O5(CLBLM_L_X56Y119_SLICE_X84Y119_AO5),
.O6(CLBLM_L_X56Y119_SLICE_X84Y119_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X56Y119_SLICE_X85Y119_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X56Y119_SLICE_X85Y119_DO5),
.O6(CLBLM_L_X56Y119_SLICE_X85Y119_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X56Y119_SLICE_X85Y119_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X56Y119_SLICE_X85Y119_CO5),
.O6(CLBLM_L_X56Y119_SLICE_X85Y119_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X56Y119_SLICE_X85Y119_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X56Y119_SLICE_X85Y119_BO5),
.O6(CLBLM_L_X56Y119_SLICE_X85Y119_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X56Y119_SLICE_X85Y119_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X56Y119_SLICE_X85Y119_AO5),
.O6(CLBLM_L_X56Y119_SLICE_X85Y119_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y110_SLICE_X2Y110_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y110_SLICE_X2Y110_DO5),
.O6(CLBLM_R_X3Y110_SLICE_X2Y110_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y110_SLICE_X2Y110_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y110_SLICE_X2Y110_CO5),
.O6(CLBLM_R_X3Y110_SLICE_X2Y110_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y110_SLICE_X2Y110_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y110_SLICE_X2Y110_BO5),
.O6(CLBLM_R_X3Y110_SLICE_X2Y110_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y110_SLICE_X2Y110_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y110_SLICE_X2Y110_AO5),
.O6(CLBLM_R_X3Y110_SLICE_X2Y110_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y110_SLICE_X3Y110_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y110_SLICE_X3Y110_DO5),
.O6(CLBLM_R_X3Y110_SLICE_X3Y110_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y110_SLICE_X3Y110_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y110_SLICE_X3Y110_CO5),
.O6(CLBLM_R_X3Y110_SLICE_X3Y110_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y110_SLICE_X3Y110_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y110_SLICE_X3Y110_BO5),
.O6(CLBLM_R_X3Y110_SLICE_X3Y110_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h5555444455505550)
  ) CLBLM_R_X3Y110_SLICE_X3Y110_ALUT (
.I0(LIOB33_X0Y95_IOB_X0Y96_I),
.I1(LIOB33_X0Y61_IOB_X0Y62_I),
.I2(LIOB33_X0Y59_IOB_X0Y59_I),
.I3(LIOB33_X0Y57_IOB_X0Y58_I),
.I4(LIOB33_X0Y59_IOB_X0Y60_I),
.I5(1'b1),
.O5(CLBLM_R_X3Y110_SLICE_X3Y110_AO5),
.O6(CLBLM_R_X3Y110_SLICE_X3Y110_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y111_SLICE_X2Y111_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y111_SLICE_X2Y111_DO5),
.O6(CLBLM_R_X3Y111_SLICE_X2Y111_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y111_SLICE_X2Y111_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y111_SLICE_X2Y111_CO5),
.O6(CLBLM_R_X3Y111_SLICE_X2Y111_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y111_SLICE_X2Y111_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y111_SLICE_X2Y111_BO5),
.O6(CLBLM_R_X3Y111_SLICE_X2Y111_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h00fa00fa33013301)
  ) CLBLM_R_X3Y111_SLICE_X2Y111_ALUT (
.I0(LIOB33_X0Y55_IOB_X0Y56_I),
.I1(LIOB33_X0Y119_IOB_X0Y120_I),
.I2(LIOB33_X0Y57_IOB_X0Y57_I),
.I3(LIOB33_X0Y95_IOB_X0Y96_I),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y111_SLICE_X2Y111_AO5),
.O6(CLBLM_R_X3Y111_SLICE_X2Y111_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hc3c3c0c0c0c0c2c0)
  ) CLBLM_R_X3Y111_SLICE_X3Y111_DLUT (
.I0(CLBLM_R_X3Y110_SLICE_X3Y110_AO6),
.I1(CLBLM_R_X3Y111_SLICE_X2Y111_AO6),
.I2(LIOB33_X0Y119_IOB_X0Y120_I),
.I3(LIOB33_X0Y115_IOB_X0Y116_I),
.I4(LIOB33_X0Y121_IOB_X0Y122_I),
.I5(CLBLM_R_X3Y110_SLICE_X3Y110_AO5),
.O5(CLBLM_R_X3Y111_SLICE_X3Y111_DO5),
.O6(CLBLM_R_X3Y111_SLICE_X3Y111_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h4444445540404050)
  ) CLBLM_R_X3Y111_SLICE_X3Y111_CLUT (
.I0(LIOB33_X0Y117_IOB_X0Y118_I),
.I1(LIOB33_X0Y95_IOB_X0Y96_I),
.I2(CLBLL_L_X4Y111_SLICE_X4Y111_BO6),
.I3(LIOB33_X0Y65_IOB_X0Y65_I),
.I4(LIOB33_X0Y63_IOB_X0Y63_I),
.I5(1'b1),
.O5(CLBLM_R_X3Y111_SLICE_X3Y111_CO5),
.O6(CLBLM_R_X3Y111_SLICE_X3Y111_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h33333300cfcfcfff)
  ) CLBLM_R_X3Y111_SLICE_X3Y111_BLUT (
.I0(1'b1),
.I1(LIOB33_X0Y95_IOB_X0Y96_I),
.I2(LIOB33_X0Y117_IOB_X0Y118_I),
.I3(LIOB33_X0Y63_IOB_X0Y63_I),
.I4(LIOB33_X0Y65_IOB_X0Y65_I),
.I5(1'b1),
.O5(CLBLM_R_X3Y111_SLICE_X3Y111_BO5),
.O6(CLBLM_R_X3Y111_SLICE_X3Y111_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000cdcd32320000)
  ) CLBLM_R_X3Y111_SLICE_X3Y111_ALUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(LIOB33_X0Y95_IOB_X0Y96_I),
.I2(LIOB33_X0Y75_IOB_X0Y75_I),
.I3(1'b1),
.I4(LIOB33_X0Y113_IOB_X0Y114_I),
.I5(1'b1),
.O5(CLBLM_R_X3Y111_SLICE_X3Y111_AO5),
.O6(CLBLM_R_X3Y111_SLICE_X3Y111_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y112_SLICE_X2Y112_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y112_SLICE_X2Y112_DO5),
.O6(CLBLM_R_X3Y112_SLICE_X2Y112_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y112_SLICE_X2Y112_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y112_SLICE_X2Y112_CO5),
.O6(CLBLM_R_X3Y112_SLICE_X2Y112_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y112_SLICE_X2Y112_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y112_SLICE_X2Y112_BO5),
.O6(CLBLM_R_X3Y112_SLICE_X2Y112_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y112_SLICE_X2Y112_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y112_SLICE_X2Y112_AO5),
.O6(CLBLM_R_X3Y112_SLICE_X2Y112_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y112_SLICE_X3Y112_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y112_SLICE_X3Y112_DO5),
.O6(CLBLM_R_X3Y112_SLICE_X3Y112_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y112_SLICE_X3Y112_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y112_SLICE_X3Y112_CO5),
.O6(CLBLM_R_X3Y112_SLICE_X3Y112_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h1100000011010000)
  ) CLBLM_R_X3Y112_SLICE_X3Y112_BLUT (
.I0(LIOB33_X0Y111_IOB_X0Y111_I),
.I1(CLBLL_L_X4Y112_SLICE_X5Y112_BO6),
.I2(LIOB33_X0Y73_IOB_X0Y74_I),
.I3(LIOB33_X0Y95_IOB_X0Y96_I),
.I4(CLBLM_R_X3Y111_SLICE_X3Y111_CO5),
.I5(LIOB33_X0Y71_IOB_X0Y72_I),
.O5(CLBLM_R_X3Y112_SLICE_X3Y112_BO5),
.O6(CLBLM_R_X3Y112_SLICE_X3Y112_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hff0fff3f0f000f03)
  ) CLBLM_R_X3Y112_SLICE_X3Y112_ALUT (
.I0(1'b1),
.I1(LIOB33_X0Y79_IOB_X0Y79_I),
.I2(LIOB33_X0Y115_IOB_X0Y115_I),
.I3(LIOB33_X0Y95_IOB_X0Y96_I),
.I4(LIOB33_X0Y77_IOB_X0Y78_I),
.I5(1'b1),
.O5(CLBLM_R_X3Y112_SLICE_X3Y112_AO5),
.O6(CLBLM_R_X3Y112_SLICE_X3Y112_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X5Y109_SLICE_X6Y109_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y109_SLICE_X6Y109_DO5),
.O6(CLBLM_R_X5Y109_SLICE_X6Y109_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X5Y109_SLICE_X6Y109_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y109_SLICE_X6Y109_CO5),
.O6(CLBLM_R_X5Y109_SLICE_X6Y109_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffff33333332)
  ) CLBLM_R_X5Y109_SLICE_X6Y109_BLUT (
.I0(LIOB33_X0Y87_IOB_X0Y88_I),
.I1(LIOB33_X0Y95_IOB_X0Y95_I),
.I2(LIOB33_X0Y85_IOB_X0Y86_I),
.I3(LIOB33_X0Y87_IOB_X0Y87_I),
.I4(LIOB33_X0Y89_IOB_X0Y90_I),
.I5(CLBLM_R_X5Y110_SLICE_X6Y110_AO6),
.O5(CLBLM_R_X5Y109_SLICE_X6Y109_BO5),
.O6(CLBLM_R_X5Y109_SLICE_X6Y109_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffeeffffffeefffe)
  ) CLBLM_R_X5Y109_SLICE_X6Y109_ALUT (
.I0(CLBLM_R_X7Y113_SLICE_X8Y113_AO6),
.I1(CLBLL_L_X4Y107_SLICE_X4Y107_AO6),
.I2(LIOB33_X0Y101_IOB_X0Y102_I),
.I3(CLBLM_R_X5Y109_SLICE_X6Y109_BO6),
.I4(LIOB33_X0Y95_IOB_X0Y95_I),
.I5(LIOB33_X0Y101_IOB_X0Y101_I),
.O5(CLBLM_R_X5Y109_SLICE_X6Y109_AO5),
.O6(CLBLM_R_X5Y109_SLICE_X6Y109_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X5Y109_SLICE_X7Y109_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y109_SLICE_X7Y109_DO5),
.O6(CLBLM_R_X5Y109_SLICE_X7Y109_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X5Y109_SLICE_X7Y109_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y109_SLICE_X7Y109_CO5),
.O6(CLBLM_R_X5Y109_SLICE_X7Y109_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X5Y109_SLICE_X7Y109_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y109_SLICE_X7Y109_BO5),
.O6(CLBLM_R_X5Y109_SLICE_X7Y109_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X5Y109_SLICE_X7Y109_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y109_SLICE_X7Y109_AO5),
.O6(CLBLM_R_X5Y109_SLICE_X7Y109_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X5Y110_SLICE_X6Y110_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y110_SLICE_X6Y110_DO5),
.O6(CLBLM_R_X5Y110_SLICE_X6Y110_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X5Y110_SLICE_X6Y110_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y110_SLICE_X6Y110_CO5),
.O6(CLBLM_R_X5Y110_SLICE_X6Y110_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X5Y110_SLICE_X6Y110_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y110_SLICE_X6Y110_BO5),
.O6(CLBLM_R_X5Y110_SLICE_X6Y110_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000fff00000aaa0)
  ) CLBLM_R_X5Y110_SLICE_X6Y110_ALUT (
.I0(LIOB33_X0Y125_IOB_X0Y125_I),
.I1(1'b1),
.I2(LIOB33_X0Y91_IOB_X0Y92_I),
.I3(LIOB33_X0Y91_IOB_X0Y91_I),
.I4(LIOB33_X0Y95_IOB_X0Y95_I),
.I5(1'b1),
.O5(CLBLM_R_X5Y110_SLICE_X6Y110_AO5),
.O6(CLBLM_R_X5Y110_SLICE_X6Y110_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X5Y110_SLICE_X7Y110_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y110_SLICE_X7Y110_DO5),
.O6(CLBLM_R_X5Y110_SLICE_X7Y110_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X5Y110_SLICE_X7Y110_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y110_SLICE_X7Y110_CO5),
.O6(CLBLM_R_X5Y110_SLICE_X7Y110_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X5Y110_SLICE_X7Y110_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y110_SLICE_X7Y110_BO5),
.O6(CLBLM_R_X5Y110_SLICE_X7Y110_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X5Y110_SLICE_X7Y110_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y110_SLICE_X7Y110_AO5),
.O6(CLBLM_R_X5Y110_SLICE_X7Y110_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffffffffffffe)
  ) CLBLM_R_X5Y111_SLICE_X6Y111_DLUT (
.I0(CLBLL_L_X4Y110_SLICE_X4Y110_BO5),
.I1(CLBLM_R_X5Y111_SLICE_X7Y111_AO5),
.I2(CLBLM_R_X5Y112_SLICE_X6Y112_BO6),
.I3(CLBLL_L_X4Y112_SLICE_X4Y112_CO6),
.I4(CLBLL_L_X4Y111_SLICE_X4Y111_AO5),
.I5(CLBLL_L_X4Y111_SLICE_X4Y111_CO6),
.O5(CLBLM_R_X5Y111_SLICE_X6Y111_DO5),
.O6(CLBLM_R_X5Y111_SLICE_X6Y111_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000001000000000)
  ) CLBLM_R_X5Y111_SLICE_X6Y111_CLUT (
.I0(CLBLL_L_X4Y111_SLICE_X5Y111_AO5),
.I1(CLBLM_R_X3Y111_SLICE_X2Y111_AO5),
.I2(LIOB33_X0Y117_IOB_X0Y118_I),
.I3(CLBLM_R_X5Y111_SLICE_X6Y111_AO5),
.I4(CLBLM_R_X5Y111_SLICE_X6Y111_DO6),
.I5(CLBLM_R_X3Y111_SLICE_X3Y111_BO6),
.O5(CLBLM_R_X5Y111_SLICE_X6Y111_CO5),
.O6(CLBLM_R_X5Y111_SLICE_X6Y111_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'ha0a0a0a0b0b0f0b0)
  ) CLBLM_R_X5Y111_SLICE_X6Y111_BLUT (
.I0(CLBLM_R_X5Y115_SLICE_X6Y115_AO5),
.I1(CLBLL_L_X4Y112_SLICE_X4Y112_BO6),
.I2(CLBLM_L_X10Y123_SLICE_X12Y123_AO6),
.I3(LIOB33_X0Y111_IOB_X0Y112_I),
.I4(CLBLL_L_X4Y111_SLICE_X5Y111_BO6),
.I5(CLBLM_R_X3Y111_SLICE_X3Y111_CO6),
.O5(CLBLM_R_X5Y111_SLICE_X6Y111_BO5),
.O6(CLBLM_R_X5Y111_SLICE_X6Y111_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h55ea55eec0c0cccc)
  ) CLBLM_R_X5Y111_SLICE_X6Y111_ALUT (
.I0(LIOB33_X0Y117_IOB_X0Y118_I),
.I1(CLBLL_L_X4Y112_SLICE_X4Y112_BO6),
.I2(CLBLL_L_X4Y111_SLICE_X5Y111_BO6),
.I3(CLBLM_R_X3Y111_SLICE_X3Y111_BO6),
.I4(LIOB33_X0Y111_IOB_X0Y112_I),
.I5(1'b1),
.O5(CLBLM_R_X5Y111_SLICE_X6Y111_AO5),
.O6(CLBLM_R_X5Y111_SLICE_X6Y111_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffffff5f5ffff)
  ) CLBLM_R_X5Y111_SLICE_X7Y111_DLUT (
.I0(LIOB33_X0Y113_IOB_X0Y114_I),
.I1(1'b1),
.I2(LIOB33_X0Y75_IOB_X0Y75_I),
.I3(1'b1),
.I4(LIOB33_X0Y109_IOB_X0Y109_I),
.I5(LIOB33_X0Y79_IOB_X0Y80_I),
.O5(CLBLM_R_X5Y111_SLICE_X7Y111_DO5),
.O6(CLBLM_R_X5Y111_SLICE_X7Y111_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h33333333ff33f733)
  ) CLBLM_R_X5Y111_SLICE_X7Y111_CLUT (
.I0(LIOB33_X0Y113_IOB_X0Y114_I),
.I1(CLBLM_L_X10Y123_SLICE_X12Y123_AO6),
.I2(LIOB33_X0Y75_IOB_X0Y75_I),
.I3(CLBLL_L_X4Y111_SLICE_X4Y111_CO6),
.I4(CLBLM_R_X5Y115_SLICE_X6Y115_AO6),
.I5(RIOB33_X105Y169_IOB_X1Y169_I),
.O5(CLBLM_R_X5Y111_SLICE_X7Y111_CO5),
.O6(CLBLM_R_X5Y111_SLICE_X7Y111_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'haabaffff00000000)
  ) CLBLM_R_X5Y111_SLICE_X7Y111_BLUT (
.I0(RIOB33_X105Y161_IOB_X1Y161_I),
.I1(LIOB33_X0Y79_IOB_X0Y80_I),
.I2(LIOB33_X0Y109_IOB_X0Y109_I),
.I3(CLBLM_R_X5Y115_SLICE_X6Y115_AO6),
.I4(CLBLL_L_X4Y110_SLICE_X4Y110_BO5),
.I5(CLBLM_L_X10Y123_SLICE_X12Y123_AO6),
.O5(CLBLM_R_X5Y111_SLICE_X7Y111_BO5),
.O6(CLBLM_R_X5Y111_SLICE_X7Y111_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0faf0f8aaffaaee)
  ) CLBLM_R_X5Y111_SLICE_X7Y111_ALUT (
.I0(LIOB33_X0Y115_IOB_X0Y116_I),
.I1(LIOB33_X0Y61_IOB_X0Y62_I),
.I2(CLBLL_L_X4Y111_SLICE_X4Y111_AO5),
.I3(LIOB33_X0Y95_IOB_X0Y96_I),
.I4(LIOB33_X0Y59_IOB_X0Y60_I),
.I5(1'b1),
.O5(CLBLM_R_X5Y111_SLICE_X7Y111_AO5),
.O6(CLBLM_R_X5Y111_SLICE_X7Y111_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X5Y112_SLICE_X6Y112_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y112_SLICE_X6Y112_DO5),
.O6(CLBLM_R_X5Y112_SLICE_X6Y112_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffdfdfffffdfdf)
  ) CLBLM_R_X5Y112_SLICE_X6Y112_CLUT (
.I0(LIOB33_X0Y139_IOB_X0Y139_I),
.I1(CLBLM_R_X3Y112_SLICE_X3Y112_AO5),
.I2(CLBLM_R_X5Y111_SLICE_X7Y111_AO5),
.I3(1'b1),
.I4(CLBLL_L_X4Y111_SLICE_X5Y111_AO5),
.I5(1'b1),
.O5(CLBLM_R_X5Y112_SLICE_X6Y112_CO5),
.O6(CLBLM_R_X5Y112_SLICE_X6Y112_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffffff30ff35b)
  ) CLBLM_R_X5Y112_SLICE_X6Y112_BLUT (
.I0(LIOB33_X0Y81_IOB_X0Y81_I),
.I1(LIOB33_X0Y111_IOB_X0Y112_I),
.I2(LIOB33_X0Y109_IOB_X0Y109_I),
.I3(LIOB33_X0Y95_IOB_X0Y96_I),
.I4(LIOB33_X0Y79_IOB_X0Y80_I),
.I5(CLBLM_R_X3Y112_SLICE_X3Y112_AO5),
.O5(CLBLM_R_X5Y112_SLICE_X6Y112_BO5),
.O6(CLBLM_R_X5Y112_SLICE_X6Y112_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaaaaaa00aa20aa)
  ) CLBLM_R_X5Y112_SLICE_X6Y112_ALUT (
.I0(CLBLM_L_X10Y123_SLICE_X12Y123_AO6),
.I1(LIOB33_X0Y77_IOB_X0Y78_I),
.I2(LIOB33_X0Y115_IOB_X0Y115_I),
.I3(CLBLM_R_X5Y112_SLICE_X6Y112_BO6),
.I4(CLBLM_R_X5Y115_SLICE_X6Y115_AO6),
.I5(RIOB33_X105Y167_IOB_X1Y168_I),
.O5(CLBLM_R_X5Y112_SLICE_X6Y112_AO5),
.O6(CLBLM_R_X5Y112_SLICE_X6Y112_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X5Y112_SLICE_X7Y112_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y112_SLICE_X7Y112_DO5),
.O6(CLBLM_R_X5Y112_SLICE_X7Y112_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X5Y112_SLICE_X7Y112_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y112_SLICE_X7Y112_CO5),
.O6(CLBLM_R_X5Y112_SLICE_X7Y112_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X5Y112_SLICE_X7Y112_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y112_SLICE_X7Y112_BO5),
.O6(CLBLM_R_X5Y112_SLICE_X7Y112_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h003000f011115555)
  ) CLBLM_R_X5Y112_SLICE_X7Y112_ALUT (
.I0(LIOB33_X0Y103_IOB_X0Y103_I),
.I1(LIOB33_X0Y67_IOB_X0Y68_I),
.I2(LIOB33_X0Y125_IOB_X0Y125_I),
.I3(LIOB33_X0Y91_IOB_X0Y91_I),
.I4(LIOB33_X0Y69_IOB_X0Y70_I),
.I5(1'b1),
.O5(CLBLM_R_X5Y112_SLICE_X7Y112_AO5),
.O6(CLBLM_R_X5Y112_SLICE_X7Y112_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaaaaaafdfdfdfd)
  ) CLBLM_R_X5Y113_SLICE_X6Y113_DLUT (
.I0(LIOB33_X0Y95_IOB_X0Y95_I),
.I1(LIOB33_X0Y129_IOB_X0Y129_I),
.I2(LIOB33_X0Y131_IOB_X0Y131_I),
.I3(1'b1),
.I4(1'b1),
.I5(LIOB33_X0Y127_IOB_X0Y127_I),
.O5(CLBLM_R_X5Y113_SLICE_X6Y113_DO5),
.O6(CLBLM_R_X5Y113_SLICE_X6Y113_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hcd00cc00ff00ff00)
  ) CLBLM_R_X5Y113_SLICE_X6Y113_CLUT (
.I0(CLBLM_R_X5Y115_SLICE_X6Y115_AO6),
.I1(RIOB33_X105Y169_IOB_X1Y170_I),
.I2(LIOB33_X0Y71_IOB_X0Y72_I),
.I3(CLBLM_L_X10Y123_SLICE_X12Y123_AO6),
.I4(LIOB33_X0Y111_IOB_X0Y111_I),
.I5(CLBLL_L_X4Y112_SLICE_X4Y112_CO6),
.O5(CLBLM_R_X5Y113_SLICE_X6Y113_CO5),
.O6(CLBLM_R_X5Y113_SLICE_X6Y113_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'haa00ba00ff00ff00)
  ) CLBLM_R_X5Y113_SLICE_X6Y113_BLUT (
.I0(LIOB33_X0Y127_IOB_X0Y128_I),
.I1(LIOB33_X0Y93_IOB_X0Y93_I),
.I2(LIOB33_X0Y125_IOB_X0Y126_I),
.I3(CLBLM_L_X10Y123_SLICE_X12Y123_AO6),
.I4(CLBLM_R_X5Y115_SLICE_X6Y115_AO6),
.I5(CLBLM_R_X5Y113_SLICE_X6Y113_AO5),
.O5(CLBLM_R_X5Y113_SLICE_X6Y113_BO5),
.O6(CLBLM_R_X5Y113_SLICE_X6Y113_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfafa0f3eafafaaab)
  ) CLBLM_R_X5Y113_SLICE_X6Y113_ALUT (
.I0(CLBLM_R_X5Y113_SLICE_X6Y113_DO6),
.I1(LIOB33_X0Y93_IOB_X0Y93_I),
.I2(LIOB33_X0Y125_IOB_X0Y126_I),
.I3(LIOB33_X0Y93_IOB_X0Y94_I),
.I4(LIOB33_X0Y95_IOB_X0Y95_I),
.I5(1'b1),
.O5(CLBLM_R_X5Y113_SLICE_X6Y113_AO5),
.O6(CLBLM_R_X5Y113_SLICE_X6Y113_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffce02ffffcc00)
  ) CLBLM_R_X5Y113_SLICE_X7Y113_DLUT (
.I0(LIOB33_X0Y125_IOB_X0Y126_I),
.I1(LIOB33_X0Y67_IOB_X0Y68_I),
.I2(LIOB33_X0Y93_IOB_X0Y93_I),
.I3(LIOB33_X0Y69_IOB_X0Y70_I),
.I4(LIOB33_X0Y103_IOB_X0Y103_I),
.I5(LIOB33_X0Y127_IOB_X0Y127_I),
.O5(CLBLM_R_X5Y113_SLICE_X7Y113_DO5),
.O6(CLBLM_R_X5Y113_SLICE_X7Y113_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffffff7ffffff)
  ) CLBLM_R_X5Y113_SLICE_X7Y113_CLUT (
.I0(LIOB33_X0Y125_IOB_X0Y126_I),
.I1(LIOB33_X0Y127_IOB_X0Y127_I),
.I2(LIOB33_SING_X0Y99_IOB_X0Y99_I),
.I3(LIOB33_X0Y129_IOB_X0Y129_I),
.I4(LIOB33_X0Y151_IOB_X0Y151_I),
.I5(LIOB33_X0Y93_IOB_X0Y93_I),
.O5(CLBLM_R_X5Y113_SLICE_X7Y113_CO5),
.O6(CLBLM_R_X5Y113_SLICE_X7Y113_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000800000808)
  ) CLBLM_R_X5Y113_SLICE_X7Y113_BLUT (
.I0(CLBLM_R_X5Y112_SLICE_X7Y112_AO6),
.I1(CLBLM_R_X7Y113_SLICE_X8Y113_BO6),
.I2(LIOB33_X0Y83_IOB_X0Y84_I),
.I3(LIOB33_X0Y65_IOB_X0Y66_I),
.I4(LIOB33_X0Y85_IOB_X0Y86_I),
.I5(LIOB33_X0Y71_IOB_X0Y71_I),
.O5(CLBLM_R_X5Y113_SLICE_X7Y113_BO5),
.O6(CLBLM_R_X5Y113_SLICE_X7Y113_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000800)
  ) CLBLM_R_X5Y113_SLICE_X7Y113_ALUT (
.I0(CLBLM_R_X5Y112_SLICE_X7Y112_AO5),
.I1(LIOB33_X0Y131_IOB_X0Y131_I),
.I2(LIOB33_X0Y101_IOB_X0Y101_I),
.I3(CLBLM_R_X5Y113_SLICE_X7Y113_BO6),
.I4(CLBLM_R_X5Y115_SLICE_X6Y115_AO6),
.I5(CLBLM_R_X5Y113_SLICE_X7Y113_CO6),
.O5(CLBLM_R_X5Y113_SLICE_X7Y113_AO5),
.O6(CLBLM_R_X5Y113_SLICE_X7Y113_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hccccccfccccccccc)
  ) CLBLM_R_X5Y114_SLICE_X6Y114_DLUT (
.I0(1'b1),
.I1(CLBLM_R_X5Y114_SLICE_X7Y114_AO5),
.I2(LIOB33_X0Y111_IOB_X0Y111_I),
.I3(LIOB33_X0Y63_IOB_X0Y63_I),
.I4(LIOB33_X0Y71_IOB_X0Y72_I),
.I5(LIOB33_X0Y117_IOB_X0Y118_I),
.O5(CLBLM_R_X5Y114_SLICE_X6Y114_DO5),
.O6(CLBLM_R_X5Y114_SLICE_X6Y114_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffffffffffffd)
  ) CLBLM_R_X5Y114_SLICE_X6Y114_CLUT (
.I0(LIOB33_X0Y121_IOB_X0Y122_I),
.I1(CLBLL_L_X4Y113_SLICE_X5Y113_AO6),
.I2(LIOB33_X0Y57_IOB_X0Y58_I),
.I3(CLBLM_R_X7Y114_SLICE_X8Y114_AO6),
.I4(CLBLM_R_X5Y114_SLICE_X6Y114_DO6),
.I5(CLBLM_R_X5Y111_SLICE_X7Y111_DO6),
.O5(CLBLM_R_X5Y114_SLICE_X6Y114_CO5),
.O6(CLBLM_R_X5Y114_SLICE_X6Y114_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffffbbbfffff)
  ) CLBLM_R_X5Y114_SLICE_X6Y114_BLUT (
.I0(LIOB33_X0Y71_IOB_X0Y72_I),
.I1(LIOB33_X0Y117_IOB_X0Y118_I),
.I2(LIOB33_SING_X0Y150_IOB_X0Y150_I),
.I3(LIOB33_X0Y151_IOB_X0Y151_I),
.I4(LIOB33_X0Y111_IOB_X0Y111_I),
.I5(LIOB33_X0Y63_IOB_X0Y63_I),
.O5(CLBLM_R_X5Y114_SLICE_X6Y114_BO5),
.O6(CLBLM_R_X5Y114_SLICE_X6Y114_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000020000)
  ) CLBLM_R_X5Y114_SLICE_X6Y114_ALUT (
.I0(CLBLM_R_X5Y114_SLICE_X7Y114_AO5),
.I1(LIOB33_X0Y57_IOB_X0Y58_I),
.I2(CLBLL_L_X4Y113_SLICE_X5Y113_AO6),
.I3(CLBLM_R_X5Y114_SLICE_X6Y114_BO6),
.I4(LIOB33_X0Y121_IOB_X0Y122_I),
.I5(CLBLM_R_X5Y111_SLICE_X7Y111_DO6),
.O5(CLBLM_R_X5Y114_SLICE_X6Y114_AO5),
.O6(CLBLM_R_X5Y114_SLICE_X6Y114_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X5Y114_SLICE_X7Y114_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y114_SLICE_X7Y114_DO5),
.O6(CLBLM_R_X5Y114_SLICE_X7Y114_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X5Y114_SLICE_X7Y114_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y114_SLICE_X7Y114_CO5),
.O6(CLBLM_R_X5Y114_SLICE_X7Y114_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X5Y114_SLICE_X7Y114_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y114_SLICE_X7Y114_BO5),
.O6(CLBLM_R_X5Y114_SLICE_X7Y114_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0d0f050f2200aa00)
  ) CLBLM_R_X5Y114_SLICE_X7Y114_ALUT (
.I0(LIOB33_X0Y119_IOB_X0Y119_I),
.I1(LIOB33_X0Y69_IOB_X0Y70_I),
.I2(RIOB33_X105Y159_IOB_X1Y159_I),
.I3(LIOB33_X0Y53_IOB_X0Y54_I),
.I4(LIOB33_X0Y67_IOB_X0Y68_I),
.I5(1'b1),
.O5(CLBLM_R_X5Y114_SLICE_X7Y114_AO5),
.O6(CLBLM_R_X5Y114_SLICE_X7Y114_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X5Y115_SLICE_X6Y115_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y115_SLICE_X6Y115_DO5),
.O6(CLBLM_R_X5Y115_SLICE_X6Y115_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X5Y115_SLICE_X6Y115_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y115_SLICE_X6Y115_CO5),
.O6(CLBLM_R_X5Y115_SLICE_X6Y115_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hccccffffbbbaaaaa)
  ) CLBLM_R_X5Y115_SLICE_X6Y115_BLUT (
.I0(LIOB33_X0Y129_IOB_X0Y130_I),
.I1(LIOB33_X0Y57_IOB_X0Y58_I),
.I2(LIOB33_SING_X0Y150_IOB_X0Y150_I),
.I3(LIOB33_X0Y151_IOB_X0Y151_I),
.I4(LIOB33_X0Y121_IOB_X0Y122_I),
.I5(1'b1),
.O5(CLBLM_R_X5Y115_SLICE_X6Y115_BO5),
.O6(CLBLM_R_X5Y115_SLICE_X6Y115_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h000f000fbbbaaaaa)
  ) CLBLM_R_X5Y115_SLICE_X6Y115_ALUT (
.I0(RIOB33_X105Y165_IOB_X1Y166_I),
.I1(LIOB33_X0Y63_IOB_X0Y63_I),
.I2(LIOB33_SING_X0Y150_IOB_X0Y150_I),
.I3(LIOB33_X0Y151_IOB_X0Y151_I),
.I4(LIOB33_X0Y117_IOB_X0Y118_I),
.I5(1'b1),
.O5(CLBLM_R_X5Y115_SLICE_X6Y115_AO5),
.O6(CLBLM_R_X5Y115_SLICE_X6Y115_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X5Y115_SLICE_X7Y115_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y115_SLICE_X7Y115_DO5),
.O6(CLBLM_R_X5Y115_SLICE_X7Y115_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X5Y115_SLICE_X7Y115_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y115_SLICE_X7Y115_CO5),
.O6(CLBLM_R_X5Y115_SLICE_X7Y115_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X5Y115_SLICE_X7Y115_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y115_SLICE_X7Y115_BO5),
.O6(CLBLM_R_X5Y115_SLICE_X7Y115_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'ha0b0a0b0a0b0f0f0)
  ) CLBLM_R_X5Y115_SLICE_X7Y115_ALUT (
.I0(LIOB33_X0Y129_IOB_X0Y130_I),
.I1(CLBLM_R_X5Y115_SLICE_X6Y115_BO6),
.I2(CLBLM_L_X10Y123_SLICE_X12Y123_AO6),
.I3(CLBLM_R_X5Y115_SLICE_X6Y115_AO6),
.I4(CLBLM_R_X5Y111_SLICE_X6Y111_AO6),
.I5(CLBLM_R_X5Y111_SLICE_X7Y111_AO6),
.O5(CLBLM_R_X5Y115_SLICE_X7Y115_AO5),
.O6(CLBLM_R_X5Y115_SLICE_X7Y115_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hff00ff00ffffff11)
  ) CLBLM_R_X7Y113_SLICE_X8Y113_DLUT (
.I0(LIOB33_X0Y87_IOB_X0Y88_I),
.I1(LIOB33_X0Y89_IOB_X0Y90_I),
.I2(1'b1),
.I3(CLBLM_R_X5Y113_SLICE_X6Y113_AO6),
.I4(LIOB33_X0Y95_IOB_X0Y95_I),
.I5(LIOB33_X0Y123_IOB_X0Y123_I),
.O5(CLBLM_R_X7Y113_SLICE_X8Y113_DO5),
.O6(CLBLM_R_X7Y113_SLICE_X8Y113_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hf1f1f1f1ff0efffe)
  ) CLBLM_R_X7Y113_SLICE_X8Y113_CLUT (
.I0(LIOB33_SING_X0Y100_IOB_X0Y100_I),
.I1(LIOB33_SING_X0Y99_IOB_X0Y99_I),
.I2(LIOB33_X0Y95_IOB_X0Y95_I),
.I3(CLBLM_R_X7Y114_SLICE_X8Y114_CO6),
.I4(LIOB33_X0Y127_IOB_X0Y127_I),
.I5(LIOB33_X0Y129_IOB_X0Y129_I),
.O5(CLBLM_R_X7Y113_SLICE_X8Y113_CO5),
.O6(CLBLM_R_X7Y113_SLICE_X8Y113_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h000050f000001030)
  ) CLBLM_R_X7Y113_SLICE_X8Y113_BLUT (
.I0(LIOB33_X0Y69_IOB_X0Y70_I),
.I1(LIOB33_X0Y85_IOB_X0Y86_I),
.I2(LIOB33_X0Y123_IOB_X0Y123_I),
.I3(LIOB33_X0Y67_IOB_X0Y68_I),
.I4(LIOB33_X0Y87_IOB_X0Y88_I),
.I5(1'b1),
.O5(CLBLM_R_X7Y113_SLICE_X8Y113_BO5),
.O6(CLBLM_R_X7Y113_SLICE_X8Y113_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0f0f0c0caafaaafb)
  ) CLBLM_R_X7Y113_SLICE_X8Y113_ALUT (
.I0(CLBLM_R_X7Y114_SLICE_X8Y114_CO6),
.I1(LIOB33_SING_X0Y99_IOB_X0Y99_I),
.I2(LIOB33_X0Y95_IOB_X0Y95_I),
.I3(LIOB33_X0Y129_IOB_X0Y129_I),
.I4(LIOB33_SING_X0Y100_IOB_X0Y100_I),
.I5(1'b1),
.O5(CLBLM_R_X7Y113_SLICE_X8Y113_AO5),
.O6(CLBLM_R_X7Y113_SLICE_X8Y113_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X7Y113_SLICE_X9Y113_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y113_SLICE_X9Y113_DO5),
.O6(CLBLM_R_X7Y113_SLICE_X9Y113_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'heaeaeaeaeaeaeaea)
  ) CLBLM_R_X7Y113_SLICE_X9Y113_CLUT (
.I0(LIOB33_X0Y83_IOB_X0Y84_I),
.I1(LIOB33_X0Y71_IOB_X0Y71_I),
.I2(LIOB33_X0Y65_IOB_X0Y66_I),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y113_SLICE_X9Y113_CO5),
.O6(CLBLM_R_X7Y113_SLICE_X9Y113_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffeffffffffff)
  ) CLBLM_R_X7Y113_SLICE_X9Y113_BLUT (
.I0(LIOB33_X0Y101_IOB_X0Y101_I),
.I1(LIOB33_X0Y159_IOB_X0Y159_I),
.I2(LIOB33_SING_X0Y99_IOB_X0Y99_I),
.I3(LIOB33_X0Y131_IOB_X0Y131_I),
.I4(LIOB33_X0Y159_IOB_X0Y160_I),
.I5(LIOB33_X0Y129_IOB_X0Y129_I),
.O5(CLBLM_R_X7Y113_SLICE_X9Y113_BO5),
.O6(CLBLM_R_X7Y113_SLICE_X9Y113_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f0f0f0f0f4f0f0)
  ) CLBLM_R_X7Y113_SLICE_X9Y113_ALUT (
.I0(CLBLM_R_X5Y113_SLICE_X7Y113_DO6),
.I1(CLBLM_R_X5Y112_SLICE_X7Y112_AO6),
.I2(CLBLL_L_X4Y141_SLICE_X4Y141_AO6),
.I3(CLBLM_R_X7Y113_SLICE_X9Y113_BO6),
.I4(CLBLM_R_X7Y113_SLICE_X8Y113_BO5),
.I5(CLBLM_R_X7Y113_SLICE_X9Y113_CO6),
.O5(CLBLM_R_X7Y113_SLICE_X9Y113_AO5),
.O6(CLBLM_R_X7Y113_SLICE_X9Y113_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X7Y114_SLICE_X8Y114_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y114_SLICE_X8Y114_DO5),
.O6(CLBLM_R_X7Y114_SLICE_X8Y114_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h33333333cccccfce)
  ) CLBLM_R_X7Y114_SLICE_X8Y114_CLUT (
.I0(LIOB33_X0Y103_IOB_X0Y103_I),
.I1(LIOB33_X0Y131_IOB_X0Y131_I),
.I2(LIOB33_X0Y95_IOB_X0Y95_I),
.I3(LIOB33_X0Y103_IOB_X0Y104_I),
.I4(LIOB33_X0Y131_IOB_X0Y132_I),
.I5(CLBLM_R_X7Y114_SLICE_X8Y114_BO6),
.O5(CLBLM_R_X7Y114_SLICE_X8Y114_CO5),
.O6(CLBLM_R_X7Y114_SLICE_X8Y114_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h5550555022232223)
  ) CLBLM_R_X7Y114_SLICE_X8Y114_BLUT (
.I0(LIOB33_X0Y95_IOB_X0Y95_I),
.I1(LIOB33_X0Y131_IOB_X0Y131_I),
.I2(LIOB33_X0Y101_IOB_X0Y102_I),
.I3(LIOB33_X0Y101_IOB_X0Y101_I),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y114_SLICE_X8Y114_BO5),
.O6(CLBLM_R_X7Y114_SLICE_X8Y114_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaa0000ccdcccfc)
  ) CLBLM_R_X7Y114_SLICE_X8Y114_ALUT (
.I0(LIOB33_X0Y69_IOB_X0Y70_I),
.I1(RIOB33_X105Y159_IOB_X1Y160_I),
.I2(LIOB33_X0Y123_IOB_X0Y123_I),
.I3(LIOB33_X0Y87_IOB_X0Y88_I),
.I4(LIOB33_X0Y67_IOB_X0Y68_I),
.I5(1'b1),
.O5(CLBLM_R_X7Y114_SLICE_X8Y114_AO5),
.O6(CLBLM_R_X7Y114_SLICE_X8Y114_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X7Y114_SLICE_X9Y114_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y114_SLICE_X9Y114_DO5),
.O6(CLBLM_R_X7Y114_SLICE_X9Y114_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X7Y114_SLICE_X9Y114_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y114_SLICE_X9Y114_CO5),
.O6(CLBLM_R_X7Y114_SLICE_X9Y114_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X7Y114_SLICE_X9Y114_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y114_SLICE_X9Y114_BO5),
.O6(CLBLM_R_X7Y114_SLICE_X9Y114_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h2222222222002200)
  ) CLBLM_R_X7Y114_SLICE_X9Y114_ALUT (
.I0(LIOB33_X0Y131_IOB_X0Y131_I),
.I1(LIOB33_X0Y101_IOB_X0Y101_I),
.I2(1'b1),
.I3(LIOB33_X0Y151_IOB_X0Y151_I),
.I4(1'b1),
.I5(LIOB33_SING_X0Y150_IOB_X0Y150_I),
.O5(CLBLM_R_X7Y114_SLICE_X9Y114_AO5),
.O6(CLBLM_R_X7Y114_SLICE_X9Y114_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X7Y121_SLICE_X8Y121_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y121_SLICE_X8Y121_DO5),
.O6(CLBLM_R_X7Y121_SLICE_X8Y121_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X7Y121_SLICE_X8Y121_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y121_SLICE_X8Y121_CO5),
.O6(CLBLM_R_X7Y121_SLICE_X8Y121_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0a0a0f0f0a0a0a0e)
  ) CLBLM_R_X7Y121_SLICE_X8Y121_BLUT (
.I0(LIOB33_X0Y159_IOB_X0Y160_I),
.I1(CLBLM_R_X5Y114_SLICE_X6Y114_CO6),
.I2(CLBLM_R_X7Y121_SLICE_X9Y121_AO5),
.I3(CLBLL_L_X4Y112_SLICE_X5Y112_CO6),
.I4(LIOB33_X0Y177_IOB_X0Y177_I),
.I5(LIOB33_X0Y159_IOB_X0Y159_I),
.O5(CLBLM_R_X7Y121_SLICE_X8Y121_BO5),
.O6(CLBLM_R_X7Y121_SLICE_X8Y121_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0a0a0f0a0a0a0f0e)
  ) CLBLM_R_X7Y121_SLICE_X8Y121_ALUT (
.I0(LIOB33_X0Y159_IOB_X0Y160_I),
.I1(CLBLM_R_X5Y114_SLICE_X6Y114_CO6),
.I2(CLBLM_R_X7Y121_SLICE_X9Y121_AO6),
.I3(LIOB33_X0Y159_IOB_X0Y159_I),
.I4(LIOB33_X0Y177_IOB_X0Y177_I),
.I5(CLBLL_L_X4Y112_SLICE_X5Y112_CO6),
.O5(CLBLM_R_X7Y121_SLICE_X8Y121_AO5),
.O6(CLBLM_R_X7Y121_SLICE_X8Y121_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X7Y121_SLICE_X9Y121_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y121_SLICE_X9Y121_DO5),
.O6(CLBLM_R_X7Y121_SLICE_X9Y121_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X7Y121_SLICE_X9Y121_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y121_SLICE_X9Y121_CO5),
.O6(CLBLM_R_X7Y121_SLICE_X9Y121_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X7Y121_SLICE_X9Y121_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y121_SLICE_X9Y121_BO5),
.O6(CLBLM_R_X7Y121_SLICE_X9Y121_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffafaffeeffee)
  ) CLBLM_R_X7Y121_SLICE_X9Y121_ALUT (
.I0(CLBLM_R_X7Y113_SLICE_X9Y113_AO6),
.I1(RIOB33_X105Y119_IOB_X1Y120_I),
.I2(LIOB33_X0Y161_IOB_X0Y162_I),
.I3(RIOB33_X105Y121_IOB_X1Y121_I),
.I4(RIOB33_X105Y105_IOB_X1Y105_I),
.I5(1'b1),
.O5(CLBLM_R_X7Y121_SLICE_X9Y121_AO5),
.O6(CLBLM_R_X7Y121_SLICE_X9Y121_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X25Y115_SLICE_X36Y115_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X25Y115_SLICE_X36Y115_DO5),
.O6(CLBLM_R_X25Y115_SLICE_X36Y115_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X25Y115_SLICE_X36Y115_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X25Y115_SLICE_X36Y115_CO5),
.O6(CLBLM_R_X25Y115_SLICE_X36Y115_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h888a888a888aaaaa)
  ) CLBLM_R_X25Y115_SLICE_X36Y115_BLUT (
.I0(CLBLM_L_X10Y123_SLICE_X12Y123_AO6),
.I1(RIOB33_X105Y157_IOB_X1Y157_I),
.I2(CLBLM_R_X5Y111_SLICE_X6Y111_AO6),
.I3(CLBLM_R_X5Y111_SLICE_X7Y111_AO5),
.I4(CLBLM_R_X25Y115_SLICE_X36Y115_AO6),
.I5(CLBLM_R_X5Y115_SLICE_X6Y115_AO6),
.O5(CLBLM_R_X25Y115_SLICE_X36Y115_BO5),
.O6(CLBLM_R_X25Y115_SLICE_X36Y115_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaaffffdddccccc)
  ) CLBLM_R_X25Y115_SLICE_X36Y115_ALUT (
.I0(LIOB33_X0Y59_IOB_X0Y60_I),
.I1(RIOB33_X105Y157_IOB_X1Y157_I),
.I2(LIOB33_SING_X0Y150_IOB_X0Y150_I),
.I3(LIOB33_X0Y151_IOB_X0Y151_I),
.I4(LIOB33_X0Y115_IOB_X0Y116_I),
.I5(1'b1),
.O5(CLBLM_R_X25Y115_SLICE_X36Y115_AO5),
.O6(CLBLM_R_X25Y115_SLICE_X36Y115_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X25Y115_SLICE_X37Y115_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X25Y115_SLICE_X37Y115_DO5),
.O6(CLBLM_R_X25Y115_SLICE_X37Y115_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X25Y115_SLICE_X37Y115_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X25Y115_SLICE_X37Y115_CO5),
.O6(CLBLM_R_X25Y115_SLICE_X37Y115_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X25Y115_SLICE_X37Y115_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X25Y115_SLICE_X37Y115_BO5),
.O6(CLBLM_R_X25Y115_SLICE_X37Y115_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X25Y115_SLICE_X37Y115_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X25Y115_SLICE_X37Y115_AO5),
.O6(CLBLM_R_X25Y115_SLICE_X37Y115_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X25Y116_SLICE_X36Y116_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X25Y116_SLICE_X36Y116_DO5),
.O6(CLBLM_R_X25Y116_SLICE_X36Y116_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X25Y116_SLICE_X36Y116_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X25Y116_SLICE_X36Y116_CO5),
.O6(CLBLM_R_X25Y116_SLICE_X36Y116_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'ha0a0a2a2a0aaa2aa)
  ) CLBLM_R_X25Y116_SLICE_X36Y116_BLUT (
.I0(CLBLM_L_X10Y123_SLICE_X12Y123_AO6),
.I1(CLBLM_R_X5Y115_SLICE_X6Y115_AO6),
.I2(RIOB33_X105Y157_IOB_X1Y158_I),
.I3(CLBLM_R_X5Y111_SLICE_X6Y111_AO6),
.I4(CLBLM_R_X25Y116_SLICE_X36Y116_AO6),
.I5(CLBLM_R_X3Y111_SLICE_X2Y111_AO5),
.O5(CLBLM_R_X25Y116_SLICE_X36Y116_BO5),
.O6(CLBLM_R_X25Y116_SLICE_X36Y116_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hff00fffff0fef0f0)
  ) CLBLM_R_X25Y116_SLICE_X36Y116_ALUT (
.I0(LIOB33_SING_X0Y150_IOB_X0Y150_I),
.I1(LIOB33_X0Y151_IOB_X0Y151_I),
.I2(RIOB33_X105Y157_IOB_X1Y158_I),
.I3(LIOB33_X0Y55_IOB_X0Y56_I),
.I4(LIOB33_X0Y119_IOB_X0Y120_I),
.I5(1'b1),
.O5(CLBLM_R_X25Y116_SLICE_X36Y116_AO5),
.O6(CLBLM_R_X25Y116_SLICE_X36Y116_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X25Y116_SLICE_X37Y116_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X25Y116_SLICE_X37Y116_DO5),
.O6(CLBLM_R_X25Y116_SLICE_X37Y116_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X25Y116_SLICE_X37Y116_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X25Y116_SLICE_X37Y116_CO5),
.O6(CLBLM_R_X25Y116_SLICE_X37Y116_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X25Y116_SLICE_X37Y116_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X25Y116_SLICE_X37Y116_BO5),
.O6(CLBLM_R_X25Y116_SLICE_X37Y116_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X25Y116_SLICE_X37Y116_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X25Y116_SLICE_X37Y116_AO5),
.O6(CLBLM_R_X25Y116_SLICE_X37Y116_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X29Y115_SLICE_X42Y115_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X29Y115_SLICE_X42Y115_DO5),
.O6(CLBLM_R_X29Y115_SLICE_X42Y115_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X29Y115_SLICE_X42Y115_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X29Y115_SLICE_X42Y115_CO5),
.O6(CLBLM_R_X29Y115_SLICE_X42Y115_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000555500005554)
  ) CLBLM_R_X29Y115_SLICE_X42Y115_BLUT (
.I0(LIOB33_X0Y157_IOB_X0Y158_I),
.I1(LIOB33_X0Y163_IOB_X0Y164_I),
.I2(CLBLM_L_X10Y114_SLICE_X12Y114_AO6),
.I3(CLBLM_R_X5Y112_SLICE_X6Y112_AO6),
.I4(LIOB33_X0Y157_IOB_X0Y157_I),
.I5(LIOB33_X0Y163_IOB_X0Y163_I),
.O5(CLBLM_R_X29Y115_SLICE_X42Y115_BO5),
.O6(CLBLM_R_X29Y115_SLICE_X42Y115_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000555500005554)
  ) CLBLM_R_X29Y115_SLICE_X42Y115_ALUT (
.I0(LIOB33_X0Y155_IOB_X0Y156_I),
.I1(LIOB33_X0Y163_IOB_X0Y164_I),
.I2(CLBLM_L_X10Y114_SLICE_X12Y114_AO6),
.I3(LIOB33_X0Y163_IOB_X0Y163_I),
.I4(LIOB33_X0Y153_IOB_X0Y154_I),
.I5(CLBLM_R_X5Y112_SLICE_X6Y112_AO6),
.O5(CLBLM_R_X29Y115_SLICE_X42Y115_AO5),
.O6(CLBLM_R_X29Y115_SLICE_X42Y115_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X29Y115_SLICE_X43Y115_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X29Y115_SLICE_X43Y115_DO5),
.O6(CLBLM_R_X29Y115_SLICE_X43Y115_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X29Y115_SLICE_X43Y115_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X29Y115_SLICE_X43Y115_CO5),
.O6(CLBLM_R_X29Y115_SLICE_X43Y115_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X29Y115_SLICE_X43Y115_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X29Y115_SLICE_X43Y115_BO5),
.O6(CLBLM_R_X29Y115_SLICE_X43Y115_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X29Y115_SLICE_X43Y115_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X29Y115_SLICE_X43Y115_AO5),
.O6(CLBLM_R_X29Y115_SLICE_X43Y115_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X49Y95_SLICE_X74Y95_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X49Y95_SLICE_X74Y95_DO5),
.O6(CLBLM_R_X49Y95_SLICE_X74Y95_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X49Y95_SLICE_X74Y95_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X49Y95_SLICE_X74Y95_CO5),
.O6(CLBLM_R_X49Y95_SLICE_X74Y95_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X49Y95_SLICE_X74Y95_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X49Y95_SLICE_X74Y95_BO5),
.O6(CLBLM_R_X49Y95_SLICE_X74Y95_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000fff033330003)
  ) CLBLM_R_X49Y95_SLICE_X74Y95_ALUT (
.I0(1'b1),
.I1(CLBLM_R_X5Y113_SLICE_X6Y113_AO6),
.I2(LIOB33_X0Y83_IOB_X0Y84_I),
.I3(LIOB33_X0Y85_IOB_X0Y85_I),
.I4(LIOB33_X0Y95_IOB_X0Y95_I),
.I5(1'b1),
.O5(CLBLM_R_X49Y95_SLICE_X74Y95_AO5),
.O6(CLBLM_R_X49Y95_SLICE_X74Y95_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X49Y95_SLICE_X75Y95_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X49Y95_SLICE_X75Y95_DO5),
.O6(CLBLM_R_X49Y95_SLICE_X75Y95_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X49Y95_SLICE_X75Y95_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X49Y95_SLICE_X75Y95_CO5),
.O6(CLBLM_R_X49Y95_SLICE_X75Y95_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X49Y95_SLICE_X75Y95_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X49Y95_SLICE_X75Y95_BO5),
.O6(CLBLM_R_X49Y95_SLICE_X75Y95_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X49Y95_SLICE_X75Y95_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X49Y95_SLICE_X75Y95_AO5),
.O6(CLBLM_R_X49Y95_SLICE_X75Y95_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X49Y101_SLICE_X74Y101_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X49Y101_SLICE_X74Y101_DO5),
.O6(CLBLM_R_X49Y101_SLICE_X74Y101_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X49Y101_SLICE_X74Y101_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X49Y101_SLICE_X74Y101_CO5),
.O6(CLBLM_R_X49Y101_SLICE_X74Y101_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X49Y101_SLICE_X74Y101_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X49Y101_SLICE_X74Y101_BO5),
.O6(CLBLM_R_X49Y101_SLICE_X74Y101_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hc3c6c3c63c39cccc)
  ) CLBLM_R_X49Y101_SLICE_X74Y101_ALUT (
.I0(LIOB33_X0Y83_IOB_X0Y84_I),
.I1(RIOB33_X105Y101_IOB_X1Y101_I),
.I2(LIOB33_X0Y95_IOB_X0Y95_I),
.I3(LIOB33_X0Y85_IOB_X0Y85_I),
.I4(CLBLM_R_X5Y113_SLICE_X6Y113_AO6),
.I5(1'b1),
.O5(CLBLM_R_X49Y101_SLICE_X74Y101_AO5),
.O6(CLBLM_R_X49Y101_SLICE_X74Y101_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X49Y101_SLICE_X75Y101_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X49Y101_SLICE_X75Y101_DO5),
.O6(CLBLM_R_X49Y101_SLICE_X75Y101_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X49Y101_SLICE_X75Y101_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X49Y101_SLICE_X75Y101_CO5),
.O6(CLBLM_R_X49Y101_SLICE_X75Y101_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X49Y101_SLICE_X75Y101_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X49Y101_SLICE_X75Y101_BO5),
.O6(CLBLM_R_X49Y101_SLICE_X75Y101_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X49Y101_SLICE_X75Y101_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X49Y101_SLICE_X75Y101_AO5),
.O6(CLBLM_R_X49Y101_SLICE_X75Y101_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X101Y116_SLICE_X158Y116_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X101Y116_SLICE_X158Y116_DO5),
.O6(CLBLM_R_X101Y116_SLICE_X158Y116_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X101Y116_SLICE_X158Y116_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X101Y116_SLICE_X158Y116_CO5),
.O6(CLBLM_R_X101Y116_SLICE_X158Y116_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X101Y116_SLICE_X158Y116_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X101Y116_SLICE_X158Y116_BO5),
.O6(CLBLM_R_X101Y116_SLICE_X158Y116_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffff0fffff1f0)
  ) CLBLM_R_X101Y116_SLICE_X158Y116_ALUT (
.I0(CLBLM_R_X7Y113_SLICE_X8Y113_DO6),
.I1(CLBLM_R_X5Y110_SLICE_X6Y110_AO5),
.I2(RIOB33_X105Y115_IOB_X1Y116_I),
.I3(CLBLM_L_X10Y123_SLICE_X12Y123_AO6),
.I4(LIOB33_SING_X0Y50_IOB_X0Y50_I),
.I5(CLBLM_R_X7Y114_SLICE_X8Y114_AO5),
.O5(CLBLM_R_X101Y116_SLICE_X158Y116_AO5),
.O6(CLBLM_R_X101Y116_SLICE_X158Y116_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X101Y116_SLICE_X159Y116_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X101Y116_SLICE_X159Y116_DO5),
.O6(CLBLM_R_X101Y116_SLICE_X159Y116_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X101Y116_SLICE_X159Y116_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X101Y116_SLICE_X159Y116_CO5),
.O6(CLBLM_R_X101Y116_SLICE_X159Y116_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X101Y116_SLICE_X159Y116_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X101Y116_SLICE_X159Y116_BO5),
.O6(CLBLM_R_X101Y116_SLICE_X159Y116_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X101Y116_SLICE_X159Y116_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X101Y116_SLICE_X159Y116_AO5),
.O6(CLBLM_R_X101Y116_SLICE_X159Y116_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X101Y117_SLICE_X158Y117_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X101Y117_SLICE_X158Y117_DO5),
.O6(CLBLM_R_X101Y117_SLICE_X158Y117_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X101Y117_SLICE_X158Y117_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X101Y117_SLICE_X158Y117_CO5),
.O6(CLBLM_R_X101Y117_SLICE_X158Y117_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X101Y117_SLICE_X158Y117_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X101Y117_SLICE_X158Y117_BO5),
.O6(CLBLM_R_X101Y117_SLICE_X158Y117_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffff0fffff1f0)
  ) CLBLM_R_X101Y117_SLICE_X158Y117_ALUT (
.I0(CLBLM_R_X7Y113_SLICE_X8Y113_DO6),
.I1(CLBLM_R_X5Y110_SLICE_X6Y110_AO5),
.I2(RIOB33_X105Y151_IOB_X1Y151_I),
.I3(CLBLM_L_X10Y123_SLICE_X12Y123_AO6),
.I4(RIOB33_X105Y151_IOB_X1Y152_I),
.I5(CLBLM_R_X7Y114_SLICE_X8Y114_AO5),
.O5(CLBLM_R_X101Y117_SLICE_X158Y117_AO5),
.O6(CLBLM_R_X101Y117_SLICE_X158Y117_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X101Y117_SLICE_X159Y117_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X101Y117_SLICE_X159Y117_DO5),
.O6(CLBLM_R_X101Y117_SLICE_X159Y117_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X101Y117_SLICE_X159Y117_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X101Y117_SLICE_X159Y117_CO5),
.O6(CLBLM_R_X101Y117_SLICE_X159Y117_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X101Y117_SLICE_X159Y117_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X101Y117_SLICE_X159Y117_BO5),
.O6(CLBLM_R_X101Y117_SLICE_X159Y117_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X101Y117_SLICE_X159Y117_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X101Y117_SLICE_X159Y117_AO5),
.O6(CLBLM_R_X101Y117_SLICE_X159Y117_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hfcfd0000cccc0000)
  ) CLBLM_R_X101Y118_SLICE_X158Y118_DLUT (
.I0(CLBLM_R_X5Y111_SLICE_X6Y111_AO6),
.I1(CLBLM_R_X101Y116_SLICE_X158Y116_AO6),
.I2(CLBLM_R_X5Y115_SLICE_X6Y115_BO5),
.I3(CLBLM_R_X5Y111_SLICE_X7Y111_AO6),
.I4(CLBLM_R_X103Y122_SLICE_X163Y122_BO5),
.I5(CLBLM_L_X10Y123_SLICE_X12Y123_AO6),
.O5(CLBLM_R_X101Y118_SLICE_X158Y118_DO5),
.O6(CLBLM_R_X101Y118_SLICE_X158Y118_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hfcfd0000cccc0000)
  ) CLBLM_R_X101Y118_SLICE_X158Y118_CLUT (
.I0(CLBLM_R_X5Y111_SLICE_X6Y111_AO6),
.I1(CLBLM_R_X101Y116_SLICE_X158Y116_AO6),
.I2(CLBLM_R_X5Y115_SLICE_X6Y115_BO5),
.I3(CLBLM_R_X5Y111_SLICE_X7Y111_AO6),
.I4(CLBLM_R_X103Y122_SLICE_X163Y122_AO5),
.I5(CLBLM_L_X10Y123_SLICE_X12Y123_AO6),
.O5(CLBLM_R_X101Y118_SLICE_X158Y118_CO5),
.O6(CLBLM_R_X101Y118_SLICE_X158Y118_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf800f800f800fc00)
  ) CLBLM_R_X101Y118_SLICE_X158Y118_BLUT (
.I0(CLBLM_R_X5Y115_SLICE_X6Y115_BO5),
.I1(CLBLM_L_X10Y123_SLICE_X12Y123_AO6),
.I2(CLBLM_R_X101Y117_SLICE_X158Y117_AO6),
.I3(CLBLL_L_X100Y123_SLICE_X156Y123_AO6),
.I4(CLBLM_R_X5Y111_SLICE_X6Y111_AO6),
.I5(CLBLM_R_X5Y111_SLICE_X7Y111_AO6),
.O5(CLBLM_R_X101Y118_SLICE_X158Y118_BO5),
.O6(CLBLM_R_X101Y118_SLICE_X158Y118_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hf800f800f800fc00)
  ) CLBLM_R_X101Y118_SLICE_X158Y118_ALUT (
.I0(CLBLM_R_X5Y115_SLICE_X6Y115_BO5),
.I1(CLBLM_L_X10Y123_SLICE_X12Y123_AO6),
.I2(CLBLM_R_X101Y117_SLICE_X158Y117_AO6),
.I3(CLBLL_L_X100Y123_SLICE_X156Y123_BO6),
.I4(CLBLM_R_X5Y111_SLICE_X6Y111_AO6),
.I5(CLBLM_R_X5Y111_SLICE_X7Y111_AO6),
.O5(CLBLM_R_X101Y118_SLICE_X158Y118_AO5),
.O6(CLBLM_R_X101Y118_SLICE_X158Y118_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X101Y118_SLICE_X159Y118_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X101Y118_SLICE_X159Y118_DO5),
.O6(CLBLM_R_X101Y118_SLICE_X159Y118_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X101Y118_SLICE_X159Y118_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X101Y118_SLICE_X159Y118_CO5),
.O6(CLBLM_R_X101Y118_SLICE_X159Y118_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X101Y118_SLICE_X159Y118_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X101Y118_SLICE_X159Y118_BO5),
.O6(CLBLM_R_X101Y118_SLICE_X159Y118_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X101Y118_SLICE_X159Y118_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X101Y118_SLICE_X159Y118_AO5),
.O6(CLBLM_R_X101Y118_SLICE_X159Y118_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hccc0c0c0ccc4c0c0)
  ) CLBLM_R_X101Y119_SLICE_X158Y119_DLUT (
.I0(CLBLM_R_X5Y111_SLICE_X7Y111_AO5),
.I1(CLBLM_R_X103Y122_SLICE_X163Y122_BO5),
.I2(CLBLM_L_X56Y119_SLICE_X84Y119_AO5),
.I3(CLBLM_R_X25Y115_SLICE_X36Y115_AO5),
.I4(CLBLM_L_X10Y123_SLICE_X12Y123_AO6),
.I5(CLBLM_R_X5Y111_SLICE_X6Y111_AO6),
.O5(CLBLM_R_X101Y119_SLICE_X158Y119_DO5),
.O6(CLBLM_R_X101Y119_SLICE_X158Y119_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hff00cd00ff000000)
  ) CLBLM_R_X101Y119_SLICE_X158Y119_CLUT (
.I0(CLBLM_R_X5Y111_SLICE_X6Y111_AO6),
.I1(CLBLM_R_X25Y115_SLICE_X36Y115_AO5),
.I2(CLBLM_R_X5Y111_SLICE_X7Y111_AO5),
.I3(CLBLM_R_X103Y122_SLICE_X163Y122_AO5),
.I4(CLBLM_L_X56Y119_SLICE_X84Y119_AO5),
.I5(CLBLM_L_X10Y123_SLICE_X12Y123_AO6),
.O5(CLBLM_R_X101Y119_SLICE_X158Y119_CO5),
.O6(CLBLM_R_X101Y119_SLICE_X158Y119_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hee00ee00aa00ae00)
  ) CLBLM_R_X101Y119_SLICE_X158Y119_BLUT (
.I0(CLBLM_L_X56Y119_SLICE_X84Y119_AO6),
.I1(CLBLM_L_X10Y123_SLICE_X12Y123_AO6),
.I2(CLBLM_R_X5Y111_SLICE_X7Y111_AO5),
.I3(CLBLL_L_X100Y123_SLICE_X156Y123_AO6),
.I4(CLBLM_R_X5Y111_SLICE_X6Y111_AO6),
.I5(CLBLM_R_X25Y115_SLICE_X36Y115_AO5),
.O5(CLBLM_R_X101Y119_SLICE_X158Y119_BO5),
.O6(CLBLM_R_X101Y119_SLICE_X158Y119_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hcc88cc88cc00cc08)
  ) CLBLM_R_X101Y119_SLICE_X158Y119_ALUT (
.I0(CLBLM_L_X10Y123_SLICE_X12Y123_AO6),
.I1(CLBLL_L_X100Y123_SLICE_X156Y123_BO6),
.I2(CLBLM_R_X5Y111_SLICE_X7Y111_AO5),
.I3(CLBLM_L_X56Y119_SLICE_X84Y119_AO6),
.I4(CLBLM_R_X5Y111_SLICE_X6Y111_AO6),
.I5(CLBLM_R_X25Y115_SLICE_X36Y115_AO5),
.O5(CLBLM_R_X101Y119_SLICE_X158Y119_AO5),
.O6(CLBLM_R_X101Y119_SLICE_X158Y119_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X101Y119_SLICE_X159Y119_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X101Y119_SLICE_X159Y119_DO5),
.O6(CLBLM_R_X101Y119_SLICE_X159Y119_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X101Y119_SLICE_X159Y119_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X101Y119_SLICE_X159Y119_CO5),
.O6(CLBLM_R_X101Y119_SLICE_X159Y119_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X101Y119_SLICE_X159Y119_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X101Y119_SLICE_X159Y119_BO5),
.O6(CLBLM_R_X101Y119_SLICE_X159Y119_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X101Y119_SLICE_X159Y119_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X101Y119_SLICE_X159Y119_AO5),
.O6(CLBLM_R_X101Y119_SLICE_X159Y119_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X101Y123_SLICE_X158Y123_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X101Y123_SLICE_X158Y123_DO5),
.O6(CLBLM_R_X101Y123_SLICE_X158Y123_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'heeaa0000eeae0000)
  ) CLBLM_R_X101Y123_SLICE_X158Y123_CLUT (
.I0(CLBLM_R_X101Y123_SLICE_X158Y123_AO6),
.I1(CLBLM_L_X10Y123_SLICE_X12Y123_AO6),
.I2(CLBLM_R_X5Y111_SLICE_X6Y111_AO6),
.I3(CLBLM_R_X25Y116_SLICE_X36Y116_AO5),
.I4(CLBLL_L_X100Y123_SLICE_X156Y123_AO6),
.I5(CLBLM_R_X3Y111_SLICE_X2Y111_AO5),
.O5(CLBLM_R_X101Y123_SLICE_X158Y123_CO5),
.O6(CLBLM_R_X101Y123_SLICE_X158Y123_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f0c0c0f0f00040)
  ) CLBLM_R_X101Y123_SLICE_X158Y123_BLUT (
.I0(CLBLM_R_X5Y111_SLICE_X6Y111_AO6),
.I1(CLBLM_L_X10Y123_SLICE_X12Y123_AO6),
.I2(CLBLL_L_X100Y123_SLICE_X156Y123_BO6),
.I3(CLBLM_R_X3Y111_SLICE_X2Y111_AO5),
.I4(CLBLM_R_X101Y123_SLICE_X158Y123_AO6),
.I5(CLBLM_R_X25Y116_SLICE_X36Y116_AO5),
.O5(CLBLM_R_X101Y123_SLICE_X158Y123_BO5),
.O6(CLBLM_R_X101Y123_SLICE_X158Y123_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffafffaffffffcc)
  ) CLBLM_R_X101Y123_SLICE_X158Y123_ALUT (
.I0(LIOB33_X0Y123_IOB_X0Y124_I),
.I1(RIOB33_X105Y115_IOB_X1Y115_I),
.I2(LIOB33_X0Y121_IOB_X0Y121_I),
.I3(CLBLM_L_X10Y113_SLICE_X12Y113_CO6),
.I4(RIOB33_X105Y125_IOB_X1Y126_I),
.I5(1'b1),
.O5(CLBLM_R_X101Y123_SLICE_X158Y123_AO5),
.O6(CLBLM_R_X101Y123_SLICE_X158Y123_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X101Y123_SLICE_X159Y123_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X101Y123_SLICE_X159Y123_DO5),
.O6(CLBLM_R_X101Y123_SLICE_X159Y123_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X101Y123_SLICE_X159Y123_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X101Y123_SLICE_X159Y123_CO5),
.O6(CLBLM_R_X101Y123_SLICE_X159Y123_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0c0f000f0c0f040)
  ) CLBLM_R_X101Y123_SLICE_X159Y123_BLUT (
.I0(CLBLM_R_X5Y111_SLICE_X6Y111_AO6),
.I1(CLBLM_L_X10Y123_SLICE_X12Y123_AO6),
.I2(CLBLM_R_X103Y122_SLICE_X163Y122_BO5),
.I3(CLBLM_R_X101Y123_SLICE_X158Y123_AO5),
.I4(CLBLM_R_X25Y116_SLICE_X36Y116_AO5),
.I5(CLBLM_R_X3Y111_SLICE_X2Y111_AO5),
.O5(CLBLM_R_X101Y123_SLICE_X159Y123_BO5),
.O6(CLBLM_R_X101Y123_SLICE_X159Y123_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hccc0c0c0ccc0c4c0)
  ) CLBLM_R_X101Y123_SLICE_X159Y123_ALUT (
.I0(CLBLM_R_X5Y111_SLICE_X6Y111_AO6),
.I1(CLBLM_R_X103Y122_SLICE_X163Y122_AO5),
.I2(CLBLM_R_X101Y123_SLICE_X158Y123_AO5),
.I3(CLBLM_L_X10Y123_SLICE_X12Y123_AO6),
.I4(CLBLM_R_X25Y116_SLICE_X36Y116_AO5),
.I5(CLBLM_R_X3Y111_SLICE_X2Y111_AO5),
.O5(CLBLM_R_X101Y123_SLICE_X159Y123_AO5),
.O6(CLBLM_R_X101Y123_SLICE_X159Y123_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y97_SLICE_X162Y97_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y97_SLICE_X162Y97_DO5),
.O6(CLBLM_R_X103Y97_SLICE_X162Y97_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y97_SLICE_X162Y97_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y97_SLICE_X162Y97_CO5),
.O6(CLBLM_R_X103Y97_SLICE_X162Y97_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y97_SLICE_X162Y97_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y97_SLICE_X162Y97_BO5),
.O6(CLBLM_R_X103Y97_SLICE_X162Y97_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y97_SLICE_X162Y97_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y97_SLICE_X162Y97_AO5),
.O6(CLBLM_R_X103Y97_SLICE_X162Y97_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y97_SLICE_X163Y97_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y97_SLICE_X163Y97_DO5),
.O6(CLBLM_R_X103Y97_SLICE_X163Y97_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y97_SLICE_X163Y97_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y97_SLICE_X163Y97_CO5),
.O6(CLBLM_R_X103Y97_SLICE_X163Y97_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaaaaaaaaaaaaa0)
  ) CLBLM_R_X103Y97_SLICE_X163Y97_BLUT (
.I0(CLBLM_R_X103Y122_SLICE_X163Y122_BO5),
.I1(1'b1),
.I2(RIOB33_X105Y117_IOB_X1Y118_I),
.I3(CLBLM_R_X5Y113_SLICE_X6Y113_BO6),
.I4(CLBLM_R_X5Y111_SLICE_X6Y111_BO6),
.I5(LIOB33_X0Y51_IOB_X0Y52_I),
.O5(CLBLM_R_X103Y97_SLICE_X163Y97_BO5),
.O6(CLBLM_R_X103Y97_SLICE_X163Y97_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffffc00000000)
  ) CLBLM_R_X103Y97_SLICE_X163Y97_ALUT (
.I0(1'b1),
.I1(CLBLM_R_X5Y113_SLICE_X6Y113_BO6),
.I2(RIOB33_X105Y117_IOB_X1Y118_I),
.I3(CLBLM_R_X5Y111_SLICE_X6Y111_BO6),
.I4(LIOB33_X0Y51_IOB_X0Y52_I),
.I5(CLBLM_R_X103Y122_SLICE_X163Y122_AO5),
.O5(CLBLM_R_X103Y97_SLICE_X163Y97_AO5),
.O6(CLBLM_R_X103Y97_SLICE_X163Y97_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y102_SLICE_X162Y102_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y102_SLICE_X162Y102_DO5),
.O6(CLBLM_R_X103Y102_SLICE_X162Y102_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y102_SLICE_X162Y102_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y102_SLICE_X162Y102_CO5),
.O6(CLBLM_R_X103Y102_SLICE_X162Y102_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y102_SLICE_X162Y102_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y102_SLICE_X162Y102_BO5),
.O6(CLBLM_R_X103Y102_SLICE_X162Y102_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y102_SLICE_X162Y102_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y102_SLICE_X162Y102_AO5),
.O6(CLBLM_R_X103Y102_SLICE_X162Y102_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y102_SLICE_X163Y102_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y102_SLICE_X163Y102_DO5),
.O6(CLBLM_R_X103Y102_SLICE_X163Y102_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y102_SLICE_X163Y102_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y102_SLICE_X163Y102_CO5),
.O6(CLBLM_R_X103Y102_SLICE_X163Y102_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff0000ffee0000)
  ) CLBLM_R_X103Y102_SLICE_X163Y102_BLUT (
.I0(CLBLM_R_X5Y113_SLICE_X6Y113_CO6),
.I1(CLBLM_L_X10Y113_SLICE_X12Y113_BO6),
.I2(1'b1),
.I3(RIOB33_X105Y109_IOB_X1Y110_I),
.I4(CLBLM_R_X103Y122_SLICE_X163Y122_BO5),
.I5(RIOB33_X105Y109_IOB_X1Y109_I),
.O5(CLBLM_R_X103Y102_SLICE_X163Y102_BO5),
.O6(CLBLM_R_X103Y102_SLICE_X163Y102_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f0f0f0f0e0f0e0)
  ) CLBLM_R_X103Y102_SLICE_X163Y102_ALUT (
.I0(CLBLM_R_X5Y113_SLICE_X6Y113_CO6),
.I1(CLBLM_L_X10Y113_SLICE_X12Y113_BO6),
.I2(CLBLM_R_X103Y122_SLICE_X163Y122_AO5),
.I3(RIOB33_X105Y109_IOB_X1Y110_I),
.I4(1'b1),
.I5(RIOB33_X105Y109_IOB_X1Y109_I),
.O5(CLBLM_R_X103Y102_SLICE_X163Y102_AO5),
.O6(CLBLM_R_X103Y102_SLICE_X163Y102_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y107_SLICE_X162Y107_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y107_SLICE_X162Y107_DO5),
.O6(CLBLM_R_X103Y107_SLICE_X162Y107_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y107_SLICE_X162Y107_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y107_SLICE_X162Y107_CO5),
.O6(CLBLM_R_X103Y107_SLICE_X162Y107_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y107_SLICE_X162Y107_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y107_SLICE_X162Y107_BO5),
.O6(CLBLM_R_X103Y107_SLICE_X162Y107_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y107_SLICE_X162Y107_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y107_SLICE_X162Y107_AO5),
.O6(CLBLM_R_X103Y107_SLICE_X162Y107_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y107_SLICE_X163Y107_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y107_SLICE_X163Y107_DO5),
.O6(CLBLM_R_X103Y107_SLICE_X163Y107_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y107_SLICE_X163Y107_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y107_SLICE_X163Y107_CO5),
.O6(CLBLM_R_X103Y107_SLICE_X163Y107_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffaff00000000)
  ) CLBLM_R_X103Y107_SLICE_X163Y107_BLUT (
.I0(RIOB33_X105Y111_IOB_X1Y111_I),
.I1(1'b1),
.I2(CLBLM_L_X8Y113_SLICE_X11Y113_BO6),
.I3(CLBLM_R_X5Y111_SLICE_X7Y111_CO6),
.I4(RIOB33_X105Y111_IOB_X1Y112_I),
.I5(CLBLM_R_X103Y122_SLICE_X163Y122_AO5),
.O5(CLBLM_R_X103Y107_SLICE_X163Y107_BO5),
.O6(CLBLM_R_X103Y107_SLICE_X163Y107_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hccccc8cc00ff00ff)
  ) CLBLM_R_X103Y107_SLICE_X163Y107_ALUT (
.I0(RIOB33_X105Y111_IOB_X1Y111_I),
.I1(CLBLM_R_X103Y122_SLICE_X163Y122_BO5),
.I2(CLBLM_L_X8Y113_SLICE_X11Y113_BO6),
.I3(CLBLM_R_X5Y111_SLICE_X7Y111_CO6),
.I4(RIOB33_X105Y111_IOB_X1Y112_I),
.I5(1'b1),
.O5(CLBLM_R_X103Y107_SLICE_X163Y107_AO5),
.O6(CLBLM_R_X103Y107_SLICE_X163Y107_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y108_SLICE_X162Y108_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y108_SLICE_X162Y108_DO5),
.O6(CLBLM_R_X103Y108_SLICE_X162Y108_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y108_SLICE_X162Y108_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y108_SLICE_X162Y108_CO5),
.O6(CLBLM_R_X103Y108_SLICE_X162Y108_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y108_SLICE_X162Y108_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y108_SLICE_X162Y108_BO5),
.O6(CLBLM_R_X103Y108_SLICE_X162Y108_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y108_SLICE_X162Y108_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y108_SLICE_X162Y108_AO5),
.O6(CLBLM_R_X103Y108_SLICE_X162Y108_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y108_SLICE_X163Y108_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y108_SLICE_X163Y108_DO5),
.O6(CLBLM_R_X103Y108_SLICE_X163Y108_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y108_SLICE_X163Y108_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y108_SLICE_X163Y108_CO5),
.O6(CLBLM_R_X103Y108_SLICE_X163Y108_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y108_SLICE_X163Y108_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y108_SLICE_X163Y108_BO5),
.O6(CLBLM_R_X103Y108_SLICE_X163Y108_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h33333333cc00cc00)
  ) CLBLM_R_X103Y108_SLICE_X163Y108_ALUT (
.I0(1'b1),
.I1(RIOB33_X105Y107_IOB_X1Y107_I),
.I2(1'b1),
.I3(RIOB33_X105Y107_IOB_X1Y108_I),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y108_SLICE_X163Y108_AO5),
.O6(CLBLM_R_X103Y108_SLICE_X163Y108_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y115_SLICE_X162Y115_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y115_SLICE_X162Y115_DO5),
.O6(CLBLM_R_X103Y115_SLICE_X162Y115_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y115_SLICE_X162Y115_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y115_SLICE_X162Y115_CO5),
.O6(CLBLM_R_X103Y115_SLICE_X162Y115_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y115_SLICE_X162Y115_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y115_SLICE_X162Y115_BO5),
.O6(CLBLM_R_X103Y115_SLICE_X162Y115_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y115_SLICE_X162Y115_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y115_SLICE_X162Y115_AO5),
.O6(CLBLM_R_X103Y115_SLICE_X162Y115_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y115_SLICE_X163Y115_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y115_SLICE_X163Y115_DO5),
.O6(CLBLM_R_X103Y115_SLICE_X163Y115_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y115_SLICE_X163Y115_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y115_SLICE_X163Y115_CO5),
.O6(CLBLM_R_X103Y115_SLICE_X163Y115_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y115_SLICE_X163Y115_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y115_SLICE_X163Y115_BO5),
.O6(CLBLM_R_X103Y115_SLICE_X163Y115_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000500000005)
  ) CLBLM_R_X103Y115_SLICE_X163Y115_ALUT (
.I0(RIOB33_X105Y123_IOB_X1Y124_I),
.I1(1'b1),
.I2(CLBLM_R_X5Y112_SLICE_X6Y112_AO6),
.I3(RIOB33_X105Y113_IOB_X1Y113_I),
.I4(CLBLM_L_X10Y114_SLICE_X12Y114_AO6),
.I5(1'b1),
.O5(CLBLM_R_X103Y115_SLICE_X163Y115_AO5),
.O6(CLBLM_R_X103Y115_SLICE_X163Y115_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y122_SLICE_X162Y122_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y122_SLICE_X162Y122_DO5),
.O6(CLBLM_R_X103Y122_SLICE_X162Y122_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y122_SLICE_X162Y122_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y122_SLICE_X162Y122_CO5),
.O6(CLBLM_R_X103Y122_SLICE_X162Y122_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y122_SLICE_X162Y122_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y122_SLICE_X162Y122_BO5),
.O6(CLBLM_R_X103Y122_SLICE_X162Y122_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffefefffffefe)
  ) CLBLM_R_X103Y122_SLICE_X162Y122_ALUT (
.I0(RIOB33_X105Y123_IOB_X1Y123_I),
.I1(RIOB33_X105Y121_IOB_X1Y122_I),
.I2(CLBLM_L_X10Y113_SLICE_X12Y113_AO6),
.I3(1'b1),
.I4(CLBLM_R_X5Y111_SLICE_X7Y111_BO6),
.I5(1'b1),
.O5(CLBLM_R_X103Y122_SLICE_X162Y122_AO5),
.O6(CLBLM_R_X103Y122_SLICE_X162Y122_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000050000000300)
  ) CLBLM_R_X103Y122_SLICE_X163Y122_DLUT (
.I0(CLBLM_R_X103Y115_SLICE_X163Y115_AO6),
.I1(CLBLM_R_X7Y121_SLICE_X8Y121_BO6),
.I2(LIOB33_X0Y141_IOB_X0Y142_I),
.I3(RIOB33_X105Y103_IOB_X1Y104_I),
.I4(LIOB33_X0Y143_IOB_X0Y143_I),
.I5(1'b1),
.O5(CLBLM_R_X103Y122_SLICE_X163Y122_DO5),
.O6(CLBLM_R_X103Y122_SLICE_X163Y122_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0101000000030000)
  ) CLBLM_R_X103Y122_SLICE_X163Y122_CLUT (
.I0(CLBLM_R_X103Y115_SLICE_X163Y115_AO6),
.I1(LIOB33_X0Y141_IOB_X0Y141_I),
.I2(LIOB33_X0Y139_IOB_X0Y140_I),
.I3(CLBLM_R_X7Y121_SLICE_X8Y121_BO6),
.I4(RIOB33_X105Y103_IOB_X1Y104_I),
.I5(1'b1),
.O5(CLBLM_R_X103Y122_SLICE_X163Y122_CO5),
.O6(CLBLM_R_X103Y122_SLICE_X163Y122_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0020002000220022)
  ) CLBLM_R_X103Y122_SLICE_X163Y122_BLUT (
.I0(RIOB33_X105Y103_IOB_X1Y104_I),
.I1(LIOB33_X0Y141_IOB_X0Y142_I),
.I2(CLBLM_R_X103Y122_SLICE_X162Y122_AO6),
.I3(LIOB33_X0Y143_IOB_X0Y143_I),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y122_SLICE_X163Y122_BO5),
.O6(CLBLM_R_X103Y122_SLICE_X163Y122_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0050000000550000)
  ) CLBLM_R_X103Y122_SLICE_X163Y122_ALUT (
.I0(LIOB33_X0Y139_IOB_X0Y140_I),
.I1(1'b1),
.I2(CLBLM_R_X103Y122_SLICE_X162Y122_AO6),
.I3(LIOB33_X0Y141_IOB_X0Y141_I),
.I4(RIOB33_X105Y103_IOB_X1Y104_I),
.I5(1'b1),
.O5(CLBLM_R_X103Y122_SLICE_X163Y122_AO5),
.O6(CLBLM_R_X103Y122_SLICE_X163Y122_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hdd00df00cc00cc00)
  ) CLBLM_R_X103Y123_SLICE_X162Y123_DLUT (
.I0(CLBLM_R_X5Y114_SLICE_X7Y114_AO6),
.I1(CLBLM_R_X103Y123_SLICE_X163Y123_AO5),
.I2(CLBLL_L_X4Y111_SLICE_X5Y111_AO5),
.I3(CLBLM_R_X103Y122_SLICE_X163Y122_BO5),
.I4(CLBLM_R_X5Y111_SLICE_X6Y111_AO6),
.I5(CLBLM_L_X10Y123_SLICE_X12Y123_AO6),
.O5(CLBLM_R_X103Y123_SLICE_X162Y123_DO5),
.O6(CLBLM_R_X103Y123_SLICE_X162Y123_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hdd00df00cc00cc00)
  ) CLBLM_R_X103Y123_SLICE_X162Y123_CLUT (
.I0(CLBLM_R_X5Y114_SLICE_X7Y114_AO6),
.I1(CLBLM_R_X103Y123_SLICE_X163Y123_AO5),
.I2(CLBLL_L_X4Y111_SLICE_X5Y111_AO5),
.I3(CLBLM_R_X103Y122_SLICE_X163Y122_AO5),
.I4(CLBLM_R_X5Y111_SLICE_X6Y111_AO6),
.I5(CLBLM_L_X10Y123_SLICE_X12Y123_AO6),
.O5(CLBLM_R_X103Y123_SLICE_X162Y123_CO5),
.O6(CLBLM_R_X103Y123_SLICE_X162Y123_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f4fcfc00000000)
  ) CLBLM_R_X103Y123_SLICE_X162Y123_BLUT (
.I0(CLBLL_L_X4Y111_SLICE_X5Y111_AO5),
.I1(CLBLM_L_X10Y123_SLICE_X12Y123_AO6),
.I2(CLBLM_R_X103Y123_SLICE_X163Y123_AO6),
.I3(CLBLM_R_X5Y111_SLICE_X6Y111_AO6),
.I4(CLBLM_R_X5Y114_SLICE_X7Y114_AO6),
.I5(CLBLL_L_X100Y123_SLICE_X156Y123_BO6),
.O5(CLBLM_R_X103Y123_SLICE_X162Y123_BO5),
.O6(CLBLM_R_X103Y123_SLICE_X162Y123_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f4fcfc00000000)
  ) CLBLM_R_X103Y123_SLICE_X162Y123_ALUT (
.I0(CLBLL_L_X4Y111_SLICE_X5Y111_AO5),
.I1(CLBLM_L_X10Y123_SLICE_X12Y123_AO6),
.I2(CLBLM_R_X103Y123_SLICE_X163Y123_AO6),
.I3(CLBLM_R_X5Y111_SLICE_X6Y111_AO6),
.I4(CLBLM_R_X5Y114_SLICE_X7Y114_AO6),
.I5(CLBLL_L_X100Y123_SLICE_X156Y123_AO6),
.O5(CLBLM_R_X103Y123_SLICE_X162Y123_AO5),
.O6(CLBLM_R_X103Y123_SLICE_X162Y123_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y123_SLICE_X163Y123_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y123_SLICE_X163Y123_DO5),
.O6(CLBLM_R_X103Y123_SLICE_X163Y123_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y123_SLICE_X163Y123_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y123_SLICE_X163Y123_CO5),
.O6(CLBLM_R_X103Y123_SLICE_X163Y123_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y123_SLICE_X163Y123_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y123_SLICE_X163Y123_BO5),
.O6(CLBLM_R_X103Y123_SLICE_X163Y123_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffeeeefffafffa)
  ) CLBLM_R_X103Y123_SLICE_X163Y123_ALUT (
.I0(CLBLM_L_X8Y113_SLICE_X10Y113_DO6),
.I1(RIOB33_X105Y153_IOB_X1Y154_I),
.I2(RIOB33_X105Y113_IOB_X1Y114_I),
.I3(RIOB33_X105Y125_IOB_X1Y125_I),
.I4(RIOB33_X105Y153_IOB_X1Y153_I),
.I5(1'b1),
.O5(CLBLM_R_X103Y123_SLICE_X163Y123_AO5),
.O6(CLBLM_R_X103Y123_SLICE_X163Y123_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y147_SLICE_X162Y147_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y147_SLICE_X162Y147_DO5),
.O6(CLBLM_R_X103Y147_SLICE_X162Y147_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y147_SLICE_X162Y147_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y147_SLICE_X162Y147_CO5),
.O6(CLBLM_R_X103Y147_SLICE_X162Y147_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y147_SLICE_X162Y147_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y147_SLICE_X162Y147_BO5),
.O6(CLBLM_R_X103Y147_SLICE_X162Y147_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y147_SLICE_X162Y147_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y147_SLICE_X162Y147_AO5),
.O6(CLBLM_R_X103Y147_SLICE_X162Y147_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y147_SLICE_X163Y147_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y147_SLICE_X163Y147_DO5),
.O6(CLBLM_R_X103Y147_SLICE_X163Y147_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y147_SLICE_X163Y147_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y147_SLICE_X163Y147_CO5),
.O6(CLBLM_R_X103Y147_SLICE_X163Y147_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y147_SLICE_X163Y147_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y147_SLICE_X163Y147_BO5),
.O6(CLBLM_R_X103Y147_SLICE_X163Y147_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'ha0a0a0a00f0f0f0f)
  ) CLBLM_R_X103Y147_SLICE_X163Y147_ALUT (
.I0(RIOB33_X105Y103_IOB_X1Y103_I),
.I1(1'b1),
.I2(LIOB33_X0Y147_IOB_X0Y147_I),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y147_SLICE_X163Y147_AO5),
.O6(CLBLM_R_X103Y147_SLICE_X163Y147_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y177_SLICE_X162Y177_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y177_SLICE_X162Y177_DO5),
.O6(CLBLM_R_X103Y177_SLICE_X162Y177_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y177_SLICE_X162Y177_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y177_SLICE_X162Y177_CO5),
.O6(CLBLM_R_X103Y177_SLICE_X162Y177_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y177_SLICE_X162Y177_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y177_SLICE_X162Y177_BO5),
.O6(CLBLM_R_X103Y177_SLICE_X162Y177_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y177_SLICE_X162Y177_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y177_SLICE_X162Y177_AO5),
.O6(CLBLM_R_X103Y177_SLICE_X162Y177_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y177_SLICE_X163Y177_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y177_SLICE_X163Y177_DO5),
.O6(CLBLM_R_X103Y177_SLICE_X163Y177_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y177_SLICE_X163Y177_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y177_SLICE_X163Y177_CO5),
.O6(CLBLM_R_X103Y177_SLICE_X163Y177_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y177_SLICE_X163Y177_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y177_SLICE_X163Y177_BO5),
.O6(CLBLM_R_X103Y177_SLICE_X163Y177_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h5f5f5f5f55555555)
  ) CLBLM_R_X103Y177_SLICE_X163Y177_ALUT (
.I0(RIOB33_SING_X105Y150_IOB_X1Y150_I),
.I1(1'b1),
.I2(LIOB33_X0Y107_IOB_X0Y108_I),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y177_SLICE_X163Y177_AO5),
.O6(CLBLM_R_X103Y177_SLICE_X163Y177_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y185_SLICE_X162Y185_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y185_SLICE_X162Y185_DO5),
.O6(CLBLM_R_X103Y185_SLICE_X162Y185_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y185_SLICE_X162Y185_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y185_SLICE_X162Y185_CO5),
.O6(CLBLM_R_X103Y185_SLICE_X162Y185_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y185_SLICE_X162Y185_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y185_SLICE_X162Y185_BO5),
.O6(CLBLM_R_X103Y185_SLICE_X162Y185_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y185_SLICE_X162Y185_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y185_SLICE_X162Y185_AO5),
.O6(CLBLM_R_X103Y185_SLICE_X162Y185_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y185_SLICE_X163Y185_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y185_SLICE_X163Y185_DO5),
.O6(CLBLM_R_X103Y185_SLICE_X163Y185_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y185_SLICE_X163Y185_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y185_SLICE_X163Y185_CO5),
.O6(CLBLM_R_X103Y185_SLICE_X163Y185_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y185_SLICE_X163Y185_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y185_SLICE_X163Y185_BO5),
.O6(CLBLM_R_X103Y185_SLICE_X163Y185_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h5555555555555555)
  ) CLBLM_R_X103Y185_SLICE_X163Y185_ALUT (
.I0(LIOB33_X0Y133_IOB_X0Y134_I),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y185_SLICE_X163Y185_AO5),
.O6(CLBLM_R_X103Y185_SLICE_X163Y185_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y193_SLICE_X162Y193_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y193_SLICE_X162Y193_DO5),
.O6(CLBLM_R_X103Y193_SLICE_X162Y193_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y193_SLICE_X162Y193_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y193_SLICE_X162Y193_CO5),
.O6(CLBLM_R_X103Y193_SLICE_X162Y193_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y193_SLICE_X162Y193_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y193_SLICE_X162Y193_BO5),
.O6(CLBLM_R_X103Y193_SLICE_X162Y193_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y193_SLICE_X162Y193_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y193_SLICE_X162Y193_AO5),
.O6(CLBLM_R_X103Y193_SLICE_X162Y193_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y193_SLICE_X163Y193_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y193_SLICE_X163Y193_DO5),
.O6(CLBLM_R_X103Y193_SLICE_X163Y193_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y193_SLICE_X163Y193_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y193_SLICE_X163Y193_CO5),
.O6(CLBLM_R_X103Y193_SLICE_X163Y193_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y193_SLICE_X163Y193_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y193_SLICE_X163Y193_BO5),
.O6(CLBLM_R_X103Y193_SLICE_X163Y193_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h00ff00ff00ff00ff)
  ) CLBLM_R_X103Y193_SLICE_X163Y193_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(LIOB33_X0Y85_IOB_X0Y85_I),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y193_SLICE_X163Y193_AO5),
.O6(CLBLM_R_X103Y193_SLICE_X163Y193_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y51_IOB_X0Y51_IBUF (
.I(LIOB33_X0Y51_IOB_X0Y51_IPAD),
.O(LIOB33_X0Y51_IOB_X0Y51_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y51_IOB_X0Y52_IBUF (
.I(LIOB33_X0Y51_IOB_X0Y52_IPAD),
.O(LIOB33_X0Y51_IOB_X0Y52_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y53_IOB_X0Y53_IBUF (
.I(LIOB33_X0Y53_IOB_X0Y53_IPAD),
.O(LIOB33_X0Y53_IOB_X0Y53_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y53_IOB_X0Y54_IBUF (
.I(LIOB33_X0Y53_IOB_X0Y54_IPAD),
.O(LIOB33_X0Y53_IOB_X0Y54_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y55_IOB_X0Y55_IBUF (
.I(LIOB33_X0Y55_IOB_X0Y55_IPAD),
.O(LIOB33_X0Y55_IOB_X0Y55_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y55_IOB_X0Y56_IBUF (
.I(LIOB33_X0Y55_IOB_X0Y56_IPAD),
.O(LIOB33_X0Y55_IOB_X0Y56_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y57_IOB_X0Y57_IBUF (
.I(LIOB33_X0Y57_IOB_X0Y57_IPAD),
.O(LIOB33_X0Y57_IOB_X0Y57_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y57_IOB_X0Y58_IBUF (
.I(LIOB33_X0Y57_IOB_X0Y58_IPAD),
.O(LIOB33_X0Y57_IOB_X0Y58_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y59_IOB_X0Y59_IBUF (
.I(LIOB33_X0Y59_IOB_X0Y59_IPAD),
.O(LIOB33_X0Y59_IOB_X0Y59_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y59_IOB_X0Y60_IBUF (
.I(LIOB33_X0Y59_IOB_X0Y60_IPAD),
.O(LIOB33_X0Y59_IOB_X0Y60_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y61_IOB_X0Y61_IBUF (
.I(LIOB33_X0Y61_IOB_X0Y61_IPAD),
.O(LIOB33_X0Y61_IOB_X0Y61_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y61_IOB_X0Y62_IBUF (
.I(LIOB33_X0Y61_IOB_X0Y62_IPAD),
.O(LIOB33_X0Y61_IOB_X0Y62_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y63_IOB_X0Y63_IBUF (
.I(LIOB33_X0Y63_IOB_X0Y63_IPAD),
.O(LIOB33_X0Y63_IOB_X0Y63_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y63_IOB_X0Y64_IBUF (
.I(LIOB33_X0Y63_IOB_X0Y64_IPAD),
.O(LIOB33_X0Y63_IOB_X0Y64_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y65_IOB_X0Y65_IBUF (
.I(LIOB33_X0Y65_IOB_X0Y65_IPAD),
.O(LIOB33_X0Y65_IOB_X0Y65_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y65_IOB_X0Y66_IBUF (
.I(LIOB33_X0Y65_IOB_X0Y66_IPAD),
.O(LIOB33_X0Y65_IOB_X0Y66_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y67_IOB_X0Y67_IBUF (
.I(LIOB33_X0Y67_IOB_X0Y67_IPAD),
.O(LIOB33_X0Y67_IOB_X0Y67_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y67_IOB_X0Y68_IBUF (
.I(LIOB33_X0Y67_IOB_X0Y68_IPAD),
.O(LIOB33_X0Y67_IOB_X0Y68_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y69_IOB_X0Y69_IBUF (
.I(LIOB33_X0Y69_IOB_X0Y69_IPAD),
.O(LIOB33_X0Y69_IOB_X0Y69_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y69_IOB_X0Y70_IBUF (
.I(LIOB33_X0Y69_IOB_X0Y70_IPAD),
.O(LIOB33_X0Y69_IOB_X0Y70_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y71_IOB_X0Y71_IBUF (
.I(LIOB33_X0Y71_IOB_X0Y71_IPAD),
.O(LIOB33_X0Y71_IOB_X0Y71_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y71_IOB_X0Y72_IBUF (
.I(LIOB33_X0Y71_IOB_X0Y72_IPAD),
.O(LIOB33_X0Y71_IOB_X0Y72_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y73_IOB_X0Y73_IBUF (
.I(LIOB33_X0Y73_IOB_X0Y73_IPAD),
.O(LIOB33_X0Y73_IOB_X0Y73_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y73_IOB_X0Y74_IBUF (
.I(LIOB33_X0Y73_IOB_X0Y74_IPAD),
.O(LIOB33_X0Y73_IOB_X0Y74_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y75_IOB_X0Y75_IBUF (
.I(LIOB33_X0Y75_IOB_X0Y75_IPAD),
.O(LIOB33_X0Y75_IOB_X0Y75_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y75_IOB_X0Y76_IBUF (
.I(LIOB33_X0Y75_IOB_X0Y76_IPAD),
.O(LIOB33_X0Y75_IOB_X0Y76_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y77_IOB_X0Y77_IBUF (
.I(LIOB33_X0Y77_IOB_X0Y77_IPAD),
.O(LIOB33_X0Y77_IOB_X0Y77_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y77_IOB_X0Y78_IBUF (
.I(LIOB33_X0Y77_IOB_X0Y78_IPAD),
.O(LIOB33_X0Y77_IOB_X0Y78_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y79_IOB_X0Y79_IBUF (
.I(LIOB33_X0Y79_IOB_X0Y79_IPAD),
.O(LIOB33_X0Y79_IOB_X0Y79_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y79_IOB_X0Y80_IBUF (
.I(LIOB33_X0Y79_IOB_X0Y80_IPAD),
.O(LIOB33_X0Y79_IOB_X0Y80_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y81_IOB_X0Y81_IBUF (
.I(LIOB33_X0Y81_IOB_X0Y81_IPAD),
.O(LIOB33_X0Y81_IOB_X0Y81_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y81_IOB_X0Y82_IBUF (
.I(LIOB33_X0Y81_IOB_X0Y82_IPAD),
.O(LIOB33_X0Y81_IOB_X0Y82_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y83_IOB_X0Y83_IBUF (
.I(LIOB33_X0Y83_IOB_X0Y83_IPAD),
.O(LIOB33_X0Y83_IOB_X0Y83_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y83_IOB_X0Y84_IBUF (
.I(LIOB33_X0Y83_IOB_X0Y84_IPAD),
.O(LIOB33_X0Y83_IOB_X0Y84_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y85_IOB_X0Y85_IBUF (
.I(LIOB33_X0Y85_IOB_X0Y85_IPAD),
.O(LIOB33_X0Y85_IOB_X0Y85_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y85_IOB_X0Y86_IBUF (
.I(LIOB33_X0Y85_IOB_X0Y86_IPAD),
.O(LIOB33_X0Y85_IOB_X0Y86_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y87_IOB_X0Y87_IBUF (
.I(LIOB33_X0Y87_IOB_X0Y87_IPAD),
.O(LIOB33_X0Y87_IOB_X0Y87_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y87_IOB_X0Y88_IBUF (
.I(LIOB33_X0Y87_IOB_X0Y88_IPAD),
.O(LIOB33_X0Y87_IOB_X0Y88_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y89_IOB_X0Y89_IBUF (
.I(LIOB33_X0Y89_IOB_X0Y89_IPAD),
.O(LIOB33_X0Y89_IOB_X0Y89_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y89_IOB_X0Y90_IBUF (
.I(LIOB33_X0Y89_IOB_X0Y90_IPAD),
.O(LIOB33_X0Y89_IOB_X0Y90_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y91_IOB_X0Y91_IBUF (
.I(LIOB33_X0Y91_IOB_X0Y91_IPAD),
.O(LIOB33_X0Y91_IOB_X0Y91_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y91_IOB_X0Y92_IBUF (
.I(LIOB33_X0Y91_IOB_X0Y92_IPAD),
.O(LIOB33_X0Y91_IOB_X0Y92_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y93_IOB_X0Y93_IBUF (
.I(LIOB33_X0Y93_IOB_X0Y93_IPAD),
.O(LIOB33_X0Y93_IOB_X0Y93_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y93_IOB_X0Y94_IBUF (
.I(LIOB33_X0Y93_IOB_X0Y94_IPAD),
.O(LIOB33_X0Y93_IOB_X0Y94_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y95_IOB_X0Y95_IBUF (
.I(LIOB33_X0Y95_IOB_X0Y95_IPAD),
.O(LIOB33_X0Y95_IOB_X0Y95_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y95_IOB_X0Y96_IBUF (
.I(LIOB33_X0Y95_IOB_X0Y96_IPAD),
.O(LIOB33_X0Y95_IOB_X0Y96_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y97_IOB_X0Y97_IBUF (
.I(LIOB33_X0Y97_IOB_X0Y97_IPAD),
.O(LIOB33_X0Y97_IOB_X0Y97_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y97_IOB_X0Y98_IBUF (
.I(LIOB33_X0Y97_IOB_X0Y98_IPAD),
.O(LIOB33_X0Y97_IOB_X0Y98_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y101_IOB_X0Y101_IBUF (
.I(LIOB33_X0Y101_IOB_X0Y101_IPAD),
.O(LIOB33_X0Y101_IOB_X0Y101_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y101_IOB_X0Y102_IBUF (
.I(LIOB33_X0Y101_IOB_X0Y102_IPAD),
.O(LIOB33_X0Y101_IOB_X0Y102_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y103_IOB_X0Y103_IBUF (
.I(LIOB33_X0Y103_IOB_X0Y103_IPAD),
.O(LIOB33_X0Y103_IOB_X0Y103_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y103_IOB_X0Y104_IBUF (
.I(LIOB33_X0Y103_IOB_X0Y104_IPAD),
.O(LIOB33_X0Y103_IOB_X0Y104_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y105_IOB_X0Y105_IBUF (
.I(LIOB33_X0Y105_IOB_X0Y105_IPAD),
.O(LIOB33_X0Y105_IOB_X0Y105_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y105_IOB_X0Y106_IBUF (
.I(LIOB33_X0Y105_IOB_X0Y106_IPAD),
.O(LIOB33_X0Y105_IOB_X0Y106_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y107_IOB_X0Y107_IBUF (
.I(LIOB33_X0Y107_IOB_X0Y107_IPAD),
.O(LIOB33_X0Y107_IOB_X0Y107_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y107_IOB_X0Y108_IBUF (
.I(LIOB33_X0Y107_IOB_X0Y108_IPAD),
.O(LIOB33_X0Y107_IOB_X0Y108_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y109_IOB_X0Y109_IBUF (
.I(LIOB33_X0Y109_IOB_X0Y109_IPAD),
.O(LIOB33_X0Y109_IOB_X0Y109_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y109_IOB_X0Y110_IBUF (
.I(LIOB33_X0Y109_IOB_X0Y110_IPAD),
.O(LIOB33_X0Y109_IOB_X0Y110_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y111_IOB_X0Y111_IBUF (
.I(LIOB33_X0Y111_IOB_X0Y111_IPAD),
.O(LIOB33_X0Y111_IOB_X0Y111_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y111_IOB_X0Y112_IBUF (
.I(LIOB33_X0Y111_IOB_X0Y112_IPAD),
.O(LIOB33_X0Y111_IOB_X0Y112_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y113_IOB_X0Y113_IBUF (
.I(LIOB33_X0Y113_IOB_X0Y113_IPAD),
.O(LIOB33_X0Y113_IOB_X0Y113_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y113_IOB_X0Y114_IBUF (
.I(LIOB33_X0Y113_IOB_X0Y114_IPAD),
.O(LIOB33_X0Y113_IOB_X0Y114_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y115_IOB_X0Y115_IBUF (
.I(LIOB33_X0Y115_IOB_X0Y115_IPAD),
.O(LIOB33_X0Y115_IOB_X0Y115_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y115_IOB_X0Y116_IBUF (
.I(LIOB33_X0Y115_IOB_X0Y116_IPAD),
.O(LIOB33_X0Y115_IOB_X0Y116_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y117_IOB_X0Y117_IBUF (
.I(LIOB33_X0Y117_IOB_X0Y117_IPAD),
.O(LIOB33_X0Y117_IOB_X0Y117_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y117_IOB_X0Y118_IBUF (
.I(LIOB33_X0Y117_IOB_X0Y118_IPAD),
.O(LIOB33_X0Y117_IOB_X0Y118_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y119_IOB_X0Y119_IBUF (
.I(LIOB33_X0Y119_IOB_X0Y119_IPAD),
.O(LIOB33_X0Y119_IOB_X0Y119_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y119_IOB_X0Y120_IBUF (
.I(LIOB33_X0Y119_IOB_X0Y120_IPAD),
.O(LIOB33_X0Y119_IOB_X0Y120_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y121_IOB_X0Y121_IBUF (
.I(LIOB33_X0Y121_IOB_X0Y121_IPAD),
.O(LIOB33_X0Y121_IOB_X0Y121_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y121_IOB_X0Y122_IBUF (
.I(LIOB33_X0Y121_IOB_X0Y122_IPAD),
.O(LIOB33_X0Y121_IOB_X0Y122_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y123_IOB_X0Y123_IBUF (
.I(LIOB33_X0Y123_IOB_X0Y123_IPAD),
.O(LIOB33_X0Y123_IOB_X0Y123_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y123_IOB_X0Y124_IBUF (
.I(LIOB33_X0Y123_IOB_X0Y124_IPAD),
.O(LIOB33_X0Y123_IOB_X0Y124_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y125_IOB_X0Y125_IBUF (
.I(LIOB33_X0Y125_IOB_X0Y125_IPAD),
.O(LIOB33_X0Y125_IOB_X0Y125_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y125_IOB_X0Y126_IBUF (
.I(LIOB33_X0Y125_IOB_X0Y126_IPAD),
.O(LIOB33_X0Y125_IOB_X0Y126_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y127_IOB_X0Y127_IBUF (
.I(LIOB33_X0Y127_IOB_X0Y127_IPAD),
.O(LIOB33_X0Y127_IOB_X0Y127_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y127_IOB_X0Y128_IBUF (
.I(LIOB33_X0Y127_IOB_X0Y128_IPAD),
.O(LIOB33_X0Y127_IOB_X0Y128_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y129_IOB_X0Y129_IBUF (
.I(LIOB33_X0Y129_IOB_X0Y129_IPAD),
.O(LIOB33_X0Y129_IOB_X0Y129_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y129_IOB_X0Y130_IBUF (
.I(LIOB33_X0Y129_IOB_X0Y130_IPAD),
.O(LIOB33_X0Y129_IOB_X0Y130_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y131_IOB_X0Y131_IBUF (
.I(LIOB33_X0Y131_IOB_X0Y131_IPAD),
.O(LIOB33_X0Y131_IOB_X0Y131_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y131_IOB_X0Y132_IBUF (
.I(LIOB33_X0Y131_IOB_X0Y132_IPAD),
.O(LIOB33_X0Y131_IOB_X0Y132_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y133_IOB_X0Y133_IBUF (
.I(LIOB33_X0Y133_IOB_X0Y133_IPAD),
.O(LIOB33_X0Y133_IOB_X0Y133_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y133_IOB_X0Y134_IBUF (
.I(LIOB33_X0Y133_IOB_X0Y134_IPAD),
.O(LIOB33_X0Y133_IOB_X0Y134_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y135_IOB_X0Y135_IBUF (
.I(LIOB33_X0Y135_IOB_X0Y135_IPAD),
.O(LIOB33_X0Y135_IOB_X0Y135_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y135_IOB_X0Y136_IBUF (
.I(LIOB33_X0Y135_IOB_X0Y136_IPAD),
.O(LIOB33_X0Y135_IOB_X0Y136_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y137_IOB_X0Y137_IBUF (
.I(LIOB33_X0Y137_IOB_X0Y137_IPAD),
.O(LIOB33_X0Y137_IOB_X0Y137_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y137_IOB_X0Y138_IBUF (
.I(LIOB33_X0Y137_IOB_X0Y138_IPAD),
.O(LIOB33_X0Y137_IOB_X0Y138_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y139_IOB_X0Y139_IBUF (
.I(LIOB33_X0Y139_IOB_X0Y139_IPAD),
.O(LIOB33_X0Y139_IOB_X0Y139_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y139_IOB_X0Y140_IBUF (
.I(LIOB33_X0Y139_IOB_X0Y140_IPAD),
.O(LIOB33_X0Y139_IOB_X0Y140_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y141_IOB_X0Y141_IBUF (
.I(LIOB33_X0Y141_IOB_X0Y141_IPAD),
.O(LIOB33_X0Y141_IOB_X0Y141_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y141_IOB_X0Y142_IBUF (
.I(LIOB33_X0Y141_IOB_X0Y142_IPAD),
.O(LIOB33_X0Y141_IOB_X0Y142_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y143_IOB_X0Y143_IBUF (
.I(LIOB33_X0Y143_IOB_X0Y143_IPAD),
.O(LIOB33_X0Y143_IOB_X0Y143_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y145_IOB_X0Y145_IBUF (
.I(LIOB33_X0Y145_IOB_X0Y145_IPAD),
.O(LIOB33_X0Y145_IOB_X0Y145_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y145_IOB_X0Y146_IBUF (
.I(LIOB33_X0Y145_IOB_X0Y146_IPAD),
.O(LIOB33_X0Y145_IOB_X0Y146_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y147_IOB_X0Y147_IBUF (
.I(LIOB33_X0Y147_IOB_X0Y147_IPAD),
.O(LIOB33_X0Y147_IOB_X0Y147_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y147_IOB_X0Y148_IBUF (
.I(LIOB33_X0Y147_IOB_X0Y148_IPAD),
.O(LIOB33_X0Y147_IOB_X0Y148_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y151_IOB_X0Y151_IBUF (
.I(LIOB33_X0Y151_IOB_X0Y151_IPAD),
.O(LIOB33_X0Y151_IOB_X0Y151_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y151_IOB_X0Y152_IBUF (
.I(LIOB33_X0Y151_IOB_X0Y152_IPAD),
.O(LIOB33_X0Y151_IOB_X0Y152_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y153_IOB_X0Y153_IBUF (
.I(LIOB33_X0Y153_IOB_X0Y153_IPAD),
.O(LIOB33_X0Y153_IOB_X0Y153_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y153_IOB_X0Y154_IBUF (
.I(LIOB33_X0Y153_IOB_X0Y154_IPAD),
.O(LIOB33_X0Y153_IOB_X0Y154_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y155_IOB_X0Y155_IBUF (
.I(LIOB33_X0Y155_IOB_X0Y155_IPAD),
.O(LIOB33_X0Y155_IOB_X0Y155_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y155_IOB_X0Y156_IBUF (
.I(LIOB33_X0Y155_IOB_X0Y156_IPAD),
.O(LIOB33_X0Y155_IOB_X0Y156_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y157_IOB_X0Y157_IBUF (
.I(LIOB33_X0Y157_IOB_X0Y157_IPAD),
.O(LIOB33_X0Y157_IOB_X0Y157_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y157_IOB_X0Y158_IBUF (
.I(LIOB33_X0Y157_IOB_X0Y158_IPAD),
.O(LIOB33_X0Y157_IOB_X0Y158_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y159_IOB_X0Y159_IBUF (
.I(LIOB33_X0Y159_IOB_X0Y159_IPAD),
.O(LIOB33_X0Y159_IOB_X0Y159_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y159_IOB_X0Y160_IBUF (
.I(LIOB33_X0Y159_IOB_X0Y160_IPAD),
.O(LIOB33_X0Y159_IOB_X0Y160_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y161_IOB_X0Y161_IBUF (
.I(LIOB33_X0Y161_IOB_X0Y161_IPAD),
.O(LIOB33_X0Y161_IOB_X0Y161_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y161_IOB_X0Y162_IBUF (
.I(LIOB33_X0Y161_IOB_X0Y162_IPAD),
.O(LIOB33_X0Y161_IOB_X0Y162_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y163_IOB_X0Y163_IBUF (
.I(LIOB33_X0Y163_IOB_X0Y163_IPAD),
.O(LIOB33_X0Y163_IOB_X0Y163_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y163_IOB_X0Y164_IBUF (
.I(LIOB33_X0Y163_IOB_X0Y164_IPAD),
.O(LIOB33_X0Y163_IOB_X0Y164_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y165_IOB_X0Y165_IBUF (
.I(LIOB33_X0Y165_IOB_X0Y165_IPAD),
.O(LIOB33_X0Y165_IOB_X0Y165_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y165_IOB_X0Y166_IBUF (
.I(LIOB33_X0Y165_IOB_X0Y166_IPAD),
.O(LIOB33_X0Y165_IOB_X0Y166_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y167_IOB_X0Y167_IBUF (
.I(LIOB33_X0Y167_IOB_X0Y167_IPAD),
.O(LIOB33_X0Y167_IOB_X0Y167_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y167_IOB_X0Y168_IBUF (
.I(LIOB33_X0Y167_IOB_X0Y168_IPAD),
.O(LIOB33_X0Y167_IOB_X0Y168_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y169_IOB_X0Y169_IBUF (
.I(LIOB33_X0Y169_IOB_X0Y169_IPAD),
.O(LIOB33_X0Y169_IOB_X0Y169_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y169_IOB_X0Y170_IBUF (
.I(LIOB33_X0Y169_IOB_X0Y170_IPAD),
.O(LIOB33_X0Y169_IOB_X0Y170_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y171_IOB_X0Y171_IBUF (
.I(LIOB33_X0Y171_IOB_X0Y171_IPAD),
.O(LIOB33_X0Y171_IOB_X0Y171_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y171_IOB_X0Y172_IBUF (
.I(LIOB33_X0Y171_IOB_X0Y172_IPAD),
.O(LIOB33_X0Y171_IOB_X0Y172_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y173_IOB_X0Y173_IBUF (
.I(LIOB33_X0Y173_IOB_X0Y173_IPAD),
.O(LIOB33_X0Y173_IOB_X0Y173_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y173_IOB_X0Y174_IBUF (
.I(LIOB33_X0Y173_IOB_X0Y174_IPAD),
.O(LIOB33_X0Y173_IOB_X0Y174_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y175_IOB_X0Y175_IBUF (
.I(LIOB33_X0Y175_IOB_X0Y175_IPAD),
.O(LIOB33_X0Y175_IOB_X0Y175_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y175_IOB_X0Y176_IBUF (
.I(LIOB33_X0Y175_IOB_X0Y176_IPAD),
.O(LIOB33_X0Y175_IOB_X0Y176_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y177_IOB_X0Y177_IBUF (
.I(LIOB33_X0Y177_IOB_X0Y177_IPAD),
.O(LIOB33_X0Y177_IOB_X0Y177_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y177_IOB_X0Y178_OBUF (
.I(CLBLL_L_X2Y175_SLICE_X0Y175_AO6),
.O(LIOB33_X0Y177_IOB_X0Y178_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y179_IOB_X0Y179_OBUF (
.I(LIOB33_X0Y133_IOB_X0Y134_I),
.O(LIOB33_X0Y179_IOB_X0Y179_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y179_IOB_X0Y180_OBUF (
.I(LIOB33_X0Y133_IOB_X0Y133_I),
.O(LIOB33_X0Y179_IOB_X0Y180_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y181_IOB_X0Y181_OBUF (
.I(LIOB33_X0Y133_IOB_X0Y133_I),
.O(LIOB33_X0Y181_IOB_X0Y181_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y181_IOB_X0Y182_OBUF (
.I(LIOB33_X0Y97_IOB_X0Y97_I),
.O(LIOB33_X0Y181_IOB_X0Y182_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y183_IOB_X0Y183_OBUF (
.I(LIOB33_X0Y101_IOB_X0Y102_I),
.O(LIOB33_X0Y183_IOB_X0Y183_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y183_IOB_X0Y184_OBUF (
.I(CLBLM_R_X103Y108_SLICE_X163Y108_AO5),
.O(LIOB33_X0Y183_IOB_X0Y184_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y185_IOB_X0Y185_OBUF (
.I(LIOB33_X0Y67_IOB_X0Y67_I),
.O(LIOB33_X0Y185_IOB_X0Y185_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y185_IOB_X0Y186_OBUF (
.I(LIOB33_X0Y135_IOB_X0Y135_I),
.O(LIOB33_X0Y185_IOB_X0Y186_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y187_IOB_X0Y187_OBUF (
.I(CLBLL_L_X2Y173_SLICE_X1Y173_BO6),
.O(LIOB33_X0Y187_IOB_X0Y187_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y187_IOB_X0Y188_OBUF (
.I(CLBLL_L_X2Y173_SLICE_X1Y173_BO6),
.O(LIOB33_X0Y187_IOB_X0Y188_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y189_IOB_X0Y189_OBUF (
.I(CLBLL_L_X2Y173_SLICE_X1Y173_BO6),
.O(LIOB33_X0Y189_IOB_X0Y189_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y189_IOB_X0Y190_OBUF (
.I(CLBLL_L_X2Y173_SLICE_X1Y173_BO6),
.O(LIOB33_X0Y189_IOB_X0Y190_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y191_IOB_X0Y191_OBUF (
.I(CLBLM_R_X5Y113_SLICE_X7Y113_AO6),
.O(LIOB33_X0Y191_IOB_X0Y191_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y191_IOB_X0Y192_OBUF (
.I(CLBLM_R_X5Y114_SLICE_X6Y114_AO6),
.O(LIOB33_X0Y191_IOB_X0Y192_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y193_IOB_X0Y193_OBUF (
.I(CLBLM_R_X3Y112_SLICE_X3Y112_BO6),
.O(LIOB33_X0Y193_IOB_X0Y193_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y193_IOB_X0Y194_OBUF (
.I(1'b0),
.O(LIOB33_X0Y193_IOB_X0Y194_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y195_IOB_X0Y195_OBUF (
.I(1'b0),
.O(LIOB33_X0Y195_IOB_X0Y195_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y195_IOB_X0Y196_OBUF (
.I(CLBLM_R_X3Y112_SLICE_X3Y112_BO6),
.O(LIOB33_X0Y195_IOB_X0Y196_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y197_IOB_X0Y197_OBUF (
.I(CLBLL_L_X4Y110_SLICE_X4Y110_CO5),
.O(LIOB33_X0Y197_IOB_X0Y197_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y197_IOB_X0Y198_OBUF (
.I(CLBLL_L_X2Y102_SLICE_X0Y102_BO6),
.O(LIOB33_X0Y197_IOB_X0Y198_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_SING_X0Y50_IOB_X0Y50_IBUF (
.I(LIOB33_SING_X0Y50_IOB_X0Y50_IPAD),
.O(LIOB33_SING_X0Y50_IOB_X0Y50_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_SING_X0Y99_IOB_X0Y99_IBUF (
.I(LIOB33_SING_X0Y99_IOB_X0Y99_IPAD),
.O(LIOB33_SING_X0Y99_IOB_X0Y99_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_SING_X0Y100_IOB_X0Y100_IBUF (
.I(LIOB33_SING_X0Y100_IOB_X0Y100_IPAD),
.O(LIOB33_SING_X0Y100_IOB_X0Y100_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_SING_X0Y149_IOB_X0Y149_IBUF (
.I(LIOB33_SING_X0Y149_IOB_X0Y149_IPAD),
.O(LIOB33_SING_X0Y149_IOB_X0Y149_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_SING_X0Y150_IOB_X0Y150_IBUF (
.I(LIOB33_SING_X0Y150_IOB_X0Y150_IPAD),
.O(LIOB33_SING_X0Y150_IOB_X0Y150_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_SING_X0Y199_IOB_X0Y199_OBUF (
.I(CLBLL_L_X4Y111_SLICE_X5Y111_CO6),
.O(LIOB33_SING_X0Y199_IOB_X0Y199_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_SING_X0Y200_IOB_X0Y200_OBUF (
.I(LIOB33_SING_X0Y100_IOB_X0Y100_I),
.O(LIOB33_SING_X0Y200_IOB_X0Y200_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y51_IOB_X1Y51_OBUF (
.I(CLBLL_L_X4Y111_SLICE_X5Y111_CO6),
.O(RIOB33_X105Y51_IOB_X1Y51_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y51_IOB_X1Y52_OBUF (
.I(CLBLM_R_X49Y95_SLICE_X74Y95_AO6),
.O(RIOB33_X105Y51_IOB_X1Y52_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y53_IOB_X1Y53_OBUF (
.I(CLBLM_L_X10Y113_SLICE_X12Y113_AO6),
.O(RIOB33_X105Y53_IOB_X1Y53_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y53_IOB_X1Y54_OBUF (
.I(CLBLM_R_X103Y108_SLICE_X163Y108_AO6),
.O(RIOB33_X105Y53_IOB_X1Y54_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y55_IOB_X1Y55_OBUF (
.I(CLBLM_L_X10Y114_SLICE_X12Y114_AO6),
.O(RIOB33_X105Y55_IOB_X1Y55_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y55_IOB_X1Y56_OBUF (
.I(CLBLM_R_X5Y111_SLICE_X7Y111_BO6),
.O(RIOB33_X105Y55_IOB_X1Y56_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y57_IOB_X1Y57_OBUF (
.I(CLBLM_R_X49Y95_SLICE_X74Y95_AO5),
.O(RIOB33_X105Y57_IOB_X1Y57_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y57_IOB_X1Y58_OBUF (
.I(CLBLL_L_X100Y121_SLICE_X156Y121_AO6),
.O(RIOB33_X105Y57_IOB_X1Y58_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y59_IOB_X1Y59_OBUF (
.I(CLBLM_R_X5Y113_SLICE_X6Y113_BO6),
.O(RIOB33_X105Y59_IOB_X1Y59_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y59_IOB_X1Y60_OBUF (
.I(CLBLM_L_X10Y113_SLICE_X12Y113_BO6),
.O(RIOB33_X105Y59_IOB_X1Y60_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y61_IOB_X1Y61_OBUF (
.I(CLBLM_L_X8Y113_SLICE_X11Y113_BO6),
.O(RIOB33_X105Y61_IOB_X1Y61_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y61_IOB_X1Y62_OBUF (
.I(CLBLL_L_X100Y121_SLICE_X156Y121_BO6),
.O(RIOB33_X105Y61_IOB_X1Y62_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y63_IOB_X1Y63_OBUF (
.I(CLBLM_R_X5Y111_SLICE_X6Y111_BO6),
.O(RIOB33_X105Y63_IOB_X1Y63_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y63_IOB_X1Y64_OBUF (
.I(CLBLM_R_X5Y113_SLICE_X6Y113_CO6),
.O(RIOB33_X105Y63_IOB_X1Y64_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y65_IOB_X1Y65_OBUF (
.I(CLBLM_R_X103Y107_SLICE_X163Y107_AO5),
.O(RIOB33_X105Y65_IOB_X1Y65_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y65_IOB_X1Y66_OBUF (
.I(CLBLM_R_X5Y112_SLICE_X6Y112_AO6),
.O(RIOB33_X105Y65_IOB_X1Y66_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y67_IOB_X1Y67_OBUF (
.I(CLBLM_R_X5Y109_SLICE_X6Y109_AO6),
.O(RIOB33_X105Y67_IOB_X1Y67_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y67_IOB_X1Y68_OBUF (
.I(CLBLL_L_X4Y109_SLICE_X4Y109_AO6),
.O(RIOB33_X105Y67_IOB_X1Y68_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y69_IOB_X1Y69_OBUF (
.I(CLBLM_R_X5Y111_SLICE_X6Y111_CO6),
.O(RIOB33_X105Y69_IOB_X1Y69_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y69_IOB_X1Y70_OBUF (
.I(CLBLM_L_X8Y113_SLICE_X11Y113_CO6),
.O(RIOB33_X105Y69_IOB_X1Y70_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y71_IOB_X1Y71_OBUF (
.I(CLBLM_R_X103Y122_SLICE_X163Y122_AO6),
.O(RIOB33_X105Y71_IOB_X1Y71_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y71_IOB_X1Y72_OBUF (
.I(CLBLM_R_X103Y122_SLICE_X163Y122_BO6),
.O(RIOB33_X105Y71_IOB_X1Y72_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y73_IOB_X1Y73_OBUF (
.I(CLBLL_L_X36Y113_SLICE_X54Y113_AO6),
.O(RIOB33_X105Y73_IOB_X1Y73_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y73_IOB_X1Y74_OBUF (
.I(CLBLL_L_X100Y113_SLICE_X156Y113_AO6),
.O(RIOB33_X105Y73_IOB_X1Y74_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y75_IOB_X1Y75_OBUF (
.I(CLBLM_R_X29Y115_SLICE_X42Y115_AO6),
.O(RIOB33_X105Y75_IOB_X1Y75_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y75_IOB_X1Y76_OBUF (
.I(CLBLL_R_X57Y113_SLICE_X86Y113_BO6),
.O(RIOB33_X105Y75_IOB_X1Y76_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y77_IOB_X1Y77_OBUF (
.I(CLBLL_L_X36Y113_SLICE_X54Y113_BO6),
.O(RIOB33_X105Y77_IOB_X1Y77_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y77_IOB_X1Y78_OBUF (
.I(CLBLL_L_X100Y113_SLICE_X156Y113_BO6),
.O(RIOB33_X105Y77_IOB_X1Y78_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y79_IOB_X1Y79_OBUF (
.I(CLBLM_R_X29Y115_SLICE_X42Y115_BO6),
.O(RIOB33_X105Y79_IOB_X1Y79_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y79_IOB_X1Y80_OBUF (
.I(CLBLM_R_X103Y97_SLICE_X163Y97_AO6),
.O(RIOB33_X105Y79_IOB_X1Y80_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y81_IOB_X1Y81_OBUF (
.I(CLBLM_R_X103Y122_SLICE_X163Y122_CO6),
.O(RIOB33_X105Y81_IOB_X1Y81_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y81_IOB_X1Y82_OBUF (
.I(CLBLM_R_X103Y107_SLICE_X163Y107_BO6),
.O(RIOB33_X105Y81_IOB_X1Y82_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y83_IOB_X1Y83_OBUF (
.I(CLBLM_R_X103Y102_SLICE_X163Y102_AO6),
.O(RIOB33_X105Y83_IOB_X1Y83_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y83_IOB_X1Y84_OBUF (
.I(CLBLM_R_X103Y97_SLICE_X163Y97_BO6),
.O(RIOB33_X105Y83_IOB_X1Y84_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y85_IOB_X1Y85_OBUF (
.I(CLBLM_R_X103Y122_SLICE_X163Y122_DO6),
.O(RIOB33_X105Y85_IOB_X1Y85_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y85_IOB_X1Y86_OBUF (
.I(CLBLM_R_X103Y107_SLICE_X163Y107_AO6),
.O(RIOB33_X105Y85_IOB_X1Y86_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y87_IOB_X1Y87_OBUF (
.I(CLBLM_R_X103Y102_SLICE_X163Y102_BO6),
.O(RIOB33_X105Y87_IOB_X1Y87_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y87_IOB_X1Y88_OBUF (
.I(CLBLM_L_X8Y113_SLICE_X10Y113_BO6),
.O(RIOB33_X105Y87_IOB_X1Y88_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y89_IOB_X1Y89_OBUF (
.I(CLBLM_R_X49Y101_SLICE_X74Y101_AO5),
.O(RIOB33_X105Y89_IOB_X1Y89_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y89_IOB_X1Y90_OBUF (
.I(CLBLM_L_X8Y113_SLICE_X10Y113_DO6),
.O(RIOB33_X105Y89_IOB_X1Y90_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y91_IOB_X1Y91_OBUF (
.I(CLBLM_L_X10Y113_SLICE_X12Y113_CO6),
.O(RIOB33_X105Y91_IOB_X1Y91_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y91_IOB_X1Y92_OBUF (
.I(CLBLM_L_X10Y113_SLICE_X13Y113_AO6),
.O(RIOB33_X105Y91_IOB_X1Y92_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y93_IOB_X1Y93_OBUF (
.I(CLBLM_L_X10Y113_SLICE_X13Y113_BO6),
.O(RIOB33_X105Y93_IOB_X1Y93_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y93_IOB_X1Y94_OBUF (
.I(CLBLL_L_X4Y109_SLICE_X4Y109_AO5),
.O(RIOB33_X105Y93_IOB_X1Y94_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y95_IOB_X1Y95_OBUF (
.I(CLBLM_L_X10Y114_SLICE_X12Y114_BO6),
.O(RIOB33_X105Y95_IOB_X1Y95_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y95_IOB_X1Y96_OBUF (
.I(CLBLM_R_X25Y116_SLICE_X36Y116_BO6),
.O(RIOB33_X105Y95_IOB_X1Y96_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y97_IOB_X1Y97_OBUF (
.I(CLBLM_R_X5Y115_SLICE_X7Y115_AO6),
.O(RIOB33_X105Y97_IOB_X1Y97_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y97_IOB_X1Y98_OBUF (
.I(CLBLM_R_X25Y115_SLICE_X36Y115_BO6),
.O(RIOB33_X105Y97_IOB_X1Y98_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y101_IOB_X1Y101_IBUF (
.I(RIOB33_X105Y101_IOB_X1Y101_IPAD),
.O(RIOB33_X105Y101_IOB_X1Y101_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y101_IOB_X1Y102_IBUF (
.I(RIOB33_X105Y101_IOB_X1Y102_IPAD),
.O(RIOB33_X105Y101_IOB_X1Y102_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y103_IOB_X1Y103_IBUF (
.I(RIOB33_X105Y103_IOB_X1Y103_IPAD),
.O(RIOB33_X105Y103_IOB_X1Y103_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y103_IOB_X1Y104_IBUF (
.I(RIOB33_X105Y103_IOB_X1Y104_IPAD),
.O(RIOB33_X105Y103_IOB_X1Y104_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y105_IOB_X1Y105_IBUF (
.I(RIOB33_X105Y105_IOB_X1Y105_IPAD),
.O(RIOB33_X105Y105_IOB_X1Y105_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y105_IOB_X1Y106_IBUF (
.I(RIOB33_X105Y105_IOB_X1Y106_IPAD),
.O(RIOB33_X105Y105_IOB_X1Y106_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y107_IOB_X1Y107_IBUF (
.I(RIOB33_X105Y107_IOB_X1Y107_IPAD),
.O(RIOB33_X105Y107_IOB_X1Y107_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y107_IOB_X1Y108_IBUF (
.I(RIOB33_X105Y107_IOB_X1Y108_IPAD),
.O(RIOB33_X105Y107_IOB_X1Y108_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y109_IOB_X1Y109_IBUF (
.I(RIOB33_X105Y109_IOB_X1Y109_IPAD),
.O(RIOB33_X105Y109_IOB_X1Y109_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y109_IOB_X1Y110_IBUF (
.I(RIOB33_X105Y109_IOB_X1Y110_IPAD),
.O(RIOB33_X105Y109_IOB_X1Y110_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y111_IOB_X1Y111_IBUF (
.I(RIOB33_X105Y111_IOB_X1Y111_IPAD),
.O(RIOB33_X105Y111_IOB_X1Y111_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y111_IOB_X1Y112_IBUF (
.I(RIOB33_X105Y111_IOB_X1Y112_IPAD),
.O(RIOB33_X105Y111_IOB_X1Y112_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y113_IOB_X1Y113_IBUF (
.I(RIOB33_X105Y113_IOB_X1Y113_IPAD),
.O(RIOB33_X105Y113_IOB_X1Y113_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y113_IOB_X1Y114_IBUF (
.I(RIOB33_X105Y113_IOB_X1Y114_IPAD),
.O(RIOB33_X105Y113_IOB_X1Y114_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y115_IOB_X1Y115_IBUF (
.I(RIOB33_X105Y115_IOB_X1Y115_IPAD),
.O(RIOB33_X105Y115_IOB_X1Y115_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y115_IOB_X1Y116_IBUF (
.I(RIOB33_X105Y115_IOB_X1Y116_IPAD),
.O(RIOB33_X105Y115_IOB_X1Y116_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y117_IOB_X1Y117_IBUF (
.I(RIOB33_X105Y117_IOB_X1Y117_IPAD),
.O(RIOB33_X105Y117_IOB_X1Y117_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y117_IOB_X1Y118_IBUF (
.I(RIOB33_X105Y117_IOB_X1Y118_IPAD),
.O(RIOB33_X105Y117_IOB_X1Y118_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y119_IOB_X1Y119_IBUF (
.I(RIOB33_X105Y119_IOB_X1Y119_IPAD),
.O(RIOB33_X105Y119_IOB_X1Y119_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y119_IOB_X1Y120_IBUF (
.I(RIOB33_X105Y119_IOB_X1Y120_IPAD),
.O(RIOB33_X105Y119_IOB_X1Y120_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y121_IOB_X1Y121_IBUF (
.I(RIOB33_X105Y121_IOB_X1Y121_IPAD),
.O(RIOB33_X105Y121_IOB_X1Y121_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y121_IOB_X1Y122_IBUF (
.I(RIOB33_X105Y121_IOB_X1Y122_IPAD),
.O(RIOB33_X105Y121_IOB_X1Y122_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y123_IOB_X1Y123_IBUF (
.I(RIOB33_X105Y123_IOB_X1Y123_IPAD),
.O(RIOB33_X105Y123_IOB_X1Y123_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y123_IOB_X1Y124_IBUF (
.I(RIOB33_X105Y123_IOB_X1Y124_IPAD),
.O(RIOB33_X105Y123_IOB_X1Y124_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y125_IOB_X1Y125_IBUF (
.I(RIOB33_X105Y125_IOB_X1Y125_IPAD),
.O(RIOB33_X105Y125_IOB_X1Y125_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y125_IOB_X1Y126_IBUF (
.I(RIOB33_X105Y125_IOB_X1Y126_IPAD),
.O(RIOB33_X105Y125_IOB_X1Y126_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y127_IOB_X1Y127_OBUF (
.I(CLBLL_R_X57Y113_SLICE_X86Y113_AO6),
.O(RIOB33_X105Y127_IOB_X1Y127_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y127_IOB_X1Y128_OBUF (
.I(CLBLM_R_X103Y123_SLICE_X162Y123_AO6),
.O(RIOB33_X105Y127_IOB_X1Y128_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y129_IOB_X1Y129_OBUF (
.I(CLBLM_R_X103Y123_SLICE_X162Y123_BO6),
.O(RIOB33_X105Y129_IOB_X1Y129_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y129_IOB_X1Y130_OBUF (
.I(CLBLM_R_X101Y123_SLICE_X158Y123_BO6),
.O(RIOB33_X105Y129_IOB_X1Y130_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y131_IOB_X1Y131_OBUF (
.I(CLBLM_R_X101Y118_SLICE_X158Y118_AO6),
.O(RIOB33_X105Y131_IOB_X1Y131_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y131_IOB_X1Y132_OBUF (
.I(CLBLM_R_X101Y119_SLICE_X158Y119_AO6),
.O(RIOB33_X105Y131_IOB_X1Y132_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y133_IOB_X1Y133_OBUF (
.I(CLBLM_R_X101Y123_SLICE_X158Y123_CO6),
.O(RIOB33_X105Y133_IOB_X1Y133_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y133_IOB_X1Y134_OBUF (
.I(CLBLM_R_X101Y118_SLICE_X158Y118_BO6),
.O(RIOB33_X105Y133_IOB_X1Y134_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y135_IOB_X1Y135_OBUF (
.I(CLBLM_R_X101Y119_SLICE_X158Y119_CO6),
.O(RIOB33_X105Y135_IOB_X1Y135_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y135_IOB_X1Y136_OBUF (
.I(CLBLM_R_X101Y118_SLICE_X158Y118_CO6),
.O(RIOB33_X105Y135_IOB_X1Y136_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y137_IOB_X1Y137_OBUF (
.I(CLBLM_R_X101Y123_SLICE_X159Y123_AO6),
.O(RIOB33_X105Y137_IOB_X1Y137_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y137_IOB_X1Y138_OBUF (
.I(CLBLM_R_X103Y123_SLICE_X162Y123_CO6),
.O(RIOB33_X105Y137_IOB_X1Y138_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y139_IOB_X1Y139_OBUF (
.I(CLBLM_R_X101Y119_SLICE_X158Y119_DO6),
.O(RIOB33_X105Y139_IOB_X1Y139_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y139_IOB_X1Y140_OBUF (
.I(CLBLM_R_X101Y118_SLICE_X158Y118_DO6),
.O(RIOB33_X105Y139_IOB_X1Y140_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y141_IOB_X1Y141_OBUF (
.I(CLBLM_R_X101Y123_SLICE_X159Y123_BO6),
.O(RIOB33_X105Y141_IOB_X1Y141_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y141_IOB_X1Y142_OBUF (
.I(CLBLM_R_X103Y123_SLICE_X162Y123_DO6),
.O(RIOB33_X105Y141_IOB_X1Y142_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y143_IOB_X1Y143_OBUF (
.I(CLBLM_L_X10Y123_SLICE_X12Y123_AO6),
.O(RIOB33_X105Y143_IOB_X1Y143_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y143_IOB_X1Y144_OBUF (
.I(CLBLM_L_X10Y123_SLICE_X12Y123_AO6),
.O(RIOB33_X105Y143_IOB_X1Y144_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y145_IOB_X1Y145_OBUF (
.I(CLBLL_L_X100Y123_SLICE_X156Y123_BO5),
.O(RIOB33_X105Y145_IOB_X1Y145_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y145_IOB_X1Y146_OBUF (
.I(CLBLL_L_X100Y123_SLICE_X156Y123_AO5),
.O(RIOB33_X105Y145_IOB_X1Y146_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y147_IOB_X1Y147_OBUF (
.I(CLBLM_R_X103Y122_SLICE_X163Y122_CO5),
.O(RIOB33_X105Y147_IOB_X1Y147_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y147_IOB_X1Y148_OBUF (
.I(CLBLM_R_X103Y122_SLICE_X163Y122_DO5),
.O(RIOB33_X105Y147_IOB_X1Y148_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y151_IOB_X1Y151_IBUF (
.I(RIOB33_X105Y151_IOB_X1Y151_IPAD),
.O(RIOB33_X105Y151_IOB_X1Y151_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y151_IOB_X1Y152_IBUF (
.I(RIOB33_X105Y151_IOB_X1Y152_IPAD),
.O(RIOB33_X105Y151_IOB_X1Y152_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y153_IOB_X1Y153_IBUF (
.I(RIOB33_X105Y153_IOB_X1Y153_IPAD),
.O(RIOB33_X105Y153_IOB_X1Y153_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y153_IOB_X1Y154_IBUF (
.I(RIOB33_X105Y153_IOB_X1Y154_IPAD),
.O(RIOB33_X105Y153_IOB_X1Y154_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y155_IOB_X1Y155_IBUF (
.I(RIOB33_X105Y155_IOB_X1Y155_IPAD),
.O(RIOB33_X105Y155_IOB_X1Y155_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y155_IOB_X1Y156_IBUF (
.I(RIOB33_X105Y155_IOB_X1Y156_IPAD),
.O(RIOB33_X105Y155_IOB_X1Y156_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y157_IOB_X1Y157_IBUF (
.I(RIOB33_X105Y157_IOB_X1Y157_IPAD),
.O(RIOB33_X105Y157_IOB_X1Y157_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y157_IOB_X1Y158_IBUF (
.I(RIOB33_X105Y157_IOB_X1Y158_IPAD),
.O(RIOB33_X105Y157_IOB_X1Y158_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y159_IOB_X1Y159_IBUF (
.I(RIOB33_X105Y159_IOB_X1Y159_IPAD),
.O(RIOB33_X105Y159_IOB_X1Y159_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y159_IOB_X1Y160_IBUF (
.I(RIOB33_X105Y159_IOB_X1Y160_IPAD),
.O(RIOB33_X105Y159_IOB_X1Y160_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y161_IOB_X1Y161_IBUF (
.I(RIOB33_X105Y161_IOB_X1Y161_IPAD),
.O(RIOB33_X105Y161_IOB_X1Y161_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y161_IOB_X1Y162_IBUF (
.I(RIOB33_X105Y161_IOB_X1Y162_IPAD),
.O(RIOB33_X105Y161_IOB_X1Y162_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y163_IOB_X1Y163_IBUF (
.I(RIOB33_X105Y163_IOB_X1Y163_IPAD),
.O(RIOB33_X105Y163_IOB_X1Y163_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y163_IOB_X1Y164_IBUF (
.I(RIOB33_X105Y163_IOB_X1Y164_IPAD),
.O(RIOB33_X105Y163_IOB_X1Y164_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y165_IOB_X1Y165_IBUF (
.I(RIOB33_X105Y165_IOB_X1Y165_IPAD),
.O(RIOB33_X105Y165_IOB_X1Y165_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y165_IOB_X1Y166_IBUF (
.I(RIOB33_X105Y165_IOB_X1Y166_IPAD),
.O(RIOB33_X105Y165_IOB_X1Y166_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y167_IOB_X1Y167_IBUF (
.I(RIOB33_X105Y167_IOB_X1Y167_IPAD),
.O(RIOB33_X105Y167_IOB_X1Y167_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y167_IOB_X1Y168_IBUF (
.I(RIOB33_X105Y167_IOB_X1Y168_IPAD),
.O(RIOB33_X105Y167_IOB_X1Y168_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y169_IOB_X1Y169_IBUF (
.I(RIOB33_X105Y169_IOB_X1Y169_IPAD),
.O(RIOB33_X105Y169_IOB_X1Y169_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y169_IOB_X1Y170_IBUF (
.I(RIOB33_X105Y169_IOB_X1Y170_IPAD),
.O(RIOB33_X105Y169_IOB_X1Y170_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y171_IOB_X1Y171_IBUF (
.I(RIOB33_X105Y171_IOB_X1Y171_IPAD),
.O(RIOB33_X105Y171_IOB_X1Y171_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y171_IOB_X1Y172_IBUF (
.I(RIOB33_X105Y171_IOB_X1Y172_IPAD),
.O(RIOB33_X105Y171_IOB_X1Y172_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y173_IOB_X1Y173_OBUF (
.I(CLBLM_R_X103Y147_SLICE_X163Y147_AO5),
.O(RIOB33_X105Y173_IOB_X1Y173_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y173_IOB_X1Y174_OBUF (
.I(LIOB33_X0Y133_IOB_X0Y133_I),
.O(RIOB33_X105Y173_IOB_X1Y174_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y175_IOB_X1Y175_OBUF (
.I(LIOB33_X0Y103_IOB_X0Y104_I),
.O(RIOB33_X105Y175_IOB_X1Y175_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y175_IOB_X1Y176_OBUF (
.I(LIOB33_X0Y137_IOB_X0Y138_I),
.O(RIOB33_X105Y175_IOB_X1Y176_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y177_IOB_X1Y177_OBUF (
.I(LIOB33_X0Y137_IOB_X0Y137_I),
.O(RIOB33_X105Y177_IOB_X1Y177_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y177_IOB_X1Y178_OBUF (
.I(CLBLM_R_X103Y177_SLICE_X163Y177_AO6),
.O(RIOB33_X105Y177_IOB_X1Y178_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y179_IOB_X1Y179_OBUF (
.I(CLBLM_R_X103Y147_SLICE_X163Y147_AO6),
.O(RIOB33_X105Y179_IOB_X1Y179_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y179_IOB_X1Y180_OBUF (
.I(CLBLL_L_X2Y146_SLICE_X1Y146_AO5),
.O(RIOB33_X105Y179_IOB_X1Y180_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y181_IOB_X1Y181_OBUF (
.I(CLBLL_L_X2Y136_SLICE_X0Y136_BO6),
.O(RIOB33_X105Y181_IOB_X1Y181_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y181_IOB_X1Y182_OBUF (
.I(RIOB33_X105Y103_IOB_X1Y104_I),
.O(RIOB33_X105Y181_IOB_X1Y182_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y183_IOB_X1Y183_OBUF (
.I(RIOB33_X105Y107_IOB_X1Y107_I),
.O(RIOB33_X105Y183_IOB_X1Y183_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y183_IOB_X1Y184_OBUF (
.I(RIOB33_SING_X105Y150_IOB_X1Y150_I),
.O(RIOB33_X105Y183_IOB_X1Y184_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y185_IOB_X1Y185_OBUF (
.I(LIOB33_X0Y133_IOB_X0Y134_I),
.O(RIOB33_X105Y185_IOB_X1Y185_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y185_IOB_X1Y186_OBUF (
.I(LIOB33_X0Y85_IOB_X0Y85_I),
.O(RIOB33_X105Y185_IOB_X1Y186_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y187_IOB_X1Y187_OBUF (
.I(CLBLM_R_X103Y185_SLICE_X163Y185_AO6),
.O(RIOB33_X105Y187_IOB_X1Y187_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y187_IOB_X1Y188_OBUF (
.I(CLBLL_L_X2Y146_SLICE_X1Y146_AO6),
.O(RIOB33_X105Y187_IOB_X1Y188_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y189_IOB_X1Y189_OBUF (
.I(CLBLL_L_X2Y173_SLICE_X1Y173_AO5),
.O(RIOB33_X105Y189_IOB_X1Y189_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y189_IOB_X1Y190_OBUF (
.I(CLBLM_R_X103Y177_SLICE_X163Y177_AO5),
.O(RIOB33_X105Y189_IOB_X1Y190_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y191_IOB_X1Y191_OBUF (
.I(CLBLM_R_X103Y177_SLICE_X163Y177_AO5),
.O(RIOB33_X105Y191_IOB_X1Y191_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y191_IOB_X1Y192_OBUF (
.I(CLBLM_R_X103Y177_SLICE_X163Y177_AO5),
.O(RIOB33_X105Y191_IOB_X1Y192_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y193_IOB_X1Y193_OBUF (
.I(CLBLM_R_X103Y177_SLICE_X163Y177_AO5),
.O(RIOB33_X105Y193_IOB_X1Y193_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y193_IOB_X1Y194_OBUF (
.I(CLBLM_R_X103Y193_SLICE_X163Y193_AO6),
.O(RIOB33_X105Y193_IOB_X1Y194_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y195_IOB_X1Y195_OBUF (
.I(LIOB33_X0Y85_IOB_X0Y85_I),
.O(RIOB33_X105Y195_IOB_X1Y195_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y195_IOB_X1Y196_OBUF (
.I(CLBLL_L_X2Y173_SLICE_X0Y173_AO6),
.O(RIOB33_X105Y195_IOB_X1Y196_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y197_IOB_X1Y197_OBUF (
.I(CLBLL_L_X2Y173_SLICE_X1Y173_AO6),
.O(RIOB33_X105Y197_IOB_X1Y197_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y197_IOB_X1Y198_OBUF (
.I(CLBLL_L_X2Y173_SLICE_X1Y173_AO6),
.O(RIOB33_X105Y197_IOB_X1Y198_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_SING_X105Y50_IOB_X1Y50_OBUF (
.I(CLBLM_R_X49Y95_SLICE_X74Y95_AO6),
.O(RIOB33_SING_X105Y50_IOB_X1Y50_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_SING_X105Y99_IOB_X1Y99_OBUF (
.I(CLBLM_R_X101Y119_SLICE_X158Y119_BO6),
.O(RIOB33_SING_X105Y99_IOB_X1Y99_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_SING_X105Y100_IOB_X1Y100_IBUF (
.I(RIOB33_SING_X105Y100_IOB_X1Y100_IPAD),
.O(RIOB33_SING_X105Y100_IOB_X1Y100_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_SING_X105Y149_IOB_X1Y149_OBUF (
.I(CLBLL_L_X4Y110_SLICE_X4Y110_CO6),
.O(RIOB33_SING_X105Y149_IOB_X1Y149_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_SING_X105Y150_IOB_X1Y150_IBUF (
.I(RIOB33_SING_X105Y150_IOB_X1Y150_IPAD),
.O(RIOB33_SING_X105Y150_IOB_X1Y150_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_SING_X105Y199_IOB_X1Y199_OBUF (
.I(CLBLL_L_X2Y173_SLICE_X1Y173_BO5),
.O(RIOB33_SING_X105Y199_IOB_X1Y199_OPAD)
  );
  assign CLBLL_L_X2Y98_SLICE_X0Y98_A = CLBLL_L_X2Y98_SLICE_X0Y98_AO6;
  assign CLBLL_L_X2Y98_SLICE_X0Y98_B = CLBLL_L_X2Y98_SLICE_X0Y98_BO6;
  assign CLBLL_L_X2Y98_SLICE_X0Y98_C = CLBLL_L_X2Y98_SLICE_X0Y98_CO6;
  assign CLBLL_L_X2Y98_SLICE_X0Y98_D = CLBLL_L_X2Y98_SLICE_X0Y98_DO6;
  assign CLBLL_L_X2Y98_SLICE_X1Y98_A = CLBLL_L_X2Y98_SLICE_X1Y98_AO6;
  assign CLBLL_L_X2Y98_SLICE_X1Y98_B = CLBLL_L_X2Y98_SLICE_X1Y98_BO6;
  assign CLBLL_L_X2Y98_SLICE_X1Y98_C = CLBLL_L_X2Y98_SLICE_X1Y98_CO6;
  assign CLBLL_L_X2Y98_SLICE_X1Y98_D = CLBLL_L_X2Y98_SLICE_X1Y98_DO6;
  assign CLBLL_L_X2Y102_SLICE_X0Y102_A = CLBLL_L_X2Y102_SLICE_X0Y102_AO6;
  assign CLBLL_L_X2Y102_SLICE_X0Y102_B = CLBLL_L_X2Y102_SLICE_X0Y102_BO6;
  assign CLBLL_L_X2Y102_SLICE_X0Y102_C = CLBLL_L_X2Y102_SLICE_X0Y102_CO6;
  assign CLBLL_L_X2Y102_SLICE_X0Y102_D = CLBLL_L_X2Y102_SLICE_X0Y102_DO6;
  assign CLBLL_L_X2Y102_SLICE_X1Y102_A = CLBLL_L_X2Y102_SLICE_X1Y102_AO6;
  assign CLBLL_L_X2Y102_SLICE_X1Y102_B = CLBLL_L_X2Y102_SLICE_X1Y102_BO6;
  assign CLBLL_L_X2Y102_SLICE_X1Y102_C = CLBLL_L_X2Y102_SLICE_X1Y102_CO6;
  assign CLBLL_L_X2Y102_SLICE_X1Y102_D = CLBLL_L_X2Y102_SLICE_X1Y102_DO6;
  assign CLBLL_L_X2Y136_SLICE_X0Y136_A = CLBLL_L_X2Y136_SLICE_X0Y136_AO6;
  assign CLBLL_L_X2Y136_SLICE_X0Y136_B = CLBLL_L_X2Y136_SLICE_X0Y136_BO6;
  assign CLBLL_L_X2Y136_SLICE_X0Y136_C = CLBLL_L_X2Y136_SLICE_X0Y136_CO6;
  assign CLBLL_L_X2Y136_SLICE_X0Y136_D = CLBLL_L_X2Y136_SLICE_X0Y136_DO6;
  assign CLBLL_L_X2Y136_SLICE_X1Y136_A = CLBLL_L_X2Y136_SLICE_X1Y136_AO6;
  assign CLBLL_L_X2Y136_SLICE_X1Y136_B = CLBLL_L_X2Y136_SLICE_X1Y136_BO6;
  assign CLBLL_L_X2Y136_SLICE_X1Y136_C = CLBLL_L_X2Y136_SLICE_X1Y136_CO6;
  assign CLBLL_L_X2Y136_SLICE_X1Y136_D = CLBLL_L_X2Y136_SLICE_X1Y136_DO6;
  assign CLBLL_L_X2Y146_SLICE_X0Y146_A = CLBLL_L_X2Y146_SLICE_X0Y146_AO6;
  assign CLBLL_L_X2Y146_SLICE_X0Y146_B = CLBLL_L_X2Y146_SLICE_X0Y146_BO6;
  assign CLBLL_L_X2Y146_SLICE_X0Y146_C = CLBLL_L_X2Y146_SLICE_X0Y146_CO6;
  assign CLBLL_L_X2Y146_SLICE_X0Y146_D = CLBLL_L_X2Y146_SLICE_X0Y146_DO6;
  assign CLBLL_L_X2Y146_SLICE_X1Y146_A = CLBLL_L_X2Y146_SLICE_X1Y146_AO6;
  assign CLBLL_L_X2Y146_SLICE_X1Y146_B = CLBLL_L_X2Y146_SLICE_X1Y146_BO6;
  assign CLBLL_L_X2Y146_SLICE_X1Y146_C = CLBLL_L_X2Y146_SLICE_X1Y146_CO6;
  assign CLBLL_L_X2Y146_SLICE_X1Y146_D = CLBLL_L_X2Y146_SLICE_X1Y146_DO6;
  assign CLBLL_L_X2Y146_SLICE_X1Y146_AMUX = CLBLL_L_X2Y146_SLICE_X1Y146_AO5;
  assign CLBLL_L_X2Y173_SLICE_X0Y173_A = CLBLL_L_X2Y173_SLICE_X0Y173_AO6;
  assign CLBLL_L_X2Y173_SLICE_X0Y173_B = CLBLL_L_X2Y173_SLICE_X0Y173_BO6;
  assign CLBLL_L_X2Y173_SLICE_X0Y173_C = CLBLL_L_X2Y173_SLICE_X0Y173_CO6;
  assign CLBLL_L_X2Y173_SLICE_X0Y173_D = CLBLL_L_X2Y173_SLICE_X0Y173_DO6;
  assign CLBLL_L_X2Y173_SLICE_X1Y173_A = CLBLL_L_X2Y173_SLICE_X1Y173_AO6;
  assign CLBLL_L_X2Y173_SLICE_X1Y173_B = CLBLL_L_X2Y173_SLICE_X1Y173_BO6;
  assign CLBLL_L_X2Y173_SLICE_X1Y173_C = CLBLL_L_X2Y173_SLICE_X1Y173_CO6;
  assign CLBLL_L_X2Y173_SLICE_X1Y173_D = CLBLL_L_X2Y173_SLICE_X1Y173_DO6;
  assign CLBLL_L_X2Y173_SLICE_X1Y173_AMUX = CLBLL_L_X2Y173_SLICE_X1Y173_AO5;
  assign CLBLL_L_X2Y173_SLICE_X1Y173_BMUX = CLBLL_L_X2Y173_SLICE_X1Y173_BO5;
  assign CLBLL_L_X2Y175_SLICE_X0Y175_A = CLBLL_L_X2Y175_SLICE_X0Y175_AO6;
  assign CLBLL_L_X2Y175_SLICE_X0Y175_B = CLBLL_L_X2Y175_SLICE_X0Y175_BO6;
  assign CLBLL_L_X2Y175_SLICE_X0Y175_C = CLBLL_L_X2Y175_SLICE_X0Y175_CO6;
  assign CLBLL_L_X2Y175_SLICE_X0Y175_D = CLBLL_L_X2Y175_SLICE_X0Y175_DO6;
  assign CLBLL_L_X2Y175_SLICE_X1Y175_A = CLBLL_L_X2Y175_SLICE_X1Y175_AO6;
  assign CLBLL_L_X2Y175_SLICE_X1Y175_B = CLBLL_L_X2Y175_SLICE_X1Y175_BO6;
  assign CLBLL_L_X2Y175_SLICE_X1Y175_C = CLBLL_L_X2Y175_SLICE_X1Y175_CO6;
  assign CLBLL_L_X2Y175_SLICE_X1Y175_D = CLBLL_L_X2Y175_SLICE_X1Y175_DO6;
  assign CLBLL_L_X4Y107_SLICE_X4Y107_A = CLBLL_L_X4Y107_SLICE_X4Y107_AO6;
  assign CLBLL_L_X4Y107_SLICE_X4Y107_B = CLBLL_L_X4Y107_SLICE_X4Y107_BO6;
  assign CLBLL_L_X4Y107_SLICE_X4Y107_C = CLBLL_L_X4Y107_SLICE_X4Y107_CO6;
  assign CLBLL_L_X4Y107_SLICE_X4Y107_D = CLBLL_L_X4Y107_SLICE_X4Y107_DO6;
  assign CLBLL_L_X4Y107_SLICE_X5Y107_A = CLBLL_L_X4Y107_SLICE_X5Y107_AO6;
  assign CLBLL_L_X4Y107_SLICE_X5Y107_B = CLBLL_L_X4Y107_SLICE_X5Y107_BO6;
  assign CLBLL_L_X4Y107_SLICE_X5Y107_C = CLBLL_L_X4Y107_SLICE_X5Y107_CO6;
  assign CLBLL_L_X4Y107_SLICE_X5Y107_D = CLBLL_L_X4Y107_SLICE_X5Y107_DO6;
  assign CLBLL_L_X4Y109_SLICE_X4Y109_A = CLBLL_L_X4Y109_SLICE_X4Y109_AO6;
  assign CLBLL_L_X4Y109_SLICE_X4Y109_B = CLBLL_L_X4Y109_SLICE_X4Y109_BO6;
  assign CLBLL_L_X4Y109_SLICE_X4Y109_C = CLBLL_L_X4Y109_SLICE_X4Y109_CO6;
  assign CLBLL_L_X4Y109_SLICE_X4Y109_D = CLBLL_L_X4Y109_SLICE_X4Y109_DO6;
  assign CLBLL_L_X4Y109_SLICE_X4Y109_AMUX = CLBLL_L_X4Y109_SLICE_X4Y109_AO5;
  assign CLBLL_L_X4Y109_SLICE_X4Y109_BMUX = CLBLL_L_X4Y109_SLICE_X4Y109_BO5;
  assign CLBLL_L_X4Y109_SLICE_X5Y109_A = CLBLL_L_X4Y109_SLICE_X5Y109_AO6;
  assign CLBLL_L_X4Y109_SLICE_X5Y109_B = CLBLL_L_X4Y109_SLICE_X5Y109_BO6;
  assign CLBLL_L_X4Y109_SLICE_X5Y109_C = CLBLL_L_X4Y109_SLICE_X5Y109_CO6;
  assign CLBLL_L_X4Y109_SLICE_X5Y109_D = CLBLL_L_X4Y109_SLICE_X5Y109_DO6;
  assign CLBLL_L_X4Y110_SLICE_X4Y110_A = CLBLL_L_X4Y110_SLICE_X4Y110_AO6;
  assign CLBLL_L_X4Y110_SLICE_X4Y110_B = CLBLL_L_X4Y110_SLICE_X4Y110_BO6;
  assign CLBLL_L_X4Y110_SLICE_X4Y110_C = CLBLL_L_X4Y110_SLICE_X4Y110_CO6;
  assign CLBLL_L_X4Y110_SLICE_X4Y110_D = CLBLL_L_X4Y110_SLICE_X4Y110_DO6;
  assign CLBLL_L_X4Y110_SLICE_X4Y110_AMUX = CLBLL_L_X4Y110_SLICE_X4Y110_AO5;
  assign CLBLL_L_X4Y110_SLICE_X4Y110_BMUX = CLBLL_L_X4Y110_SLICE_X4Y110_BO5;
  assign CLBLL_L_X4Y110_SLICE_X4Y110_CMUX = CLBLL_L_X4Y110_SLICE_X4Y110_CO5;
  assign CLBLL_L_X4Y110_SLICE_X5Y110_A = CLBLL_L_X4Y110_SLICE_X5Y110_AO6;
  assign CLBLL_L_X4Y110_SLICE_X5Y110_B = CLBLL_L_X4Y110_SLICE_X5Y110_BO6;
  assign CLBLL_L_X4Y110_SLICE_X5Y110_C = CLBLL_L_X4Y110_SLICE_X5Y110_CO6;
  assign CLBLL_L_X4Y110_SLICE_X5Y110_D = CLBLL_L_X4Y110_SLICE_X5Y110_DO6;
  assign CLBLL_L_X4Y111_SLICE_X4Y111_A = CLBLL_L_X4Y111_SLICE_X4Y111_AO6;
  assign CLBLL_L_X4Y111_SLICE_X4Y111_B = CLBLL_L_X4Y111_SLICE_X4Y111_BO6;
  assign CLBLL_L_X4Y111_SLICE_X4Y111_C = CLBLL_L_X4Y111_SLICE_X4Y111_CO6;
  assign CLBLL_L_X4Y111_SLICE_X4Y111_D = CLBLL_L_X4Y111_SLICE_X4Y111_DO6;
  assign CLBLL_L_X4Y111_SLICE_X4Y111_AMUX = CLBLL_L_X4Y111_SLICE_X4Y111_AO5;
  assign CLBLL_L_X4Y111_SLICE_X4Y111_BMUX = CLBLL_L_X4Y111_SLICE_X4Y111_BO6;
  assign CLBLL_L_X4Y111_SLICE_X5Y111_A = CLBLL_L_X4Y111_SLICE_X5Y111_AO6;
  assign CLBLL_L_X4Y111_SLICE_X5Y111_B = CLBLL_L_X4Y111_SLICE_X5Y111_BO6;
  assign CLBLL_L_X4Y111_SLICE_X5Y111_C = CLBLL_L_X4Y111_SLICE_X5Y111_CO6;
  assign CLBLL_L_X4Y111_SLICE_X5Y111_D = CLBLL_L_X4Y111_SLICE_X5Y111_DO6;
  assign CLBLL_L_X4Y111_SLICE_X5Y111_AMUX = CLBLL_L_X4Y111_SLICE_X5Y111_AO5;
  assign CLBLL_L_X4Y111_SLICE_X5Y111_BMUX = CLBLL_L_X4Y111_SLICE_X5Y111_BO5;
  assign CLBLL_L_X4Y112_SLICE_X4Y112_A = CLBLL_L_X4Y112_SLICE_X4Y112_AO6;
  assign CLBLL_L_X4Y112_SLICE_X4Y112_B = CLBLL_L_X4Y112_SLICE_X4Y112_BO6;
  assign CLBLL_L_X4Y112_SLICE_X4Y112_C = CLBLL_L_X4Y112_SLICE_X4Y112_CO6;
  assign CLBLL_L_X4Y112_SLICE_X4Y112_D = CLBLL_L_X4Y112_SLICE_X4Y112_DO6;
  assign CLBLL_L_X4Y112_SLICE_X4Y112_AMUX = CLBLL_L_X4Y112_SLICE_X4Y112_AO5;
  assign CLBLL_L_X4Y112_SLICE_X5Y112_A = CLBLL_L_X4Y112_SLICE_X5Y112_AO6;
  assign CLBLL_L_X4Y112_SLICE_X5Y112_B = CLBLL_L_X4Y112_SLICE_X5Y112_BO6;
  assign CLBLL_L_X4Y112_SLICE_X5Y112_C = CLBLL_L_X4Y112_SLICE_X5Y112_CO6;
  assign CLBLL_L_X4Y112_SLICE_X5Y112_D = CLBLL_L_X4Y112_SLICE_X5Y112_DO6;
  assign CLBLL_L_X4Y112_SLICE_X5Y112_AMUX = CLBLL_L_X4Y112_SLICE_X5Y112_AO5;
  assign CLBLL_L_X4Y112_SLICE_X5Y112_BMUX = CLBLL_L_X4Y112_SLICE_X5Y112_BO6;
  assign CLBLL_L_X4Y113_SLICE_X4Y113_A = CLBLL_L_X4Y113_SLICE_X4Y113_AO6;
  assign CLBLL_L_X4Y113_SLICE_X4Y113_B = CLBLL_L_X4Y113_SLICE_X4Y113_BO6;
  assign CLBLL_L_X4Y113_SLICE_X4Y113_C = CLBLL_L_X4Y113_SLICE_X4Y113_CO6;
  assign CLBLL_L_X4Y113_SLICE_X4Y113_D = CLBLL_L_X4Y113_SLICE_X4Y113_DO6;
  assign CLBLL_L_X4Y113_SLICE_X5Y113_A = CLBLL_L_X4Y113_SLICE_X5Y113_AO6;
  assign CLBLL_L_X4Y113_SLICE_X5Y113_B = CLBLL_L_X4Y113_SLICE_X5Y113_BO6;
  assign CLBLL_L_X4Y113_SLICE_X5Y113_C = CLBLL_L_X4Y113_SLICE_X5Y113_CO6;
  assign CLBLL_L_X4Y113_SLICE_X5Y113_D = CLBLL_L_X4Y113_SLICE_X5Y113_DO6;
  assign CLBLL_L_X4Y141_SLICE_X4Y141_A = CLBLL_L_X4Y141_SLICE_X4Y141_AO6;
  assign CLBLL_L_X4Y141_SLICE_X4Y141_B = CLBLL_L_X4Y141_SLICE_X4Y141_BO6;
  assign CLBLL_L_X4Y141_SLICE_X4Y141_C = CLBLL_L_X4Y141_SLICE_X4Y141_CO6;
  assign CLBLL_L_X4Y141_SLICE_X4Y141_D = CLBLL_L_X4Y141_SLICE_X4Y141_DO6;
  assign CLBLL_L_X4Y141_SLICE_X5Y141_A = CLBLL_L_X4Y141_SLICE_X5Y141_AO6;
  assign CLBLL_L_X4Y141_SLICE_X5Y141_B = CLBLL_L_X4Y141_SLICE_X5Y141_BO6;
  assign CLBLL_L_X4Y141_SLICE_X5Y141_C = CLBLL_L_X4Y141_SLICE_X5Y141_CO6;
  assign CLBLL_L_X4Y141_SLICE_X5Y141_D = CLBLL_L_X4Y141_SLICE_X5Y141_DO6;
  assign CLBLL_L_X36Y113_SLICE_X54Y113_A = CLBLL_L_X36Y113_SLICE_X54Y113_AO6;
  assign CLBLL_L_X36Y113_SLICE_X54Y113_B = CLBLL_L_X36Y113_SLICE_X54Y113_BO6;
  assign CLBLL_L_X36Y113_SLICE_X54Y113_C = CLBLL_L_X36Y113_SLICE_X54Y113_CO6;
  assign CLBLL_L_X36Y113_SLICE_X54Y113_D = CLBLL_L_X36Y113_SLICE_X54Y113_DO6;
  assign CLBLL_L_X36Y113_SLICE_X55Y113_A = CLBLL_L_X36Y113_SLICE_X55Y113_AO6;
  assign CLBLL_L_X36Y113_SLICE_X55Y113_B = CLBLL_L_X36Y113_SLICE_X55Y113_BO6;
  assign CLBLL_L_X36Y113_SLICE_X55Y113_C = CLBLL_L_X36Y113_SLICE_X55Y113_CO6;
  assign CLBLL_L_X36Y113_SLICE_X55Y113_D = CLBLL_L_X36Y113_SLICE_X55Y113_DO6;
  assign CLBLL_L_X100Y113_SLICE_X156Y113_A = CLBLL_L_X100Y113_SLICE_X156Y113_AO6;
  assign CLBLL_L_X100Y113_SLICE_X156Y113_B = CLBLL_L_X100Y113_SLICE_X156Y113_BO6;
  assign CLBLL_L_X100Y113_SLICE_X156Y113_C = CLBLL_L_X100Y113_SLICE_X156Y113_CO6;
  assign CLBLL_L_X100Y113_SLICE_X156Y113_D = CLBLL_L_X100Y113_SLICE_X156Y113_DO6;
  assign CLBLL_L_X100Y113_SLICE_X157Y113_A = CLBLL_L_X100Y113_SLICE_X157Y113_AO6;
  assign CLBLL_L_X100Y113_SLICE_X157Y113_B = CLBLL_L_X100Y113_SLICE_X157Y113_BO6;
  assign CLBLL_L_X100Y113_SLICE_X157Y113_C = CLBLL_L_X100Y113_SLICE_X157Y113_CO6;
  assign CLBLL_L_X100Y113_SLICE_X157Y113_D = CLBLL_L_X100Y113_SLICE_X157Y113_DO6;
  assign CLBLL_L_X100Y121_SLICE_X156Y121_A = CLBLL_L_X100Y121_SLICE_X156Y121_AO6;
  assign CLBLL_L_X100Y121_SLICE_X156Y121_B = CLBLL_L_X100Y121_SLICE_X156Y121_BO6;
  assign CLBLL_L_X100Y121_SLICE_X156Y121_C = CLBLL_L_X100Y121_SLICE_X156Y121_CO6;
  assign CLBLL_L_X100Y121_SLICE_X156Y121_D = CLBLL_L_X100Y121_SLICE_X156Y121_DO6;
  assign CLBLL_L_X100Y121_SLICE_X157Y121_A = CLBLL_L_X100Y121_SLICE_X157Y121_AO6;
  assign CLBLL_L_X100Y121_SLICE_X157Y121_B = CLBLL_L_X100Y121_SLICE_X157Y121_BO6;
  assign CLBLL_L_X100Y121_SLICE_X157Y121_C = CLBLL_L_X100Y121_SLICE_X157Y121_CO6;
  assign CLBLL_L_X100Y121_SLICE_X157Y121_D = CLBLL_L_X100Y121_SLICE_X157Y121_DO6;
  assign CLBLL_L_X100Y123_SLICE_X156Y123_A = CLBLL_L_X100Y123_SLICE_X156Y123_AO6;
  assign CLBLL_L_X100Y123_SLICE_X156Y123_B = CLBLL_L_X100Y123_SLICE_X156Y123_BO6;
  assign CLBLL_L_X100Y123_SLICE_X156Y123_C = CLBLL_L_X100Y123_SLICE_X156Y123_CO6;
  assign CLBLL_L_X100Y123_SLICE_X156Y123_D = CLBLL_L_X100Y123_SLICE_X156Y123_DO6;
  assign CLBLL_L_X100Y123_SLICE_X156Y123_AMUX = CLBLL_L_X100Y123_SLICE_X156Y123_AO5;
  assign CLBLL_L_X100Y123_SLICE_X156Y123_BMUX = CLBLL_L_X100Y123_SLICE_X156Y123_BO5;
  assign CLBLL_L_X100Y123_SLICE_X157Y123_A = CLBLL_L_X100Y123_SLICE_X157Y123_AO6;
  assign CLBLL_L_X100Y123_SLICE_X157Y123_B = CLBLL_L_X100Y123_SLICE_X157Y123_BO6;
  assign CLBLL_L_X100Y123_SLICE_X157Y123_C = CLBLL_L_X100Y123_SLICE_X157Y123_CO6;
  assign CLBLL_L_X100Y123_SLICE_X157Y123_D = CLBLL_L_X100Y123_SLICE_X157Y123_DO6;
  assign CLBLL_R_X57Y113_SLICE_X86Y113_A = CLBLL_R_X57Y113_SLICE_X86Y113_AO6;
  assign CLBLL_R_X57Y113_SLICE_X86Y113_B = CLBLL_R_X57Y113_SLICE_X86Y113_BO6;
  assign CLBLL_R_X57Y113_SLICE_X86Y113_C = CLBLL_R_X57Y113_SLICE_X86Y113_CO6;
  assign CLBLL_R_X57Y113_SLICE_X86Y113_D = CLBLL_R_X57Y113_SLICE_X86Y113_DO6;
  assign CLBLL_R_X57Y113_SLICE_X87Y113_A = CLBLL_R_X57Y113_SLICE_X87Y113_AO6;
  assign CLBLL_R_X57Y113_SLICE_X87Y113_B = CLBLL_R_X57Y113_SLICE_X87Y113_BO6;
  assign CLBLL_R_X57Y113_SLICE_X87Y113_C = CLBLL_R_X57Y113_SLICE_X87Y113_CO6;
  assign CLBLL_R_X57Y113_SLICE_X87Y113_D = CLBLL_R_X57Y113_SLICE_X87Y113_DO6;
  assign CLBLM_L_X8Y113_SLICE_X10Y113_A = CLBLM_L_X8Y113_SLICE_X10Y113_AO6;
  assign CLBLM_L_X8Y113_SLICE_X10Y113_B = CLBLM_L_X8Y113_SLICE_X10Y113_BO6;
  assign CLBLM_L_X8Y113_SLICE_X10Y113_C = CLBLM_L_X8Y113_SLICE_X10Y113_CO6;
  assign CLBLM_L_X8Y113_SLICE_X10Y113_D = CLBLM_L_X8Y113_SLICE_X10Y113_DO6;
  assign CLBLM_L_X8Y113_SLICE_X10Y113_AMUX = CLBLM_L_X8Y113_SLICE_X10Y113_AO5;
  assign CLBLM_L_X8Y113_SLICE_X11Y113_A = CLBLM_L_X8Y113_SLICE_X11Y113_AO6;
  assign CLBLM_L_X8Y113_SLICE_X11Y113_B = CLBLM_L_X8Y113_SLICE_X11Y113_BO6;
  assign CLBLM_L_X8Y113_SLICE_X11Y113_C = CLBLM_L_X8Y113_SLICE_X11Y113_CO6;
  assign CLBLM_L_X8Y113_SLICE_X11Y113_D = CLBLM_L_X8Y113_SLICE_X11Y113_DO6;
  assign CLBLM_L_X8Y113_SLICE_X11Y113_AMUX = CLBLM_L_X8Y113_SLICE_X11Y113_AO5;
  assign CLBLM_L_X10Y113_SLICE_X12Y113_A = CLBLM_L_X10Y113_SLICE_X12Y113_AO6;
  assign CLBLM_L_X10Y113_SLICE_X12Y113_B = CLBLM_L_X10Y113_SLICE_X12Y113_BO6;
  assign CLBLM_L_X10Y113_SLICE_X12Y113_C = CLBLM_L_X10Y113_SLICE_X12Y113_CO6;
  assign CLBLM_L_X10Y113_SLICE_X12Y113_D = CLBLM_L_X10Y113_SLICE_X12Y113_DO6;
  assign CLBLM_L_X10Y113_SLICE_X13Y113_A = CLBLM_L_X10Y113_SLICE_X13Y113_AO6;
  assign CLBLM_L_X10Y113_SLICE_X13Y113_B = CLBLM_L_X10Y113_SLICE_X13Y113_BO6;
  assign CLBLM_L_X10Y113_SLICE_X13Y113_C = CLBLM_L_X10Y113_SLICE_X13Y113_CO6;
  assign CLBLM_L_X10Y113_SLICE_X13Y113_D = CLBLM_L_X10Y113_SLICE_X13Y113_DO6;
  assign CLBLM_L_X10Y114_SLICE_X12Y114_A = CLBLM_L_X10Y114_SLICE_X12Y114_AO6;
  assign CLBLM_L_X10Y114_SLICE_X12Y114_B = CLBLM_L_X10Y114_SLICE_X12Y114_BO6;
  assign CLBLM_L_X10Y114_SLICE_X12Y114_C = CLBLM_L_X10Y114_SLICE_X12Y114_CO6;
  assign CLBLM_L_X10Y114_SLICE_X12Y114_D = CLBLM_L_X10Y114_SLICE_X12Y114_DO6;
  assign CLBLM_L_X10Y114_SLICE_X13Y114_A = CLBLM_L_X10Y114_SLICE_X13Y114_AO6;
  assign CLBLM_L_X10Y114_SLICE_X13Y114_B = CLBLM_L_X10Y114_SLICE_X13Y114_BO6;
  assign CLBLM_L_X10Y114_SLICE_X13Y114_C = CLBLM_L_X10Y114_SLICE_X13Y114_CO6;
  assign CLBLM_L_X10Y114_SLICE_X13Y114_D = CLBLM_L_X10Y114_SLICE_X13Y114_DO6;
  assign CLBLM_L_X10Y123_SLICE_X12Y123_A = CLBLM_L_X10Y123_SLICE_X12Y123_AO6;
  assign CLBLM_L_X10Y123_SLICE_X12Y123_B = CLBLM_L_X10Y123_SLICE_X12Y123_BO6;
  assign CLBLM_L_X10Y123_SLICE_X12Y123_C = CLBLM_L_X10Y123_SLICE_X12Y123_CO6;
  assign CLBLM_L_X10Y123_SLICE_X12Y123_D = CLBLM_L_X10Y123_SLICE_X12Y123_DO6;
  assign CLBLM_L_X10Y123_SLICE_X13Y123_A = CLBLM_L_X10Y123_SLICE_X13Y123_AO6;
  assign CLBLM_L_X10Y123_SLICE_X13Y123_B = CLBLM_L_X10Y123_SLICE_X13Y123_BO6;
  assign CLBLM_L_X10Y123_SLICE_X13Y123_C = CLBLM_L_X10Y123_SLICE_X13Y123_CO6;
  assign CLBLM_L_X10Y123_SLICE_X13Y123_D = CLBLM_L_X10Y123_SLICE_X13Y123_DO6;
  assign CLBLM_L_X56Y119_SLICE_X84Y119_A = CLBLM_L_X56Y119_SLICE_X84Y119_AO6;
  assign CLBLM_L_X56Y119_SLICE_X84Y119_B = CLBLM_L_X56Y119_SLICE_X84Y119_BO6;
  assign CLBLM_L_X56Y119_SLICE_X84Y119_C = CLBLM_L_X56Y119_SLICE_X84Y119_CO6;
  assign CLBLM_L_X56Y119_SLICE_X84Y119_D = CLBLM_L_X56Y119_SLICE_X84Y119_DO6;
  assign CLBLM_L_X56Y119_SLICE_X84Y119_AMUX = CLBLM_L_X56Y119_SLICE_X84Y119_AO5;
  assign CLBLM_L_X56Y119_SLICE_X85Y119_A = CLBLM_L_X56Y119_SLICE_X85Y119_AO6;
  assign CLBLM_L_X56Y119_SLICE_X85Y119_B = CLBLM_L_X56Y119_SLICE_X85Y119_BO6;
  assign CLBLM_L_X56Y119_SLICE_X85Y119_C = CLBLM_L_X56Y119_SLICE_X85Y119_CO6;
  assign CLBLM_L_X56Y119_SLICE_X85Y119_D = CLBLM_L_X56Y119_SLICE_X85Y119_DO6;
  assign CLBLM_R_X3Y110_SLICE_X2Y110_A = CLBLM_R_X3Y110_SLICE_X2Y110_AO6;
  assign CLBLM_R_X3Y110_SLICE_X2Y110_B = CLBLM_R_X3Y110_SLICE_X2Y110_BO6;
  assign CLBLM_R_X3Y110_SLICE_X2Y110_C = CLBLM_R_X3Y110_SLICE_X2Y110_CO6;
  assign CLBLM_R_X3Y110_SLICE_X2Y110_D = CLBLM_R_X3Y110_SLICE_X2Y110_DO6;
  assign CLBLM_R_X3Y110_SLICE_X3Y110_A = CLBLM_R_X3Y110_SLICE_X3Y110_AO6;
  assign CLBLM_R_X3Y110_SLICE_X3Y110_B = CLBLM_R_X3Y110_SLICE_X3Y110_BO6;
  assign CLBLM_R_X3Y110_SLICE_X3Y110_C = CLBLM_R_X3Y110_SLICE_X3Y110_CO6;
  assign CLBLM_R_X3Y110_SLICE_X3Y110_D = CLBLM_R_X3Y110_SLICE_X3Y110_DO6;
  assign CLBLM_R_X3Y110_SLICE_X3Y110_AMUX = CLBLM_R_X3Y110_SLICE_X3Y110_AO5;
  assign CLBLM_R_X3Y111_SLICE_X2Y111_A = CLBLM_R_X3Y111_SLICE_X2Y111_AO6;
  assign CLBLM_R_X3Y111_SLICE_X2Y111_B = CLBLM_R_X3Y111_SLICE_X2Y111_BO6;
  assign CLBLM_R_X3Y111_SLICE_X2Y111_C = CLBLM_R_X3Y111_SLICE_X2Y111_CO6;
  assign CLBLM_R_X3Y111_SLICE_X2Y111_D = CLBLM_R_X3Y111_SLICE_X2Y111_DO6;
  assign CLBLM_R_X3Y111_SLICE_X2Y111_AMUX = CLBLM_R_X3Y111_SLICE_X2Y111_AO5;
  assign CLBLM_R_X3Y111_SLICE_X3Y111_A = CLBLM_R_X3Y111_SLICE_X3Y111_AO6;
  assign CLBLM_R_X3Y111_SLICE_X3Y111_B = CLBLM_R_X3Y111_SLICE_X3Y111_BO6;
  assign CLBLM_R_X3Y111_SLICE_X3Y111_C = CLBLM_R_X3Y111_SLICE_X3Y111_CO6;
  assign CLBLM_R_X3Y111_SLICE_X3Y111_D = CLBLM_R_X3Y111_SLICE_X3Y111_DO6;
  assign CLBLM_R_X3Y111_SLICE_X3Y111_AMUX = CLBLM_R_X3Y111_SLICE_X3Y111_AO5;
  assign CLBLM_R_X3Y111_SLICE_X3Y111_BMUX = CLBLM_R_X3Y111_SLICE_X3Y111_BO5;
  assign CLBLM_R_X3Y111_SLICE_X3Y111_CMUX = CLBLM_R_X3Y111_SLICE_X3Y111_CO5;
  assign CLBLM_R_X3Y111_SLICE_X3Y111_DMUX = CLBLM_R_X3Y111_SLICE_X3Y111_DO6;
  assign CLBLM_R_X3Y112_SLICE_X2Y112_A = CLBLM_R_X3Y112_SLICE_X2Y112_AO6;
  assign CLBLM_R_X3Y112_SLICE_X2Y112_B = CLBLM_R_X3Y112_SLICE_X2Y112_BO6;
  assign CLBLM_R_X3Y112_SLICE_X2Y112_C = CLBLM_R_X3Y112_SLICE_X2Y112_CO6;
  assign CLBLM_R_X3Y112_SLICE_X2Y112_D = CLBLM_R_X3Y112_SLICE_X2Y112_DO6;
  assign CLBLM_R_X3Y112_SLICE_X3Y112_A = CLBLM_R_X3Y112_SLICE_X3Y112_AO6;
  assign CLBLM_R_X3Y112_SLICE_X3Y112_B = CLBLM_R_X3Y112_SLICE_X3Y112_BO6;
  assign CLBLM_R_X3Y112_SLICE_X3Y112_C = CLBLM_R_X3Y112_SLICE_X3Y112_CO6;
  assign CLBLM_R_X3Y112_SLICE_X3Y112_D = CLBLM_R_X3Y112_SLICE_X3Y112_DO6;
  assign CLBLM_R_X3Y112_SLICE_X3Y112_AMUX = CLBLM_R_X3Y112_SLICE_X3Y112_AO5;
  assign CLBLM_R_X5Y109_SLICE_X6Y109_A = CLBLM_R_X5Y109_SLICE_X6Y109_AO6;
  assign CLBLM_R_X5Y109_SLICE_X6Y109_B = CLBLM_R_X5Y109_SLICE_X6Y109_BO6;
  assign CLBLM_R_X5Y109_SLICE_X6Y109_C = CLBLM_R_X5Y109_SLICE_X6Y109_CO6;
  assign CLBLM_R_X5Y109_SLICE_X6Y109_D = CLBLM_R_X5Y109_SLICE_X6Y109_DO6;
  assign CLBLM_R_X5Y109_SLICE_X7Y109_A = CLBLM_R_X5Y109_SLICE_X7Y109_AO6;
  assign CLBLM_R_X5Y109_SLICE_X7Y109_B = CLBLM_R_X5Y109_SLICE_X7Y109_BO6;
  assign CLBLM_R_X5Y109_SLICE_X7Y109_C = CLBLM_R_X5Y109_SLICE_X7Y109_CO6;
  assign CLBLM_R_X5Y109_SLICE_X7Y109_D = CLBLM_R_X5Y109_SLICE_X7Y109_DO6;
  assign CLBLM_R_X5Y110_SLICE_X6Y110_A = CLBLM_R_X5Y110_SLICE_X6Y110_AO6;
  assign CLBLM_R_X5Y110_SLICE_X6Y110_B = CLBLM_R_X5Y110_SLICE_X6Y110_BO6;
  assign CLBLM_R_X5Y110_SLICE_X6Y110_C = CLBLM_R_X5Y110_SLICE_X6Y110_CO6;
  assign CLBLM_R_X5Y110_SLICE_X6Y110_D = CLBLM_R_X5Y110_SLICE_X6Y110_DO6;
  assign CLBLM_R_X5Y110_SLICE_X6Y110_AMUX = CLBLM_R_X5Y110_SLICE_X6Y110_AO5;
  assign CLBLM_R_X5Y110_SLICE_X7Y110_A = CLBLM_R_X5Y110_SLICE_X7Y110_AO6;
  assign CLBLM_R_X5Y110_SLICE_X7Y110_B = CLBLM_R_X5Y110_SLICE_X7Y110_BO6;
  assign CLBLM_R_X5Y110_SLICE_X7Y110_C = CLBLM_R_X5Y110_SLICE_X7Y110_CO6;
  assign CLBLM_R_X5Y110_SLICE_X7Y110_D = CLBLM_R_X5Y110_SLICE_X7Y110_DO6;
  assign CLBLM_R_X5Y111_SLICE_X6Y111_A = CLBLM_R_X5Y111_SLICE_X6Y111_AO6;
  assign CLBLM_R_X5Y111_SLICE_X6Y111_B = CLBLM_R_X5Y111_SLICE_X6Y111_BO6;
  assign CLBLM_R_X5Y111_SLICE_X6Y111_C = CLBLM_R_X5Y111_SLICE_X6Y111_CO6;
  assign CLBLM_R_X5Y111_SLICE_X6Y111_D = CLBLM_R_X5Y111_SLICE_X6Y111_DO6;
  assign CLBLM_R_X5Y111_SLICE_X6Y111_AMUX = CLBLM_R_X5Y111_SLICE_X6Y111_AO5;
  assign CLBLM_R_X5Y111_SLICE_X7Y111_A = CLBLM_R_X5Y111_SLICE_X7Y111_AO6;
  assign CLBLM_R_X5Y111_SLICE_X7Y111_B = CLBLM_R_X5Y111_SLICE_X7Y111_BO6;
  assign CLBLM_R_X5Y111_SLICE_X7Y111_C = CLBLM_R_X5Y111_SLICE_X7Y111_CO6;
  assign CLBLM_R_X5Y111_SLICE_X7Y111_D = CLBLM_R_X5Y111_SLICE_X7Y111_DO6;
  assign CLBLM_R_X5Y111_SLICE_X7Y111_AMUX = CLBLM_R_X5Y111_SLICE_X7Y111_AO5;
  assign CLBLM_R_X5Y112_SLICE_X6Y112_A = CLBLM_R_X5Y112_SLICE_X6Y112_AO6;
  assign CLBLM_R_X5Y112_SLICE_X6Y112_B = CLBLM_R_X5Y112_SLICE_X6Y112_BO6;
  assign CLBLM_R_X5Y112_SLICE_X6Y112_C = CLBLM_R_X5Y112_SLICE_X6Y112_CO6;
  assign CLBLM_R_X5Y112_SLICE_X6Y112_D = CLBLM_R_X5Y112_SLICE_X6Y112_DO6;
  assign CLBLM_R_X5Y112_SLICE_X7Y112_A = CLBLM_R_X5Y112_SLICE_X7Y112_AO6;
  assign CLBLM_R_X5Y112_SLICE_X7Y112_B = CLBLM_R_X5Y112_SLICE_X7Y112_BO6;
  assign CLBLM_R_X5Y112_SLICE_X7Y112_C = CLBLM_R_X5Y112_SLICE_X7Y112_CO6;
  assign CLBLM_R_X5Y112_SLICE_X7Y112_D = CLBLM_R_X5Y112_SLICE_X7Y112_DO6;
  assign CLBLM_R_X5Y112_SLICE_X7Y112_AMUX = CLBLM_R_X5Y112_SLICE_X7Y112_AO5;
  assign CLBLM_R_X5Y113_SLICE_X6Y113_A = CLBLM_R_X5Y113_SLICE_X6Y113_AO6;
  assign CLBLM_R_X5Y113_SLICE_X6Y113_B = CLBLM_R_X5Y113_SLICE_X6Y113_BO6;
  assign CLBLM_R_X5Y113_SLICE_X6Y113_C = CLBLM_R_X5Y113_SLICE_X6Y113_CO6;
  assign CLBLM_R_X5Y113_SLICE_X6Y113_D = CLBLM_R_X5Y113_SLICE_X6Y113_DO6;
  assign CLBLM_R_X5Y113_SLICE_X6Y113_AMUX = CLBLM_R_X5Y113_SLICE_X6Y113_AO5;
  assign CLBLM_R_X5Y113_SLICE_X7Y113_A = CLBLM_R_X5Y113_SLICE_X7Y113_AO6;
  assign CLBLM_R_X5Y113_SLICE_X7Y113_B = CLBLM_R_X5Y113_SLICE_X7Y113_BO6;
  assign CLBLM_R_X5Y113_SLICE_X7Y113_C = CLBLM_R_X5Y113_SLICE_X7Y113_CO6;
  assign CLBLM_R_X5Y113_SLICE_X7Y113_D = CLBLM_R_X5Y113_SLICE_X7Y113_DO6;
  assign CLBLM_R_X5Y114_SLICE_X6Y114_A = CLBLM_R_X5Y114_SLICE_X6Y114_AO6;
  assign CLBLM_R_X5Y114_SLICE_X6Y114_B = CLBLM_R_X5Y114_SLICE_X6Y114_BO6;
  assign CLBLM_R_X5Y114_SLICE_X6Y114_C = CLBLM_R_X5Y114_SLICE_X6Y114_CO6;
  assign CLBLM_R_X5Y114_SLICE_X6Y114_D = CLBLM_R_X5Y114_SLICE_X6Y114_DO6;
  assign CLBLM_R_X5Y114_SLICE_X7Y114_A = CLBLM_R_X5Y114_SLICE_X7Y114_AO6;
  assign CLBLM_R_X5Y114_SLICE_X7Y114_B = CLBLM_R_X5Y114_SLICE_X7Y114_BO6;
  assign CLBLM_R_X5Y114_SLICE_X7Y114_C = CLBLM_R_X5Y114_SLICE_X7Y114_CO6;
  assign CLBLM_R_X5Y114_SLICE_X7Y114_D = CLBLM_R_X5Y114_SLICE_X7Y114_DO6;
  assign CLBLM_R_X5Y114_SLICE_X7Y114_AMUX = CLBLM_R_X5Y114_SLICE_X7Y114_AO5;
  assign CLBLM_R_X5Y115_SLICE_X6Y115_A = CLBLM_R_X5Y115_SLICE_X6Y115_AO6;
  assign CLBLM_R_X5Y115_SLICE_X6Y115_B = CLBLM_R_X5Y115_SLICE_X6Y115_BO6;
  assign CLBLM_R_X5Y115_SLICE_X6Y115_C = CLBLM_R_X5Y115_SLICE_X6Y115_CO6;
  assign CLBLM_R_X5Y115_SLICE_X6Y115_D = CLBLM_R_X5Y115_SLICE_X6Y115_DO6;
  assign CLBLM_R_X5Y115_SLICE_X6Y115_AMUX = CLBLM_R_X5Y115_SLICE_X6Y115_AO5;
  assign CLBLM_R_X5Y115_SLICE_X6Y115_BMUX = CLBLM_R_X5Y115_SLICE_X6Y115_BO5;
  assign CLBLM_R_X5Y115_SLICE_X7Y115_A = CLBLM_R_X5Y115_SLICE_X7Y115_AO6;
  assign CLBLM_R_X5Y115_SLICE_X7Y115_B = CLBLM_R_X5Y115_SLICE_X7Y115_BO6;
  assign CLBLM_R_X5Y115_SLICE_X7Y115_C = CLBLM_R_X5Y115_SLICE_X7Y115_CO6;
  assign CLBLM_R_X5Y115_SLICE_X7Y115_D = CLBLM_R_X5Y115_SLICE_X7Y115_DO6;
  assign CLBLM_R_X7Y113_SLICE_X8Y113_A = CLBLM_R_X7Y113_SLICE_X8Y113_AO6;
  assign CLBLM_R_X7Y113_SLICE_X8Y113_B = CLBLM_R_X7Y113_SLICE_X8Y113_BO6;
  assign CLBLM_R_X7Y113_SLICE_X8Y113_C = CLBLM_R_X7Y113_SLICE_X8Y113_CO6;
  assign CLBLM_R_X7Y113_SLICE_X8Y113_D = CLBLM_R_X7Y113_SLICE_X8Y113_DO6;
  assign CLBLM_R_X7Y113_SLICE_X8Y113_AMUX = CLBLM_R_X7Y113_SLICE_X8Y113_AO5;
  assign CLBLM_R_X7Y113_SLICE_X8Y113_BMUX = CLBLM_R_X7Y113_SLICE_X8Y113_BO5;
  assign CLBLM_R_X7Y113_SLICE_X9Y113_A = CLBLM_R_X7Y113_SLICE_X9Y113_AO6;
  assign CLBLM_R_X7Y113_SLICE_X9Y113_B = CLBLM_R_X7Y113_SLICE_X9Y113_BO6;
  assign CLBLM_R_X7Y113_SLICE_X9Y113_C = CLBLM_R_X7Y113_SLICE_X9Y113_CO6;
  assign CLBLM_R_X7Y113_SLICE_X9Y113_D = CLBLM_R_X7Y113_SLICE_X9Y113_DO6;
  assign CLBLM_R_X7Y114_SLICE_X8Y114_A = CLBLM_R_X7Y114_SLICE_X8Y114_AO6;
  assign CLBLM_R_X7Y114_SLICE_X8Y114_B = CLBLM_R_X7Y114_SLICE_X8Y114_BO6;
  assign CLBLM_R_X7Y114_SLICE_X8Y114_C = CLBLM_R_X7Y114_SLICE_X8Y114_CO6;
  assign CLBLM_R_X7Y114_SLICE_X8Y114_D = CLBLM_R_X7Y114_SLICE_X8Y114_DO6;
  assign CLBLM_R_X7Y114_SLICE_X8Y114_AMUX = CLBLM_R_X7Y114_SLICE_X8Y114_AO5;
  assign CLBLM_R_X7Y114_SLICE_X8Y114_BMUX = CLBLM_R_X7Y114_SLICE_X8Y114_BO5;
  assign CLBLM_R_X7Y114_SLICE_X9Y114_A = CLBLM_R_X7Y114_SLICE_X9Y114_AO6;
  assign CLBLM_R_X7Y114_SLICE_X9Y114_B = CLBLM_R_X7Y114_SLICE_X9Y114_BO6;
  assign CLBLM_R_X7Y114_SLICE_X9Y114_C = CLBLM_R_X7Y114_SLICE_X9Y114_CO6;
  assign CLBLM_R_X7Y114_SLICE_X9Y114_D = CLBLM_R_X7Y114_SLICE_X9Y114_DO6;
  assign CLBLM_R_X7Y121_SLICE_X8Y121_A = CLBLM_R_X7Y121_SLICE_X8Y121_AO6;
  assign CLBLM_R_X7Y121_SLICE_X8Y121_B = CLBLM_R_X7Y121_SLICE_X8Y121_BO6;
  assign CLBLM_R_X7Y121_SLICE_X8Y121_C = CLBLM_R_X7Y121_SLICE_X8Y121_CO6;
  assign CLBLM_R_X7Y121_SLICE_X8Y121_D = CLBLM_R_X7Y121_SLICE_X8Y121_DO6;
  assign CLBLM_R_X7Y121_SLICE_X9Y121_A = CLBLM_R_X7Y121_SLICE_X9Y121_AO6;
  assign CLBLM_R_X7Y121_SLICE_X9Y121_B = CLBLM_R_X7Y121_SLICE_X9Y121_BO6;
  assign CLBLM_R_X7Y121_SLICE_X9Y121_C = CLBLM_R_X7Y121_SLICE_X9Y121_CO6;
  assign CLBLM_R_X7Y121_SLICE_X9Y121_D = CLBLM_R_X7Y121_SLICE_X9Y121_DO6;
  assign CLBLM_R_X7Y121_SLICE_X9Y121_AMUX = CLBLM_R_X7Y121_SLICE_X9Y121_AO5;
  assign CLBLM_R_X25Y115_SLICE_X36Y115_A = CLBLM_R_X25Y115_SLICE_X36Y115_AO6;
  assign CLBLM_R_X25Y115_SLICE_X36Y115_B = CLBLM_R_X25Y115_SLICE_X36Y115_BO6;
  assign CLBLM_R_X25Y115_SLICE_X36Y115_C = CLBLM_R_X25Y115_SLICE_X36Y115_CO6;
  assign CLBLM_R_X25Y115_SLICE_X36Y115_D = CLBLM_R_X25Y115_SLICE_X36Y115_DO6;
  assign CLBLM_R_X25Y115_SLICE_X36Y115_AMUX = CLBLM_R_X25Y115_SLICE_X36Y115_AO5;
  assign CLBLM_R_X25Y115_SLICE_X37Y115_A = CLBLM_R_X25Y115_SLICE_X37Y115_AO6;
  assign CLBLM_R_X25Y115_SLICE_X37Y115_B = CLBLM_R_X25Y115_SLICE_X37Y115_BO6;
  assign CLBLM_R_X25Y115_SLICE_X37Y115_C = CLBLM_R_X25Y115_SLICE_X37Y115_CO6;
  assign CLBLM_R_X25Y115_SLICE_X37Y115_D = CLBLM_R_X25Y115_SLICE_X37Y115_DO6;
  assign CLBLM_R_X25Y116_SLICE_X36Y116_A = CLBLM_R_X25Y116_SLICE_X36Y116_AO6;
  assign CLBLM_R_X25Y116_SLICE_X36Y116_B = CLBLM_R_X25Y116_SLICE_X36Y116_BO6;
  assign CLBLM_R_X25Y116_SLICE_X36Y116_C = CLBLM_R_X25Y116_SLICE_X36Y116_CO6;
  assign CLBLM_R_X25Y116_SLICE_X36Y116_D = CLBLM_R_X25Y116_SLICE_X36Y116_DO6;
  assign CLBLM_R_X25Y116_SLICE_X36Y116_AMUX = CLBLM_R_X25Y116_SLICE_X36Y116_AO5;
  assign CLBLM_R_X25Y116_SLICE_X37Y116_A = CLBLM_R_X25Y116_SLICE_X37Y116_AO6;
  assign CLBLM_R_X25Y116_SLICE_X37Y116_B = CLBLM_R_X25Y116_SLICE_X37Y116_BO6;
  assign CLBLM_R_X25Y116_SLICE_X37Y116_C = CLBLM_R_X25Y116_SLICE_X37Y116_CO6;
  assign CLBLM_R_X25Y116_SLICE_X37Y116_D = CLBLM_R_X25Y116_SLICE_X37Y116_DO6;
  assign CLBLM_R_X29Y115_SLICE_X42Y115_A = CLBLM_R_X29Y115_SLICE_X42Y115_AO6;
  assign CLBLM_R_X29Y115_SLICE_X42Y115_B = CLBLM_R_X29Y115_SLICE_X42Y115_BO6;
  assign CLBLM_R_X29Y115_SLICE_X42Y115_C = CLBLM_R_X29Y115_SLICE_X42Y115_CO6;
  assign CLBLM_R_X29Y115_SLICE_X42Y115_D = CLBLM_R_X29Y115_SLICE_X42Y115_DO6;
  assign CLBLM_R_X29Y115_SLICE_X43Y115_A = CLBLM_R_X29Y115_SLICE_X43Y115_AO6;
  assign CLBLM_R_X29Y115_SLICE_X43Y115_B = CLBLM_R_X29Y115_SLICE_X43Y115_BO6;
  assign CLBLM_R_X29Y115_SLICE_X43Y115_C = CLBLM_R_X29Y115_SLICE_X43Y115_CO6;
  assign CLBLM_R_X29Y115_SLICE_X43Y115_D = CLBLM_R_X29Y115_SLICE_X43Y115_DO6;
  assign CLBLM_R_X49Y95_SLICE_X74Y95_A = CLBLM_R_X49Y95_SLICE_X74Y95_AO6;
  assign CLBLM_R_X49Y95_SLICE_X74Y95_B = CLBLM_R_X49Y95_SLICE_X74Y95_BO6;
  assign CLBLM_R_X49Y95_SLICE_X74Y95_C = CLBLM_R_X49Y95_SLICE_X74Y95_CO6;
  assign CLBLM_R_X49Y95_SLICE_X74Y95_D = CLBLM_R_X49Y95_SLICE_X74Y95_DO6;
  assign CLBLM_R_X49Y95_SLICE_X74Y95_AMUX = CLBLM_R_X49Y95_SLICE_X74Y95_AO5;
  assign CLBLM_R_X49Y95_SLICE_X75Y95_A = CLBLM_R_X49Y95_SLICE_X75Y95_AO6;
  assign CLBLM_R_X49Y95_SLICE_X75Y95_B = CLBLM_R_X49Y95_SLICE_X75Y95_BO6;
  assign CLBLM_R_X49Y95_SLICE_X75Y95_C = CLBLM_R_X49Y95_SLICE_X75Y95_CO6;
  assign CLBLM_R_X49Y95_SLICE_X75Y95_D = CLBLM_R_X49Y95_SLICE_X75Y95_DO6;
  assign CLBLM_R_X49Y101_SLICE_X74Y101_A = CLBLM_R_X49Y101_SLICE_X74Y101_AO6;
  assign CLBLM_R_X49Y101_SLICE_X74Y101_B = CLBLM_R_X49Y101_SLICE_X74Y101_BO6;
  assign CLBLM_R_X49Y101_SLICE_X74Y101_C = CLBLM_R_X49Y101_SLICE_X74Y101_CO6;
  assign CLBLM_R_X49Y101_SLICE_X74Y101_D = CLBLM_R_X49Y101_SLICE_X74Y101_DO6;
  assign CLBLM_R_X49Y101_SLICE_X74Y101_AMUX = CLBLM_R_X49Y101_SLICE_X74Y101_AO5;
  assign CLBLM_R_X49Y101_SLICE_X75Y101_A = CLBLM_R_X49Y101_SLICE_X75Y101_AO6;
  assign CLBLM_R_X49Y101_SLICE_X75Y101_B = CLBLM_R_X49Y101_SLICE_X75Y101_BO6;
  assign CLBLM_R_X49Y101_SLICE_X75Y101_C = CLBLM_R_X49Y101_SLICE_X75Y101_CO6;
  assign CLBLM_R_X49Y101_SLICE_X75Y101_D = CLBLM_R_X49Y101_SLICE_X75Y101_DO6;
  assign CLBLM_R_X101Y116_SLICE_X158Y116_A = CLBLM_R_X101Y116_SLICE_X158Y116_AO6;
  assign CLBLM_R_X101Y116_SLICE_X158Y116_B = CLBLM_R_X101Y116_SLICE_X158Y116_BO6;
  assign CLBLM_R_X101Y116_SLICE_X158Y116_C = CLBLM_R_X101Y116_SLICE_X158Y116_CO6;
  assign CLBLM_R_X101Y116_SLICE_X158Y116_D = CLBLM_R_X101Y116_SLICE_X158Y116_DO6;
  assign CLBLM_R_X101Y116_SLICE_X159Y116_A = CLBLM_R_X101Y116_SLICE_X159Y116_AO6;
  assign CLBLM_R_X101Y116_SLICE_X159Y116_B = CLBLM_R_X101Y116_SLICE_X159Y116_BO6;
  assign CLBLM_R_X101Y116_SLICE_X159Y116_C = CLBLM_R_X101Y116_SLICE_X159Y116_CO6;
  assign CLBLM_R_X101Y116_SLICE_X159Y116_D = CLBLM_R_X101Y116_SLICE_X159Y116_DO6;
  assign CLBLM_R_X101Y117_SLICE_X158Y117_A = CLBLM_R_X101Y117_SLICE_X158Y117_AO6;
  assign CLBLM_R_X101Y117_SLICE_X158Y117_B = CLBLM_R_X101Y117_SLICE_X158Y117_BO6;
  assign CLBLM_R_X101Y117_SLICE_X158Y117_C = CLBLM_R_X101Y117_SLICE_X158Y117_CO6;
  assign CLBLM_R_X101Y117_SLICE_X158Y117_D = CLBLM_R_X101Y117_SLICE_X158Y117_DO6;
  assign CLBLM_R_X101Y117_SLICE_X159Y117_A = CLBLM_R_X101Y117_SLICE_X159Y117_AO6;
  assign CLBLM_R_X101Y117_SLICE_X159Y117_B = CLBLM_R_X101Y117_SLICE_X159Y117_BO6;
  assign CLBLM_R_X101Y117_SLICE_X159Y117_C = CLBLM_R_X101Y117_SLICE_X159Y117_CO6;
  assign CLBLM_R_X101Y117_SLICE_X159Y117_D = CLBLM_R_X101Y117_SLICE_X159Y117_DO6;
  assign CLBLM_R_X101Y118_SLICE_X158Y118_A = CLBLM_R_X101Y118_SLICE_X158Y118_AO6;
  assign CLBLM_R_X101Y118_SLICE_X158Y118_B = CLBLM_R_X101Y118_SLICE_X158Y118_BO6;
  assign CLBLM_R_X101Y118_SLICE_X158Y118_C = CLBLM_R_X101Y118_SLICE_X158Y118_CO6;
  assign CLBLM_R_X101Y118_SLICE_X158Y118_D = CLBLM_R_X101Y118_SLICE_X158Y118_DO6;
  assign CLBLM_R_X101Y118_SLICE_X159Y118_A = CLBLM_R_X101Y118_SLICE_X159Y118_AO6;
  assign CLBLM_R_X101Y118_SLICE_X159Y118_B = CLBLM_R_X101Y118_SLICE_X159Y118_BO6;
  assign CLBLM_R_X101Y118_SLICE_X159Y118_C = CLBLM_R_X101Y118_SLICE_X159Y118_CO6;
  assign CLBLM_R_X101Y118_SLICE_X159Y118_D = CLBLM_R_X101Y118_SLICE_X159Y118_DO6;
  assign CLBLM_R_X101Y119_SLICE_X158Y119_A = CLBLM_R_X101Y119_SLICE_X158Y119_AO6;
  assign CLBLM_R_X101Y119_SLICE_X158Y119_B = CLBLM_R_X101Y119_SLICE_X158Y119_BO6;
  assign CLBLM_R_X101Y119_SLICE_X158Y119_C = CLBLM_R_X101Y119_SLICE_X158Y119_CO6;
  assign CLBLM_R_X101Y119_SLICE_X158Y119_D = CLBLM_R_X101Y119_SLICE_X158Y119_DO6;
  assign CLBLM_R_X101Y119_SLICE_X159Y119_A = CLBLM_R_X101Y119_SLICE_X159Y119_AO6;
  assign CLBLM_R_X101Y119_SLICE_X159Y119_B = CLBLM_R_X101Y119_SLICE_X159Y119_BO6;
  assign CLBLM_R_X101Y119_SLICE_X159Y119_C = CLBLM_R_X101Y119_SLICE_X159Y119_CO6;
  assign CLBLM_R_X101Y119_SLICE_X159Y119_D = CLBLM_R_X101Y119_SLICE_X159Y119_DO6;
  assign CLBLM_R_X101Y123_SLICE_X158Y123_A = CLBLM_R_X101Y123_SLICE_X158Y123_AO6;
  assign CLBLM_R_X101Y123_SLICE_X158Y123_B = CLBLM_R_X101Y123_SLICE_X158Y123_BO6;
  assign CLBLM_R_X101Y123_SLICE_X158Y123_C = CLBLM_R_X101Y123_SLICE_X158Y123_CO6;
  assign CLBLM_R_X101Y123_SLICE_X158Y123_D = CLBLM_R_X101Y123_SLICE_X158Y123_DO6;
  assign CLBLM_R_X101Y123_SLICE_X158Y123_AMUX = CLBLM_R_X101Y123_SLICE_X158Y123_AO5;
  assign CLBLM_R_X101Y123_SLICE_X159Y123_A = CLBLM_R_X101Y123_SLICE_X159Y123_AO6;
  assign CLBLM_R_X101Y123_SLICE_X159Y123_B = CLBLM_R_X101Y123_SLICE_X159Y123_BO6;
  assign CLBLM_R_X101Y123_SLICE_X159Y123_C = CLBLM_R_X101Y123_SLICE_X159Y123_CO6;
  assign CLBLM_R_X101Y123_SLICE_X159Y123_D = CLBLM_R_X101Y123_SLICE_X159Y123_DO6;
  assign CLBLM_R_X103Y97_SLICE_X162Y97_A = CLBLM_R_X103Y97_SLICE_X162Y97_AO6;
  assign CLBLM_R_X103Y97_SLICE_X162Y97_B = CLBLM_R_X103Y97_SLICE_X162Y97_BO6;
  assign CLBLM_R_X103Y97_SLICE_X162Y97_C = CLBLM_R_X103Y97_SLICE_X162Y97_CO6;
  assign CLBLM_R_X103Y97_SLICE_X162Y97_D = CLBLM_R_X103Y97_SLICE_X162Y97_DO6;
  assign CLBLM_R_X103Y97_SLICE_X163Y97_A = CLBLM_R_X103Y97_SLICE_X163Y97_AO6;
  assign CLBLM_R_X103Y97_SLICE_X163Y97_B = CLBLM_R_X103Y97_SLICE_X163Y97_BO6;
  assign CLBLM_R_X103Y97_SLICE_X163Y97_C = CLBLM_R_X103Y97_SLICE_X163Y97_CO6;
  assign CLBLM_R_X103Y97_SLICE_X163Y97_D = CLBLM_R_X103Y97_SLICE_X163Y97_DO6;
  assign CLBLM_R_X103Y102_SLICE_X162Y102_A = CLBLM_R_X103Y102_SLICE_X162Y102_AO6;
  assign CLBLM_R_X103Y102_SLICE_X162Y102_B = CLBLM_R_X103Y102_SLICE_X162Y102_BO6;
  assign CLBLM_R_X103Y102_SLICE_X162Y102_C = CLBLM_R_X103Y102_SLICE_X162Y102_CO6;
  assign CLBLM_R_X103Y102_SLICE_X162Y102_D = CLBLM_R_X103Y102_SLICE_X162Y102_DO6;
  assign CLBLM_R_X103Y102_SLICE_X163Y102_A = CLBLM_R_X103Y102_SLICE_X163Y102_AO6;
  assign CLBLM_R_X103Y102_SLICE_X163Y102_B = CLBLM_R_X103Y102_SLICE_X163Y102_BO6;
  assign CLBLM_R_X103Y102_SLICE_X163Y102_C = CLBLM_R_X103Y102_SLICE_X163Y102_CO6;
  assign CLBLM_R_X103Y102_SLICE_X163Y102_D = CLBLM_R_X103Y102_SLICE_X163Y102_DO6;
  assign CLBLM_R_X103Y107_SLICE_X162Y107_A = CLBLM_R_X103Y107_SLICE_X162Y107_AO6;
  assign CLBLM_R_X103Y107_SLICE_X162Y107_B = CLBLM_R_X103Y107_SLICE_X162Y107_BO6;
  assign CLBLM_R_X103Y107_SLICE_X162Y107_C = CLBLM_R_X103Y107_SLICE_X162Y107_CO6;
  assign CLBLM_R_X103Y107_SLICE_X162Y107_D = CLBLM_R_X103Y107_SLICE_X162Y107_DO6;
  assign CLBLM_R_X103Y107_SLICE_X163Y107_A = CLBLM_R_X103Y107_SLICE_X163Y107_AO6;
  assign CLBLM_R_X103Y107_SLICE_X163Y107_B = CLBLM_R_X103Y107_SLICE_X163Y107_BO6;
  assign CLBLM_R_X103Y107_SLICE_X163Y107_C = CLBLM_R_X103Y107_SLICE_X163Y107_CO6;
  assign CLBLM_R_X103Y107_SLICE_X163Y107_D = CLBLM_R_X103Y107_SLICE_X163Y107_DO6;
  assign CLBLM_R_X103Y107_SLICE_X163Y107_AMUX = CLBLM_R_X103Y107_SLICE_X163Y107_AO5;
  assign CLBLM_R_X103Y108_SLICE_X162Y108_A = CLBLM_R_X103Y108_SLICE_X162Y108_AO6;
  assign CLBLM_R_X103Y108_SLICE_X162Y108_B = CLBLM_R_X103Y108_SLICE_X162Y108_BO6;
  assign CLBLM_R_X103Y108_SLICE_X162Y108_C = CLBLM_R_X103Y108_SLICE_X162Y108_CO6;
  assign CLBLM_R_X103Y108_SLICE_X162Y108_D = CLBLM_R_X103Y108_SLICE_X162Y108_DO6;
  assign CLBLM_R_X103Y108_SLICE_X163Y108_A = CLBLM_R_X103Y108_SLICE_X163Y108_AO6;
  assign CLBLM_R_X103Y108_SLICE_X163Y108_B = CLBLM_R_X103Y108_SLICE_X163Y108_BO6;
  assign CLBLM_R_X103Y108_SLICE_X163Y108_C = CLBLM_R_X103Y108_SLICE_X163Y108_CO6;
  assign CLBLM_R_X103Y108_SLICE_X163Y108_D = CLBLM_R_X103Y108_SLICE_X163Y108_DO6;
  assign CLBLM_R_X103Y108_SLICE_X163Y108_AMUX = CLBLM_R_X103Y108_SLICE_X163Y108_AO5;
  assign CLBLM_R_X103Y115_SLICE_X162Y115_A = CLBLM_R_X103Y115_SLICE_X162Y115_AO6;
  assign CLBLM_R_X103Y115_SLICE_X162Y115_B = CLBLM_R_X103Y115_SLICE_X162Y115_BO6;
  assign CLBLM_R_X103Y115_SLICE_X162Y115_C = CLBLM_R_X103Y115_SLICE_X162Y115_CO6;
  assign CLBLM_R_X103Y115_SLICE_X162Y115_D = CLBLM_R_X103Y115_SLICE_X162Y115_DO6;
  assign CLBLM_R_X103Y115_SLICE_X163Y115_A = CLBLM_R_X103Y115_SLICE_X163Y115_AO6;
  assign CLBLM_R_X103Y115_SLICE_X163Y115_B = CLBLM_R_X103Y115_SLICE_X163Y115_BO6;
  assign CLBLM_R_X103Y115_SLICE_X163Y115_C = CLBLM_R_X103Y115_SLICE_X163Y115_CO6;
  assign CLBLM_R_X103Y115_SLICE_X163Y115_D = CLBLM_R_X103Y115_SLICE_X163Y115_DO6;
  assign CLBLM_R_X103Y122_SLICE_X162Y122_A = CLBLM_R_X103Y122_SLICE_X162Y122_AO6;
  assign CLBLM_R_X103Y122_SLICE_X162Y122_B = CLBLM_R_X103Y122_SLICE_X162Y122_BO6;
  assign CLBLM_R_X103Y122_SLICE_X162Y122_C = CLBLM_R_X103Y122_SLICE_X162Y122_CO6;
  assign CLBLM_R_X103Y122_SLICE_X162Y122_D = CLBLM_R_X103Y122_SLICE_X162Y122_DO6;
  assign CLBLM_R_X103Y122_SLICE_X163Y122_A = CLBLM_R_X103Y122_SLICE_X163Y122_AO6;
  assign CLBLM_R_X103Y122_SLICE_X163Y122_B = CLBLM_R_X103Y122_SLICE_X163Y122_BO6;
  assign CLBLM_R_X103Y122_SLICE_X163Y122_C = CLBLM_R_X103Y122_SLICE_X163Y122_CO6;
  assign CLBLM_R_X103Y122_SLICE_X163Y122_D = CLBLM_R_X103Y122_SLICE_X163Y122_DO6;
  assign CLBLM_R_X103Y122_SLICE_X163Y122_AMUX = CLBLM_R_X103Y122_SLICE_X163Y122_AO5;
  assign CLBLM_R_X103Y122_SLICE_X163Y122_BMUX = CLBLM_R_X103Y122_SLICE_X163Y122_BO5;
  assign CLBLM_R_X103Y122_SLICE_X163Y122_CMUX = CLBLM_R_X103Y122_SLICE_X163Y122_CO5;
  assign CLBLM_R_X103Y122_SLICE_X163Y122_DMUX = CLBLM_R_X103Y122_SLICE_X163Y122_DO5;
  assign CLBLM_R_X103Y123_SLICE_X162Y123_A = CLBLM_R_X103Y123_SLICE_X162Y123_AO6;
  assign CLBLM_R_X103Y123_SLICE_X162Y123_B = CLBLM_R_X103Y123_SLICE_X162Y123_BO6;
  assign CLBLM_R_X103Y123_SLICE_X162Y123_C = CLBLM_R_X103Y123_SLICE_X162Y123_CO6;
  assign CLBLM_R_X103Y123_SLICE_X162Y123_D = CLBLM_R_X103Y123_SLICE_X162Y123_DO6;
  assign CLBLM_R_X103Y123_SLICE_X163Y123_A = CLBLM_R_X103Y123_SLICE_X163Y123_AO6;
  assign CLBLM_R_X103Y123_SLICE_X163Y123_B = CLBLM_R_X103Y123_SLICE_X163Y123_BO6;
  assign CLBLM_R_X103Y123_SLICE_X163Y123_C = CLBLM_R_X103Y123_SLICE_X163Y123_CO6;
  assign CLBLM_R_X103Y123_SLICE_X163Y123_D = CLBLM_R_X103Y123_SLICE_X163Y123_DO6;
  assign CLBLM_R_X103Y123_SLICE_X163Y123_AMUX = CLBLM_R_X103Y123_SLICE_X163Y123_AO5;
  assign CLBLM_R_X103Y147_SLICE_X162Y147_A = CLBLM_R_X103Y147_SLICE_X162Y147_AO6;
  assign CLBLM_R_X103Y147_SLICE_X162Y147_B = CLBLM_R_X103Y147_SLICE_X162Y147_BO6;
  assign CLBLM_R_X103Y147_SLICE_X162Y147_C = CLBLM_R_X103Y147_SLICE_X162Y147_CO6;
  assign CLBLM_R_X103Y147_SLICE_X162Y147_D = CLBLM_R_X103Y147_SLICE_X162Y147_DO6;
  assign CLBLM_R_X103Y147_SLICE_X163Y147_A = CLBLM_R_X103Y147_SLICE_X163Y147_AO6;
  assign CLBLM_R_X103Y147_SLICE_X163Y147_B = CLBLM_R_X103Y147_SLICE_X163Y147_BO6;
  assign CLBLM_R_X103Y147_SLICE_X163Y147_C = CLBLM_R_X103Y147_SLICE_X163Y147_CO6;
  assign CLBLM_R_X103Y147_SLICE_X163Y147_D = CLBLM_R_X103Y147_SLICE_X163Y147_DO6;
  assign CLBLM_R_X103Y147_SLICE_X163Y147_AMUX = CLBLM_R_X103Y147_SLICE_X163Y147_AO5;
  assign CLBLM_R_X103Y177_SLICE_X162Y177_A = CLBLM_R_X103Y177_SLICE_X162Y177_AO6;
  assign CLBLM_R_X103Y177_SLICE_X162Y177_B = CLBLM_R_X103Y177_SLICE_X162Y177_BO6;
  assign CLBLM_R_X103Y177_SLICE_X162Y177_C = CLBLM_R_X103Y177_SLICE_X162Y177_CO6;
  assign CLBLM_R_X103Y177_SLICE_X162Y177_D = CLBLM_R_X103Y177_SLICE_X162Y177_DO6;
  assign CLBLM_R_X103Y177_SLICE_X163Y177_A = CLBLM_R_X103Y177_SLICE_X163Y177_AO6;
  assign CLBLM_R_X103Y177_SLICE_X163Y177_B = CLBLM_R_X103Y177_SLICE_X163Y177_BO6;
  assign CLBLM_R_X103Y177_SLICE_X163Y177_C = CLBLM_R_X103Y177_SLICE_X163Y177_CO6;
  assign CLBLM_R_X103Y177_SLICE_X163Y177_D = CLBLM_R_X103Y177_SLICE_X163Y177_DO6;
  assign CLBLM_R_X103Y177_SLICE_X163Y177_AMUX = CLBLM_R_X103Y177_SLICE_X163Y177_AO5;
  assign CLBLM_R_X103Y185_SLICE_X162Y185_A = CLBLM_R_X103Y185_SLICE_X162Y185_AO6;
  assign CLBLM_R_X103Y185_SLICE_X162Y185_B = CLBLM_R_X103Y185_SLICE_X162Y185_BO6;
  assign CLBLM_R_X103Y185_SLICE_X162Y185_C = CLBLM_R_X103Y185_SLICE_X162Y185_CO6;
  assign CLBLM_R_X103Y185_SLICE_X162Y185_D = CLBLM_R_X103Y185_SLICE_X162Y185_DO6;
  assign CLBLM_R_X103Y185_SLICE_X163Y185_A = CLBLM_R_X103Y185_SLICE_X163Y185_AO6;
  assign CLBLM_R_X103Y185_SLICE_X163Y185_B = CLBLM_R_X103Y185_SLICE_X163Y185_BO6;
  assign CLBLM_R_X103Y185_SLICE_X163Y185_C = CLBLM_R_X103Y185_SLICE_X163Y185_CO6;
  assign CLBLM_R_X103Y185_SLICE_X163Y185_D = CLBLM_R_X103Y185_SLICE_X163Y185_DO6;
  assign CLBLM_R_X103Y193_SLICE_X162Y193_A = CLBLM_R_X103Y193_SLICE_X162Y193_AO6;
  assign CLBLM_R_X103Y193_SLICE_X162Y193_B = CLBLM_R_X103Y193_SLICE_X162Y193_BO6;
  assign CLBLM_R_X103Y193_SLICE_X162Y193_C = CLBLM_R_X103Y193_SLICE_X162Y193_CO6;
  assign CLBLM_R_X103Y193_SLICE_X162Y193_D = CLBLM_R_X103Y193_SLICE_X162Y193_DO6;
  assign CLBLM_R_X103Y193_SLICE_X163Y193_A = CLBLM_R_X103Y193_SLICE_X163Y193_AO6;
  assign CLBLM_R_X103Y193_SLICE_X163Y193_B = CLBLM_R_X103Y193_SLICE_X163Y193_BO6;
  assign CLBLM_R_X103Y193_SLICE_X163Y193_C = CLBLM_R_X103Y193_SLICE_X163Y193_CO6;
  assign CLBLM_R_X103Y193_SLICE_X163Y193_D = CLBLM_R_X103Y193_SLICE_X163Y193_DO6;
  assign LIOI3_X0Y51_ILOGIC_X0Y52_O = LIOB33_X0Y51_IOB_X0Y52_I;
  assign LIOI3_X0Y51_ILOGIC_X0Y51_O = LIOB33_X0Y51_IOB_X0Y51_I;
  assign LIOI3_X0Y53_ILOGIC_X0Y54_O = LIOB33_X0Y53_IOB_X0Y54_I;
  assign LIOI3_X0Y53_ILOGIC_X0Y53_O = LIOB33_X0Y53_IOB_X0Y53_I;
  assign LIOI3_X0Y55_ILOGIC_X0Y56_O = LIOB33_X0Y55_IOB_X0Y56_I;
  assign LIOI3_X0Y55_ILOGIC_X0Y55_O = LIOB33_X0Y55_IOB_X0Y55_I;
  assign LIOI3_X0Y59_ILOGIC_X0Y60_O = LIOB33_X0Y59_IOB_X0Y60_I;
  assign LIOI3_X0Y59_ILOGIC_X0Y59_O = LIOB33_X0Y59_IOB_X0Y59_I;
  assign LIOI3_X0Y61_ILOGIC_X0Y62_O = LIOB33_X0Y61_IOB_X0Y62_I;
  assign LIOI3_X0Y65_ILOGIC_X0Y66_O = LIOB33_X0Y65_IOB_X0Y66_I;
  assign LIOI3_X0Y65_ILOGIC_X0Y65_O = LIOB33_X0Y65_IOB_X0Y65_I;
  assign LIOI3_X0Y67_ILOGIC_X0Y68_O = LIOB33_X0Y67_IOB_X0Y68_I;
  assign LIOI3_X0Y67_ILOGIC_X0Y67_O = LIOB33_X0Y67_IOB_X0Y67_I;
  assign LIOI3_X0Y71_ILOGIC_X0Y72_O = LIOB33_X0Y71_IOB_X0Y72_I;
  assign LIOI3_X0Y71_ILOGIC_X0Y71_O = LIOB33_X0Y71_IOB_X0Y71_I;
  assign LIOI3_X0Y73_ILOGIC_X0Y74_O = LIOB33_X0Y73_IOB_X0Y74_I;
  assign LIOI3_X0Y75_ILOGIC_X0Y76_O = LIOB33_X0Y75_IOB_X0Y76_I;
  assign LIOI3_X0Y75_ILOGIC_X0Y75_O = LIOB33_X0Y75_IOB_X0Y75_I;
  assign LIOI3_X0Y77_ILOGIC_X0Y78_O = LIOB33_X0Y77_IOB_X0Y78_I;
  assign LIOI3_X0Y77_ILOGIC_X0Y77_O = LIOB33_X0Y77_IOB_X0Y77_I;
  assign LIOI3_X0Y79_ILOGIC_X0Y80_O = LIOB33_X0Y79_IOB_X0Y80_I;
  assign LIOI3_X0Y79_ILOGIC_X0Y79_O = LIOB33_X0Y79_IOB_X0Y79_I;
  assign LIOI3_X0Y83_ILOGIC_X0Y84_O = LIOB33_X0Y83_IOB_X0Y84_I;
  assign LIOI3_X0Y83_ILOGIC_X0Y83_O = LIOB33_X0Y83_IOB_X0Y83_I;
  assign LIOI3_X0Y85_ILOGIC_X0Y86_O = LIOB33_X0Y85_IOB_X0Y86_I;
  assign LIOI3_X0Y85_ILOGIC_X0Y85_O = LIOB33_X0Y85_IOB_X0Y85_I;
  assign LIOI3_X0Y89_ILOGIC_X0Y90_O = LIOB33_X0Y89_IOB_X0Y90_I;
  assign LIOI3_X0Y89_ILOGIC_X0Y89_O = LIOB33_X0Y89_IOB_X0Y89_I;
  assign LIOI3_X0Y91_ILOGIC_X0Y92_O = LIOB33_X0Y91_IOB_X0Y92_I;
  assign LIOI3_X0Y91_ILOGIC_X0Y91_O = LIOB33_X0Y91_IOB_X0Y91_I;
  assign LIOI3_X0Y95_ILOGIC_X0Y96_O = LIOB33_X0Y95_IOB_X0Y96_I;
  assign LIOI3_X0Y95_ILOGIC_X0Y95_O = LIOB33_X0Y95_IOB_X0Y95_I;
  assign LIOI3_X0Y97_ILOGIC_X0Y98_O = LIOB33_X0Y97_IOB_X0Y98_I;
  assign LIOI3_X0Y97_ILOGIC_X0Y97_O = LIOB33_X0Y97_IOB_X0Y97_I;
  assign LIOI3_X0Y101_ILOGIC_X0Y102_O = LIOB33_X0Y101_IOB_X0Y102_I;
  assign LIOI3_X0Y101_ILOGIC_X0Y101_O = LIOB33_X0Y101_IOB_X0Y101_I;
  assign LIOI3_X0Y103_ILOGIC_X0Y104_O = LIOB33_X0Y103_IOB_X0Y104_I;
  assign LIOI3_X0Y103_ILOGIC_X0Y103_O = LIOB33_X0Y103_IOB_X0Y103_I;
  assign LIOI3_X0Y105_ILOGIC_X0Y106_O = LIOB33_X0Y105_IOB_X0Y106_I;
  assign LIOI3_X0Y105_ILOGIC_X0Y105_O = LIOB33_X0Y105_IOB_X0Y105_I;
  assign LIOI3_X0Y109_ILOGIC_X0Y110_O = LIOB33_X0Y109_IOB_X0Y110_I;
  assign LIOI3_X0Y109_ILOGIC_X0Y109_O = LIOB33_X0Y109_IOB_X0Y109_I;
  assign LIOI3_X0Y111_ILOGIC_X0Y112_O = LIOB33_X0Y111_IOB_X0Y112_I;
  assign LIOI3_X0Y111_ILOGIC_X0Y111_O = LIOB33_X0Y111_IOB_X0Y111_I;
  assign LIOI3_X0Y115_ILOGIC_X0Y116_O = LIOB33_X0Y115_IOB_X0Y116_I;
  assign LIOI3_X0Y115_ILOGIC_X0Y115_O = LIOB33_X0Y115_IOB_X0Y115_I;
  assign LIOI3_X0Y117_ILOGIC_X0Y118_O = LIOB33_X0Y117_IOB_X0Y118_I;
  assign LIOI3_X0Y117_ILOGIC_X0Y117_O = LIOB33_X0Y117_IOB_X0Y117_I;
  assign LIOI3_X0Y121_ILOGIC_X0Y122_O = LIOB33_X0Y121_IOB_X0Y122_I;
  assign LIOI3_X0Y121_ILOGIC_X0Y121_O = LIOB33_X0Y121_IOB_X0Y121_I;
  assign LIOI3_X0Y123_ILOGIC_X0Y124_O = LIOB33_X0Y123_IOB_X0Y124_I;
  assign LIOI3_X0Y123_ILOGIC_X0Y123_O = LIOB33_X0Y123_IOB_X0Y123_I;
  assign LIOI3_X0Y125_ILOGIC_X0Y126_O = LIOB33_X0Y125_IOB_X0Y126_I;
  assign LIOI3_X0Y125_ILOGIC_X0Y125_O = LIOB33_X0Y125_IOB_X0Y125_I;
  assign LIOI3_X0Y127_ILOGIC_X0Y128_O = LIOB33_X0Y127_IOB_X0Y128_I;
  assign LIOI3_X0Y127_ILOGIC_X0Y127_O = LIOB33_X0Y127_IOB_X0Y127_I;
  assign LIOI3_X0Y129_ILOGIC_X0Y130_O = LIOB33_X0Y129_IOB_X0Y130_I;
  assign LIOI3_X0Y129_ILOGIC_X0Y129_O = LIOB33_X0Y129_IOB_X0Y129_I;
  assign LIOI3_X0Y133_ILOGIC_X0Y134_O = LIOB33_X0Y133_IOB_X0Y134_I;
  assign LIOI3_X0Y133_ILOGIC_X0Y133_O = LIOB33_X0Y133_IOB_X0Y133_I;
  assign LIOI3_X0Y135_ILOGIC_X0Y136_O = LIOB33_X0Y135_IOB_X0Y136_I;
  assign LIOI3_X0Y135_ILOGIC_X0Y135_O = LIOB33_X0Y135_IOB_X0Y135_I;
  assign LIOI3_X0Y139_ILOGIC_X0Y140_O = LIOB33_X0Y139_IOB_X0Y140_I;
  assign LIOI3_X0Y139_ILOGIC_X0Y139_O = LIOB33_X0Y139_IOB_X0Y139_I;
  assign LIOI3_X0Y141_ILOGIC_X0Y142_O = LIOB33_X0Y141_IOB_X0Y142_I;
  assign LIOI3_X0Y141_ILOGIC_X0Y141_O = LIOB33_X0Y141_IOB_X0Y141_I;
  assign LIOI3_X0Y145_ILOGIC_X0Y146_O = LIOB33_X0Y145_IOB_X0Y146_I;
  assign LIOI3_X0Y145_ILOGIC_X0Y145_O = LIOB33_X0Y145_IOB_X0Y145_I;
  assign LIOI3_X0Y147_ILOGIC_X0Y147_O = LIOB33_X0Y147_IOB_X0Y147_I;
  assign LIOI3_X0Y151_ILOGIC_X0Y152_O = LIOB33_X0Y151_IOB_X0Y152_I;
  assign LIOI3_X0Y151_ILOGIC_X0Y151_O = LIOB33_X0Y151_IOB_X0Y151_I;
  assign LIOI3_X0Y153_ILOGIC_X0Y154_O = LIOB33_X0Y153_IOB_X0Y154_I;
  assign LIOI3_X0Y153_ILOGIC_X0Y153_O = LIOB33_X0Y153_IOB_X0Y153_I;
  assign LIOI3_X0Y155_ILOGIC_X0Y156_O = LIOB33_X0Y155_IOB_X0Y156_I;
  assign LIOI3_X0Y155_ILOGIC_X0Y155_O = LIOB33_X0Y155_IOB_X0Y155_I;
  assign LIOI3_X0Y159_ILOGIC_X0Y160_O = LIOB33_X0Y159_IOB_X0Y160_I;
  assign LIOI3_X0Y159_ILOGIC_X0Y159_O = LIOB33_X0Y159_IOB_X0Y159_I;
  assign LIOI3_X0Y161_ILOGIC_X0Y162_O = LIOB33_X0Y161_IOB_X0Y162_I;
  assign LIOI3_X0Y161_ILOGIC_X0Y161_O = LIOB33_X0Y161_IOB_X0Y161_I;
  assign LIOI3_X0Y165_ILOGIC_X0Y166_O = LIOB33_X0Y165_IOB_X0Y166_I;
  assign LIOI3_X0Y165_ILOGIC_X0Y165_O = LIOB33_X0Y165_IOB_X0Y165_I;
  assign LIOI3_X0Y171_ILOGIC_X0Y172_O = LIOB33_X0Y171_IOB_X0Y172_I;
  assign LIOI3_X0Y171_ILOGIC_X0Y171_O = LIOB33_X0Y171_IOB_X0Y171_I;
  assign LIOI3_X0Y173_ILOGIC_X0Y174_O = LIOB33_X0Y173_IOB_X0Y174_I;
  assign LIOI3_X0Y173_ILOGIC_X0Y173_O = LIOB33_X0Y173_IOB_X0Y173_I;
  assign LIOI3_X0Y175_ILOGIC_X0Y176_O = LIOB33_X0Y175_IOB_X0Y176_I;
  assign LIOI3_X0Y175_ILOGIC_X0Y175_O = LIOB33_X0Y175_IOB_X0Y175_I;
  assign LIOI3_X0Y177_ILOGIC_X0Y177_O = LIOB33_X0Y177_IOB_X0Y177_I;
  assign LIOI3_X0Y177_OLOGIC_X0Y178_OQ = CLBLL_L_X2Y175_SLICE_X0Y175_AO6;
  assign LIOI3_X0Y177_OLOGIC_X0Y178_TQ = 1'b1;
  assign LIOI3_X0Y179_OLOGIC_X0Y180_OQ = LIOB33_X0Y133_IOB_X0Y133_I;
  assign LIOI3_X0Y179_OLOGIC_X0Y180_TQ = 1'b1;
  assign LIOI3_X0Y179_OLOGIC_X0Y179_OQ = LIOB33_X0Y133_IOB_X0Y134_I;
  assign LIOI3_X0Y179_OLOGIC_X0Y179_TQ = 1'b1;
  assign LIOI3_X0Y183_OLOGIC_X0Y184_OQ = CLBLM_R_X103Y108_SLICE_X163Y108_AO5;
  assign LIOI3_X0Y183_OLOGIC_X0Y184_TQ = 1'b1;
  assign LIOI3_X0Y183_OLOGIC_X0Y183_OQ = LIOB33_X0Y101_IOB_X0Y102_I;
  assign LIOI3_X0Y183_OLOGIC_X0Y183_TQ = 1'b1;
  assign LIOI3_X0Y185_OLOGIC_X0Y186_OQ = LIOB33_X0Y135_IOB_X0Y135_I;
  assign LIOI3_X0Y185_OLOGIC_X0Y186_TQ = 1'b1;
  assign LIOI3_X0Y185_OLOGIC_X0Y185_OQ = LIOB33_X0Y67_IOB_X0Y67_I;
  assign LIOI3_X0Y185_OLOGIC_X0Y185_TQ = 1'b1;
  assign LIOI3_X0Y189_OLOGIC_X0Y190_OQ = CLBLL_L_X2Y173_SLICE_X1Y173_BO6;
  assign LIOI3_X0Y189_OLOGIC_X0Y190_TQ = 1'b1;
  assign LIOI3_X0Y189_OLOGIC_X0Y189_OQ = CLBLL_L_X2Y173_SLICE_X1Y173_BO6;
  assign LIOI3_X0Y189_OLOGIC_X0Y189_TQ = 1'b1;
  assign LIOI3_X0Y191_OLOGIC_X0Y192_OQ = CLBLM_R_X5Y114_SLICE_X6Y114_AO6;
  assign LIOI3_X0Y191_OLOGIC_X0Y192_TQ = 1'b1;
  assign LIOI3_X0Y191_OLOGIC_X0Y191_OQ = CLBLM_R_X5Y113_SLICE_X7Y113_AO6;
  assign LIOI3_X0Y191_OLOGIC_X0Y191_TQ = 1'b1;
  assign LIOI3_X0Y195_OLOGIC_X0Y196_OQ = CLBLM_R_X3Y112_SLICE_X3Y112_BO6;
  assign LIOI3_X0Y195_OLOGIC_X0Y196_TQ = 1'b1;
  assign LIOI3_X0Y195_OLOGIC_X0Y195_OQ = 1'b0;
  assign LIOI3_X0Y195_OLOGIC_X0Y195_TQ = 1'b1;
  assign LIOI3_X0Y197_OLOGIC_X0Y198_OQ = CLBLL_L_X2Y102_SLICE_X0Y102_BO6;
  assign LIOI3_X0Y197_OLOGIC_X0Y198_TQ = 1'b1;
  assign LIOI3_X0Y197_OLOGIC_X0Y197_OQ = CLBLL_L_X4Y110_SLICE_X4Y110_CO5;
  assign LIOI3_X0Y197_OLOGIC_X0Y197_TQ = 1'b1;
  assign LIOI3_SING_X0Y50_ILOGIC_X0Y50_O = LIOB33_SING_X0Y50_IOB_X0Y50_I;
  assign LIOI3_SING_X0Y99_ILOGIC_X0Y99_O = LIOB33_SING_X0Y99_IOB_X0Y99_I;
  assign LIOI3_SING_X0Y100_ILOGIC_X0Y100_O = LIOB33_SING_X0Y100_IOB_X0Y100_I;
  assign LIOI3_SING_X0Y150_ILOGIC_X0Y150_O = LIOB33_SING_X0Y150_IOB_X0Y150_I;
  assign LIOI3_SING_X0Y199_OLOGIC_X0Y199_OQ = CLBLL_L_X4Y111_SLICE_X5Y111_CO6;
  assign LIOI3_SING_X0Y199_OLOGIC_X0Y199_TQ = 1'b1;
  assign LIOI3_SING_X0Y200_OLOGIC_X0Y200_OQ = LIOB33_SING_X0Y100_IOB_X0Y100_I;
  assign LIOI3_SING_X0Y200_OLOGIC_X0Y200_TQ = 1'b1;
  assign LIOI3_TBYTESRC_X0Y57_ILOGIC_X0Y58_O = LIOB33_X0Y57_IOB_X0Y58_I;
  assign LIOI3_TBYTESRC_X0Y57_ILOGIC_X0Y57_O = LIOB33_X0Y57_IOB_X0Y57_I;
  assign LIOI3_TBYTESRC_X0Y69_ILOGIC_X0Y70_O = LIOB33_X0Y69_IOB_X0Y70_I;
  assign LIOI3_TBYTESRC_X0Y81_ILOGIC_X0Y82_O = LIOB33_X0Y81_IOB_X0Y82_I;
  assign LIOI3_TBYTESRC_X0Y81_ILOGIC_X0Y81_O = LIOB33_X0Y81_IOB_X0Y81_I;
  assign LIOI3_TBYTESRC_X0Y93_ILOGIC_X0Y94_O = LIOB33_X0Y93_IOB_X0Y94_I;
  assign LIOI3_TBYTESRC_X0Y93_ILOGIC_X0Y93_O = LIOB33_X0Y93_IOB_X0Y93_I;
  assign LIOI3_TBYTESRC_X0Y107_ILOGIC_X0Y108_O = LIOB33_X0Y107_IOB_X0Y108_I;
  assign LIOI3_TBYTESRC_X0Y107_ILOGIC_X0Y107_O = LIOB33_X0Y107_IOB_X0Y107_I;
  assign LIOI3_TBYTESRC_X0Y119_ILOGIC_X0Y120_O = LIOB33_X0Y119_IOB_X0Y120_I;
  assign LIOI3_TBYTESRC_X0Y119_ILOGIC_X0Y119_O = LIOB33_X0Y119_IOB_X0Y119_I;
  assign LIOI3_TBYTESRC_X0Y131_ILOGIC_X0Y132_O = LIOB33_X0Y131_IOB_X0Y132_I;
  assign LIOI3_TBYTESRC_X0Y131_ILOGIC_X0Y131_O = LIOB33_X0Y131_IOB_X0Y131_I;
  assign LIOI3_TBYTESRC_X0Y143_ILOGIC_X0Y143_O = LIOB33_X0Y143_IOB_X0Y143_I;
  assign LIOI3_TBYTESRC_X0Y157_ILOGIC_X0Y158_O = LIOB33_X0Y157_IOB_X0Y158_I;
  assign LIOI3_TBYTESRC_X0Y157_ILOGIC_X0Y157_O = LIOB33_X0Y157_IOB_X0Y157_I;
  assign LIOI3_TBYTESRC_X0Y181_OLOGIC_X0Y182_OQ = LIOB33_X0Y97_IOB_X0Y97_I;
  assign LIOI3_TBYTESRC_X0Y181_OLOGIC_X0Y182_TQ = 1'b1;
  assign LIOI3_TBYTESRC_X0Y181_OLOGIC_X0Y181_OQ = LIOB33_X0Y133_IOB_X0Y133_I;
  assign LIOI3_TBYTESRC_X0Y181_OLOGIC_X0Y181_TQ = 1'b1;
  assign LIOI3_TBYTESRC_X0Y193_OLOGIC_X0Y194_OQ = 1'b0;
  assign LIOI3_TBYTESRC_X0Y193_OLOGIC_X0Y194_TQ = 1'b1;
  assign LIOI3_TBYTESRC_X0Y193_OLOGIC_X0Y193_OQ = CLBLM_R_X3Y112_SLICE_X3Y112_BO6;
  assign LIOI3_TBYTESRC_X0Y193_OLOGIC_X0Y193_TQ = 1'b1;
  assign LIOI3_TBYTETERM_X0Y63_ILOGIC_X0Y63_O = LIOB33_X0Y63_IOB_X0Y63_I;
  assign LIOI3_TBYTETERM_X0Y87_ILOGIC_X0Y88_O = LIOB33_X0Y87_IOB_X0Y88_I;
  assign LIOI3_TBYTETERM_X0Y87_ILOGIC_X0Y87_O = LIOB33_X0Y87_IOB_X0Y87_I;
  assign LIOI3_TBYTETERM_X0Y113_ILOGIC_X0Y114_O = LIOB33_X0Y113_IOB_X0Y114_I;
  assign LIOI3_TBYTETERM_X0Y113_ILOGIC_X0Y113_O = LIOB33_X0Y113_IOB_X0Y113_I;
  assign LIOI3_TBYTETERM_X0Y137_ILOGIC_X0Y138_O = LIOB33_X0Y137_IOB_X0Y138_I;
  assign LIOI3_TBYTETERM_X0Y137_ILOGIC_X0Y137_O = LIOB33_X0Y137_IOB_X0Y137_I;
  assign LIOI3_TBYTETERM_X0Y163_ILOGIC_X0Y164_O = LIOB33_X0Y163_IOB_X0Y164_I;
  assign LIOI3_TBYTETERM_X0Y163_ILOGIC_X0Y163_O = LIOB33_X0Y163_IOB_X0Y163_I;
  assign LIOI3_TBYTETERM_X0Y187_OLOGIC_X0Y188_OQ = CLBLL_L_X2Y173_SLICE_X1Y173_BO6;
  assign LIOI3_TBYTETERM_X0Y187_OLOGIC_X0Y188_TQ = 1'b1;
  assign LIOI3_TBYTETERM_X0Y187_OLOGIC_X0Y187_OQ = CLBLL_L_X2Y173_SLICE_X1Y173_BO6;
  assign LIOI3_TBYTETERM_X0Y187_OLOGIC_X0Y187_TQ = 1'b1;
  assign RIOI3_X105Y51_OLOGIC_X1Y52_OQ = CLBLM_R_X49Y95_SLICE_X74Y95_AO6;
  assign RIOI3_X105Y51_OLOGIC_X1Y52_TQ = 1'b1;
  assign RIOI3_X105Y51_OLOGIC_X1Y51_OQ = CLBLL_L_X4Y111_SLICE_X5Y111_CO6;
  assign RIOI3_X105Y51_OLOGIC_X1Y51_TQ = 1'b1;
  assign RIOI3_X105Y53_OLOGIC_X1Y54_OQ = CLBLM_R_X103Y108_SLICE_X163Y108_AO6;
  assign RIOI3_X105Y53_OLOGIC_X1Y54_TQ = 1'b1;
  assign RIOI3_X105Y53_OLOGIC_X1Y53_OQ = CLBLM_L_X10Y113_SLICE_X12Y113_AO6;
  assign RIOI3_X105Y53_OLOGIC_X1Y53_TQ = 1'b1;
  assign RIOI3_X105Y55_OLOGIC_X1Y56_OQ = CLBLM_R_X5Y111_SLICE_X7Y111_BO6;
  assign RIOI3_X105Y55_OLOGIC_X1Y56_TQ = 1'b1;
  assign RIOI3_X105Y55_OLOGIC_X1Y55_OQ = CLBLM_L_X10Y114_SLICE_X12Y114_AO6;
  assign RIOI3_X105Y55_OLOGIC_X1Y55_TQ = 1'b1;
  assign RIOI3_X105Y59_OLOGIC_X1Y60_OQ = CLBLM_L_X10Y113_SLICE_X12Y113_BO6;
  assign RIOI3_X105Y59_OLOGIC_X1Y60_TQ = 1'b1;
  assign RIOI3_X105Y59_OLOGIC_X1Y59_OQ = CLBLM_R_X5Y113_SLICE_X6Y113_BO6;
  assign RIOI3_X105Y59_OLOGIC_X1Y59_TQ = 1'b1;
  assign RIOI3_X105Y61_OLOGIC_X1Y62_OQ = CLBLL_L_X100Y121_SLICE_X156Y121_BO6;
  assign RIOI3_X105Y61_OLOGIC_X1Y62_TQ = 1'b1;
  assign RIOI3_X105Y61_OLOGIC_X1Y61_OQ = CLBLM_L_X8Y113_SLICE_X11Y113_BO6;
  assign RIOI3_X105Y61_OLOGIC_X1Y61_TQ = 1'b1;
  assign RIOI3_X105Y65_OLOGIC_X1Y66_OQ = CLBLM_R_X5Y112_SLICE_X6Y112_AO6;
  assign RIOI3_X105Y65_OLOGIC_X1Y66_TQ = 1'b1;
  assign RIOI3_X105Y65_OLOGIC_X1Y65_OQ = CLBLM_R_X103Y107_SLICE_X163Y107_AO5;
  assign RIOI3_X105Y65_OLOGIC_X1Y65_TQ = 1'b1;
  assign RIOI3_X105Y67_OLOGIC_X1Y68_OQ = CLBLL_L_X4Y109_SLICE_X4Y109_AO6;
  assign RIOI3_X105Y67_OLOGIC_X1Y68_TQ = 1'b1;
  assign RIOI3_X105Y67_OLOGIC_X1Y67_OQ = CLBLM_R_X5Y109_SLICE_X6Y109_AO6;
  assign RIOI3_X105Y67_OLOGIC_X1Y67_TQ = 1'b1;
  assign RIOI3_X105Y71_OLOGIC_X1Y72_OQ = CLBLM_R_X103Y122_SLICE_X163Y122_BO6;
  assign RIOI3_X105Y71_OLOGIC_X1Y72_TQ = 1'b1;
  assign RIOI3_X105Y71_OLOGIC_X1Y71_OQ = CLBLM_R_X103Y122_SLICE_X163Y122_AO6;
  assign RIOI3_X105Y71_OLOGIC_X1Y71_TQ = 1'b1;
  assign RIOI3_X105Y73_OLOGIC_X1Y74_OQ = CLBLL_L_X100Y113_SLICE_X156Y113_AO6;
  assign RIOI3_X105Y73_OLOGIC_X1Y74_TQ = 1'b1;
  assign RIOI3_X105Y73_OLOGIC_X1Y73_OQ = CLBLL_L_X36Y113_SLICE_X54Y113_AO6;
  assign RIOI3_X105Y73_OLOGIC_X1Y73_TQ = 1'b1;
  assign RIOI3_X105Y75_OLOGIC_X1Y76_OQ = CLBLL_R_X57Y113_SLICE_X86Y113_BO6;
  assign RIOI3_X105Y75_OLOGIC_X1Y76_TQ = 1'b1;
  assign RIOI3_X105Y75_OLOGIC_X1Y75_OQ = CLBLM_R_X29Y115_SLICE_X42Y115_AO6;
  assign RIOI3_X105Y75_OLOGIC_X1Y75_TQ = 1'b1;
  assign RIOI3_X105Y77_OLOGIC_X1Y78_OQ = CLBLL_L_X100Y113_SLICE_X156Y113_BO6;
  assign RIOI3_X105Y77_OLOGIC_X1Y78_TQ = 1'b1;
  assign RIOI3_X105Y77_OLOGIC_X1Y77_OQ = CLBLL_L_X36Y113_SLICE_X54Y113_BO6;
  assign RIOI3_X105Y77_OLOGIC_X1Y77_TQ = 1'b1;
  assign RIOI3_X105Y79_OLOGIC_X1Y80_OQ = CLBLM_R_X103Y97_SLICE_X163Y97_AO6;
  assign RIOI3_X105Y79_OLOGIC_X1Y80_TQ = 1'b1;
  assign RIOI3_X105Y79_OLOGIC_X1Y79_OQ = CLBLM_R_X29Y115_SLICE_X42Y115_BO6;
  assign RIOI3_X105Y79_OLOGIC_X1Y79_TQ = 1'b1;
  assign RIOI3_X105Y83_OLOGIC_X1Y84_OQ = CLBLM_R_X103Y97_SLICE_X163Y97_BO6;
  assign RIOI3_X105Y83_OLOGIC_X1Y84_TQ = 1'b1;
  assign RIOI3_X105Y83_OLOGIC_X1Y83_OQ = CLBLM_R_X103Y102_SLICE_X163Y102_AO6;
  assign RIOI3_X105Y83_OLOGIC_X1Y83_TQ = 1'b1;
  assign RIOI3_X105Y85_OLOGIC_X1Y86_OQ = CLBLM_R_X103Y107_SLICE_X163Y107_AO6;
  assign RIOI3_X105Y85_OLOGIC_X1Y86_TQ = 1'b1;
  assign RIOI3_X105Y85_OLOGIC_X1Y85_OQ = CLBLM_R_X103Y122_SLICE_X163Y122_DO6;
  assign RIOI3_X105Y85_OLOGIC_X1Y85_TQ = 1'b1;
  assign RIOI3_X105Y89_OLOGIC_X1Y90_OQ = CLBLM_L_X8Y113_SLICE_X10Y113_DO6;
  assign RIOI3_X105Y89_OLOGIC_X1Y90_TQ = 1'b1;
  assign RIOI3_X105Y89_OLOGIC_X1Y89_OQ = CLBLM_R_X49Y101_SLICE_X74Y101_AO5;
  assign RIOI3_X105Y89_OLOGIC_X1Y89_TQ = 1'b1;
  assign RIOI3_X105Y91_OLOGIC_X1Y92_OQ = CLBLM_L_X10Y113_SLICE_X13Y113_AO6;
  assign RIOI3_X105Y91_OLOGIC_X1Y92_TQ = 1'b1;
  assign RIOI3_X105Y91_OLOGIC_X1Y91_OQ = CLBLM_L_X10Y113_SLICE_X12Y113_CO6;
  assign RIOI3_X105Y91_OLOGIC_X1Y91_TQ = 1'b1;
  assign RIOI3_X105Y95_OLOGIC_X1Y96_OQ = CLBLM_R_X25Y116_SLICE_X36Y116_BO6;
  assign RIOI3_X105Y95_OLOGIC_X1Y96_TQ = 1'b1;
  assign RIOI3_X105Y95_OLOGIC_X1Y95_OQ = CLBLM_L_X10Y114_SLICE_X12Y114_BO6;
  assign RIOI3_X105Y95_OLOGIC_X1Y95_TQ = 1'b1;
  assign RIOI3_X105Y97_OLOGIC_X1Y98_OQ = CLBLM_R_X25Y115_SLICE_X36Y115_BO6;
  assign RIOI3_X105Y97_OLOGIC_X1Y98_TQ = 1'b1;
  assign RIOI3_X105Y97_OLOGIC_X1Y97_OQ = CLBLM_R_X5Y115_SLICE_X7Y115_AO6;
  assign RIOI3_X105Y97_OLOGIC_X1Y97_TQ = 1'b1;
  assign RIOI3_X105Y101_ILOGIC_X1Y102_O = RIOB33_X105Y101_IOB_X1Y102_I;
  assign RIOI3_X105Y101_ILOGIC_X1Y101_O = RIOB33_X105Y101_IOB_X1Y101_I;
  assign RIOI3_X105Y103_ILOGIC_X1Y104_O = RIOB33_X105Y103_IOB_X1Y104_I;
  assign RIOI3_X105Y103_ILOGIC_X1Y103_O = RIOB33_X105Y103_IOB_X1Y103_I;
  assign RIOI3_X105Y105_ILOGIC_X1Y106_O = RIOB33_X105Y105_IOB_X1Y106_I;
  assign RIOI3_X105Y105_ILOGIC_X1Y105_O = RIOB33_X105Y105_IOB_X1Y105_I;
  assign RIOI3_X105Y109_ILOGIC_X1Y110_O = RIOB33_X105Y109_IOB_X1Y110_I;
  assign RIOI3_X105Y109_ILOGIC_X1Y109_O = RIOB33_X105Y109_IOB_X1Y109_I;
  assign RIOI3_X105Y111_ILOGIC_X1Y112_O = RIOB33_X105Y111_IOB_X1Y112_I;
  assign RIOI3_X105Y111_ILOGIC_X1Y111_O = RIOB33_X105Y111_IOB_X1Y111_I;
  assign RIOI3_X105Y115_ILOGIC_X1Y116_O = RIOB33_X105Y115_IOB_X1Y116_I;
  assign RIOI3_X105Y115_ILOGIC_X1Y115_O = RIOB33_X105Y115_IOB_X1Y115_I;
  assign RIOI3_X105Y117_ILOGIC_X1Y118_O = RIOB33_X105Y117_IOB_X1Y118_I;
  assign RIOI3_X105Y117_ILOGIC_X1Y117_O = RIOB33_X105Y117_IOB_X1Y117_I;
  assign RIOI3_X105Y121_ILOGIC_X1Y122_O = RIOB33_X105Y121_IOB_X1Y122_I;
  assign RIOI3_X105Y121_ILOGIC_X1Y121_O = RIOB33_X105Y121_IOB_X1Y121_I;
  assign RIOI3_X105Y123_ILOGIC_X1Y124_O = RIOB33_X105Y123_IOB_X1Y124_I;
  assign RIOI3_X105Y123_ILOGIC_X1Y123_O = RIOB33_X105Y123_IOB_X1Y123_I;
  assign RIOI3_X105Y125_ILOGIC_X1Y126_O = RIOB33_X105Y125_IOB_X1Y126_I;
  assign RIOI3_X105Y125_ILOGIC_X1Y125_O = RIOB33_X105Y125_IOB_X1Y125_I;
  assign RIOI3_X105Y127_OLOGIC_X1Y128_OQ = CLBLM_R_X103Y123_SLICE_X162Y123_AO6;
  assign RIOI3_X105Y127_OLOGIC_X1Y128_TQ = 1'b1;
  assign RIOI3_X105Y127_OLOGIC_X1Y127_OQ = CLBLL_R_X57Y113_SLICE_X86Y113_AO6;
  assign RIOI3_X105Y127_OLOGIC_X1Y127_TQ = 1'b1;
  assign RIOI3_X105Y129_OLOGIC_X1Y130_OQ = CLBLM_R_X101Y123_SLICE_X158Y123_BO6;
  assign RIOI3_X105Y129_OLOGIC_X1Y130_TQ = 1'b1;
  assign RIOI3_X105Y129_OLOGIC_X1Y129_OQ = CLBLM_R_X103Y123_SLICE_X162Y123_BO6;
  assign RIOI3_X105Y129_OLOGIC_X1Y129_TQ = 1'b1;
  assign RIOI3_X105Y133_OLOGIC_X1Y134_OQ = CLBLM_R_X101Y118_SLICE_X158Y118_BO6;
  assign RIOI3_X105Y133_OLOGIC_X1Y134_TQ = 1'b1;
  assign RIOI3_X105Y133_OLOGIC_X1Y133_OQ = CLBLM_R_X101Y123_SLICE_X158Y123_CO6;
  assign RIOI3_X105Y133_OLOGIC_X1Y133_TQ = 1'b1;
  assign RIOI3_X105Y135_OLOGIC_X1Y136_OQ = CLBLM_R_X101Y118_SLICE_X158Y118_CO6;
  assign RIOI3_X105Y135_OLOGIC_X1Y136_TQ = 1'b1;
  assign RIOI3_X105Y135_OLOGIC_X1Y135_OQ = CLBLM_R_X101Y119_SLICE_X158Y119_CO6;
  assign RIOI3_X105Y135_OLOGIC_X1Y135_TQ = 1'b1;
  assign RIOI3_X105Y139_OLOGIC_X1Y140_OQ = CLBLM_R_X101Y118_SLICE_X158Y118_DO6;
  assign RIOI3_X105Y139_OLOGIC_X1Y140_TQ = 1'b1;
  assign RIOI3_X105Y139_OLOGIC_X1Y139_OQ = CLBLM_R_X101Y119_SLICE_X158Y119_DO6;
  assign RIOI3_X105Y139_OLOGIC_X1Y139_TQ = 1'b1;
  assign RIOI3_X105Y141_OLOGIC_X1Y142_OQ = CLBLM_R_X103Y123_SLICE_X162Y123_DO6;
  assign RIOI3_X105Y141_OLOGIC_X1Y142_TQ = 1'b1;
  assign RIOI3_X105Y141_OLOGIC_X1Y141_OQ = CLBLM_R_X101Y123_SLICE_X159Y123_BO6;
  assign RIOI3_X105Y141_OLOGIC_X1Y141_TQ = 1'b1;
  assign RIOI3_X105Y145_OLOGIC_X1Y146_OQ = CLBLL_L_X100Y123_SLICE_X156Y123_AO5;
  assign RIOI3_X105Y145_OLOGIC_X1Y146_TQ = 1'b1;
  assign RIOI3_X105Y145_OLOGIC_X1Y145_OQ = CLBLL_L_X100Y123_SLICE_X156Y123_BO5;
  assign RIOI3_X105Y145_OLOGIC_X1Y145_TQ = 1'b1;
  assign RIOI3_X105Y147_OLOGIC_X1Y148_OQ = CLBLM_R_X103Y122_SLICE_X163Y122_DO5;
  assign RIOI3_X105Y147_OLOGIC_X1Y148_TQ = 1'b1;
  assign RIOI3_X105Y147_OLOGIC_X1Y147_OQ = CLBLM_R_X103Y122_SLICE_X163Y122_CO5;
  assign RIOI3_X105Y147_OLOGIC_X1Y147_TQ = 1'b1;
  assign RIOI3_X105Y151_ILOGIC_X1Y152_O = RIOB33_X105Y151_IOB_X1Y152_I;
  assign RIOI3_X105Y151_ILOGIC_X1Y151_O = RIOB33_X105Y151_IOB_X1Y151_I;
  assign RIOI3_X105Y153_ILOGIC_X1Y154_O = RIOB33_X105Y153_IOB_X1Y154_I;
  assign RIOI3_X105Y153_ILOGIC_X1Y153_O = RIOB33_X105Y153_IOB_X1Y153_I;
  assign RIOI3_X105Y155_ILOGIC_X1Y156_O = RIOB33_X105Y155_IOB_X1Y156_I;
  assign RIOI3_X105Y155_ILOGIC_X1Y155_O = RIOB33_X105Y155_IOB_X1Y155_I;
  assign RIOI3_X105Y159_ILOGIC_X1Y160_O = RIOB33_X105Y159_IOB_X1Y160_I;
  assign RIOI3_X105Y159_ILOGIC_X1Y159_O = RIOB33_X105Y159_IOB_X1Y159_I;
  assign RIOI3_X105Y161_ILOGIC_X1Y161_O = RIOB33_X105Y161_IOB_X1Y161_I;
  assign RIOI3_X105Y165_ILOGIC_X1Y166_O = RIOB33_X105Y165_IOB_X1Y166_I;
  assign RIOI3_X105Y165_ILOGIC_X1Y165_O = RIOB33_X105Y165_IOB_X1Y165_I;
  assign RIOI3_X105Y167_ILOGIC_X1Y168_O = RIOB33_X105Y167_IOB_X1Y168_I;
  assign RIOI3_X105Y167_ILOGIC_X1Y167_O = RIOB33_X105Y167_IOB_X1Y167_I;
  assign RIOI3_X105Y171_ILOGIC_X1Y172_O = RIOB33_X105Y171_IOB_X1Y172_I;
  assign RIOI3_X105Y171_ILOGIC_X1Y171_O = RIOB33_X105Y171_IOB_X1Y171_I;
  assign RIOI3_X105Y173_OLOGIC_X1Y174_OQ = LIOB33_X0Y133_IOB_X0Y133_I;
  assign RIOI3_X105Y173_OLOGIC_X1Y174_TQ = 1'b1;
  assign RIOI3_X105Y173_OLOGIC_X1Y173_OQ = CLBLM_R_X103Y147_SLICE_X163Y147_AO5;
  assign RIOI3_X105Y173_OLOGIC_X1Y173_TQ = 1'b1;
  assign RIOI3_X105Y175_OLOGIC_X1Y176_OQ = LIOB33_X0Y137_IOB_X0Y138_I;
  assign RIOI3_X105Y175_OLOGIC_X1Y176_TQ = 1'b1;
  assign RIOI3_X105Y175_OLOGIC_X1Y175_OQ = LIOB33_X0Y103_IOB_X0Y104_I;
  assign RIOI3_X105Y175_OLOGIC_X1Y175_TQ = 1'b1;
  assign RIOI3_X105Y177_OLOGIC_X1Y178_OQ = CLBLM_R_X103Y177_SLICE_X163Y177_AO6;
  assign RIOI3_X105Y177_OLOGIC_X1Y178_TQ = 1'b1;
  assign RIOI3_X105Y177_OLOGIC_X1Y177_OQ = LIOB33_X0Y137_IOB_X0Y137_I;
  assign RIOI3_X105Y177_OLOGIC_X1Y177_TQ = 1'b1;
  assign RIOI3_X105Y179_OLOGIC_X1Y180_OQ = CLBLL_L_X2Y146_SLICE_X1Y146_AO5;
  assign RIOI3_X105Y179_OLOGIC_X1Y180_TQ = 1'b1;
  assign RIOI3_X105Y179_OLOGIC_X1Y179_OQ = CLBLM_R_X103Y147_SLICE_X163Y147_AO6;
  assign RIOI3_X105Y179_OLOGIC_X1Y179_TQ = 1'b1;
  assign RIOI3_X105Y183_OLOGIC_X1Y184_OQ = RIOB33_SING_X105Y150_IOB_X1Y150_I;
  assign RIOI3_X105Y183_OLOGIC_X1Y184_TQ = 1'b1;
  assign RIOI3_X105Y183_OLOGIC_X1Y183_OQ = RIOB33_X105Y107_IOB_X1Y107_I;
  assign RIOI3_X105Y183_OLOGIC_X1Y183_TQ = 1'b1;
  assign RIOI3_X105Y185_OLOGIC_X1Y186_OQ = LIOB33_X0Y85_IOB_X0Y85_I;
  assign RIOI3_X105Y185_OLOGIC_X1Y186_TQ = 1'b1;
  assign RIOI3_X105Y185_OLOGIC_X1Y185_OQ = LIOB33_X0Y133_IOB_X0Y134_I;
  assign RIOI3_X105Y185_OLOGIC_X1Y185_TQ = 1'b1;
  assign RIOI3_X105Y189_OLOGIC_X1Y190_OQ = CLBLM_R_X103Y177_SLICE_X163Y177_AO5;
  assign RIOI3_X105Y189_OLOGIC_X1Y190_TQ = 1'b1;
  assign RIOI3_X105Y189_OLOGIC_X1Y189_OQ = CLBLL_L_X2Y173_SLICE_X1Y173_AO5;
  assign RIOI3_X105Y189_OLOGIC_X1Y189_TQ = 1'b1;
  assign RIOI3_X105Y191_OLOGIC_X1Y192_OQ = CLBLM_R_X103Y177_SLICE_X163Y177_AO5;
  assign RIOI3_X105Y191_OLOGIC_X1Y192_TQ = 1'b1;
  assign RIOI3_X105Y191_OLOGIC_X1Y191_OQ = CLBLM_R_X103Y177_SLICE_X163Y177_AO5;
  assign RIOI3_X105Y191_OLOGIC_X1Y191_TQ = 1'b1;
  assign RIOI3_X105Y195_OLOGIC_X1Y196_OQ = CLBLL_L_X2Y173_SLICE_X0Y173_AO6;
  assign RIOI3_X105Y195_OLOGIC_X1Y196_TQ = 1'b1;
  assign RIOI3_X105Y195_OLOGIC_X1Y195_OQ = LIOB33_X0Y85_IOB_X0Y85_I;
  assign RIOI3_X105Y195_OLOGIC_X1Y195_TQ = 1'b1;
  assign RIOI3_X105Y197_OLOGIC_X1Y198_OQ = CLBLL_L_X2Y173_SLICE_X1Y173_AO6;
  assign RIOI3_X105Y197_OLOGIC_X1Y198_TQ = 1'b1;
  assign RIOI3_X105Y197_OLOGIC_X1Y197_OQ = CLBLL_L_X2Y173_SLICE_X1Y173_AO6;
  assign RIOI3_X105Y197_OLOGIC_X1Y197_TQ = 1'b1;
  assign RIOI3_SING_X105Y50_OLOGIC_X1Y50_OQ = CLBLM_R_X49Y95_SLICE_X74Y95_AO6;
  assign RIOI3_SING_X105Y50_OLOGIC_X1Y50_TQ = 1'b1;
  assign RIOI3_SING_X105Y99_OLOGIC_X1Y99_OQ = CLBLM_R_X101Y119_SLICE_X158Y119_BO6;
  assign RIOI3_SING_X105Y99_OLOGIC_X1Y99_TQ = 1'b1;
  assign RIOI3_SING_X105Y100_ILOGIC_X1Y100_O = RIOB33_SING_X105Y100_IOB_X1Y100_I;
  assign RIOI3_SING_X105Y149_OLOGIC_X1Y149_OQ = CLBLL_L_X4Y110_SLICE_X4Y110_CO6;
  assign RIOI3_SING_X105Y149_OLOGIC_X1Y149_TQ = 1'b1;
  assign RIOI3_SING_X105Y150_ILOGIC_X1Y150_O = RIOB33_SING_X105Y150_IOB_X1Y150_I;
  assign RIOI3_SING_X105Y199_OLOGIC_X1Y199_OQ = CLBLL_L_X2Y173_SLICE_X1Y173_BO5;
  assign RIOI3_SING_X105Y199_OLOGIC_X1Y199_TQ = 1'b1;
  assign RIOI3_TBYTESRC_X105Y57_OLOGIC_X1Y58_OQ = CLBLL_L_X100Y121_SLICE_X156Y121_AO6;
  assign RIOI3_TBYTESRC_X105Y57_OLOGIC_X1Y58_TQ = 1'b1;
  assign RIOI3_TBYTESRC_X105Y57_OLOGIC_X1Y57_OQ = CLBLM_R_X49Y95_SLICE_X74Y95_AO5;
  assign RIOI3_TBYTESRC_X105Y57_OLOGIC_X1Y57_TQ = 1'b1;
  assign RIOI3_TBYTESRC_X105Y69_OLOGIC_X1Y70_OQ = CLBLM_L_X8Y113_SLICE_X11Y113_CO6;
  assign RIOI3_TBYTESRC_X105Y69_OLOGIC_X1Y70_TQ = 1'b1;
  assign RIOI3_TBYTESRC_X105Y69_OLOGIC_X1Y69_OQ = CLBLM_R_X5Y111_SLICE_X6Y111_CO6;
  assign RIOI3_TBYTESRC_X105Y69_OLOGIC_X1Y69_TQ = 1'b1;
  assign RIOI3_TBYTESRC_X105Y81_OLOGIC_X1Y82_OQ = CLBLM_R_X103Y107_SLICE_X163Y107_BO6;
  assign RIOI3_TBYTESRC_X105Y81_OLOGIC_X1Y82_TQ = 1'b1;
  assign RIOI3_TBYTESRC_X105Y81_OLOGIC_X1Y81_OQ = CLBLM_R_X103Y122_SLICE_X163Y122_CO6;
  assign RIOI3_TBYTESRC_X105Y81_OLOGIC_X1Y81_TQ = 1'b1;
  assign RIOI3_TBYTESRC_X105Y93_OLOGIC_X1Y94_OQ = CLBLL_L_X4Y109_SLICE_X4Y109_AO5;
  assign RIOI3_TBYTESRC_X105Y93_OLOGIC_X1Y94_TQ = 1'b1;
  assign RIOI3_TBYTESRC_X105Y93_OLOGIC_X1Y93_OQ = CLBLM_L_X10Y113_SLICE_X13Y113_BO6;
  assign RIOI3_TBYTESRC_X105Y93_OLOGIC_X1Y93_TQ = 1'b1;
  assign RIOI3_TBYTESRC_X105Y107_ILOGIC_X1Y108_O = RIOB33_X105Y107_IOB_X1Y108_I;
  assign RIOI3_TBYTESRC_X105Y107_ILOGIC_X1Y107_O = RIOB33_X105Y107_IOB_X1Y107_I;
  assign RIOI3_TBYTESRC_X105Y119_ILOGIC_X1Y120_O = RIOB33_X105Y119_IOB_X1Y120_I;
  assign RIOI3_TBYTESRC_X105Y119_ILOGIC_X1Y119_O = RIOB33_X105Y119_IOB_X1Y119_I;
  assign RIOI3_TBYTESRC_X105Y131_OLOGIC_X1Y132_OQ = CLBLM_R_X101Y119_SLICE_X158Y119_AO6;
  assign RIOI3_TBYTESRC_X105Y131_OLOGIC_X1Y132_TQ = 1'b1;
  assign RIOI3_TBYTESRC_X105Y131_OLOGIC_X1Y131_OQ = CLBLM_R_X101Y118_SLICE_X158Y118_AO6;
  assign RIOI3_TBYTESRC_X105Y131_OLOGIC_X1Y131_TQ = 1'b1;
  assign RIOI3_TBYTESRC_X105Y143_OLOGIC_X1Y144_OQ = CLBLM_L_X10Y123_SLICE_X12Y123_AO6;
  assign RIOI3_TBYTESRC_X105Y143_OLOGIC_X1Y144_TQ = 1'b1;
  assign RIOI3_TBYTESRC_X105Y143_OLOGIC_X1Y143_OQ = CLBLM_L_X10Y123_SLICE_X12Y123_AO6;
  assign RIOI3_TBYTESRC_X105Y143_OLOGIC_X1Y143_TQ = 1'b1;
  assign RIOI3_TBYTESRC_X105Y157_ILOGIC_X1Y158_O = RIOB33_X105Y157_IOB_X1Y158_I;
  assign RIOI3_TBYTESRC_X105Y157_ILOGIC_X1Y157_O = RIOB33_X105Y157_IOB_X1Y157_I;
  assign RIOI3_TBYTESRC_X105Y169_ILOGIC_X1Y170_O = RIOB33_X105Y169_IOB_X1Y170_I;
  assign RIOI3_TBYTESRC_X105Y169_ILOGIC_X1Y169_O = RIOB33_X105Y169_IOB_X1Y169_I;
  assign RIOI3_TBYTESRC_X105Y181_OLOGIC_X1Y182_OQ = RIOB33_X105Y103_IOB_X1Y104_I;
  assign RIOI3_TBYTESRC_X105Y181_OLOGIC_X1Y182_TQ = 1'b1;
  assign RIOI3_TBYTESRC_X105Y181_OLOGIC_X1Y181_OQ = CLBLL_L_X2Y136_SLICE_X0Y136_BO6;
  assign RIOI3_TBYTESRC_X105Y181_OLOGIC_X1Y181_TQ = 1'b1;
  assign RIOI3_TBYTESRC_X105Y193_OLOGIC_X1Y194_OQ = CLBLM_R_X103Y193_SLICE_X163Y193_AO6;
  assign RIOI3_TBYTESRC_X105Y193_OLOGIC_X1Y194_TQ = 1'b1;
  assign RIOI3_TBYTESRC_X105Y193_OLOGIC_X1Y193_OQ = CLBLM_R_X103Y177_SLICE_X163Y177_AO5;
  assign RIOI3_TBYTESRC_X105Y193_OLOGIC_X1Y193_TQ = 1'b1;
  assign RIOI3_TBYTETERM_X105Y63_OLOGIC_X1Y64_OQ = CLBLM_R_X5Y113_SLICE_X6Y113_CO6;
  assign RIOI3_TBYTETERM_X105Y63_OLOGIC_X1Y64_TQ = 1'b1;
  assign RIOI3_TBYTETERM_X105Y63_OLOGIC_X1Y63_OQ = CLBLM_R_X5Y111_SLICE_X6Y111_BO6;
  assign RIOI3_TBYTETERM_X105Y63_OLOGIC_X1Y63_TQ = 1'b1;
  assign RIOI3_TBYTETERM_X105Y87_OLOGIC_X1Y88_OQ = CLBLM_L_X8Y113_SLICE_X10Y113_BO6;
  assign RIOI3_TBYTETERM_X105Y87_OLOGIC_X1Y88_TQ = 1'b1;
  assign RIOI3_TBYTETERM_X105Y87_OLOGIC_X1Y87_OQ = CLBLM_R_X103Y102_SLICE_X163Y102_BO6;
  assign RIOI3_TBYTETERM_X105Y87_OLOGIC_X1Y87_TQ = 1'b1;
  assign RIOI3_TBYTETERM_X105Y113_ILOGIC_X1Y114_O = RIOB33_X105Y113_IOB_X1Y114_I;
  assign RIOI3_TBYTETERM_X105Y113_ILOGIC_X1Y113_O = RIOB33_X105Y113_IOB_X1Y113_I;
  assign RIOI3_TBYTETERM_X105Y137_OLOGIC_X1Y138_OQ = CLBLM_R_X103Y123_SLICE_X162Y123_CO6;
  assign RIOI3_TBYTETERM_X105Y137_OLOGIC_X1Y138_TQ = 1'b1;
  assign RIOI3_TBYTETERM_X105Y137_OLOGIC_X1Y137_OQ = CLBLM_R_X101Y123_SLICE_X159Y123_AO6;
  assign RIOI3_TBYTETERM_X105Y137_OLOGIC_X1Y137_TQ = 1'b1;
  assign RIOI3_TBYTETERM_X105Y163_ILOGIC_X1Y163_O = RIOB33_X105Y163_IOB_X1Y163_I;
  assign RIOI3_TBYTETERM_X105Y187_OLOGIC_X1Y188_OQ = CLBLL_L_X2Y146_SLICE_X1Y146_AO6;
  assign RIOI3_TBYTETERM_X105Y187_OLOGIC_X1Y188_TQ = 1'b1;
  assign RIOI3_TBYTETERM_X105Y187_OLOGIC_X1Y187_OQ = CLBLM_R_X103Y185_SLICE_X163Y185_AO6;
  assign RIOI3_TBYTETERM_X105Y187_OLOGIC_X1Y187_TQ = 1'b1;
  assign CLBLM_R_X103Y102_SLICE_X162Y102_C2 = 1'b1;
  assign RIOB33_X105Y175_IOB_X1Y175_O = LIOB33_X0Y103_IOB_X0Y104_I;
  assign RIOB33_X105Y175_IOB_X1Y176_O = LIOB33_X0Y137_IOB_X0Y138_I;
  assign CLBLM_R_X103Y102_SLICE_X162Y102_C3 = 1'b1;
  assign RIOB33_SING_X105Y149_IOB_X1Y149_O = CLBLL_L_X4Y110_SLICE_X4Y110_CO6;
  assign CLBLM_R_X103Y102_SLICE_X162Y102_C4 = 1'b1;
  assign CLBLM_R_X103Y97_SLICE_X163Y97_C2 = 1'b1;
  assign CLBLM_R_X103Y97_SLICE_X163Y97_C3 = 1'b1;
  assign CLBLM_R_X103Y97_SLICE_X163Y97_C4 = 1'b1;
  assign LIOI3_SING_X0Y150_ILOGIC_X0Y150_D = LIOB33_SING_X0Y150_IOB_X0Y150_I;
  assign CLBLM_R_X103Y97_SLICE_X163Y97_C5 = 1'b1;
  assign CLBLM_R_X103Y97_SLICE_X163Y97_C6 = 1'b1;
  assign LIOI3_X0Y185_OLOGIC_X0Y186_D1 = LIOB33_X0Y135_IOB_X0Y135_I;
  assign LIOI3_X0Y185_OLOGIC_X0Y186_T1 = 1'b1;
  assign CLBLM_R_X103Y102_SLICE_X162Y102_D2 = 1'b1;
  assign CLBLM_R_X7Y113_SLICE_X9Y113_A1 = CLBLM_R_X5Y113_SLICE_X7Y113_DO6;
  assign CLBLM_R_X7Y113_SLICE_X9Y113_A2 = CLBLM_R_X5Y112_SLICE_X7Y112_AO6;
  assign CLBLM_R_X7Y113_SLICE_X9Y113_A3 = CLBLL_L_X4Y141_SLICE_X4Y141_AO6;
  assign CLBLM_R_X7Y113_SLICE_X9Y113_A4 = CLBLM_R_X7Y113_SLICE_X9Y113_BO6;
  assign CLBLM_R_X7Y113_SLICE_X9Y113_A5 = CLBLM_R_X7Y113_SLICE_X8Y113_BO5;
  assign CLBLM_R_X7Y113_SLICE_X9Y113_A6 = CLBLM_R_X7Y113_SLICE_X9Y113_CO6;
  assign CLBLM_R_X103Y97_SLICE_X163Y97_D1 = 1'b1;
  assign CLBLM_R_X7Y113_SLICE_X9Y113_B1 = LIOB33_X0Y101_IOB_X0Y101_I;
  assign CLBLM_R_X7Y113_SLICE_X9Y113_B2 = LIOB33_X0Y159_IOB_X0Y159_I;
  assign CLBLM_R_X7Y113_SLICE_X9Y113_B3 = LIOB33_SING_X0Y99_IOB_X0Y99_I;
  assign CLBLM_R_X7Y113_SLICE_X9Y113_B4 = LIOB33_X0Y131_IOB_X0Y131_I;
  assign CLBLM_R_X7Y113_SLICE_X9Y113_B5 = LIOB33_X0Y159_IOB_X0Y160_I;
  assign CLBLM_R_X7Y113_SLICE_X9Y113_B6 = LIOB33_X0Y129_IOB_X0Y129_I;
  assign CLBLM_R_X103Y97_SLICE_X163Y97_D2 = 1'b1;
  assign LIOI3_X0Y185_OLOGIC_X0Y185_D1 = LIOB33_X0Y67_IOB_X0Y67_I;
  assign CLBLM_R_X7Y113_SLICE_X9Y113_C1 = LIOB33_X0Y83_IOB_X0Y84_I;
  assign CLBLM_R_X7Y113_SLICE_X9Y113_C2 = LIOB33_X0Y71_IOB_X0Y71_I;
  assign CLBLM_R_X7Y113_SLICE_X9Y113_C3 = LIOB33_X0Y65_IOB_X0Y66_I;
  assign CLBLM_R_X7Y113_SLICE_X9Y113_C4 = 1'b1;
  assign CLBLM_R_X7Y113_SLICE_X9Y113_C5 = 1'b1;
  assign CLBLM_R_X7Y113_SLICE_X9Y113_C6 = 1'b1;
  assign CLBLM_R_X103Y97_SLICE_X163Y97_D4 = 1'b1;
  assign CLBLM_R_X103Y97_SLICE_X163Y97_D5 = 1'b1;
  assign LIOI3_X0Y185_OLOGIC_X0Y185_T1 = 1'b1;
  assign RIOI3_X105Y139_OLOGIC_X1Y140_D1 = CLBLM_R_X101Y118_SLICE_X158Y118_DO6;
  assign CLBLM_R_X103Y97_SLICE_X163Y97_D6 = 1'b1;
  assign CLBLM_R_X7Y113_SLICE_X9Y113_D1 = 1'b1;
  assign CLBLM_R_X7Y113_SLICE_X9Y113_D2 = 1'b1;
  assign CLBLM_R_X7Y113_SLICE_X9Y113_D3 = 1'b1;
  assign CLBLM_R_X7Y113_SLICE_X9Y113_D4 = 1'b1;
  assign CLBLM_R_X7Y113_SLICE_X9Y113_D5 = 1'b1;
  assign CLBLM_R_X7Y113_SLICE_X9Y113_D6 = 1'b1;
  assign RIOI3_X105Y77_OLOGIC_X1Y78_D1 = CLBLL_L_X100Y113_SLICE_X156Y113_BO6;
  assign RIOI3_X105Y139_OLOGIC_X1Y140_T1 = 1'b1;
  assign CLBLM_R_X7Y113_SLICE_X8Y113_A1 = CLBLM_R_X7Y114_SLICE_X8Y114_CO6;
  assign CLBLM_R_X7Y113_SLICE_X8Y113_A2 = LIOB33_SING_X0Y99_IOB_X0Y99_I;
  assign CLBLM_R_X7Y113_SLICE_X8Y113_A3 = LIOB33_X0Y95_IOB_X0Y95_I;
  assign CLBLM_R_X7Y113_SLICE_X8Y113_A4 = LIOB33_X0Y129_IOB_X0Y129_I;
  assign CLBLM_R_X7Y113_SLICE_X8Y113_A5 = LIOB33_SING_X0Y100_IOB_X0Y100_I;
  assign CLBLM_R_X7Y113_SLICE_X8Y113_A6 = 1'b1;
  assign RIOI3_X105Y77_OLOGIC_X1Y78_T1 = 1'b1;
  assign RIOI3_X105Y139_OLOGIC_X1Y139_D1 = CLBLM_R_X101Y119_SLICE_X158Y119_DO6;
  assign CLBLM_R_X7Y113_SLICE_X8Y113_B1 = LIOB33_X0Y69_IOB_X0Y70_I;
  assign CLBLM_R_X7Y113_SLICE_X8Y113_B2 = LIOB33_X0Y85_IOB_X0Y86_I;
  assign CLBLM_R_X7Y113_SLICE_X8Y113_B3 = LIOB33_X0Y123_IOB_X0Y123_I;
  assign CLBLM_R_X7Y113_SLICE_X8Y113_B4 = LIOB33_X0Y67_IOB_X0Y68_I;
  assign CLBLM_R_X7Y113_SLICE_X8Y113_B5 = LIOB33_X0Y87_IOB_X0Y88_I;
  assign CLBLM_R_X7Y113_SLICE_X8Y113_B6 = 1'b1;
  assign RIOI3_X105Y77_OLOGIC_X1Y77_D1 = CLBLL_L_X36Y113_SLICE_X54Y113_BO6;
  assign RIOI3_X105Y139_OLOGIC_X1Y139_T1 = 1'b1;
  assign RIOI3_TBYTETERM_X105Y137_OLOGIC_X1Y138_D1 = CLBLM_R_X103Y123_SLICE_X162Y123_CO6;
  assign CLBLM_R_X7Y113_SLICE_X8Y113_C1 = LIOB33_SING_X0Y100_IOB_X0Y100_I;
  assign CLBLM_R_X7Y113_SLICE_X8Y113_C2 = LIOB33_SING_X0Y99_IOB_X0Y99_I;
  assign CLBLM_R_X7Y113_SLICE_X8Y113_C3 = LIOB33_X0Y95_IOB_X0Y95_I;
  assign CLBLM_R_X7Y113_SLICE_X8Y113_C4 = CLBLM_R_X7Y114_SLICE_X8Y114_CO6;
  assign CLBLM_R_X7Y113_SLICE_X8Y113_C5 = LIOB33_X0Y127_IOB_X0Y127_I;
  assign CLBLM_R_X7Y113_SLICE_X8Y113_C6 = LIOB33_X0Y129_IOB_X0Y129_I;
  assign RIOI3_X105Y77_OLOGIC_X1Y77_T1 = 1'b1;
  assign RIOI3_TBYTESRC_X105Y181_OLOGIC_X1Y182_D1 = RIOB33_X105Y103_IOB_X1Y104_I;
  assign RIOI3_TBYTETERM_X105Y137_OLOGIC_X1Y138_T1 = 1'b1;
  assign CLBLM_R_X103Y185_SLICE_X163Y185_B1 = 1'b1;
  assign CLBLM_R_X103Y123_SLICE_X163Y123_D4 = 1'b1;
  assign CLBLM_R_X7Y113_SLICE_X8Y113_D1 = LIOB33_X0Y87_IOB_X0Y88_I;
  assign CLBLM_R_X7Y113_SLICE_X8Y113_D2 = LIOB33_X0Y89_IOB_X0Y90_I;
  assign CLBLM_R_X7Y113_SLICE_X8Y113_D3 = 1'b1;
  assign CLBLM_R_X7Y113_SLICE_X8Y113_D4 = CLBLM_R_X5Y113_SLICE_X6Y113_AO6;
  assign CLBLM_R_X7Y113_SLICE_X8Y113_D5 = LIOB33_X0Y95_IOB_X0Y95_I;
  assign CLBLM_R_X7Y113_SLICE_X8Y113_D6 = LIOB33_X0Y123_IOB_X0Y123_I;
  assign CLBLM_R_X103Y185_SLICE_X163Y185_B2 = 1'b1;
  assign CLBLM_R_X103Y185_SLICE_X163Y185_B3 = 1'b1;
  assign RIOI3_TBYTETERM_X105Y137_OLOGIC_X1Y137_D1 = CLBLM_R_X101Y123_SLICE_X159Y123_AO6;
  assign CLBLM_R_X103Y185_SLICE_X163Y185_B4 = 1'b1;
  assign RIOI3_TBYTESRC_X105Y181_OLOGIC_X1Y181_D1 = CLBLL_L_X2Y136_SLICE_X0Y136_BO6;
  assign CLBLM_R_X103Y123_SLICE_X163Y123_A6 = 1'b1;
  assign CLBLM_R_X103Y185_SLICE_X163Y185_B5 = 1'b1;
  assign RIOI3_TBYTETERM_X105Y137_OLOGIC_X1Y137_T1 = 1'b1;
  assign CLBLM_R_X103Y185_SLICE_X163Y185_B6 = 1'b1;
  assign RIOI3_TBYTESRC_X105Y181_OLOGIC_X1Y181_T1 = 1'b1;
  assign CLBLM_R_X103Y123_SLICE_X163Y123_D5 = 1'b1;
  assign RIOB33_X105Y57_IOB_X1Y58_O = CLBLL_L_X100Y121_SLICE_X156Y121_AO6;
  assign RIOB33_X105Y57_IOB_X1Y57_O = CLBLM_R_X49Y95_SLICE_X74Y95_AO5;
  assign CLBLM_R_X103Y123_SLICE_X163Y123_B2 = 1'b1;
  assign CLBLM_R_X103Y185_SLICE_X163Y185_C1 = 1'b1;
  assign CLBLM_R_X103Y185_SLICE_X162Y185_A1 = 1'b1;
  assign CLBLM_R_X103Y123_SLICE_X163Y123_D6 = 1'b1;
  assign CLBLM_R_X103Y123_SLICE_X163Y123_B3 = 1'b1;
  assign CLBLM_R_X103Y185_SLICE_X163Y185_C2 = 1'b1;
  assign CLBLM_R_X103Y123_SLICE_X163Y123_B4 = 1'b1;
  assign CLBLM_R_X103Y185_SLICE_X163Y185_C3 = 1'b1;
  assign CLBLM_R_X103Y123_SLICE_X163Y123_B5 = 1'b1;
  assign CLBLM_R_X103Y185_SLICE_X163Y185_C4 = 1'b1;
  assign CLBLM_R_X103Y123_SLICE_X163Y123_B6 = 1'b1;
  assign CLBLM_R_X103Y185_SLICE_X163Y185_C5 = 1'b1;
  assign CLBLM_R_X103Y185_SLICE_X163Y185_C6 = 1'b1;
  assign CLBLM_R_X103Y185_SLICE_X162Y185_A2 = 1'b1;
  assign CLBLM_R_X103Y123_SLICE_X163Y123_C1 = 1'b1;
  assign CLBLM_R_X103Y123_SLICE_X163Y123_C2 = 1'b1;
  assign CLBLM_R_X103Y185_SLICE_X162Y185_A3 = 1'b1;
  assign CLBLM_R_X103Y123_SLICE_X163Y123_C3 = 1'b1;
  assign CLBLM_R_X103Y123_SLICE_X163Y123_C4 = 1'b1;
  assign CLBLM_R_X103Y123_SLICE_X163Y123_C5 = 1'b1;
  assign LIOI3_X0Y155_ILOGIC_X0Y156_D = LIOB33_X0Y155_IOB_X0Y156_I;
  assign CLBLM_R_X103Y123_SLICE_X163Y123_C6 = 1'b1;
  assign LIOI3_X0Y155_ILOGIC_X0Y155_D = LIOB33_X0Y155_IOB_X0Y155_I;
  assign RIOB33_X105Y177_IOB_X1Y178_O = CLBLM_R_X103Y177_SLICE_X163Y177_AO6;
  assign RIOB33_X105Y177_IOB_X1Y177_O = LIOB33_X0Y137_IOB_X0Y137_I;
  assign LIOI3_X0Y125_ILOGIC_X0Y126_D = LIOB33_X0Y125_IOB_X0Y126_I;
  assign LIOI3_SING_X0Y199_OLOGIC_X0Y199_D1 = CLBLL_L_X4Y111_SLICE_X5Y111_CO6;
  assign CLBLM_R_X103Y185_SLICE_X163Y185_D1 = 1'b1;
  assign CLBLM_R_X103Y185_SLICE_X162Y185_A4 = 1'b1;
  assign LIOI3_X0Y125_ILOGIC_X0Y125_D = LIOB33_X0Y125_IOB_X0Y125_I;
  assign RIOB33_SING_X105Y199_IOB_X1Y199_O = CLBLL_L_X2Y173_SLICE_X1Y173_BO5;
  assign CLBLM_R_X103Y185_SLICE_X163Y185_D2 = 1'b1;
  assign LIOI3_X0Y95_ILOGIC_X0Y96_D = LIOB33_X0Y95_IOB_X0Y96_I;
  assign CLBLM_R_X103Y185_SLICE_X163Y185_D3 = 1'b1;
  assign LIOI3_X0Y95_ILOGIC_X0Y95_D = LIOB33_X0Y95_IOB_X0Y95_I;
  assign LIOI3_SING_X0Y199_OLOGIC_X0Y199_T1 = 1'b1;
  assign RIOI3_X105Y171_ILOGIC_X1Y172_D = RIOB33_X105Y171_IOB_X1Y172_I;
  assign LIOI3_X0Y65_ILOGIC_X0Y66_D = LIOB33_X0Y65_IOB_X0Y66_I;
  assign CLBLM_R_X103Y185_SLICE_X163Y185_D4 = 1'b1;
  assign RIOI3_X105Y171_ILOGIC_X1Y171_D = RIOB33_X105Y171_IOB_X1Y171_I;
  assign LIOI3_X0Y65_ILOGIC_X0Y65_D = LIOB33_X0Y65_IOB_X0Y65_I;
  assign CLBLM_R_X103Y185_SLICE_X163Y185_D5 = 1'b1;
  assign CLBLM_R_X103Y185_SLICE_X163Y185_D6 = 1'b1;
  assign CLBLM_R_X103Y185_SLICE_X162Y185_A5 = 1'b1;
  assign RIOI3_X105Y109_ILOGIC_X1Y110_D = RIOB33_X105Y109_IOB_X1Y110_I;
  assign CLBLM_R_X103Y185_SLICE_X163Y185_A1 = LIOB33_X0Y133_IOB_X0Y134_I;
  assign CLBLM_R_X103Y185_SLICE_X163Y185_A2 = 1'b1;
  assign CLBLM_R_X103Y185_SLICE_X163Y185_A3 = 1'b1;
  assign CLBLM_R_X103Y185_SLICE_X163Y185_A4 = 1'b1;
  assign CLBLM_R_X103Y185_SLICE_X163Y185_A5 = 1'b1;
  assign CLBLM_R_X103Y107_SLICE_X163Y107_A1 = RIOB33_X105Y111_IOB_X1Y111_I;
  assign CLBLM_R_X103Y107_SLICE_X163Y107_A2 = CLBLM_R_X103Y122_SLICE_X163Y122_BO5;
  assign CLBLM_R_X103Y107_SLICE_X163Y107_A3 = CLBLM_L_X8Y113_SLICE_X11Y113_BO6;
  assign CLBLM_R_X103Y107_SLICE_X163Y107_A4 = CLBLM_R_X5Y111_SLICE_X7Y111_CO6;
  assign CLBLM_R_X103Y107_SLICE_X163Y107_A5 = RIOB33_X105Y111_IOB_X1Y112_I;
  assign CLBLM_R_X103Y107_SLICE_X163Y107_A6 = 1'b1;
  assign CLBLM_R_X103Y123_SLICE_X163Y123_D1 = 1'b1;
  assign CLBLM_R_X103Y185_SLICE_X163Y185_A6 = 1'b1;
  assign CLBLM_R_X103Y107_SLICE_X163Y107_B1 = RIOB33_X105Y111_IOB_X1Y111_I;
  assign CLBLM_R_X103Y107_SLICE_X163Y107_B2 = 1'b1;
  assign CLBLM_R_X103Y107_SLICE_X163Y107_B3 = CLBLM_L_X8Y113_SLICE_X11Y113_BO6;
  assign CLBLM_R_X103Y107_SLICE_X163Y107_B4 = CLBLM_R_X5Y111_SLICE_X7Y111_CO6;
  assign CLBLM_R_X103Y107_SLICE_X163Y107_B5 = RIOB33_X105Y111_IOB_X1Y112_I;
  assign CLBLM_R_X103Y107_SLICE_X163Y107_B6 = CLBLM_R_X103Y122_SLICE_X163Y122_AO5;
  assign CLBLM_R_X103Y123_SLICE_X163Y123_D2 = 1'b1;
  assign CLBLM_R_X103Y123_SLICE_X163Y123_D3 = 1'b1;
  assign CLBLM_R_X101Y123_SLICE_X159Y123_A1 = CLBLM_R_X5Y111_SLICE_X6Y111_AO6;
  assign CLBLM_R_X101Y123_SLICE_X159Y123_A2 = CLBLM_R_X103Y122_SLICE_X163Y122_AO5;
  assign CLBLM_R_X101Y123_SLICE_X159Y123_A3 = CLBLM_R_X101Y123_SLICE_X158Y123_AO5;
  assign CLBLM_R_X101Y123_SLICE_X159Y123_A4 = CLBLM_L_X10Y123_SLICE_X12Y123_AO6;
  assign CLBLM_R_X101Y123_SLICE_X159Y123_A5 = CLBLM_R_X25Y116_SLICE_X36Y116_AO5;
  assign CLBLM_R_X101Y123_SLICE_X159Y123_A6 = CLBLM_R_X3Y111_SLICE_X2Y111_AO5;
  assign CLBLM_R_X103Y107_SLICE_X163Y107_C1 = 1'b1;
  assign CLBLM_R_X103Y107_SLICE_X163Y107_C2 = 1'b1;
  assign CLBLM_R_X101Y123_SLICE_X159Y123_B1 = CLBLM_R_X5Y111_SLICE_X6Y111_AO6;
  assign CLBLM_R_X101Y123_SLICE_X159Y123_B2 = CLBLM_L_X10Y123_SLICE_X12Y123_AO6;
  assign CLBLM_R_X101Y123_SLICE_X159Y123_B3 = CLBLM_R_X103Y122_SLICE_X163Y122_BO5;
  assign CLBLM_R_X101Y123_SLICE_X159Y123_B4 = CLBLM_R_X101Y123_SLICE_X158Y123_AO5;
  assign CLBLM_R_X101Y123_SLICE_X159Y123_B5 = CLBLM_R_X25Y116_SLICE_X36Y116_AO5;
  assign CLBLM_R_X101Y123_SLICE_X159Y123_B6 = CLBLM_R_X3Y111_SLICE_X2Y111_AO5;
  assign CLBLM_R_X103Y107_SLICE_X163Y107_C6 = 1'b1;
  assign CLBLM_R_X103Y97_SLICE_X162Y97_D5 = 1'b1;
  assign CLBLM_R_X101Y123_SLICE_X159Y123_C1 = 1'b1;
  assign CLBLM_R_X101Y123_SLICE_X159Y123_C2 = 1'b1;
  assign CLBLM_R_X101Y123_SLICE_X159Y123_C3 = 1'b1;
  assign CLBLM_R_X101Y123_SLICE_X159Y123_C4 = 1'b1;
  assign CLBLM_R_X101Y123_SLICE_X159Y123_C5 = 1'b1;
  assign CLBLM_R_X101Y123_SLICE_X159Y123_C6 = 1'b1;
  assign CLBLM_R_X103Y97_SLICE_X162Y97_D6 = 1'b1;
  assign CLBLM_R_X103Y107_SLICE_X163Y107_D2 = 1'b1;
  assign CLBLM_R_X103Y107_SLICE_X163Y107_D3 = 1'b1;
  assign CLBLM_R_X103Y107_SLICE_X163Y107_D4 = 1'b1;
  assign CLBLM_R_X103Y107_SLICE_X162Y107_A1 = 1'b1;
  assign CLBLM_R_X103Y107_SLICE_X162Y107_A2 = 1'b1;
  assign CLBLM_R_X103Y107_SLICE_X162Y107_A3 = 1'b1;
  assign CLBLM_R_X103Y107_SLICE_X162Y107_A4 = 1'b1;
  assign CLBLM_R_X101Y123_SLICE_X159Y123_D1 = 1'b1;
  assign CLBLM_R_X101Y123_SLICE_X159Y123_D2 = 1'b1;
  assign CLBLM_R_X101Y123_SLICE_X159Y123_D3 = 1'b1;
  assign CLBLM_R_X101Y123_SLICE_X159Y123_D4 = 1'b1;
  assign CLBLM_R_X101Y123_SLICE_X159Y123_D5 = 1'b1;
  assign CLBLM_R_X101Y123_SLICE_X159Y123_D6 = 1'b1;
  assign CLBLM_R_X103Y107_SLICE_X162Y107_A5 = 1'b1;
  assign CLBLM_R_X103Y107_SLICE_X162Y107_B1 = 1'b1;
  assign CLBLM_R_X103Y107_SLICE_X162Y107_B2 = 1'b1;
  assign CLBLM_R_X101Y123_SLICE_X158Y123_A1 = LIOB33_X0Y123_IOB_X0Y124_I;
  assign CLBLM_R_X101Y123_SLICE_X158Y123_A2 = RIOB33_X105Y115_IOB_X1Y115_I;
  assign CLBLM_R_X101Y123_SLICE_X158Y123_A3 = LIOB33_X0Y121_IOB_X0Y121_I;
  assign CLBLM_R_X7Y114_SLICE_X9Y114_A1 = LIOB33_X0Y131_IOB_X0Y131_I;
  assign CLBLM_R_X7Y114_SLICE_X9Y114_A2 = LIOB33_X0Y101_IOB_X0Y101_I;
  assign CLBLM_R_X7Y114_SLICE_X9Y114_A3 = 1'b1;
  assign CLBLM_R_X7Y114_SLICE_X9Y114_A4 = LIOB33_X0Y151_IOB_X0Y151_I;
  assign CLBLM_R_X7Y114_SLICE_X9Y114_A5 = 1'b1;
  assign CLBLM_R_X7Y114_SLICE_X9Y114_A6 = LIOB33_SING_X0Y150_IOB_X0Y150_I;
  assign CLBLM_R_X101Y123_SLICE_X158Y123_A4 = CLBLM_L_X10Y113_SLICE_X12Y113_CO6;
  assign CLBLM_R_X101Y123_SLICE_X158Y123_A5 = RIOB33_X105Y125_IOB_X1Y126_I;
  assign CLBLM_R_X101Y123_SLICE_X158Y123_A6 = 1'b1;
  assign CLBLM_R_X7Y114_SLICE_X9Y114_B1 = 1'b1;
  assign CLBLM_R_X7Y114_SLICE_X9Y114_B2 = 1'b1;
  assign CLBLM_R_X7Y114_SLICE_X9Y114_B3 = 1'b1;
  assign CLBLM_R_X7Y114_SLICE_X9Y114_B4 = 1'b1;
  assign CLBLM_R_X7Y114_SLICE_X9Y114_B5 = 1'b1;
  assign CLBLM_R_X7Y114_SLICE_X9Y114_B6 = 1'b1;
  assign CLBLM_R_X101Y123_SLICE_X158Y123_B1 = CLBLM_R_X5Y111_SLICE_X6Y111_AO6;
  assign CLBLM_R_X101Y123_SLICE_X158Y123_B2 = CLBLM_L_X10Y123_SLICE_X12Y123_AO6;
  assign CLBLM_R_X101Y123_SLICE_X158Y123_B3 = CLBLL_L_X100Y123_SLICE_X156Y123_BO6;
  assign CLBLM_R_X7Y114_SLICE_X9Y114_C1 = 1'b1;
  assign CLBLM_R_X7Y114_SLICE_X9Y114_C2 = 1'b1;
  assign CLBLM_R_X7Y114_SLICE_X9Y114_C3 = 1'b1;
  assign CLBLM_R_X7Y114_SLICE_X9Y114_C4 = 1'b1;
  assign CLBLM_R_X7Y114_SLICE_X9Y114_C5 = 1'b1;
  assign CLBLM_R_X7Y114_SLICE_X9Y114_C6 = 1'b1;
  assign CLBLM_R_X101Y123_SLICE_X158Y123_C1 = CLBLM_R_X101Y123_SLICE_X158Y123_AO6;
  assign CLBLM_R_X101Y123_SLICE_X158Y123_C2 = CLBLM_L_X10Y123_SLICE_X12Y123_AO6;
  assign CLBLM_R_X101Y123_SLICE_X158Y123_C3 = CLBLM_R_X5Y111_SLICE_X6Y111_AO6;
  assign CLBLM_R_X101Y123_SLICE_X158Y123_C4 = CLBLM_R_X25Y116_SLICE_X36Y116_AO5;
  assign CLBLM_R_X101Y123_SLICE_X158Y123_C5 = CLBLL_L_X100Y123_SLICE_X156Y123_AO6;
  assign CLBLM_R_X101Y123_SLICE_X158Y123_C6 = CLBLM_R_X3Y111_SLICE_X2Y111_AO5;
  assign CLBLM_R_X7Y114_SLICE_X9Y114_D1 = 1'b1;
  assign CLBLM_R_X7Y114_SLICE_X9Y114_D2 = 1'b1;
  assign CLBLM_R_X7Y114_SLICE_X9Y114_D3 = 1'b1;
  assign CLBLM_R_X7Y114_SLICE_X9Y114_D4 = 1'b1;
  assign CLBLM_R_X7Y114_SLICE_X9Y114_D5 = 1'b1;
  assign CLBLM_R_X7Y114_SLICE_X9Y114_D6 = 1'b1;
  assign CLBLM_R_X101Y123_SLICE_X158Y123_D1 = 1'b1;
  assign CLBLM_R_X101Y123_SLICE_X158Y123_D2 = 1'b1;
  assign CLBLM_R_X101Y123_SLICE_X158Y123_D3 = 1'b1;
  assign CLBLM_R_X101Y123_SLICE_X158Y123_D4 = 1'b1;
  assign CLBLM_R_X101Y123_SLICE_X158Y123_D5 = 1'b1;
  assign CLBLM_R_X101Y123_SLICE_X158Y123_D6 = 1'b1;
  assign CLBLM_R_X7Y114_SLICE_X8Y114_A1 = LIOB33_X0Y69_IOB_X0Y70_I;
  assign CLBLM_R_X7Y114_SLICE_X8Y114_A2 = RIOB33_X105Y159_IOB_X1Y160_I;
  assign CLBLM_R_X7Y114_SLICE_X8Y114_A3 = LIOB33_X0Y123_IOB_X0Y123_I;
  assign CLBLM_R_X7Y114_SLICE_X8Y114_A4 = LIOB33_X0Y87_IOB_X0Y88_I;
  assign CLBLM_R_X7Y114_SLICE_X8Y114_A5 = LIOB33_X0Y67_IOB_X0Y68_I;
  assign CLBLM_R_X7Y114_SLICE_X8Y114_A6 = 1'b1;
  assign CLBLM_R_X103Y123_SLICE_X162Y123_B1 = CLBLL_L_X4Y111_SLICE_X5Y111_AO5;
  assign CLBLM_R_X7Y114_SLICE_X8Y114_B1 = LIOB33_X0Y95_IOB_X0Y95_I;
  assign CLBLM_R_X7Y114_SLICE_X8Y114_B2 = LIOB33_X0Y131_IOB_X0Y131_I;
  assign CLBLM_R_X7Y114_SLICE_X8Y114_B3 = LIOB33_X0Y101_IOB_X0Y102_I;
  assign CLBLM_R_X7Y114_SLICE_X8Y114_B4 = LIOB33_X0Y101_IOB_X0Y101_I;
  assign CLBLM_R_X7Y114_SLICE_X8Y114_B5 = 1'b1;
  assign CLBLM_R_X7Y114_SLICE_X8Y114_B6 = 1'b1;
  assign CLBLM_R_X103Y123_SLICE_X162Y123_B2 = CLBLM_L_X10Y123_SLICE_X12Y123_AO6;
  assign CLBLM_R_X103Y123_SLICE_X162Y123_B3 = CLBLM_R_X103Y123_SLICE_X163Y123_AO6;
  assign CLBLM_R_X103Y123_SLICE_X162Y123_A3 = CLBLM_R_X103Y123_SLICE_X163Y123_AO6;
  assign CLBLM_R_X7Y114_SLICE_X8Y114_C1 = LIOB33_X0Y103_IOB_X0Y103_I;
  assign CLBLM_R_X7Y114_SLICE_X8Y114_C2 = LIOB33_X0Y131_IOB_X0Y131_I;
  assign CLBLM_R_X7Y114_SLICE_X8Y114_C3 = LIOB33_X0Y95_IOB_X0Y95_I;
  assign CLBLM_R_X7Y114_SLICE_X8Y114_C4 = LIOB33_X0Y103_IOB_X0Y104_I;
  assign CLBLM_R_X7Y114_SLICE_X8Y114_C5 = LIOB33_X0Y131_IOB_X0Y132_I;
  assign CLBLM_R_X7Y114_SLICE_X8Y114_C6 = CLBLM_R_X7Y114_SLICE_X8Y114_BO6;
  assign CLBLM_R_X103Y123_SLICE_X162Y123_B4 = CLBLM_R_X5Y111_SLICE_X6Y111_AO6;
  assign CLBLM_R_X103Y123_SLICE_X162Y123_B5 = CLBLM_R_X5Y114_SLICE_X7Y114_AO6;
  assign CLBLM_R_X103Y185_SLICE_X162Y185_C2 = 1'b1;
  assign CLBLM_R_X103Y185_SLICE_X162Y185_C3 = 1'b1;
  assign CLBLM_R_X103Y123_SLICE_X162Y123_B6 = CLBLL_L_X100Y123_SLICE_X156Y123_BO6;
  assign CLBLM_R_X103Y185_SLICE_X162Y185_C4 = 1'b1;
  assign RIOB33_X105Y59_IOB_X1Y59_O = CLBLM_R_X5Y113_SLICE_X6Y113_BO6;
  assign CLBLM_R_X7Y114_SLICE_X8Y114_D1 = 1'b1;
  assign CLBLM_R_X7Y114_SLICE_X8Y114_D2 = 1'b1;
  assign CLBLM_R_X7Y114_SLICE_X8Y114_D3 = 1'b1;
  assign CLBLM_R_X7Y114_SLICE_X8Y114_D4 = 1'b1;
  assign CLBLM_R_X7Y114_SLICE_X8Y114_D5 = 1'b1;
  assign CLBLM_R_X7Y114_SLICE_X8Y114_D6 = 1'b1;
  assign CLBLM_R_X5Y111_SLICE_X6Y111_B6 = CLBLM_R_X3Y111_SLICE_X3Y111_CO6;
  assign CLBLM_R_X103Y185_SLICE_X162Y185_C5 = 1'b1;
  assign CLBLM_R_X103Y123_SLICE_X162Y123_A4 = CLBLM_R_X5Y111_SLICE_X6Y111_AO6;
  assign CLBLM_R_X103Y185_SLICE_X162Y185_C6 = 1'b1;
  assign CLBLM_R_X103Y185_SLICE_X162Y185_B1 = 1'b1;
  assign CLBLM_R_X103Y123_SLICE_X162Y123_C1 = CLBLM_R_X5Y114_SLICE_X7Y114_AO6;
  assign CLBLM_R_X103Y123_SLICE_X162Y123_A5 = CLBLM_R_X5Y114_SLICE_X7Y114_AO6;
  assign CLBLM_R_X103Y185_SLICE_X162Y185_B2 = 1'b1;
  assign CLBLM_R_X103Y123_SLICE_X162Y123_C6 = CLBLM_L_X10Y123_SLICE_X12Y123_AO6;
  assign CLBLM_R_X103Y123_SLICE_X162Y123_A6 = CLBLL_L_X100Y123_SLICE_X156Y123_AO6;
  assign CLBLM_R_X103Y185_SLICE_X162Y185_B3 = 1'b1;
  assign CLBLM_R_X103Y185_SLICE_X162Y185_D1 = 1'b1;
  assign CLBLM_R_X103Y185_SLICE_X162Y185_D2 = 1'b1;
  assign CLBLM_R_X103Y185_SLICE_X162Y185_D3 = 1'b1;
  assign CLBLM_R_X103Y185_SLICE_X162Y185_D4 = 1'b1;
  assign CLBLM_R_X103Y185_SLICE_X162Y185_D5 = 1'b1;
  assign RIOB33_X105Y179_IOB_X1Y180_O = CLBLL_L_X2Y146_SLICE_X1Y146_AO5;
  assign RIOB33_X105Y179_IOB_X1Y179_O = CLBLM_R_X103Y147_SLICE_X163Y147_AO6;
  assign CLBLM_R_X103Y185_SLICE_X162Y185_B4 = 1'b1;
  assign CLBLM_R_X103Y185_SLICE_X162Y185_D6 = 1'b1;
  assign LIOB33_X0Y187_IOB_X0Y188_O = CLBLL_L_X2Y173_SLICE_X1Y173_BO6;
  assign LIOB33_X0Y187_IOB_X0Y187_O = CLBLL_L_X2Y173_SLICE_X1Y173_BO6;
  assign CLBLM_R_X103Y123_SLICE_X162Y123_D2 = CLBLM_R_X103Y123_SLICE_X163Y123_AO5;
  assign CLBLM_R_X103Y185_SLICE_X162Y185_B5 = 1'b1;
  assign CLBLM_R_X103Y123_SLICE_X162Y123_D3 = CLBLL_L_X4Y111_SLICE_X5Y111_AO5;
  assign CLBLM_R_X103Y123_SLICE_X162Y123_D4 = CLBLM_R_X103Y122_SLICE_X163Y122_BO5;
  assign CLBLM_R_X103Y123_SLICE_X162Y123_D5 = CLBLM_R_X5Y111_SLICE_X6Y111_AO6;
  assign CLBLM_R_X103Y123_SLICE_X162Y123_D6 = CLBLM_L_X10Y123_SLICE_X12Y123_AO6;
  assign CLBLM_R_X103Y185_SLICE_X162Y185_B6 = 1'b1;
  assign CLBLM_R_X103Y108_SLICE_X163Y108_A1 = 1'b1;
  assign CLBLM_R_X103Y108_SLICE_X163Y108_A2 = RIOB33_X105Y107_IOB_X1Y107_I;
  assign CLBLM_R_X103Y108_SLICE_X163Y108_A3 = 1'b1;
  assign CLBLM_R_X103Y108_SLICE_X163Y108_A4 = RIOB33_X105Y107_IOB_X1Y108_I;
  assign CLBLM_R_X103Y108_SLICE_X163Y108_A5 = 1'b1;
  assign CLBLM_R_X103Y108_SLICE_X163Y108_A6 = 1'b1;
  assign LIOI3_SING_X0Y200_OLOGIC_X0Y200_D1 = LIOB33_SING_X0Y100_IOB_X0Y100_I;
  assign CLBLM_R_X103Y108_SLICE_X163Y108_B1 = 1'b1;
  assign CLBLM_R_X103Y108_SLICE_X163Y108_B2 = 1'b1;
  assign CLBLM_R_X103Y108_SLICE_X163Y108_B3 = 1'b1;
  assign CLBLM_R_X103Y108_SLICE_X163Y108_B4 = 1'b1;
  assign CLBLM_R_X103Y108_SLICE_X163Y108_B5 = 1'b1;
  assign CLBLM_R_X103Y108_SLICE_X163Y108_B6 = 1'b1;
  assign LIOI3_SING_X0Y200_OLOGIC_X0Y200_T1 = 1'b1;
  assign CLBLM_R_X103Y108_SLICE_X163Y108_C1 = 1'b1;
  assign CLBLM_R_X103Y108_SLICE_X163Y108_C2 = 1'b1;
  assign CLBLM_R_X103Y108_SLICE_X163Y108_C3 = 1'b1;
  assign CLBLM_R_X103Y108_SLICE_X163Y108_C4 = 1'b1;
  assign CLBLM_R_X103Y108_SLICE_X163Y108_C5 = 1'b1;
  assign CLBLM_R_X103Y108_SLICE_X163Y108_C6 = 1'b1;
  assign CLBLM_R_X103Y108_SLICE_X163Y108_D1 = 1'b1;
  assign CLBLM_R_X103Y108_SLICE_X163Y108_D2 = 1'b1;
  assign CLBLM_R_X103Y108_SLICE_X163Y108_D3 = 1'b1;
  assign CLBLM_R_X103Y108_SLICE_X163Y108_D4 = 1'b1;
  assign CLBLM_R_X103Y108_SLICE_X163Y108_D5 = 1'b1;
  assign CLBLM_R_X103Y108_SLICE_X163Y108_D6 = 1'b1;
  assign CLBLM_R_X103Y108_SLICE_X162Y108_A1 = 1'b1;
  assign CLBLM_R_X103Y108_SLICE_X162Y108_A2 = 1'b1;
  assign CLBLM_R_X103Y108_SLICE_X162Y108_A3 = 1'b1;
  assign CLBLM_R_X103Y108_SLICE_X162Y108_A4 = 1'b1;
  assign CLBLM_R_X103Y108_SLICE_X162Y108_A5 = 1'b1;
  assign CLBLM_R_X103Y108_SLICE_X162Y108_A6 = 1'b1;
  assign RIOI3_X105Y67_OLOGIC_X1Y67_T1 = 1'b1;
  assign CLBLM_R_X103Y108_SLICE_X162Y108_B1 = 1'b1;
  assign CLBLM_R_X103Y108_SLICE_X162Y108_B2 = 1'b1;
  assign CLBLM_R_X103Y108_SLICE_X162Y108_B3 = 1'b1;
  assign CLBLM_R_X103Y108_SLICE_X162Y108_B4 = 1'b1;
  assign CLBLM_R_X103Y108_SLICE_X162Y108_B5 = 1'b1;
  assign CLBLM_R_X103Y108_SLICE_X162Y108_B6 = 1'b1;
  assign CLBLM_R_X103Y108_SLICE_X162Y108_C1 = 1'b1;
  assign CLBLM_R_X103Y108_SLICE_X162Y108_C2 = 1'b1;
  assign CLBLM_R_X103Y108_SLICE_X162Y108_C3 = 1'b1;
  assign CLBLM_R_X103Y108_SLICE_X162Y108_C4 = 1'b1;
  assign CLBLM_R_X103Y108_SLICE_X162Y108_C5 = 1'b1;
  assign CLBLM_R_X103Y108_SLICE_X162Y108_C6 = 1'b1;
  assign CLBLL_L_X2Y175_SLICE_X0Y175_A3 = LIOB33_X0Y137_IOB_X0Y138_I;
  assign CLBLM_R_X103Y108_SLICE_X162Y108_D1 = 1'b1;
  assign CLBLM_R_X103Y108_SLICE_X162Y108_D2 = 1'b1;
  assign CLBLM_R_X103Y108_SLICE_X162Y108_D3 = 1'b1;
  assign CLBLM_R_X103Y108_SLICE_X162Y108_D4 = 1'b1;
  assign CLBLM_R_X103Y108_SLICE_X162Y108_D5 = 1'b1;
  assign CLBLM_R_X103Y108_SLICE_X162Y108_D6 = 1'b1;
  assign CLBLL_L_X2Y175_SLICE_X0Y175_B1 = 1'b1;
  assign RIOB33_X105Y61_IOB_X1Y62_O = CLBLL_L_X100Y121_SLICE_X156Y121_BO6;
  assign RIOB33_X105Y61_IOB_X1Y61_O = CLBLM_L_X8Y113_SLICE_X11Y113_BO6;
  assign CLBLL_L_X2Y175_SLICE_X0Y175_B2 = 1'b1;
  assign CLBLM_R_X103Y185_SLICE_X162Y185_C1 = 1'b1;
  assign CLBLL_L_X2Y175_SLICE_X0Y175_B3 = 1'b1;
  assign CLBLL_L_X2Y175_SLICE_X0Y175_B4 = 1'b1;
  assign CLBLL_L_X2Y175_SLICE_X0Y175_B5 = 1'b1;
  assign RIOB33_X105Y85_IOB_X1Y86_O = CLBLM_R_X103Y107_SLICE_X163Y107_AO6;
  assign RIOB33_X105Y85_IOB_X1Y85_O = CLBLM_R_X103Y122_SLICE_X163Y122_DO6;
  assign LIOI3_X0Y189_OLOGIC_X0Y190_D1 = CLBLL_L_X2Y173_SLICE_X1Y173_BO6;
  assign LIOI3_X0Y189_OLOGIC_X0Y190_T1 = 1'b1;
  assign LIOI3_X0Y189_OLOGIC_X0Y189_D1 = CLBLL_L_X2Y173_SLICE_X1Y173_BO6;
  assign RIOI3_X105Y173_OLOGIC_X1Y174_D1 = LIOB33_X0Y133_IOB_X0Y133_I;
  assign LIOI3_X0Y189_OLOGIC_X0Y189_T1 = 1'b1;
  assign RIOI3_X105Y141_OLOGIC_X1Y142_D1 = CLBLM_R_X103Y123_SLICE_X162Y123_DO6;
  assign RIOB33_X105Y181_IOB_X1Y182_O = RIOB33_X105Y103_IOB_X1Y104_I;
  assign RIOB33_X105Y181_IOB_X1Y181_O = CLBLL_L_X2Y136_SLICE_X0Y136_BO6;
  assign RIOI3_X105Y173_OLOGIC_X1Y174_T1 = 1'b1;
  assign RIOI3_X105Y141_OLOGIC_X1Y142_T1 = 1'b1;
  assign RIOI3_X105Y79_OLOGIC_X1Y80_D1 = CLBLM_R_X103Y97_SLICE_X163Y97_AO6;
  assign RIOI3_X105Y173_OLOGIC_X1Y173_D1 = CLBLM_R_X103Y147_SLICE_X163Y147_AO5;
  assign CLBLL_L_X36Y113_SLICE_X54Y113_A1 = LIOB33_X0Y165_IOB_X0Y166_I;
  assign CLBLL_L_X36Y113_SLICE_X54Y113_A2 = CLBLM_R_X5Y113_SLICE_X6Y113_CO6;
  assign CLBLL_L_X36Y113_SLICE_X54Y113_A3 = LIOB33_X0Y51_IOB_X0Y51_I;
  assign CLBLL_L_X36Y113_SLICE_X54Y113_A4 = CLBLM_L_X10Y113_SLICE_X12Y113_BO6;
  assign CLBLL_L_X36Y113_SLICE_X54Y113_A5 = LIOB33_X0Y153_IOB_X0Y154_I;
  assign CLBLL_L_X36Y113_SLICE_X54Y113_A6 = LIOB33_X0Y155_IOB_X0Y156_I;
  assign RIOI3_X105Y51_OLOGIC_X1Y52_D1 = CLBLM_R_X49Y95_SLICE_X74Y95_AO6;
  assign RIOI3_X105Y79_OLOGIC_X1Y80_T1 = 1'b1;
  assign RIOI3_X105Y141_OLOGIC_X1Y141_D1 = CLBLM_R_X101Y123_SLICE_X159Y123_BO6;
  assign CLBLL_L_X36Y113_SLICE_X54Y113_B1 = LIOB33_X0Y157_IOB_X0Y157_I;
  assign CLBLL_L_X36Y113_SLICE_X54Y113_B2 = CLBLM_L_X10Y113_SLICE_X12Y113_BO6;
  assign CLBLL_L_X36Y113_SLICE_X54Y113_B3 = CLBLM_R_X5Y113_SLICE_X6Y113_CO6;
  assign CLBLL_L_X36Y113_SLICE_X54Y113_B4 = LIOB33_X0Y51_IOB_X0Y51_I;
  assign CLBLL_L_X36Y113_SLICE_X54Y113_B5 = LIOB33_X0Y157_IOB_X0Y158_I;
  assign CLBLL_L_X36Y113_SLICE_X54Y113_B6 = LIOB33_X0Y165_IOB_X0Y166_I;
  assign RIOI3_X105Y51_OLOGIC_X1Y52_T1 = 1'b1;
  assign RIOI3_X105Y79_OLOGIC_X1Y79_D1 = CLBLM_R_X29Y115_SLICE_X42Y115_BO6;
  assign RIOI3_X105Y141_OLOGIC_X1Y141_T1 = 1'b1;
  assign CLBLL_L_X36Y113_SLICE_X54Y113_C1 = 1'b1;
  assign CLBLL_L_X36Y113_SLICE_X54Y113_C2 = 1'b1;
  assign CLBLL_L_X36Y113_SLICE_X54Y113_C3 = 1'b1;
  assign CLBLL_L_X36Y113_SLICE_X54Y113_C4 = 1'b1;
  assign CLBLL_L_X36Y113_SLICE_X54Y113_C5 = 1'b1;
  assign CLBLL_L_X36Y113_SLICE_X54Y113_C6 = 1'b1;
  assign RIOI3_X105Y51_OLOGIC_X1Y51_D1 = CLBLL_L_X4Y111_SLICE_X5Y111_CO6;
  assign RIOI3_TBYTESRC_X105Y193_OLOGIC_X1Y194_D1 = CLBLM_R_X103Y193_SLICE_X163Y193_AO6;
  assign RIOI3_X105Y79_OLOGIC_X1Y79_T1 = 1'b1;
  assign RIOI3_TBYTESRC_X105Y57_OLOGIC_X1Y58_D1 = CLBLL_L_X100Y121_SLICE_X156Y121_AO6;
  assign CLBLL_L_X36Y113_SLICE_X54Y113_D1 = 1'b1;
  assign CLBLL_L_X36Y113_SLICE_X54Y113_D2 = 1'b1;
  assign CLBLL_L_X36Y113_SLICE_X54Y113_D3 = 1'b1;
  assign CLBLL_L_X36Y113_SLICE_X54Y113_D4 = 1'b1;
  assign CLBLL_L_X36Y113_SLICE_X54Y113_D5 = 1'b1;
  assign CLBLL_L_X36Y113_SLICE_X54Y113_D6 = 1'b1;
  assign RIOI3_X105Y51_OLOGIC_X1Y51_T1 = 1'b1;
  assign RIOI3_TBYTESRC_X105Y193_OLOGIC_X1Y194_T1 = 1'b1;
  assign RIOI3_TBYTESRC_X105Y57_OLOGIC_X1Y58_T1 = 1'b1;
  assign RIOI3_TBYTESRC_X105Y193_OLOGIC_X1Y193_D1 = CLBLM_R_X103Y177_SLICE_X163Y177_AO5;
  assign RIOI3_TBYTESRC_X105Y57_OLOGIC_X1Y57_D1 = CLBLM_R_X49Y95_SLICE_X74Y95_AO5;
  assign RIOI3_TBYTESRC_X105Y193_OLOGIC_X1Y193_T1 = 1'b1;
  assign RIOI3_TBYTESRC_X105Y57_OLOGIC_X1Y57_T1 = 1'b1;
  assign CLBLL_L_X36Y113_SLICE_X55Y113_A1 = 1'b1;
  assign CLBLL_L_X36Y113_SLICE_X55Y113_A2 = 1'b1;
  assign CLBLL_L_X36Y113_SLICE_X55Y113_A3 = 1'b1;
  assign CLBLL_L_X36Y113_SLICE_X55Y113_A4 = 1'b1;
  assign CLBLL_L_X36Y113_SLICE_X55Y113_A5 = 1'b1;
  assign CLBLL_L_X36Y113_SLICE_X55Y113_A6 = 1'b1;
  assign CLBLL_L_X36Y113_SLICE_X55Y113_B1 = 1'b1;
  assign CLBLL_L_X36Y113_SLICE_X55Y113_B2 = 1'b1;
  assign CLBLL_L_X36Y113_SLICE_X55Y113_B3 = 1'b1;
  assign CLBLL_L_X36Y113_SLICE_X55Y113_B4 = 1'b1;
  assign CLBLL_L_X36Y113_SLICE_X55Y113_B5 = 1'b1;
  assign CLBLL_L_X36Y113_SLICE_X55Y113_B6 = 1'b1;
  assign CLBLL_L_X36Y113_SLICE_X55Y113_C1 = 1'b1;
  assign CLBLL_L_X36Y113_SLICE_X55Y113_C2 = 1'b1;
  assign CLBLL_L_X36Y113_SLICE_X55Y113_C3 = 1'b1;
  assign CLBLL_L_X36Y113_SLICE_X55Y113_C4 = 1'b1;
  assign CLBLL_L_X36Y113_SLICE_X55Y113_C5 = 1'b1;
  assign CLBLL_L_X36Y113_SLICE_X55Y113_C6 = 1'b1;
  assign CLBLL_L_X36Y113_SLICE_X55Y113_D1 = 1'b1;
  assign CLBLL_L_X36Y113_SLICE_X55Y113_D2 = 1'b1;
  assign CLBLL_L_X36Y113_SLICE_X55Y113_D3 = 1'b1;
  assign CLBLL_L_X36Y113_SLICE_X55Y113_D4 = 1'b1;
  assign CLBLL_L_X36Y113_SLICE_X55Y113_D5 = 1'b1;
  assign CLBLL_L_X36Y113_SLICE_X55Y113_D6 = 1'b1;
  assign LIOI3_X0Y159_ILOGIC_X0Y160_D = LIOB33_X0Y159_IOB_X0Y160_I;
  assign LIOI3_X0Y159_ILOGIC_X0Y159_D = LIOB33_X0Y159_IOB_X0Y159_I;
  assign LIOI3_X0Y127_ILOGIC_X0Y128_D = LIOB33_X0Y127_IOB_X0Y128_I;
  assign LIOI3_X0Y127_ILOGIC_X0Y127_D = LIOB33_X0Y127_IOB_X0Y127_I;
  assign LIOI3_X0Y97_ILOGIC_X0Y98_D = LIOB33_X0Y97_IOB_X0Y98_I;
  assign LIOI3_X0Y97_ILOGIC_X0Y97_D = LIOB33_X0Y97_IOB_X0Y97_I;
  assign LIOI3_X0Y67_ILOGIC_X0Y68_D = LIOB33_X0Y67_IOB_X0Y68_I;
  assign RIOB33_X105Y63_IOB_X1Y64_O = CLBLM_R_X5Y113_SLICE_X6Y113_CO6;
  assign RIOB33_X105Y63_IOB_X1Y63_O = CLBLM_R_X5Y111_SLICE_X6Y111_BO6;
  assign RIOI3_SING_X105Y149_OLOGIC_X1Y149_T1 = 1'b1;
  assign LIOI3_X0Y67_ILOGIC_X0Y67_D = LIOB33_X0Y67_IOB_X0Y67_I;
  assign RIOI3_X105Y103_ILOGIC_X1Y104_D = RIOB33_X105Y103_IOB_X1Y104_I;
  assign RIOI3_X105Y111_ILOGIC_X1Y112_D = RIOB33_X105Y111_IOB_X1Y112_I;
  assign RIOI3_X105Y111_ILOGIC_X1Y111_D = RIOB33_X105Y111_IOB_X1Y111_I;
  assign RIOI3_X105Y103_ILOGIC_X1Y103_D = RIOB33_X105Y103_IOB_X1Y103_I;
  assign LIOI3_TBYTESRC_X0Y131_ILOGIC_X0Y132_D = LIOB33_X0Y131_IOB_X0Y132_I;
  assign CLBLM_R_X103Y147_SLICE_X163Y147_A5 = 1'b1;
  assign LIOI3_TBYTESRC_X0Y131_ILOGIC_X0Y131_D = LIOB33_X0Y131_IOB_X0Y131_I;
  assign RIOI3_TBYTETERM_X105Y163_ILOGIC_X1Y163_D = RIOB33_X105Y163_IOB_X1Y163_I;
  assign RIOB33_X105Y183_IOB_X1Y184_O = RIOB33_SING_X105Y150_IOB_X1Y150_I;
  assign RIOB33_X105Y183_IOB_X1Y183_O = RIOB33_X105Y107_IOB_X1Y107_I;
  assign CLBLM_R_X103Y147_SLICE_X163Y147_B2 = 1'b1;
  assign CLBLM_R_X103Y147_SLICE_X163Y147_B4 = 1'b1;
  assign RIOB33_X105Y65_IOB_X1Y66_O = CLBLM_R_X5Y112_SLICE_X6Y112_AO6;
  assign RIOB33_X105Y65_IOB_X1Y65_O = CLBLM_R_X103Y107_SLICE_X163Y107_AO5;
  assign RIOI3_TBYTESRC_X105Y107_ILOGIC_X1Y108_D = RIOB33_X105Y107_IOB_X1Y108_I;
  assign RIOI3_X105Y61_OLOGIC_X1Y61_T1 = 1'b1;
  assign RIOB33_X105Y185_IOB_X1Y186_O = LIOB33_X0Y85_IOB_X0Y85_I;
  assign RIOB33_X105Y185_IOB_X1Y185_O = LIOB33_X0Y133_IOB_X0Y134_I;
  assign RIOI3_X105Y165_ILOGIC_X1Y166_D = RIOB33_X105Y165_IOB_X1Y166_I;
  assign RIOI3_X105Y165_ILOGIC_X1Y165_D = RIOB33_X105Y165_IOB_X1Y165_I;
  assign LIOI3_X0Y191_OLOGIC_X0Y192_D1 = CLBLM_R_X5Y114_SLICE_X6Y114_AO6;
  assign LIOI3_X0Y191_OLOGIC_X0Y192_T1 = 1'b1;
  assign LIOI3_X0Y191_OLOGIC_X0Y191_D1 = CLBLM_R_X5Y113_SLICE_X7Y113_AO6;
  assign RIOI3_X105Y175_OLOGIC_X1Y176_D1 = LIOB33_X0Y137_IOB_X0Y138_I;
  assign LIOI3_X0Y191_OLOGIC_X0Y191_T1 = 1'b1;
  assign RIOI3_X105Y145_OLOGIC_X1Y146_D1 = CLBLL_L_X100Y123_SLICE_X156Y123_AO5;
  assign RIOI3_X105Y175_OLOGIC_X1Y176_T1 = 1'b1;
  assign RIOI3_X105Y145_OLOGIC_X1Y146_T1 = 1'b1;
  assign RIOI3_X105Y83_OLOGIC_X1Y84_D1 = CLBLM_R_X103Y97_SLICE_X163Y97_BO6;
  assign RIOI3_X105Y175_OLOGIC_X1Y175_D1 = LIOB33_X0Y103_IOB_X0Y104_I;
  assign RIOB33_X105Y67_IOB_X1Y68_O = CLBLL_L_X4Y109_SLICE_X4Y109_AO6;
  assign RIOB33_X105Y67_IOB_X1Y67_O = CLBLM_R_X5Y109_SLICE_X6Y109_AO6;
  assign RIOI3_X105Y53_OLOGIC_X1Y54_D1 = CLBLM_R_X103Y108_SLICE_X163Y108_AO6;
  assign RIOI3_X105Y145_OLOGIC_X1Y145_D1 = CLBLL_L_X100Y123_SLICE_X156Y123_BO5;
  assign RIOI3_X105Y83_OLOGIC_X1Y84_T1 = 1'b1;
  assign RIOI3_X105Y175_OLOGIC_X1Y175_T1 = 1'b1;
  assign RIOI3_X105Y53_OLOGIC_X1Y54_T1 = 1'b1;
  assign RIOI3_X105Y145_OLOGIC_X1Y145_T1 = 1'b1;
  assign RIOI3_X105Y83_OLOGIC_X1Y83_D1 = CLBLM_R_X103Y102_SLICE_X163Y102_AO6;
  assign RIOI3_TBYTETERM_X105Y187_OLOGIC_X1Y188_D1 = CLBLL_L_X2Y146_SLICE_X1Y146_AO6;
  assign RIOI3_X105Y53_OLOGIC_X1Y53_D1 = CLBLM_L_X10Y113_SLICE_X12Y113_AO6;
  assign RIOI3_X105Y83_OLOGIC_X1Y83_T1 = 1'b1;
  assign RIOI3_TBYTETERM_X105Y187_OLOGIC_X1Y188_T1 = 1'b1;
  assign RIOI3_TBYTESRC_X105Y69_OLOGIC_X1Y70_D1 = CLBLM_L_X8Y113_SLICE_X11Y113_CO6;
  assign RIOI3_X105Y53_OLOGIC_X1Y53_T1 = 1'b1;
  assign RIOI3_TBYTETERM_X105Y187_OLOGIC_X1Y187_D1 = CLBLM_R_X103Y185_SLICE_X163Y185_AO6;
  assign RIOB33_X105Y127_IOB_X1Y128_O = CLBLM_R_X103Y123_SLICE_X162Y123_AO6;
  assign RIOB33_X105Y127_IOB_X1Y127_O = CLBLL_R_X57Y113_SLICE_X86Y113_AO6;
  assign RIOI3_TBYTESRC_X105Y69_OLOGIC_X1Y70_T1 = 1'b1;
  assign RIOI3_TBYTETERM_X105Y187_OLOGIC_X1Y187_T1 = 1'b1;
  assign RIOI3_TBYTESRC_X105Y69_OLOGIC_X1Y69_D1 = CLBLM_R_X5Y111_SLICE_X6Y111_CO6;
  assign RIOI3_TBYTESRC_X105Y69_OLOGIC_X1Y69_T1 = 1'b1;
  assign RIOB33_X105Y187_IOB_X1Y188_O = CLBLL_L_X2Y146_SLICE_X1Y146_AO6;
  assign RIOB33_X105Y187_IOB_X1Y187_O = CLBLM_R_X103Y185_SLICE_X163Y185_AO6;
  assign CLBLM_R_X49Y101_SLICE_X75Y101_A1 = 1'b1;
  assign CLBLM_R_X49Y101_SLICE_X75Y101_A2 = 1'b1;
  assign CLBLM_R_X49Y101_SLICE_X75Y101_A3 = 1'b1;
  assign CLBLM_R_X49Y101_SLICE_X75Y101_A4 = 1'b1;
  assign CLBLM_R_X49Y101_SLICE_X75Y101_A5 = 1'b1;
  assign CLBLM_R_X49Y101_SLICE_X75Y101_A6 = 1'b1;
  assign LIOI3_X0Y161_ILOGIC_X0Y162_D = LIOB33_X0Y161_IOB_X0Y162_I;
  assign CLBLM_R_X49Y101_SLICE_X75Y101_B1 = 1'b1;
  assign CLBLM_R_X49Y101_SLICE_X75Y101_B2 = 1'b1;
  assign CLBLM_R_X49Y101_SLICE_X75Y101_B3 = 1'b1;
  assign CLBLM_R_X49Y101_SLICE_X75Y101_B4 = 1'b1;
  assign CLBLM_R_X49Y101_SLICE_X75Y101_B5 = 1'b1;
  assign CLBLM_R_X49Y101_SLICE_X75Y101_B6 = 1'b1;
  assign LIOI3_X0Y161_ILOGIC_X0Y161_D = LIOB33_X0Y161_IOB_X0Y161_I;
  assign LIOI3_X0Y129_ILOGIC_X0Y130_D = LIOB33_X0Y129_IOB_X0Y130_I;
  assign CLBLM_R_X49Y101_SLICE_X75Y101_C1 = 1'b1;
  assign CLBLM_R_X49Y101_SLICE_X75Y101_C2 = 1'b1;
  assign CLBLM_R_X49Y101_SLICE_X75Y101_C3 = 1'b1;
  assign CLBLM_R_X49Y101_SLICE_X75Y101_C4 = 1'b1;
  assign CLBLM_R_X49Y101_SLICE_X75Y101_C5 = 1'b1;
  assign CLBLM_R_X49Y101_SLICE_X75Y101_C6 = 1'b1;
  assign LIOI3_X0Y101_ILOGIC_X0Y102_D = LIOB33_X0Y101_IOB_X0Y102_I;
  assign LIOI3_X0Y129_ILOGIC_X0Y129_D = LIOB33_X0Y129_IOB_X0Y129_I;
  assign LIOI3_X0Y101_ILOGIC_X0Y101_D = LIOB33_X0Y101_IOB_X0Y101_I;
  assign CLBLL_R_X57Y113_SLICE_X86Y113_A4 = CLBLM_R_X5Y111_SLICE_X6Y111_BO6;
  assign CLBLM_R_X49Y101_SLICE_X75Y101_D1 = 1'b1;
  assign CLBLM_R_X49Y101_SLICE_X75Y101_D2 = 1'b1;
  assign CLBLM_R_X49Y101_SLICE_X75Y101_D3 = 1'b1;
  assign CLBLM_R_X49Y101_SLICE_X75Y101_D4 = 1'b1;
  assign CLBLM_R_X49Y101_SLICE_X75Y101_D5 = 1'b1;
  assign CLBLM_R_X49Y101_SLICE_X75Y101_D6 = 1'b1;
  assign LIOI3_X0Y71_ILOGIC_X0Y72_D = LIOB33_X0Y71_IOB_X0Y72_I;
  assign LIOI3_X0Y71_ILOGIC_X0Y71_D = LIOB33_X0Y71_IOB_X0Y71_I;
  assign CLBLM_R_X49Y101_SLICE_X74Y101_A1 = LIOB33_X0Y83_IOB_X0Y84_I;
  assign CLBLM_R_X49Y101_SLICE_X74Y101_A2 = RIOB33_X105Y101_IOB_X1Y101_I;
  assign CLBLM_R_X49Y101_SLICE_X74Y101_A3 = LIOB33_X0Y95_IOB_X0Y95_I;
  assign CLBLM_R_X49Y101_SLICE_X74Y101_A4 = LIOB33_X0Y85_IOB_X0Y85_I;
  assign CLBLM_R_X49Y101_SLICE_X74Y101_A5 = CLBLM_R_X5Y113_SLICE_X6Y113_AO6;
  assign CLBLM_R_X49Y101_SLICE_X74Y101_A6 = 1'b1;
  assign RIOI3_X105Y115_ILOGIC_X1Y116_D = RIOB33_X105Y115_IOB_X1Y116_I;
  assign RIOI3_X105Y115_ILOGIC_X1Y115_D = RIOB33_X105Y115_IOB_X1Y115_I;
  assign CLBLM_R_X49Y101_SLICE_X74Y101_B1 = 1'b1;
  assign CLBLM_R_X49Y101_SLICE_X74Y101_B2 = 1'b1;
  assign CLBLM_R_X49Y101_SLICE_X74Y101_B3 = 1'b1;
  assign CLBLM_R_X49Y101_SLICE_X74Y101_B4 = 1'b1;
  assign CLBLM_R_X49Y101_SLICE_X74Y101_B5 = 1'b1;
  assign CLBLM_R_X49Y101_SLICE_X74Y101_B6 = 1'b1;
  assign LIOI3_TBYTETERM_X0Y63_ILOGIC_X0Y63_D = LIOB33_X0Y63_IOB_X0Y63_I;
  assign LIOI3_TBYTESRC_X0Y143_ILOGIC_X0Y143_D = LIOB33_X0Y143_IOB_X0Y143_I;
  assign CLBLL_R_X57Y113_SLICE_X86Y113_B1 = LIOB33_X0Y157_IOB_X0Y158_I;
  assign CLBLM_R_X49Y101_SLICE_X74Y101_C1 = 1'b1;
  assign CLBLM_R_X49Y101_SLICE_X74Y101_C2 = 1'b1;
  assign CLBLM_R_X49Y101_SLICE_X74Y101_C3 = 1'b1;
  assign CLBLM_R_X49Y101_SLICE_X74Y101_C4 = 1'b1;
  assign CLBLL_R_X57Y113_SLICE_X86Y113_B2 = CLBLM_R_X5Y111_SLICE_X6Y111_BO6;
  assign CLBLM_R_X49Y101_SLICE_X74Y101_C5 = 1'b1;
  assign CLBLM_R_X49Y101_SLICE_X74Y101_C6 = 1'b1;
  assign CLBLM_R_X49Y101_SLICE_X74Y101_D1 = 1'b1;
  assign CLBLM_R_X49Y101_SLICE_X74Y101_D2 = 1'b1;
  assign CLBLM_R_X49Y101_SLICE_X74Y101_D3 = 1'b1;
  assign CLBLM_R_X49Y101_SLICE_X74Y101_D4 = 1'b1;
  assign CLBLL_R_X57Y113_SLICE_X86Y113_B5 = LIOB33_X0Y157_IOB_X0Y157_I;
  assign CLBLM_R_X49Y101_SLICE_X74Y101_D5 = 1'b1;
  assign CLBLM_R_X49Y101_SLICE_X74Y101_D6 = 1'b1;
  assign RIOB33_X105Y69_IOB_X1Y70_O = CLBLM_L_X8Y113_SLICE_X11Y113_CO6;
  assign RIOB33_X105Y69_IOB_X1Y69_O = CLBLM_R_X5Y111_SLICE_X6Y111_CO6;
  assign CLBLM_R_X103Y185_SLICE_X162Y185_A6 = 1'b1;
  assign RIOB33_X105Y129_IOB_X1Y130_O = CLBLM_R_X101Y123_SLICE_X158Y123_BO6;
  assign RIOB33_X105Y129_IOB_X1Y129_O = CLBLM_R_X103Y123_SLICE_X162Y123_BO6;
  assign RIOB33_X105Y189_IOB_X1Y190_O = CLBLM_R_X103Y177_SLICE_X163Y177_AO5;
  assign RIOB33_X105Y189_IOB_X1Y189_O = CLBLL_L_X2Y173_SLICE_X1Y173_AO5;
  assign CLBLM_R_X5Y109_SLICE_X7Y109_A1 = 1'b1;
  assign CLBLM_R_X5Y109_SLICE_X7Y109_A2 = 1'b1;
  assign CLBLM_R_X5Y109_SLICE_X7Y109_A3 = 1'b1;
  assign CLBLM_R_X5Y109_SLICE_X7Y109_A4 = 1'b1;
  assign CLBLM_R_X5Y109_SLICE_X7Y109_A5 = 1'b1;
  assign CLBLM_R_X5Y109_SLICE_X7Y109_A6 = 1'b1;
  assign CLBLM_R_X5Y109_SLICE_X7Y109_B1 = 1'b1;
  assign CLBLM_R_X5Y109_SLICE_X7Y109_B2 = 1'b1;
  assign CLBLM_R_X5Y109_SLICE_X7Y109_B3 = 1'b1;
  assign CLBLM_R_X5Y109_SLICE_X7Y109_B4 = 1'b1;
  assign CLBLM_R_X5Y109_SLICE_X7Y109_B5 = 1'b1;
  assign CLBLM_R_X5Y109_SLICE_X7Y109_B6 = 1'b1;
  assign LIOI3_X0Y59_ILOGIC_X0Y60_D = LIOB33_X0Y59_IOB_X0Y60_I;
  assign CLBLM_R_X5Y109_SLICE_X7Y109_C1 = 1'b1;
  assign CLBLM_R_X5Y109_SLICE_X7Y109_C2 = 1'b1;
  assign CLBLM_R_X5Y109_SLICE_X7Y109_C3 = 1'b1;
  assign CLBLM_R_X5Y109_SLICE_X7Y109_C4 = 1'b1;
  assign CLBLM_R_X5Y109_SLICE_X7Y109_C5 = 1'b1;
  assign CLBLM_R_X5Y109_SLICE_X7Y109_C6 = 1'b1;
  assign LIOI3_X0Y59_ILOGIC_X0Y59_D = LIOB33_X0Y59_IOB_X0Y59_I;
  assign CLBLM_R_X5Y109_SLICE_X7Y109_D1 = 1'b1;
  assign CLBLM_R_X5Y109_SLICE_X7Y109_D2 = 1'b1;
  assign CLBLM_R_X5Y109_SLICE_X7Y109_D3 = 1'b1;
  assign CLBLM_R_X5Y109_SLICE_X7Y109_D4 = 1'b1;
  assign CLBLM_R_X5Y109_SLICE_X7Y109_D5 = 1'b1;
  assign CLBLM_R_X5Y109_SLICE_X7Y109_D6 = 1'b1;
  assign CLBLM_R_X5Y109_SLICE_X6Y109_A1 = CLBLM_R_X7Y113_SLICE_X8Y113_AO6;
  assign CLBLM_R_X5Y109_SLICE_X6Y109_A2 = CLBLL_L_X4Y107_SLICE_X4Y107_AO6;
  assign CLBLM_R_X5Y109_SLICE_X6Y109_A3 = LIOB33_X0Y101_IOB_X0Y102_I;
  assign CLBLM_R_X5Y109_SLICE_X6Y109_A4 = CLBLM_R_X5Y109_SLICE_X6Y109_BO6;
  assign CLBLM_R_X5Y109_SLICE_X6Y109_A5 = LIOB33_X0Y95_IOB_X0Y95_I;
  assign CLBLM_R_X5Y109_SLICE_X6Y109_A6 = LIOB33_X0Y101_IOB_X0Y101_I;
  assign CLBLM_R_X5Y109_SLICE_X6Y109_B1 = LIOB33_X0Y87_IOB_X0Y88_I;
  assign CLBLM_R_X5Y109_SLICE_X6Y109_B2 = LIOB33_X0Y95_IOB_X0Y95_I;
  assign CLBLM_R_X5Y109_SLICE_X6Y109_B3 = LIOB33_X0Y85_IOB_X0Y86_I;
  assign CLBLM_R_X5Y109_SLICE_X6Y109_B4 = LIOB33_X0Y87_IOB_X0Y87_I;
  assign CLBLM_R_X5Y109_SLICE_X6Y109_B5 = LIOB33_X0Y89_IOB_X0Y90_I;
  assign CLBLM_R_X5Y109_SLICE_X6Y109_B6 = CLBLM_R_X5Y110_SLICE_X6Y110_AO6;
  assign CLBLM_R_X5Y109_SLICE_X6Y109_C1 = 1'b1;
  assign CLBLM_R_X5Y109_SLICE_X6Y109_C2 = 1'b1;
  assign CLBLM_R_X5Y109_SLICE_X6Y109_C3 = 1'b1;
  assign CLBLM_R_X5Y109_SLICE_X6Y109_C4 = 1'b1;
  assign CLBLM_R_X5Y109_SLICE_X6Y109_C5 = 1'b1;
  assign CLBLM_R_X5Y109_SLICE_X6Y109_C6 = 1'b1;
  assign CLBLM_R_X5Y109_SLICE_X6Y109_D1 = 1'b1;
  assign CLBLM_R_X5Y109_SLICE_X6Y109_D2 = 1'b1;
  assign CLBLM_R_X5Y109_SLICE_X6Y109_D3 = 1'b1;
  assign CLBLM_R_X5Y109_SLICE_X6Y109_D4 = 1'b1;
  assign CLBLM_R_X5Y109_SLICE_X6Y109_D5 = 1'b1;
  assign CLBLM_R_X5Y109_SLICE_X6Y109_D6 = 1'b1;
  assign RIOB33_X105Y71_IOB_X1Y72_O = CLBLM_R_X103Y122_SLICE_X163Y122_BO6;
  assign RIOB33_X105Y71_IOB_X1Y71_O = CLBLM_R_X103Y122_SLICE_X163Y122_AO6;
  assign RIOI3_X105Y183_OLOGIC_X1Y183_D1 = RIOB33_X105Y107_IOB_X1Y107_I;
  assign LIOI3_X0Y89_ILOGIC_X0Y90_D = LIOB33_X0Y89_IOB_X0Y90_I;
  assign RIOB33_X105Y87_IOB_X1Y88_O = CLBLM_L_X8Y113_SLICE_X10Y113_BO6;
  assign RIOB33_X105Y131_IOB_X1Y132_O = CLBLM_R_X101Y119_SLICE_X158Y119_AO6;
  assign RIOB33_X105Y87_IOB_X1Y87_O = CLBLM_R_X103Y102_SLICE_X163Y102_BO6;
  assign RIOB33_X105Y131_IOB_X1Y131_O = CLBLM_R_X101Y118_SLICE_X158Y118_AO6;
  assign LIOI3_X0Y89_ILOGIC_X0Y89_D = LIOB33_X0Y89_IOB_X0Y89_I;
  assign CLBLM_L_X10Y123_SLICE_X13Y123_C4 = 1'b1;
  assign CLBLM_L_X10Y123_SLICE_X13Y123_C5 = 1'b1;
  assign CLBLM_L_X10Y123_SLICE_X13Y123_C6 = 1'b1;
  assign RIOB33_X105Y191_IOB_X1Y192_O = CLBLM_R_X103Y177_SLICE_X163Y177_AO5;
  assign RIOB33_X105Y191_IOB_X1Y191_O = CLBLM_R_X103Y177_SLICE_X163Y177_AO5;
  assign LIOI3_X0Y195_OLOGIC_X0Y196_D1 = CLBLM_R_X3Y112_SLICE_X3Y112_BO6;
  assign CLBLM_R_X5Y110_SLICE_X7Y110_A1 = 1'b1;
  assign CLBLM_R_X5Y110_SLICE_X7Y110_A2 = 1'b1;
  assign CLBLM_R_X5Y110_SLICE_X7Y110_A3 = 1'b1;
  assign CLBLM_R_X5Y110_SLICE_X7Y110_A4 = 1'b1;
  assign CLBLM_R_X5Y110_SLICE_X7Y110_A5 = 1'b1;
  assign CLBLM_R_X5Y110_SLICE_X7Y110_A6 = 1'b1;
  assign LIOI3_X0Y195_OLOGIC_X0Y196_T1 = 1'b1;
  assign CLBLM_R_X103Y123_SLICE_X162Y123_A1 = CLBLL_L_X4Y111_SLICE_X5Y111_AO5;
  assign CLBLM_R_X5Y110_SLICE_X7Y110_B1 = 1'b1;
  assign CLBLM_R_X5Y110_SLICE_X7Y110_B2 = 1'b1;
  assign CLBLM_R_X5Y110_SLICE_X7Y110_B3 = 1'b1;
  assign CLBLM_R_X5Y110_SLICE_X7Y110_B4 = 1'b1;
  assign CLBLM_R_X5Y110_SLICE_X7Y110_B5 = 1'b1;
  assign CLBLM_R_X5Y110_SLICE_X7Y110_B6 = 1'b1;
  assign LIOI3_X0Y195_OLOGIC_X0Y195_D1 = 1'b0;
  assign CLBLM_L_X10Y123_SLICE_X13Y123_D5 = 1'b1;
  assign CLBLM_R_X5Y110_SLICE_X7Y110_C1 = 1'b1;
  assign CLBLM_R_X5Y110_SLICE_X7Y110_C2 = 1'b1;
  assign CLBLM_R_X5Y110_SLICE_X7Y110_C3 = 1'b1;
  assign CLBLM_L_X10Y123_SLICE_X13Y123_D6 = 1'b1;
  assign CLBLM_R_X5Y110_SLICE_X7Y110_C4 = 1'b1;
  assign CLBLM_R_X5Y110_SLICE_X7Y110_C5 = 1'b1;
  assign CLBLM_R_X5Y110_SLICE_X7Y110_C6 = 1'b1;
  assign RIOI3_X105Y177_OLOGIC_X1Y178_D1 = CLBLM_R_X103Y177_SLICE_X163Y177_AO6;
  assign LIOI3_X0Y195_OLOGIC_X0Y195_T1 = 1'b1;
  assign RIOI3_X105Y147_OLOGIC_X1Y148_D1 = CLBLM_R_X103Y122_SLICE_X163Y122_DO5;
  assign CLBLM_R_X5Y110_SLICE_X7Y110_D1 = 1'b1;
  assign CLBLM_R_X5Y110_SLICE_X7Y110_D2 = 1'b1;
  assign CLBLM_R_X5Y110_SLICE_X7Y110_D3 = 1'b1;
  assign CLBLM_R_X5Y110_SLICE_X7Y110_D4 = 1'b1;
  assign CLBLM_R_X5Y110_SLICE_X7Y110_D5 = 1'b1;
  assign CLBLM_R_X5Y110_SLICE_X7Y110_D6 = 1'b1;
  assign RIOI3_X105Y177_OLOGIC_X1Y178_T1 = 1'b1;
  assign RIOI3_X105Y147_OLOGIC_X1Y148_T1 = 1'b1;
  assign RIOI3_X105Y85_OLOGIC_X1Y86_D1 = CLBLM_R_X103Y107_SLICE_X163Y107_AO6;
  assign CLBLM_R_X5Y110_SLICE_X6Y110_A1 = LIOB33_X0Y125_IOB_X0Y125_I;
  assign CLBLM_R_X5Y110_SLICE_X6Y110_A2 = 1'b1;
  assign CLBLM_R_X5Y110_SLICE_X6Y110_A3 = LIOB33_X0Y91_IOB_X0Y92_I;
  assign CLBLM_R_X5Y110_SLICE_X6Y110_A4 = LIOB33_X0Y91_IOB_X0Y91_I;
  assign CLBLM_R_X5Y110_SLICE_X6Y110_A5 = LIOB33_X0Y95_IOB_X0Y95_I;
  assign CLBLM_R_X5Y110_SLICE_X6Y110_A6 = 1'b1;
  assign RIOI3_X105Y177_OLOGIC_X1Y177_D1 = LIOB33_X0Y137_IOB_X0Y137_I;
  assign RIOI3_X105Y55_OLOGIC_X1Y56_D1 = CLBLM_R_X5Y111_SLICE_X7Y111_BO6;
  assign RIOI3_X105Y147_OLOGIC_X1Y147_D1 = CLBLM_R_X103Y122_SLICE_X163Y122_CO5;
  assign CLBLM_R_X5Y110_SLICE_X6Y110_B1 = 1'b1;
  assign CLBLM_R_X5Y110_SLICE_X6Y110_B2 = 1'b1;
  assign CLBLM_R_X5Y110_SLICE_X6Y110_B3 = 1'b1;
  assign CLBLM_R_X5Y110_SLICE_X6Y110_B4 = 1'b1;
  assign CLBLM_R_X5Y110_SLICE_X6Y110_B5 = 1'b1;
  assign CLBLM_R_X5Y110_SLICE_X6Y110_B6 = 1'b1;
  assign RIOI3_X105Y85_OLOGIC_X1Y86_T1 = 1'b1;
  assign RIOI3_X105Y177_OLOGIC_X1Y177_T1 = 1'b1;
  assign RIOI3_X105Y55_OLOGIC_X1Y56_T1 = 1'b1;
  assign RIOI3_X105Y147_OLOGIC_X1Y147_T1 = 1'b1;
  assign CLBLM_R_X5Y110_SLICE_X6Y110_C1 = 1'b1;
  assign CLBLM_R_X5Y110_SLICE_X6Y110_C2 = 1'b1;
  assign CLBLM_R_X5Y110_SLICE_X6Y110_C3 = 1'b1;
  assign CLBLM_R_X5Y110_SLICE_X6Y110_C4 = 1'b1;
  assign CLBLM_R_X5Y110_SLICE_X6Y110_C5 = 1'b1;
  assign CLBLM_R_X5Y110_SLICE_X6Y110_C6 = 1'b1;
  assign RIOI3_X105Y85_OLOGIC_X1Y85_D1 = CLBLM_R_X103Y122_SLICE_X163Y122_DO6;
  assign RIOI3_X105Y55_OLOGIC_X1Y55_D1 = CLBLM_L_X10Y114_SLICE_X12Y114_AO6;
  assign RIOI3_X105Y85_OLOGIC_X1Y85_T1 = 1'b1;
  assign CLBLM_R_X5Y110_SLICE_X6Y110_D1 = 1'b1;
  assign CLBLM_R_X5Y110_SLICE_X6Y110_D2 = 1'b1;
  assign CLBLM_R_X5Y110_SLICE_X6Y110_D3 = 1'b1;
  assign CLBLM_R_X5Y110_SLICE_X6Y110_D4 = 1'b1;
  assign CLBLM_R_X5Y110_SLICE_X6Y110_D5 = 1'b1;
  assign CLBLM_R_X5Y110_SLICE_X6Y110_D6 = 1'b1;
  assign RIOI3_X105Y55_OLOGIC_X1Y55_T1 = 1'b1;
  assign RIOI3_TBYTESRC_X105Y81_OLOGIC_X1Y82_D1 = CLBLM_R_X103Y107_SLICE_X163Y107_BO6;
  assign RIOI3_TBYTESRC_X105Y81_OLOGIC_X1Y82_T1 = 1'b1;
  assign RIOI3_TBYTESRC_X105Y81_OLOGIC_X1Y81_D1 = CLBLM_R_X103Y122_SLICE_X163Y122_CO6;
  assign RIOI3_TBYTESRC_X105Y81_OLOGIC_X1Y81_T1 = 1'b1;
  assign LIOI3_X0Y121_ILOGIC_X0Y122_D = LIOB33_X0Y121_IOB_X0Y122_I;
  assign CLBLM_R_X103Y123_SLICE_X162Y123_A2 = CLBLM_L_X10Y123_SLICE_X12Y123_AO6;
  assign LIOI3_X0Y121_ILOGIC_X0Y121_D = LIOB33_X0Y121_IOB_X0Y121_I;
  assign RIOB33_X105Y73_IOB_X1Y74_O = CLBLL_L_X100Y113_SLICE_X156Y113_AO6;
  assign RIOB33_X105Y73_IOB_X1Y73_O = CLBLL_L_X36Y113_SLICE_X54Y113_AO6;
  assign CLBLM_L_X10Y123_SLICE_X12Y123_C2 = 1'b1;
  assign CLBLM_L_X10Y123_SLICE_X12Y123_C3 = 1'b1;
  assign CLBLM_L_X10Y123_SLICE_X12Y123_C4 = 1'b1;
  assign LIOI3_X0Y165_ILOGIC_X0Y166_D = LIOB33_X0Y165_IOB_X0Y166_I;
  assign RIOB33_X105Y133_IOB_X1Y134_O = CLBLM_R_X101Y118_SLICE_X158Y118_BO6;
  assign RIOB33_X105Y133_IOB_X1Y133_O = CLBLM_R_X101Y123_SLICE_X158Y123_CO6;
  assign LIOI3_X0Y165_ILOGIC_X0Y165_D = LIOB33_X0Y165_IOB_X0Y165_I;
  assign CLBLL_L_X4Y107_SLICE_X4Y107_A1 = LIOB33_X0Y83_IOB_X0Y84_I;
  assign CLBLL_L_X4Y107_SLICE_X4Y107_A2 = LIOB33_X0Y105_IOB_X0Y105_I;
  assign CLBLL_L_X4Y107_SLICE_X4Y107_A3 = LIOB33_X0Y95_IOB_X0Y95_I;
  assign CLBLL_L_X4Y107_SLICE_X4Y107_A4 = CLBLL_L_X4Y107_SLICE_X4Y107_BO6;
  assign CLBLL_L_X4Y107_SLICE_X4Y107_A5 = LIOB33_X0Y85_IOB_X0Y85_I;
  assign CLBLL_L_X4Y107_SLICE_X4Y107_A6 = LIOB33_X0Y107_IOB_X0Y107_I;
  assign LIOI3_X0Y133_ILOGIC_X0Y134_D = LIOB33_X0Y133_IOB_X0Y134_I;
  assign LIOI3_X0Y133_ILOGIC_X0Y133_D = LIOB33_X0Y133_IOB_X0Y133_I;
  assign LIOI3_X0Y103_ILOGIC_X0Y104_D = LIOB33_X0Y103_IOB_X0Y104_I;
  assign CLBLL_L_X4Y107_SLICE_X4Y107_B1 = 1'b1;
  assign CLBLL_L_X4Y107_SLICE_X4Y107_B2 = 1'b1;
  assign CLBLL_L_X4Y107_SLICE_X4Y107_B3 = LIOB33_X0Y103_IOB_X0Y103_I;
  assign CLBLL_L_X4Y107_SLICE_X4Y107_B4 = LIOB33_X0Y103_IOB_X0Y104_I;
  assign CLBLL_L_X4Y107_SLICE_X4Y107_B5 = 1'b1;
  assign CLBLL_L_X4Y107_SLICE_X4Y107_B6 = 1'b1;
  assign LIOI3_X0Y73_ILOGIC_X0Y74_D = LIOB33_X0Y73_IOB_X0Y74_I;
  assign LIOI3_X0Y103_ILOGIC_X0Y103_D = LIOB33_X0Y103_IOB_X0Y103_I;
  assign CLBLL_L_X4Y107_SLICE_X4Y107_C1 = 1'b1;
  assign CLBLL_L_X4Y107_SLICE_X4Y107_C2 = 1'b1;
  assign CLBLL_L_X4Y107_SLICE_X4Y107_C3 = 1'b1;
  assign CLBLL_L_X4Y107_SLICE_X4Y107_C4 = 1'b1;
  assign CLBLL_L_X4Y107_SLICE_X4Y107_C5 = 1'b1;
  assign CLBLL_L_X4Y107_SLICE_X4Y107_C6 = 1'b1;
  assign LIOI3_X0Y151_ILOGIC_X0Y152_D = LIOB33_X0Y151_IOB_X0Y152_I;
  assign CLBLL_L_X4Y110_SLICE_X4Y110_A4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign RIOI3_X105Y117_ILOGIC_X1Y118_D = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLL_L_X4Y107_SLICE_X4Y107_D1 = 1'b1;
  assign CLBLL_L_X4Y107_SLICE_X4Y107_D2 = 1'b1;
  assign CLBLL_L_X4Y107_SLICE_X4Y107_D3 = 1'b1;
  assign CLBLL_L_X4Y107_SLICE_X4Y107_D4 = 1'b1;
  assign CLBLL_L_X4Y107_SLICE_X4Y107_D5 = 1'b1;
  assign CLBLL_L_X4Y107_SLICE_X4Y107_D6 = 1'b1;
  assign CLBLL_L_X4Y110_SLICE_X4Y110_A6 = 1'b1;
  assign LIOI3_TBYTETERM_X0Y87_ILOGIC_X0Y88_D = LIOB33_X0Y87_IOB_X0Y88_I;
  assign LIOI3_TBYTETERM_X0Y87_ILOGIC_X0Y87_D = LIOB33_X0Y87_IOB_X0Y87_I;
  assign RIOB33_X105Y193_IOB_X1Y193_O = CLBLM_R_X103Y177_SLICE_X163Y177_AO5;
  assign RIOB33_X105Y193_IOB_X1Y194_O = CLBLM_R_X103Y193_SLICE_X163Y193_AO6;
  assign LIOI3_TBYTESRC_X0Y157_ILOGIC_X0Y158_D = LIOB33_X0Y157_IOB_X0Y158_I;
  assign LIOI3_TBYTESRC_X0Y157_ILOGIC_X0Y157_D = LIOB33_X0Y157_IOB_X0Y157_I;
  assign CLBLL_L_X4Y110_SLICE_X4Y110_B1 = LIOB33_X0Y81_IOB_X0Y81_I;
  assign CLBLL_L_X4Y107_SLICE_X5Y107_A1 = 1'b1;
  assign CLBLL_L_X4Y107_SLICE_X5Y107_A2 = 1'b1;
  assign CLBLL_L_X4Y107_SLICE_X5Y107_A3 = 1'b1;
  assign CLBLL_L_X4Y107_SLICE_X5Y107_A4 = 1'b1;
  assign CLBLL_L_X4Y107_SLICE_X5Y107_A5 = 1'b1;
  assign CLBLL_L_X4Y107_SLICE_X5Y107_A6 = 1'b1;
  assign CLBLL_L_X4Y107_SLICE_X5Y107_B1 = 1'b1;
  assign CLBLL_L_X4Y107_SLICE_X5Y107_B2 = 1'b1;
  assign CLBLL_L_X4Y107_SLICE_X5Y107_B3 = 1'b1;
  assign CLBLM_R_X7Y121_SLICE_X9Y121_A1 = CLBLM_R_X7Y113_SLICE_X9Y113_AO6;
  assign CLBLM_R_X7Y121_SLICE_X9Y121_A2 = RIOB33_X105Y119_IOB_X1Y120_I;
  assign CLBLM_R_X7Y121_SLICE_X9Y121_A3 = LIOB33_X0Y161_IOB_X0Y162_I;
  assign CLBLM_R_X7Y121_SLICE_X9Y121_A4 = RIOB33_X105Y121_IOB_X1Y121_I;
  assign CLBLM_R_X7Y121_SLICE_X9Y121_A5 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X7Y121_SLICE_X9Y121_A6 = 1'b1;
  assign CLBLL_L_X4Y107_SLICE_X5Y107_B4 = 1'b1;
  assign CLBLL_L_X4Y107_SLICE_X5Y107_B5 = 1'b1;
  assign CLBLL_L_X4Y107_SLICE_X5Y107_B6 = 1'b1;
  assign CLBLM_R_X7Y121_SLICE_X9Y121_B1 = 1'b1;
  assign CLBLM_R_X7Y121_SLICE_X9Y121_B2 = 1'b1;
  assign CLBLM_R_X7Y121_SLICE_X9Y121_B3 = 1'b1;
  assign CLBLM_R_X7Y121_SLICE_X9Y121_B4 = 1'b1;
  assign CLBLL_L_X4Y107_SLICE_X5Y107_C1 = 1'b1;
  assign CLBLL_L_X4Y107_SLICE_X5Y107_C2 = 1'b1;
  assign CLBLL_L_X4Y107_SLICE_X5Y107_C3 = 1'b1;
  assign CLBLL_L_X4Y107_SLICE_X5Y107_C4 = 1'b1;
  assign CLBLL_L_X4Y107_SLICE_X5Y107_C5 = 1'b1;
  assign CLBLM_R_X5Y111_SLICE_X7Y111_A1 = LIOB33_X0Y115_IOB_X0Y116_I;
  assign CLBLM_R_X5Y111_SLICE_X7Y111_A2 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X5Y111_SLICE_X7Y111_A3 = CLBLL_L_X4Y111_SLICE_X4Y111_AO5;
  assign CLBLM_R_X5Y111_SLICE_X7Y111_A4 = LIOB33_X0Y95_IOB_X0Y96_I;
  assign CLBLM_R_X5Y111_SLICE_X7Y111_A5 = LIOB33_X0Y59_IOB_X0Y60_I;
  assign CLBLM_R_X5Y111_SLICE_X7Y111_A6 = 1'b1;
  assign CLBLL_L_X4Y107_SLICE_X5Y107_D1 = 1'b1;
  assign CLBLL_L_X4Y107_SLICE_X5Y107_D2 = 1'b1;
  assign CLBLM_R_X5Y111_SLICE_X7Y111_B1 = RIOB33_X105Y161_IOB_X1Y161_I;
  assign CLBLM_R_X5Y111_SLICE_X7Y111_B2 = LIOB33_X0Y79_IOB_X0Y80_I;
  assign CLBLM_R_X5Y111_SLICE_X7Y111_B3 = LIOB33_X0Y109_IOB_X0Y109_I;
  assign CLBLM_R_X5Y111_SLICE_X7Y111_B4 = CLBLM_R_X5Y115_SLICE_X6Y115_AO6;
  assign CLBLM_R_X5Y111_SLICE_X7Y111_B5 = CLBLL_L_X4Y110_SLICE_X4Y110_BO5;
  assign CLBLM_R_X5Y111_SLICE_X7Y111_B6 = CLBLM_L_X10Y123_SLICE_X12Y123_AO6;
  assign CLBLL_L_X4Y107_SLICE_X5Y107_D6 = 1'b1;
  assign CLBLM_R_X5Y111_SLICE_X7Y111_C1 = LIOB33_X0Y113_IOB_X0Y114_I;
  assign CLBLM_R_X5Y111_SLICE_X7Y111_C2 = CLBLM_L_X10Y123_SLICE_X12Y123_AO6;
  assign CLBLM_R_X5Y111_SLICE_X7Y111_C3 = LIOB33_X0Y75_IOB_X0Y75_I;
  assign CLBLM_R_X5Y111_SLICE_X7Y111_C4 = CLBLL_L_X4Y111_SLICE_X4Y111_CO6;
  assign CLBLM_R_X5Y111_SLICE_X7Y111_C5 = CLBLM_R_X5Y115_SLICE_X6Y115_AO6;
  assign CLBLM_R_X5Y111_SLICE_X7Y111_C6 = RIOB33_X105Y169_IOB_X1Y169_I;
  assign CLBLL_L_X2Y146_SLICE_X0Y146_A1 = 1'b1;
  assign CLBLL_L_X2Y146_SLICE_X0Y146_A2 = 1'b1;
  assign CLBLL_L_X2Y146_SLICE_X0Y146_A3 = 1'b1;
  assign CLBLL_L_X2Y146_SLICE_X0Y146_A4 = 1'b1;
  assign CLBLL_L_X2Y146_SLICE_X0Y146_A5 = 1'b1;
  assign CLBLL_L_X2Y146_SLICE_X0Y146_A6 = 1'b1;
  assign CLBLL_L_X2Y146_SLICE_X0Y146_B1 = 1'b1;
  assign CLBLM_R_X5Y111_SLICE_X7Y111_D1 = LIOB33_X0Y113_IOB_X0Y114_I;
  assign CLBLM_R_X5Y111_SLICE_X7Y111_D2 = 1'b1;
  assign CLBLM_R_X5Y111_SLICE_X7Y111_D3 = LIOB33_X0Y75_IOB_X0Y75_I;
  assign CLBLM_R_X5Y111_SLICE_X7Y111_D4 = 1'b1;
  assign CLBLM_R_X5Y111_SLICE_X7Y111_D5 = LIOB33_X0Y109_IOB_X0Y109_I;
  assign CLBLM_R_X5Y111_SLICE_X7Y111_D6 = LIOB33_X0Y79_IOB_X0Y80_I;
  assign CLBLL_L_X2Y146_SLICE_X0Y146_B2 = 1'b1;
  assign CLBLL_L_X2Y146_SLICE_X0Y146_B3 = 1'b1;
  assign CLBLL_L_X2Y146_SLICE_X0Y146_B4 = 1'b1;
  assign CLBLL_L_X2Y146_SLICE_X0Y146_B5 = 1'b1;
  assign CLBLL_L_X2Y146_SLICE_X0Y146_B6 = 1'b1;
  assign CLBLL_L_X2Y146_SLICE_X0Y146_C1 = 1'b1;
  assign CLBLM_R_X5Y111_SLICE_X6Y111_A1 = LIOB33_X0Y117_IOB_X0Y118_I;
  assign CLBLM_R_X5Y111_SLICE_X6Y111_A2 = CLBLL_L_X4Y112_SLICE_X4Y112_BO6;
  assign CLBLM_R_X5Y111_SLICE_X6Y111_A3 = CLBLL_L_X4Y111_SLICE_X5Y111_BO6;
  assign CLBLM_R_X5Y111_SLICE_X6Y111_A4 = CLBLM_R_X3Y111_SLICE_X3Y111_BO6;
  assign CLBLM_R_X5Y111_SLICE_X6Y111_A5 = LIOB33_X0Y111_IOB_X0Y112_I;
  assign CLBLM_R_X5Y111_SLICE_X6Y111_A6 = 1'b1;
  assign CLBLL_L_X2Y146_SLICE_X0Y146_C3 = 1'b1;
  assign CLBLL_L_X2Y146_SLICE_X0Y146_C4 = 1'b1;
  assign CLBLL_L_X2Y146_SLICE_X0Y146_C5 = 1'b1;
  assign CLBLM_R_X5Y111_SLICE_X6Y111_B1 = CLBLM_R_X5Y115_SLICE_X6Y115_AO5;
  assign CLBLM_R_X5Y111_SLICE_X6Y111_B2 = CLBLL_L_X4Y112_SLICE_X4Y112_BO6;
  assign CLBLM_R_X5Y111_SLICE_X6Y111_B3 = CLBLM_L_X10Y123_SLICE_X12Y123_AO6;
  assign CLBLM_R_X5Y111_SLICE_X6Y111_B4 = LIOB33_X0Y111_IOB_X0Y112_I;
  assign CLBLM_R_X5Y111_SLICE_X6Y111_B5 = CLBLL_L_X4Y111_SLICE_X5Y111_BO6;
  assign CLBLL_L_X2Y146_SLICE_X0Y146_D1 = 1'b1;
  assign CLBLL_L_X2Y146_SLICE_X0Y146_D2 = 1'b1;
  assign CLBLL_L_X2Y146_SLICE_X0Y146_D3 = 1'b1;
  assign CLBLL_L_X2Y146_SLICE_X0Y146_D4 = 1'b1;
  assign CLBLL_L_X2Y146_SLICE_X0Y146_D5 = 1'b1;
  assign CLBLL_L_X2Y146_SLICE_X0Y146_D6 = 1'b1;
  assign CLBLM_R_X7Y121_SLICE_X8Y121_D5 = 1'b1;
  assign CLBLM_R_X7Y121_SLICE_X8Y121_D6 = 1'b1;
  assign CLBLM_R_X5Y111_SLICE_X6Y111_C3 = LIOB33_X0Y117_IOB_X0Y118_I;
  assign CLBLM_R_X5Y111_SLICE_X6Y111_C4 = CLBLM_R_X5Y111_SLICE_X6Y111_AO5;
  assign CLBLM_R_X5Y111_SLICE_X6Y111_C5 = CLBLM_R_X5Y111_SLICE_X6Y111_DO6;
  assign CLBLM_R_X5Y111_SLICE_X6Y111_C1 = CLBLL_L_X4Y111_SLICE_X5Y111_AO5;
  assign CLBLM_R_X5Y111_SLICE_X6Y111_C2 = CLBLM_R_X3Y111_SLICE_X2Y111_AO5;
  assign CLBLM_R_X5Y111_SLICE_X6Y111_C6 = CLBLM_R_X3Y111_SLICE_X3Y111_BO6;
  assign CLBLM_R_X7Y121_SLICE_X9Y121_B5 = 1'b1;
  assign CLBLM_R_X7Y121_SLICE_X9Y121_B6 = 1'b1;
  assign RIOB33_X105Y147_IOB_X1Y148_O = CLBLM_R_X103Y122_SLICE_X163Y122_DO5;
  assign RIOB33_X105Y147_IOB_X1Y147_O = CLBLM_R_X103Y122_SLICE_X163Y122_CO5;
  assign CLBLM_R_X5Y111_SLICE_X6Y111_D1 = CLBLL_L_X4Y110_SLICE_X4Y110_BO5;
  assign CLBLM_R_X5Y111_SLICE_X6Y111_D2 = CLBLM_R_X5Y111_SLICE_X7Y111_AO5;
  assign CLBLM_R_X5Y111_SLICE_X6Y111_D3 = CLBLM_R_X5Y112_SLICE_X6Y112_BO6;
  assign CLBLM_R_X5Y111_SLICE_X6Y111_D4 = CLBLL_L_X4Y112_SLICE_X4Y112_CO6;
  assign CLBLM_R_X5Y111_SLICE_X6Y111_D5 = CLBLL_L_X4Y111_SLICE_X4Y111_AO5;
  assign CLBLM_R_X5Y111_SLICE_X6Y111_D6 = CLBLL_L_X4Y111_SLICE_X4Y111_CO6;
  assign CLBLL_L_X2Y146_SLICE_X1Y146_A1 = LIOB33_X0Y75_IOB_X0Y76_I;
  assign CLBLL_L_X2Y146_SLICE_X1Y146_A2 = 1'b1;
  assign CLBLL_L_X2Y146_SLICE_X1Y146_A3 = LIOB33_X0Y89_IOB_X0Y89_I;
  assign CLBLL_L_X2Y146_SLICE_X1Y146_A4 = RIOB33_X105Y105_IOB_X1Y106_I;
  assign CLBLL_L_X2Y146_SLICE_X1Y146_A5 = LIOB33_X0Y145_IOB_X0Y146_I;
  assign CLBLL_L_X2Y146_SLICE_X1Y146_A6 = 1'b1;
  assign CLBLL_L_X2Y146_SLICE_X1Y146_B1 = 1'b1;
  assign CLBLL_L_X2Y146_SLICE_X1Y146_B2 = 1'b1;
  assign CLBLL_L_X2Y146_SLICE_X1Y146_B3 = 1'b1;
  assign CLBLL_L_X2Y146_SLICE_X1Y146_B4 = 1'b1;
  assign CLBLL_L_X2Y146_SLICE_X1Y146_B5 = 1'b1;
  assign CLBLL_L_X2Y146_SLICE_X1Y146_B6 = 1'b1;
  assign CLBLM_R_X7Y121_SLICE_X9Y121_C1 = 1'b1;
  assign CLBLM_R_X7Y121_SLICE_X9Y121_C2 = 1'b1;
  assign CLBLL_L_X2Y146_SLICE_X1Y146_C1 = 1'b1;
  assign CLBLL_L_X2Y146_SLICE_X1Y146_C2 = 1'b1;
  assign CLBLL_L_X2Y146_SLICE_X1Y146_C3 = 1'b1;
  assign CLBLL_L_X2Y146_SLICE_X1Y146_C4 = 1'b1;
  assign CLBLL_L_X2Y146_SLICE_X1Y146_C5 = 1'b1;
  assign CLBLL_L_X2Y146_SLICE_X1Y146_C6 = 1'b1;
  assign CLBLM_R_X7Y121_SLICE_X9Y121_C3 = 1'b1;
  assign CLBLM_R_X7Y121_SLICE_X9Y121_C4 = 1'b1;
  assign CLBLM_R_X7Y121_SLICE_X9Y121_C5 = 1'b1;
  assign CLBLL_L_X2Y146_SLICE_X1Y146_D1 = 1'b1;
  assign CLBLL_L_X2Y146_SLICE_X1Y146_D2 = 1'b1;
  assign CLBLL_L_X2Y146_SLICE_X1Y146_D3 = 1'b1;
  assign CLBLL_L_X2Y146_SLICE_X1Y146_D4 = 1'b1;
  assign CLBLL_L_X2Y146_SLICE_X1Y146_D5 = 1'b1;
  assign CLBLL_L_X2Y146_SLICE_X1Y146_D6 = 1'b1;
  assign CLBLM_R_X7Y121_SLICE_X9Y121_C6 = 1'b1;
  assign RIOB33_X105Y75_IOB_X1Y75_O = CLBLM_R_X29Y115_SLICE_X42Y115_AO6;
  assign RIOB33_X105Y75_IOB_X1Y76_O = CLBLL_R_X57Y113_SLICE_X86Y113_BO6;
  assign RIOB33_X105Y135_IOB_X1Y136_O = CLBLM_R_X101Y118_SLICE_X158Y118_CO6;
  assign RIOB33_X105Y135_IOB_X1Y135_O = CLBLM_R_X101Y119_SLICE_X158Y119_CO6;
  assign RIOB33_X105Y195_IOB_X1Y196_O = CLBLL_L_X2Y173_SLICE_X0Y173_AO6;
  assign CLBLM_R_X7Y121_SLICE_X9Y121_D1 = 1'b1;
  assign RIOB33_X105Y195_IOB_X1Y195_O = LIOB33_X0Y85_IOB_X0Y85_I;
  assign CLBLM_R_X7Y121_SLICE_X9Y121_D2 = 1'b1;
  assign CLBLM_R_X7Y121_SLICE_X9Y121_D3 = 1'b1;
  assign CLBLM_R_X7Y121_SLICE_X9Y121_D4 = 1'b1;
  assign CLBLM_R_X7Y121_SLICE_X9Y121_D5 = 1'b1;
  assign CLBLL_L_X2Y173_SLICE_X0Y173_A1 = LIOB33_X0Y145_IOB_X0Y145_I;
  assign CLBLL_L_X2Y173_SLICE_X0Y173_A2 = 1'b1;
  assign CLBLL_L_X2Y173_SLICE_X0Y173_A3 = LIOB33_X0Y171_IOB_X0Y172_I;
  assign CLBLL_L_X2Y173_SLICE_X0Y173_A4 = LIOB33_X0Y75_IOB_X0Y76_I;
  assign CLBLL_L_X2Y173_SLICE_X0Y173_A5 = LIOB33_X0Y173_IOB_X0Y173_I;
  assign CLBLL_L_X2Y173_SLICE_X0Y173_A6 = LIOB33_X0Y89_IOB_X0Y89_I;
  assign CLBLM_R_X7Y121_SLICE_X9Y121_D6 = 1'b1;
  assign CLBLL_L_X2Y173_SLICE_X0Y173_B1 = 1'b1;
  assign CLBLL_L_X2Y173_SLICE_X0Y173_B2 = 1'b1;
  assign CLBLL_L_X2Y173_SLICE_X0Y173_B3 = 1'b1;
  assign CLBLL_L_X2Y173_SLICE_X0Y173_B4 = 1'b1;
  assign CLBLL_L_X2Y173_SLICE_X0Y173_B5 = 1'b1;
  assign CLBLL_L_X2Y173_SLICE_X0Y173_B6 = 1'b1;
  assign CLBLM_R_X103Y115_SLICE_X162Y115_B1 = 1'b1;
  assign CLBLM_R_X103Y193_SLICE_X163Y193_A1 = 1'b1;
  assign CLBLL_L_X2Y173_SLICE_X0Y173_C1 = 1'b1;
  assign CLBLL_L_X2Y173_SLICE_X0Y173_C2 = 1'b1;
  assign CLBLL_L_X2Y173_SLICE_X0Y173_C3 = 1'b1;
  assign CLBLL_L_X2Y173_SLICE_X0Y173_C4 = 1'b1;
  assign CLBLL_L_X2Y173_SLICE_X0Y173_C5 = 1'b1;
  assign CLBLL_L_X2Y173_SLICE_X0Y173_C6 = 1'b1;
  assign CLBLM_R_X103Y115_SLICE_X163Y115_A1 = RIOB33_X105Y123_IOB_X1Y124_I;
  assign CLBLM_R_X103Y115_SLICE_X163Y115_A2 = 1'b1;
  assign CLBLM_R_X103Y115_SLICE_X163Y115_A3 = CLBLM_R_X5Y112_SLICE_X6Y112_AO6;
  assign CLBLM_R_X103Y115_SLICE_X163Y115_A4 = RIOB33_X105Y113_IOB_X1Y113_I;
  assign CLBLM_R_X103Y115_SLICE_X163Y115_A5 = CLBLM_L_X10Y114_SLICE_X12Y114_AO6;
  assign CLBLM_R_X103Y115_SLICE_X163Y115_A6 = 1'b1;
  assign CLBLM_R_X103Y193_SLICE_X163Y193_A5 = 1'b1;
  assign CLBLL_L_X2Y173_SLICE_X0Y173_D1 = 1'b1;
  assign CLBLL_L_X2Y173_SLICE_X0Y173_D2 = 1'b1;
  assign CLBLL_L_X2Y173_SLICE_X0Y173_D3 = 1'b1;
  assign CLBLL_L_X2Y173_SLICE_X0Y173_D4 = 1'b1;
  assign CLBLL_L_X2Y173_SLICE_X0Y173_D5 = 1'b1;
  assign CLBLL_L_X2Y173_SLICE_X0Y173_D6 = 1'b1;
  assign CLBLM_R_X103Y115_SLICE_X162Y115_B2 = 1'b1;
  assign CLBLM_R_X103Y115_SLICE_X163Y115_B1 = 1'b1;
  assign CLBLM_R_X7Y121_SLICE_X8Y121_A1 = LIOB33_X0Y159_IOB_X0Y160_I;
  assign CLBLM_R_X103Y115_SLICE_X163Y115_B2 = 1'b1;
  assign CLBLM_R_X103Y115_SLICE_X163Y115_B3 = 1'b1;
  assign CLBLM_R_X103Y115_SLICE_X163Y115_B4 = 1'b1;
  assign CLBLM_R_X7Y121_SLICE_X8Y121_A2 = CLBLM_R_X5Y114_SLICE_X6Y114_CO6;
  assign CLBLM_R_X103Y115_SLICE_X163Y115_B6 = 1'b1;
  assign CLBLM_R_X103Y115_SLICE_X163Y115_C1 = 1'b1;
  assign CLBLM_R_X103Y115_SLICE_X163Y115_C2 = 1'b1;
  assign CLBLM_R_X7Y121_SLICE_X8Y121_A3 = CLBLM_R_X7Y121_SLICE_X9Y121_AO6;
  assign CLBLM_R_X103Y115_SLICE_X163Y115_C3 = 1'b1;
  assign CLBLM_R_X103Y115_SLICE_X163Y115_C4 = 1'b1;
  assign CLBLM_R_X103Y115_SLICE_X163Y115_C5 = 1'b1;
  assign CLBLM_R_X103Y115_SLICE_X163Y115_C6 = 1'b1;
  assign CLBLM_R_X7Y121_SLICE_X8Y121_A4 = LIOB33_X0Y159_IOB_X0Y159_I;
  assign CLBLM_R_X103Y115_SLICE_X163Y115_D1 = 1'b1;
  assign CLBLM_R_X103Y115_SLICE_X162Y115_B3 = 1'b1;
  assign CLBLM_R_X103Y115_SLICE_X163Y115_D2 = 1'b1;
  assign CLBLM_R_X7Y121_SLICE_X8Y121_A5 = LIOB33_X0Y177_IOB_X0Y177_I;
  assign CLBLM_R_X103Y115_SLICE_X163Y115_D3 = 1'b1;
  assign CLBLM_R_X103Y115_SLICE_X163Y115_D4 = 1'b1;
  assign CLBLM_R_X103Y115_SLICE_X163Y115_D5 = 1'b1;
  assign CLBLM_R_X103Y115_SLICE_X163Y115_D6 = 1'b1;
  assign CLBLM_R_X7Y121_SLICE_X8Y121_A6 = CLBLL_L_X4Y112_SLICE_X5Y112_CO6;
  assign CLBLL_L_X2Y173_SLICE_X1Y173_A1 = LIOB33_X0Y145_IOB_X0Y145_I;
  assign CLBLL_L_X2Y173_SLICE_X1Y173_A2 = LIOB33_X0Y75_IOB_X0Y76_I;
  assign CLBLL_L_X2Y173_SLICE_X1Y173_A3 = LIOB33_X0Y173_IOB_X0Y174_I;
  assign CLBLL_L_X2Y173_SLICE_X1Y173_A4 = LIOB33_X0Y89_IOB_X0Y89_I;
  assign CLBLL_L_X2Y173_SLICE_X1Y173_A5 = LIOB33_X0Y97_IOB_X0Y98_I;
  assign CLBLL_L_X2Y173_SLICE_X1Y173_A6 = 1'b1;
  assign CLBLM_R_X103Y115_SLICE_X162Y115_A1 = 1'b1;
  assign CLBLM_R_X103Y115_SLICE_X162Y115_A2 = 1'b1;
  assign CLBLM_R_X103Y115_SLICE_X162Y115_A3 = 1'b1;
  assign CLBLL_L_X2Y173_SLICE_X1Y173_B1 = LIOB33_X0Y145_IOB_X0Y145_I;
  assign CLBLL_L_X2Y173_SLICE_X1Y173_B2 = LIOB33_X0Y75_IOB_X0Y76_I;
  assign CLBLL_L_X2Y173_SLICE_X1Y173_B3 = RIOB33_X105Y107_IOB_X1Y107_I;
  assign CLBLL_L_X2Y173_SLICE_X1Y173_B4 = LIOB33_X0Y89_IOB_X0Y89_I;
  assign CLBLL_L_X2Y173_SLICE_X1Y173_B5 = LIOB33_X0Y171_IOB_X0Y171_I;
  assign CLBLL_L_X2Y173_SLICE_X1Y173_B6 = 1'b1;
  assign CLBLM_R_X103Y115_SLICE_X162Y115_A5 = 1'b1;
  assign CLBLM_R_X103Y115_SLICE_X162Y115_A6 = 1'b1;
  assign CLBLL_L_X2Y173_SLICE_X1Y173_C1 = 1'b1;
  assign CLBLL_L_X2Y173_SLICE_X1Y173_C2 = 1'b1;
  assign CLBLL_L_X2Y173_SLICE_X1Y173_C3 = 1'b1;
  assign CLBLL_L_X2Y173_SLICE_X1Y173_C4 = 1'b1;
  assign CLBLL_L_X2Y173_SLICE_X1Y173_C5 = 1'b1;
  assign CLBLL_L_X2Y173_SLICE_X1Y173_C6 = 1'b1;
  assign CLBLM_R_X103Y115_SLICE_X162Y115_B4 = 1'b1;
  assign CLBLM_R_X103Y115_SLICE_X162Y115_B5 = 1'b1;
  assign CLBLM_R_X7Y121_SLICE_X8Y121_B1 = LIOB33_X0Y159_IOB_X0Y160_I;
  assign CLBLM_R_X103Y115_SLICE_X162Y115_C1 = 1'b1;
  assign CLBLM_R_X103Y115_SLICE_X162Y115_C2 = 1'b1;
  assign CLBLM_R_X103Y115_SLICE_X162Y115_C3 = 1'b1;
  assign CLBLM_R_X7Y121_SLICE_X8Y121_B2 = CLBLM_R_X5Y114_SLICE_X6Y114_CO6;
  assign CLBLL_L_X2Y173_SLICE_X1Y173_D1 = 1'b1;
  assign CLBLL_L_X2Y173_SLICE_X1Y173_D2 = 1'b1;
  assign CLBLL_L_X2Y173_SLICE_X1Y173_D3 = 1'b1;
  assign CLBLL_L_X2Y173_SLICE_X1Y173_D4 = 1'b1;
  assign CLBLL_L_X2Y173_SLICE_X1Y173_D5 = 1'b1;
  assign CLBLL_L_X2Y173_SLICE_X1Y173_D6 = 1'b1;
  assign CLBLM_R_X7Y121_SLICE_X8Y121_B3 = CLBLM_R_X7Y121_SLICE_X9Y121_AO5;
  assign CLBLM_R_X5Y112_SLICE_X7Y112_A1 = LIOB33_X0Y103_IOB_X0Y103_I;
  assign CLBLM_R_X5Y112_SLICE_X7Y112_A2 = LIOB33_X0Y67_IOB_X0Y68_I;
  assign CLBLM_R_X5Y112_SLICE_X7Y112_A3 = LIOB33_X0Y125_IOB_X0Y125_I;
  assign CLBLM_R_X5Y112_SLICE_X7Y112_A4 = LIOB33_X0Y91_IOB_X0Y91_I;
  assign CLBLM_R_X5Y112_SLICE_X7Y112_A5 = LIOB33_X0Y69_IOB_X0Y70_I;
  assign CLBLM_R_X5Y112_SLICE_X7Y112_A6 = 1'b1;
  assign CLBLM_R_X7Y121_SLICE_X8Y121_B4 = CLBLL_L_X4Y112_SLICE_X5Y112_CO6;
  assign CLBLM_R_X7Y121_SLICE_X8Y121_B5 = LIOB33_X0Y177_IOB_X0Y177_I;
  assign CLBLM_R_X7Y121_SLICE_X8Y121_B6 = LIOB33_X0Y159_IOB_X0Y159_I;
  assign CLBLM_R_X5Y112_SLICE_X7Y112_B1 = 1'b1;
  assign CLBLM_R_X5Y112_SLICE_X7Y112_B2 = 1'b1;
  assign CLBLM_R_X5Y112_SLICE_X7Y112_B3 = 1'b1;
  assign CLBLM_R_X5Y112_SLICE_X7Y112_B4 = 1'b1;
  assign CLBLM_R_X5Y112_SLICE_X7Y112_B5 = 1'b1;
  assign CLBLM_R_X5Y112_SLICE_X7Y112_B6 = 1'b1;
  assign CLBLL_L_X4Y110_SLICE_X5Y110_B5 = 1'b1;
  assign CLBLM_R_X5Y112_SLICE_X7Y112_C1 = 1'b1;
  assign CLBLM_R_X5Y112_SLICE_X7Y112_C2 = 1'b1;
  assign CLBLM_R_X5Y112_SLICE_X7Y112_C3 = 1'b1;
  assign CLBLM_R_X5Y112_SLICE_X7Y112_C4 = 1'b1;
  assign CLBLM_R_X5Y112_SLICE_X7Y112_C5 = 1'b1;
  assign CLBLM_R_X5Y112_SLICE_X7Y112_C6 = 1'b1;
  assign CLBLM_R_X5Y112_SLICE_X7Y112_D1 = 1'b1;
  assign CLBLM_R_X5Y112_SLICE_X7Y112_D2 = 1'b1;
  assign CLBLM_R_X5Y112_SLICE_X7Y112_D3 = 1'b1;
  assign CLBLM_R_X5Y112_SLICE_X7Y112_D4 = 1'b1;
  assign CLBLM_R_X5Y112_SLICE_X7Y112_D5 = 1'b1;
  assign CLBLM_R_X5Y112_SLICE_X7Y112_D6 = 1'b1;
  assign CLBLM_R_X7Y121_SLICE_X8Y121_C1 = 1'b1;
  assign CLBLM_R_X7Y121_SLICE_X8Y121_C2 = 1'b1;
  assign RIOI3_SING_X105Y50_OLOGIC_X1Y50_T1 = 1'b1;
  assign CLBLM_R_X5Y112_SLICE_X6Y112_A1 = CLBLM_L_X10Y123_SLICE_X12Y123_AO6;
  assign CLBLM_R_X5Y112_SLICE_X6Y112_A2 = LIOB33_X0Y77_IOB_X0Y78_I;
  assign CLBLM_R_X5Y112_SLICE_X6Y112_A3 = LIOB33_X0Y115_IOB_X0Y115_I;
  assign CLBLM_R_X5Y112_SLICE_X6Y112_A4 = CLBLM_R_X5Y112_SLICE_X6Y112_BO6;
  assign CLBLM_R_X5Y112_SLICE_X6Y112_A5 = CLBLM_R_X5Y115_SLICE_X6Y115_AO6;
  assign CLBLM_R_X5Y112_SLICE_X6Y112_A6 = RIOB33_X105Y167_IOB_X1Y168_I;
  assign CLBLM_R_X7Y121_SLICE_X8Y121_C3 = 1'b1;
  assign CLBLM_R_X7Y121_SLICE_X8Y121_C4 = 1'b1;
  assign CLBLM_R_X5Y112_SLICE_X6Y112_B1 = LIOB33_X0Y81_IOB_X0Y81_I;
  assign CLBLM_R_X5Y112_SLICE_X6Y112_B2 = LIOB33_X0Y111_IOB_X0Y112_I;
  assign CLBLM_R_X5Y112_SLICE_X6Y112_B3 = LIOB33_X0Y109_IOB_X0Y109_I;
  assign CLBLM_R_X5Y112_SLICE_X6Y112_B4 = LIOB33_X0Y95_IOB_X0Y96_I;
  assign CLBLM_R_X5Y112_SLICE_X6Y112_B5 = LIOB33_X0Y79_IOB_X0Y80_I;
  assign CLBLM_R_X5Y112_SLICE_X6Y112_B6 = CLBLM_R_X3Y112_SLICE_X3Y112_AO5;
  assign CLBLM_R_X7Y121_SLICE_X8Y121_C5 = 1'b1;
  assign CLBLM_R_X7Y121_SLICE_X8Y121_C6 = 1'b1;
  assign CLBLM_R_X5Y112_SLICE_X6Y112_C1 = LIOB33_X0Y139_IOB_X0Y139_I;
  assign CLBLM_R_X5Y112_SLICE_X6Y112_C2 = CLBLM_R_X3Y112_SLICE_X3Y112_AO5;
  assign CLBLM_R_X5Y112_SLICE_X6Y112_C3 = CLBLM_R_X5Y111_SLICE_X7Y111_AO5;
  assign CLBLM_R_X5Y112_SLICE_X6Y112_C4 = 1'b1;
  assign CLBLM_R_X5Y112_SLICE_X6Y112_C5 = CLBLL_L_X4Y111_SLICE_X5Y111_AO5;
  assign CLBLM_R_X5Y112_SLICE_X6Y112_C6 = 1'b1;
  assign CLBLM_R_X5Y112_SLICE_X6Y112_D1 = 1'b1;
  assign CLBLM_R_X5Y112_SLICE_X6Y112_D2 = 1'b1;
  assign CLBLM_R_X5Y112_SLICE_X6Y112_D3 = 1'b1;
  assign CLBLM_R_X5Y112_SLICE_X6Y112_D4 = 1'b1;
  assign CLBLM_R_X5Y112_SLICE_X6Y112_D5 = 1'b1;
  assign CLBLM_R_X5Y112_SLICE_X6Y112_D6 = 1'b1;
  assign RIOB33_X105Y77_IOB_X1Y78_O = CLBLL_L_X100Y113_SLICE_X156Y113_BO6;
  assign RIOB33_X105Y77_IOB_X1Y77_O = CLBLL_L_X36Y113_SLICE_X54Y113_BO6;
  assign LIOI3_X0Y197_OLOGIC_X0Y198_D1 = CLBLL_L_X2Y102_SLICE_X0Y102_BO6;
  assign LIOI3_X0Y197_OLOGIC_X0Y198_T1 = 1'b1;
  assign CLBLM_R_X7Y121_SLICE_X8Y121_D1 = 1'b1;
  assign CLBLM_R_X7Y121_SLICE_X8Y121_D2 = 1'b1;
  assign CLBLM_R_X7Y121_SLICE_X8Y121_D3 = 1'b1;
  assign CLBLM_L_X10Y113_SLICE_X13Y113_A1 = CLBLM_R_X5Y110_SLICE_X6Y110_AO6;
  assign CLBLM_L_X10Y113_SLICE_X13Y113_A2 = CLBLM_L_X10Y123_SLICE_X12Y123_AO6;
  assign CLBLM_L_X10Y113_SLICE_X13Y113_A3 = LIOB33_X0Y125_IOB_X0Y125_I;
  assign CLBLM_L_X10Y113_SLICE_X13Y113_A4 = RIOB33_X105Y159_IOB_X1Y160_I;
  assign CLBLM_L_X10Y113_SLICE_X13Y113_A5 = CLBLM_R_X7Y113_SLICE_X8Y113_BO6;
  assign CLBLM_L_X10Y113_SLICE_X13Y113_A6 = CLBLM_R_X7Y113_SLICE_X8Y113_DO6;
  assign CLBLM_R_X7Y121_SLICE_X8Y121_D4 = 1'b1;
  assign LIOI3_X0Y197_OLOGIC_X0Y197_D1 = CLBLL_L_X4Y110_SLICE_X4Y110_CO5;
  assign RIOI3_X105Y179_OLOGIC_X1Y180_D1 = CLBLL_L_X2Y146_SLICE_X1Y146_AO5;
  assign CLBLM_L_X10Y113_SLICE_X13Y113_B1 = CLBLM_R_X5Y110_SLICE_X6Y110_AO6;
  assign CLBLM_L_X10Y113_SLICE_X13Y113_B2 = CLBLM_R_X5Y113_SLICE_X6Y113_AO6;
  assign CLBLM_L_X10Y113_SLICE_X13Y113_B3 = CLBLM_L_X10Y123_SLICE_X12Y123_AO6;
  assign CLBLM_L_X10Y113_SLICE_X13Y113_B4 = RIOB33_X105Y155_IOB_X1Y156_I;
  assign CLBLM_L_X10Y113_SLICE_X13Y113_B5 = LIOB33_X0Y125_IOB_X0Y125_I;
  assign CLBLM_L_X10Y113_SLICE_X13Y113_B6 = CLBLM_R_X5Y112_SLICE_X7Y112_AO6;
  assign LIOI3_X0Y197_OLOGIC_X0Y197_T1 = 1'b1;
  assign RIOB33_X105Y137_IOB_X1Y137_O = CLBLM_R_X101Y123_SLICE_X159Y123_AO6;
  assign RIOB33_X105Y137_IOB_X1Y138_O = CLBLM_R_X103Y123_SLICE_X162Y123_CO6;
  assign CLBLM_L_X10Y113_SLICE_X13Y113_C1 = 1'b1;
  assign CLBLM_L_X10Y113_SLICE_X13Y113_C2 = 1'b1;
  assign CLBLM_L_X10Y113_SLICE_X13Y113_C3 = 1'b1;
  assign CLBLM_L_X10Y113_SLICE_X13Y113_C4 = 1'b1;
  assign CLBLM_L_X10Y113_SLICE_X13Y113_C5 = 1'b1;
  assign CLBLM_L_X10Y113_SLICE_X13Y113_C6 = 1'b1;
  assign RIOI3_X105Y89_OLOGIC_X1Y90_D1 = CLBLM_L_X8Y113_SLICE_X10Y113_DO6;
  assign RIOI3_X105Y179_OLOGIC_X1Y179_D1 = CLBLM_R_X103Y147_SLICE_X163Y147_AO6;
  assign CLBLM_L_X10Y113_SLICE_X13Y113_D1 = 1'b1;
  assign CLBLM_L_X10Y113_SLICE_X13Y113_D2 = 1'b1;
  assign CLBLM_L_X10Y113_SLICE_X13Y113_D3 = 1'b1;
  assign CLBLM_L_X10Y113_SLICE_X13Y113_D4 = 1'b1;
  assign CLBLM_L_X10Y113_SLICE_X13Y113_D5 = 1'b1;
  assign CLBLM_L_X10Y113_SLICE_X13Y113_D6 = 1'b1;
  assign RIOI3_X105Y59_OLOGIC_X1Y60_D1 = CLBLM_L_X10Y113_SLICE_X12Y113_BO6;
  assign RIOI3_X105Y89_OLOGIC_X1Y90_T1 = 1'b1;
  assign RIOI3_X105Y179_OLOGIC_X1Y179_T1 = 1'b1;
  assign CLBLM_L_X10Y113_SLICE_X12Y113_A1 = CLBLM_R_X7Y114_SLICE_X8Y114_AO6;
  assign CLBLM_L_X10Y113_SLICE_X12Y113_A2 = CLBLM_L_X8Y113_SLICE_X11Y113_AO6;
  assign CLBLM_L_X10Y113_SLICE_X12Y113_A3 = RIOB33_SING_X105Y100_IOB_X1Y100_I;
  assign CLBLM_L_X10Y113_SLICE_X12Y113_A4 = LIOB33_X0Y103_IOB_X0Y103_I;
  assign CLBLM_L_X10Y113_SLICE_X12Y113_A5 = CLBLM_L_X10Y123_SLICE_X12Y123_AO6;
  assign CLBLM_L_X10Y113_SLICE_X12Y113_A6 = LIOB33_X0Y131_IOB_X0Y132_I;
  assign CLBLM_L_X10Y113_SLICE_X12Y113_D5 = 1'b1;
  assign CLBLM_L_X10Y113_SLICE_X12Y113_D6 = 1'b1;
  assign RIOB33_X105Y197_IOB_X1Y198_O = CLBLL_L_X2Y173_SLICE_X1Y173_AO6;
  assign RIOB33_X105Y197_IOB_X1Y197_O = CLBLL_L_X2Y173_SLICE_X1Y173_AO6;
  assign CLBLM_L_X10Y113_SLICE_X12Y113_B1 = CLBLM_R_X7Y113_SLICE_X8Y113_CO6;
  assign CLBLM_L_X10Y113_SLICE_X12Y113_B2 = LIOB33_X0Y159_IOB_X0Y160_I;
  assign CLBLM_L_X10Y113_SLICE_X12Y113_B3 = RIOB33_X105Y171_IOB_X1Y172_I;
  assign CLBLM_L_X10Y113_SLICE_X12Y113_B4 = LIOB33_X0Y151_IOB_X0Y151_I;
  assign CLBLM_L_X10Y113_SLICE_X12Y113_B5 = LIOB33_X0Y127_IOB_X0Y127_I;
  assign CLBLM_L_X10Y113_SLICE_X12Y113_B6 = LIOB33_X0Y159_IOB_X0Y159_I;
  assign RIOI3_X105Y59_OLOGIC_X1Y59_D1 = CLBLM_R_X5Y113_SLICE_X6Y113_BO6;
  assign RIOI3_X105Y89_OLOGIC_X1Y89_T1 = 1'b1;
  assign CLBLM_L_X10Y113_SLICE_X12Y113_C1 = CLBLM_L_X10Y123_SLICE_X12Y123_AO6;
  assign CLBLL_L_X4Y109_SLICE_X4Y109_A1 = CLBLL_L_X4Y110_SLICE_X4Y110_DO6;
  assign CLBLL_L_X4Y109_SLICE_X4Y109_A2 = CLBLM_R_X5Y109_SLICE_X6Y109_AO6;
  assign CLBLL_L_X4Y109_SLICE_X4Y109_A3 = CLBLL_L_X2Y136_SLICE_X0Y136_AO6;
  assign CLBLM_L_X10Y113_SLICE_X12Y113_C5 = LIOB33_X0Y85_IOB_X0Y86_I;
  assign CLBLM_L_X10Y113_SLICE_X12Y113_C6 = CLBLM_R_X5Y113_SLICE_X6Y113_AO6;
  assign CLBLL_L_X4Y109_SLICE_X4Y109_A4 = CLBLL_L_X4Y110_SLICE_X4Y110_CO5;
  assign CLBLL_L_X4Y109_SLICE_X4Y109_A5 = CLBLL_L_X2Y102_SLICE_X0Y102_BO6;
  assign CLBLL_L_X4Y109_SLICE_X4Y109_A6 = 1'b1;
  assign CLBLM_L_X10Y113_SLICE_X12Y113_C2 = CLBLM_L_X8Y113_SLICE_X10Y113_AO5;
  assign CLBLM_L_X10Y113_SLICE_X12Y113_C3 = CLBLM_R_X7Y114_SLICE_X8Y114_AO6;
  assign CLBLM_L_X10Y113_SLICE_X12Y113_C4 = RIOB33_X105Y165_IOB_X1Y165_I;
  assign CLBLL_L_X4Y109_SLICE_X4Y109_B1 = LIOB33_X0Y81_IOB_X0Y81_I;
  assign CLBLL_L_X4Y109_SLICE_X4Y109_B2 = LIOB33_X0Y79_IOB_X0Y80_I;
  assign CLBLL_L_X4Y109_SLICE_X4Y109_B3 = LIOB33_X0Y77_IOB_X0Y78_I;
  assign CLBLL_L_X4Y109_SLICE_X4Y109_B4 = LIOB33_X0Y95_IOB_X0Y96_I;
  assign CLBLL_L_X4Y109_SLICE_X4Y109_B5 = LIOB33_X0Y79_IOB_X0Y79_I;
  assign CLBLM_L_X10Y113_SLICE_X12Y113_D3 = 1'b1;
  assign CLBLM_L_X10Y113_SLICE_X12Y113_D4 = 1'b1;
  assign CLBLL_L_X4Y109_SLICE_X4Y109_B6 = 1'b1;
  assign CLBLM_L_X10Y113_SLICE_X12Y113_D1 = 1'b1;
  assign CLBLM_L_X10Y113_SLICE_X12Y113_D2 = 1'b1;
  assign CLBLL_L_X4Y109_SLICE_X4Y109_C1 = LIOB33_X0Y75_IOB_X0Y75_I;
  assign CLBLL_L_X4Y109_SLICE_X4Y109_C2 = CLBLL_L_X4Y110_SLICE_X4Y110_AO5;
  assign CLBLL_L_X4Y109_SLICE_X4Y109_C3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLL_L_X4Y109_SLICE_X4Y109_C4 = LIOB33_X0Y95_IOB_X0Y96_I;
  assign CLBLL_L_X4Y109_SLICE_X4Y109_C5 = CLBLL_L_X4Y109_SLICE_X4Y109_BO5;
  assign CLBLL_L_X4Y109_SLICE_X4Y109_C6 = CLBLL_L_X4Y109_SLICE_X4Y109_BO6;
  assign RIOI3_TBYTESRC_X105Y93_OLOGIC_X1Y93_D1 = CLBLM_L_X10Y113_SLICE_X13Y113_BO6;
  assign CLBLL_L_X4Y109_SLICE_X4Y109_D1 = LIOB33_X0Y103_IOB_X0Y103_I;
  assign CLBLL_L_X4Y109_SLICE_X4Y109_D2 = LIOB33_X0Y93_IOB_X0Y93_I;
  assign CLBLL_L_X4Y109_SLICE_X4Y109_D3 = LIOB33_SING_X0Y99_IOB_X0Y99_I;
  assign CLBLL_L_X4Y109_SLICE_X4Y109_D4 = 1'b1;
  assign CLBLL_L_X4Y109_SLICE_X4Y109_D5 = LIOB33_X0Y101_IOB_X0Y101_I;
  assign CLBLL_L_X4Y109_SLICE_X4Y109_D6 = LIOB33_X0Y105_IOB_X0Y105_I;
  assign RIOI3_TBYTESRC_X105Y93_OLOGIC_X1Y93_T1 = 1'b1;
  assign CLBLL_L_X4Y109_SLICE_X5Y109_A1 = 1'b1;
  assign CLBLL_L_X4Y109_SLICE_X5Y109_A2 = 1'b1;
  assign CLBLL_L_X4Y109_SLICE_X5Y109_A3 = 1'b1;
  assign CLBLL_L_X4Y109_SLICE_X5Y109_A4 = 1'b1;
  assign CLBLL_L_X4Y109_SLICE_X5Y109_A5 = 1'b1;
  assign CLBLL_L_X4Y109_SLICE_X5Y109_A6 = 1'b1;
  assign CLBLL_L_X4Y109_SLICE_X5Y109_B1 = 1'b1;
  assign CLBLL_L_X4Y109_SLICE_X5Y109_B2 = 1'b1;
  assign CLBLL_L_X4Y109_SLICE_X5Y109_B3 = 1'b1;
  assign CLBLL_L_X4Y109_SLICE_X5Y109_B4 = 1'b1;
  assign CLBLL_L_X4Y109_SLICE_X5Y109_B5 = 1'b1;
  assign CLBLL_L_X4Y109_SLICE_X5Y109_B6 = 1'b1;
  assign CLBLL_L_X4Y109_SLICE_X5Y109_C1 = 1'b1;
  assign CLBLL_L_X4Y109_SLICE_X5Y109_C2 = 1'b1;
  assign CLBLL_L_X4Y109_SLICE_X5Y109_C3 = 1'b1;
  assign CLBLL_L_X4Y109_SLICE_X5Y109_C4 = 1'b1;
  assign CLBLL_L_X4Y109_SLICE_X5Y109_C5 = 1'b1;
  assign CLBLL_L_X4Y109_SLICE_X5Y109_C6 = 1'b1;
  assign CLBLL_L_X4Y109_SLICE_X5Y109_D1 = 1'b1;
  assign CLBLL_L_X4Y109_SLICE_X5Y109_D2 = 1'b1;
  assign CLBLL_L_X4Y109_SLICE_X5Y109_D3 = 1'b1;
  assign CLBLL_L_X4Y109_SLICE_X5Y109_D4 = 1'b1;
  assign CLBLL_L_X4Y109_SLICE_X5Y109_D5 = 1'b1;
  assign CLBLL_L_X4Y109_SLICE_X5Y109_D6 = 1'b1;
  assign CLBLM_R_X5Y113_SLICE_X7Y113_A1 = CLBLM_R_X5Y112_SLICE_X7Y112_AO5;
  assign CLBLM_R_X5Y113_SLICE_X7Y113_A2 = LIOB33_X0Y131_IOB_X0Y131_I;
  assign CLBLM_R_X5Y113_SLICE_X7Y113_A3 = LIOB33_X0Y101_IOB_X0Y101_I;
  assign CLBLM_R_X5Y113_SLICE_X7Y113_A4 = CLBLM_R_X5Y113_SLICE_X7Y113_BO6;
  assign CLBLM_R_X5Y113_SLICE_X7Y113_A5 = CLBLM_R_X5Y115_SLICE_X6Y115_AO6;
  assign CLBLM_R_X5Y113_SLICE_X7Y113_A6 = CLBLM_R_X5Y113_SLICE_X7Y113_CO6;
  assign CLBLM_R_X5Y113_SLICE_X7Y113_B1 = CLBLM_R_X5Y112_SLICE_X7Y112_AO6;
  assign CLBLM_R_X5Y113_SLICE_X7Y113_B2 = CLBLM_R_X7Y113_SLICE_X8Y113_BO6;
  assign CLBLM_R_X5Y113_SLICE_X7Y113_B3 = LIOB33_X0Y83_IOB_X0Y84_I;
  assign CLBLM_R_X5Y113_SLICE_X7Y113_B4 = LIOB33_X0Y65_IOB_X0Y66_I;
  assign CLBLM_R_X5Y113_SLICE_X7Y113_B5 = LIOB33_X0Y85_IOB_X0Y86_I;
  assign CLBLM_R_X5Y113_SLICE_X7Y113_B6 = LIOB33_X0Y71_IOB_X0Y71_I;
  assign LIOI3_X0Y135_ILOGIC_X0Y136_D = LIOB33_X0Y135_IOB_X0Y136_I;
  assign LIOI3_X0Y135_ILOGIC_X0Y135_D = LIOB33_X0Y135_IOB_X0Y135_I;
  assign LIOI3_X0Y105_ILOGIC_X0Y106_D = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLM_R_X5Y113_SLICE_X7Y113_C1 = LIOB33_X0Y125_IOB_X0Y126_I;
  assign CLBLM_R_X5Y113_SLICE_X7Y113_C2 = LIOB33_X0Y127_IOB_X0Y127_I;
  assign CLBLM_R_X5Y113_SLICE_X7Y113_C3 = LIOB33_SING_X0Y99_IOB_X0Y99_I;
  assign CLBLM_R_X5Y113_SLICE_X7Y113_C4 = LIOB33_X0Y129_IOB_X0Y129_I;
  assign CLBLM_R_X5Y113_SLICE_X7Y113_C5 = LIOB33_X0Y151_IOB_X0Y151_I;
  assign CLBLM_R_X5Y113_SLICE_X7Y113_C6 = LIOB33_X0Y93_IOB_X0Y93_I;
  assign LIOI3_X0Y105_ILOGIC_X0Y105_D = LIOB33_X0Y105_IOB_X0Y105_I;
  assign LIOI3_X0Y75_ILOGIC_X0Y76_D = LIOB33_X0Y75_IOB_X0Y76_I;
  assign LIOI3_X0Y75_ILOGIC_X0Y75_D = LIOB33_X0Y75_IOB_X0Y75_I;
  assign RIOI3_X105Y151_ILOGIC_X1Y152_D = RIOB33_X105Y151_IOB_X1Y152_I;
  assign CLBLM_R_X5Y113_SLICE_X7Y113_D1 = LIOB33_X0Y125_IOB_X0Y126_I;
  assign CLBLM_R_X5Y113_SLICE_X7Y113_D2 = LIOB33_X0Y67_IOB_X0Y68_I;
  assign CLBLM_R_X5Y113_SLICE_X7Y113_D3 = LIOB33_X0Y93_IOB_X0Y93_I;
  assign CLBLM_R_X5Y113_SLICE_X7Y113_D4 = LIOB33_X0Y69_IOB_X0Y70_I;
  assign CLBLM_R_X5Y113_SLICE_X7Y113_D5 = LIOB33_X0Y103_IOB_X0Y103_I;
  assign CLBLM_R_X5Y113_SLICE_X7Y113_D6 = LIOB33_X0Y127_IOB_X0Y127_I;
  assign RIOI3_X105Y151_ILOGIC_X1Y151_D = RIOB33_X105Y151_IOB_X1Y151_I;
  assign RIOI3_X105Y121_ILOGIC_X1Y122_D = RIOB33_X105Y121_IOB_X1Y122_I;
  assign RIOI3_X105Y121_ILOGIC_X1Y121_D = RIOB33_X105Y121_IOB_X1Y121_I;
  assign CLBLM_R_X5Y113_SLICE_X6Y113_A1 = CLBLM_R_X5Y113_SLICE_X6Y113_DO6;
  assign CLBLM_R_X5Y113_SLICE_X6Y113_A2 = LIOB33_X0Y93_IOB_X0Y93_I;
  assign CLBLM_R_X5Y113_SLICE_X6Y113_A3 = LIOB33_X0Y125_IOB_X0Y126_I;
  assign CLBLM_R_X5Y113_SLICE_X6Y113_A4 = LIOB33_X0Y93_IOB_X0Y94_I;
  assign CLBLM_R_X5Y113_SLICE_X6Y113_A5 = LIOB33_X0Y95_IOB_X0Y95_I;
  assign CLBLM_R_X5Y113_SLICE_X6Y113_A6 = 1'b1;
  assign LIOI3_TBYTETERM_X0Y113_ILOGIC_X0Y114_D = LIOB33_X0Y113_IOB_X0Y114_I;
  assign LIOI3_TBYTETERM_X0Y113_ILOGIC_X0Y113_D = LIOB33_X0Y113_IOB_X0Y113_I;
  assign CLBLM_R_X5Y113_SLICE_X6Y113_B1 = LIOB33_X0Y127_IOB_X0Y128_I;
  assign CLBLM_R_X5Y113_SLICE_X6Y113_B2 = LIOB33_X0Y93_IOB_X0Y93_I;
  assign CLBLM_R_X5Y113_SLICE_X6Y113_B3 = LIOB33_X0Y125_IOB_X0Y126_I;
  assign CLBLM_R_X5Y113_SLICE_X6Y113_B4 = CLBLM_L_X10Y123_SLICE_X12Y123_AO6;
  assign CLBLM_R_X5Y113_SLICE_X6Y113_B5 = CLBLM_R_X5Y115_SLICE_X6Y115_AO6;
  assign CLBLM_R_X5Y113_SLICE_X6Y113_B6 = CLBLM_R_X5Y113_SLICE_X6Y113_AO5;
  assign RIOB33_X105Y79_IOB_X1Y79_O = CLBLM_R_X29Y115_SLICE_X42Y115_BO6;
  assign CLBLM_R_X5Y113_SLICE_X6Y113_C1 = CLBLM_R_X5Y115_SLICE_X6Y115_AO6;
  assign CLBLM_R_X5Y113_SLICE_X6Y113_C2 = RIOB33_X105Y169_IOB_X1Y170_I;
  assign CLBLM_R_X5Y113_SLICE_X6Y113_C3 = LIOB33_X0Y71_IOB_X0Y72_I;
  assign CLBLM_R_X5Y113_SLICE_X6Y113_C4 = CLBLM_L_X10Y123_SLICE_X12Y123_AO6;
  assign CLBLM_R_X5Y113_SLICE_X6Y113_C5 = LIOB33_X0Y111_IOB_X0Y111_I;
  assign CLBLM_R_X5Y113_SLICE_X6Y113_C6 = CLBLL_L_X4Y112_SLICE_X4Y112_CO6;
  assign RIOB33_X105Y79_IOB_X1Y80_O = CLBLM_R_X103Y97_SLICE_X163Y97_AO6;
  assign RIOI3_SING_X105Y99_OLOGIC_X1Y99_D1 = CLBLM_R_X101Y119_SLICE_X158Y119_BO6;
  assign CLBLM_R_X5Y113_SLICE_X6Y113_D1 = LIOB33_X0Y95_IOB_X0Y95_I;
  assign CLBLM_R_X5Y113_SLICE_X6Y113_D2 = LIOB33_X0Y129_IOB_X0Y129_I;
  assign CLBLM_R_X5Y113_SLICE_X6Y113_D3 = LIOB33_X0Y131_IOB_X0Y131_I;
  assign CLBLM_R_X5Y113_SLICE_X6Y113_D4 = 1'b1;
  assign CLBLM_R_X5Y113_SLICE_X6Y113_D5 = 1'b1;
  assign CLBLM_R_X5Y113_SLICE_X6Y113_D6 = LIOB33_X0Y127_IOB_X0Y127_I;
  assign RIOI3_SING_X105Y99_OLOGIC_X1Y99_T1 = 1'b1;
  assign LIOI3_X0Y145_ILOGIC_X0Y146_D = LIOB33_X0Y145_IOB_X0Y146_I;
  assign RIOB33_X105Y139_IOB_X1Y140_O = CLBLM_R_X101Y118_SLICE_X158Y118_DO6;
  assign RIOB33_X105Y139_IOB_X1Y139_O = CLBLM_R_X101Y119_SLICE_X158Y119_DO6;
  assign LIOI3_X0Y145_ILOGIC_X0Y145_D = LIOB33_X0Y145_IOB_X0Y145_I;
  assign CLBLM_L_X10Y114_SLICE_X13Y114_A1 = 1'b1;
  assign CLBLM_L_X10Y114_SLICE_X13Y114_A2 = 1'b1;
  assign CLBLM_L_X10Y114_SLICE_X13Y114_A3 = 1'b1;
  assign CLBLM_L_X10Y114_SLICE_X13Y114_A4 = 1'b1;
  assign CLBLM_L_X10Y114_SLICE_X13Y114_A5 = 1'b1;
  assign CLBLM_L_X10Y114_SLICE_X13Y114_A6 = 1'b1;
  assign CLBLM_L_X10Y114_SLICE_X13Y114_B1 = 1'b1;
  assign CLBLM_L_X10Y114_SLICE_X13Y114_B2 = 1'b1;
  assign CLBLM_L_X10Y114_SLICE_X13Y114_B3 = 1'b1;
  assign CLBLM_L_X10Y114_SLICE_X13Y114_B4 = 1'b1;
  assign CLBLM_L_X10Y114_SLICE_X13Y114_B5 = 1'b1;
  assign CLBLM_L_X10Y114_SLICE_X13Y114_B6 = 1'b1;
  assign CLBLM_L_X10Y114_SLICE_X13Y114_C1 = 1'b1;
  assign CLBLM_L_X10Y114_SLICE_X13Y114_C2 = 1'b1;
  assign CLBLM_L_X10Y114_SLICE_X13Y114_C3 = 1'b1;
  assign CLBLM_L_X10Y114_SLICE_X13Y114_C4 = 1'b1;
  assign CLBLM_L_X10Y114_SLICE_X13Y114_C5 = 1'b1;
  assign CLBLM_L_X10Y114_SLICE_X13Y114_C6 = 1'b1;
  assign RIOI3_X105Y117_ILOGIC_X1Y117_D = RIOB33_X105Y117_IOB_X1Y117_I;
  assign CLBLM_L_X10Y114_SLICE_X13Y114_D1 = 1'b1;
  assign CLBLM_L_X10Y114_SLICE_X13Y114_D2 = 1'b1;
  assign CLBLM_L_X10Y114_SLICE_X13Y114_D3 = 1'b1;
  assign CLBLM_L_X10Y114_SLICE_X13Y114_D4 = 1'b1;
  assign CLBLM_L_X10Y114_SLICE_X13Y114_D5 = 1'b1;
  assign CLBLM_L_X10Y114_SLICE_X13Y114_D6 = 1'b1;
  assign CLBLM_L_X10Y114_SLICE_X12Y114_A1 = RIOB33_X105Y171_IOB_X1Y171_I;
  assign CLBLM_L_X10Y114_SLICE_X12Y114_A2 = LIOB33_X0Y131_IOB_X0Y132_I;
  assign CLBLM_L_X10Y114_SLICE_X12Y114_A3 = CLBLM_L_X10Y123_SLICE_X12Y123_AO6;
  assign CLBLM_L_X10Y114_SLICE_X12Y114_A4 = CLBLM_R_X7Y114_SLICE_X9Y114_AO6;
  assign CLBLM_L_X10Y114_SLICE_X12Y114_A5 = CLBLM_L_X8Y113_SLICE_X11Y113_AO6;
  assign CLBLM_L_X10Y114_SLICE_X12Y114_A6 = CLBLM_R_X7Y114_SLICE_X8Y114_BO5;
  assign CLBLM_L_X10Y114_SLICE_X12Y114_B1 = CLBLL_L_X4Y111_SLICE_X5Y111_AO5;
  assign CLBLL_L_X2Y175_SLICE_X0Y175_A1 = 1'b1;
  assign CLBLL_L_X2Y175_SLICE_X0Y175_A2 = 1'b1;
  assign CLBLM_L_X10Y114_SLICE_X12Y114_B2 = CLBLM_R_X5Y114_SLICE_X7Y114_AO5;
  assign CLBLM_L_X10Y114_SLICE_X12Y114_B3 = RIOB33_X105Y159_IOB_X1Y159_I;
  assign CLBLM_L_X10Y114_SLICE_X12Y114_B6 = LIOB33_X0Y159_IOB_X0Y159_I;
  assign CLBLL_L_X2Y175_SLICE_X0Y175_A5 = LIOB33_X0Y135_IOB_X0Y135_I;
  assign CLBLL_L_X2Y175_SLICE_X0Y175_A6 = 1'b1;
  assign CLBLM_L_X10Y114_SLICE_X12Y114_B4 = LIOB33_X0Y159_IOB_X0Y160_I;
  assign CLBLL_L_X4Y110_SLICE_X4Y110_A3 = LIOB33_X0Y95_IOB_X0Y96_I;
  assign CLBLL_L_X4Y110_SLICE_X4Y110_A5 = LIOB33_X0Y75_IOB_X0Y75_I;
  assign CLBLM_L_X10Y114_SLICE_X12Y114_B5 = CLBLM_R_X5Y111_SLICE_X6Y111_AO6;
  assign CLBLL_L_X2Y175_SLICE_X0Y175_A4 = 1'b1;
  assign CLBLL_L_X4Y110_SLICE_X4Y110_A1 = LIOB33_X0Y73_IOB_X0Y74_I;
  assign CLBLL_L_X4Y110_SLICE_X4Y110_A2 = LIOB33_X0Y71_IOB_X0Y72_I;
  assign CLBLL_L_X2Y175_SLICE_X0Y175_B6 = 1'b1;
  assign CLBLL_L_X4Y110_SLICE_X4Y110_B2 = LIOB33_X0Y79_IOB_X0Y80_I;
  assign CLBLL_L_X4Y110_SLICE_X4Y110_B3 = LIOB33_X0Y109_IOB_X0Y109_I;
  assign CLBLL_L_X4Y110_SLICE_X4Y110_B4 = LIOB33_X0Y95_IOB_X0Y96_I;
  assign CLBLL_L_X2Y175_SLICE_X0Y175_C1 = 1'b1;
  assign CLBLL_L_X2Y175_SLICE_X0Y175_C2 = 1'b1;
  assign CLBLL_L_X2Y175_SLICE_X0Y175_C3 = 1'b1;
  assign CLBLL_L_X2Y175_SLICE_X0Y175_C4 = 1'b1;
  assign CLBLL_L_X2Y175_SLICE_X0Y175_C5 = 1'b1;
  assign CLBLL_L_X2Y175_SLICE_X0Y175_C6 = 1'b1;
  assign CLBLL_L_X4Y110_SLICE_X4Y110_B5 = LIOB33_X0Y111_IOB_X0Y112_I;
  assign CLBLL_L_X4Y110_SLICE_X4Y110_B6 = 1'b1;
  assign CLBLL_L_X4Y110_SLICE_X4Y110_C1 = LIOB33_X0Y91_IOB_X0Y91_I;
  assign CLBLM_L_X10Y114_SLICE_X12Y114_D1 = 1'b1;
  assign CLBLL_L_X4Y110_SLICE_X4Y110_C2 = LIOB33_X0Y83_IOB_X0Y84_I;
  assign CLBLM_L_X10Y114_SLICE_X12Y114_D3 = 1'b1;
  assign CLBLM_L_X10Y114_SLICE_X12Y114_D4 = 1'b1;
  assign CLBLM_L_X10Y114_SLICE_X12Y114_D2 = 1'b1;
  assign CLBLL_L_X4Y110_SLICE_X4Y110_C3 = LIOB33_X0Y87_IOB_X0Y88_I;
  assign CLBLL_L_X4Y110_SLICE_X4Y110_C5 = LIOB33_X0Y85_IOB_X0Y86_I;
  assign CLBLL_L_X4Y110_SLICE_X4Y110_C6 = 1'b1;
  assign CLBLM_L_X10Y114_SLICE_X12Y114_D6 = 1'b1;
  assign CLBLL_L_X2Y175_SLICE_X0Y175_D1 = 1'b1;
  assign CLBLL_L_X2Y175_SLICE_X0Y175_D2 = 1'b1;
  assign CLBLL_L_X2Y175_SLICE_X0Y175_D3 = 1'b1;
  assign CLBLL_L_X2Y175_SLICE_X0Y175_D4 = 1'b1;
  assign CLBLL_L_X2Y175_SLICE_X0Y175_D5 = 1'b1;
  assign CLBLL_L_X2Y175_SLICE_X0Y175_D6 = 1'b1;
  assign CLBLL_L_X4Y110_SLICE_X4Y110_D1 = CLBLM_R_X3Y111_SLICE_X2Y111_AO6;
  assign CLBLL_L_X4Y110_SLICE_X4Y110_D2 = CLBLL_L_X2Y98_SLICE_X0Y98_AO6;
  assign CLBLL_L_X4Y110_SLICE_X4Y110_D3 = CLBLM_R_X3Y111_SLICE_X3Y111_BO6;
  assign CLBLL_L_X4Y110_SLICE_X4Y110_D4 = CLBLL_L_X4Y109_SLICE_X4Y109_CO6;
  assign CLBLL_L_X4Y110_SLICE_X4Y110_D5 = CLBLM_R_X3Y110_SLICE_X3Y110_AO5;
  assign CLBLL_L_X4Y110_SLICE_X4Y110_D6 = CLBLM_R_X3Y110_SLICE_X3Y110_AO6;
  assign CLBLL_L_X2Y175_SLICE_X1Y175_A1 = 1'b1;
  assign CLBLL_L_X2Y175_SLICE_X1Y175_A2 = 1'b1;
  assign CLBLL_L_X2Y175_SLICE_X1Y175_A3 = 1'b1;
  assign CLBLL_L_X2Y175_SLICE_X1Y175_A4 = 1'b1;
  assign CLBLL_L_X2Y175_SLICE_X1Y175_A5 = 1'b1;
  assign CLBLL_L_X2Y175_SLICE_X1Y175_A6 = 1'b1;
  assign CLBLL_L_X4Y110_SLICE_X5Y110_A1 = 1'b1;
  assign CLBLL_L_X4Y110_SLICE_X5Y110_A2 = 1'b1;
  assign CLBLL_L_X4Y110_SLICE_X5Y110_A4 = 1'b1;
  assign CLBLL_L_X4Y110_SLICE_X5Y110_A5 = 1'b1;
  assign CLBLL_L_X4Y110_SLICE_X5Y110_A3 = 1'b1;
  assign CLBLL_L_X4Y110_SLICE_X5Y110_A6 = 1'b1;
  assign CLBLL_L_X2Y175_SLICE_X1Y175_B1 = 1'b1;
  assign CLBLL_L_X2Y175_SLICE_X1Y175_B2 = 1'b1;
  assign CLBLL_L_X2Y175_SLICE_X1Y175_B3 = 1'b1;
  assign CLBLL_L_X4Y110_SLICE_X5Y110_B1 = 1'b1;
  assign CLBLL_L_X2Y175_SLICE_X1Y175_B4 = 1'b1;
  assign CLBLL_L_X4Y110_SLICE_X5Y110_B4 = 1'b1;
  assign CLBLL_L_X2Y175_SLICE_X1Y175_B5 = 1'b1;
  assign CLBLL_L_X4Y110_SLICE_X5Y110_B6 = 1'b1;
  assign CLBLL_L_X2Y175_SLICE_X1Y175_B6 = 1'b1;
  assign CLBLL_L_X4Y110_SLICE_X5Y110_B2 = 1'b1;
  assign CLBLL_L_X4Y110_SLICE_X5Y110_B3 = 1'b1;
  assign CLBLL_L_X2Y175_SLICE_X1Y175_C1 = 1'b1;
  assign CLBLL_L_X2Y175_SLICE_X1Y175_C2 = 1'b1;
  assign CLBLL_L_X2Y175_SLICE_X1Y175_C3 = 1'b1;
  assign CLBLL_L_X2Y175_SLICE_X1Y175_C4 = 1'b1;
  assign CLBLL_L_X2Y175_SLICE_X1Y175_C5 = 1'b1;
  assign CLBLL_L_X2Y175_SLICE_X1Y175_C6 = 1'b1;
  assign CLBLL_L_X4Y110_SLICE_X5Y110_C5 = 1'b1;
  assign CLBLL_L_X4Y110_SLICE_X5Y110_C6 = 1'b1;
  assign CLBLL_L_X4Y110_SLICE_X5Y110_C1 = 1'b1;
  assign CLBLL_L_X4Y110_SLICE_X5Y110_C2 = 1'b1;
  assign CLBLL_L_X4Y110_SLICE_X5Y110_C3 = 1'b1;
  assign CLBLL_L_X4Y110_SLICE_X5Y110_C4 = 1'b1;
  assign CLBLL_L_X2Y175_SLICE_X1Y175_D1 = 1'b1;
  assign CLBLL_L_X2Y175_SLICE_X1Y175_D2 = 1'b1;
  assign CLBLL_L_X4Y110_SLICE_X5Y110_D1 = 1'b1;
  assign CLBLL_L_X2Y175_SLICE_X1Y175_D3 = 1'b1;
  assign CLBLL_L_X2Y175_SLICE_X1Y175_D4 = 1'b1;
  assign CLBLL_L_X2Y175_SLICE_X1Y175_D5 = 1'b1;
  assign CLBLL_L_X2Y175_SLICE_X1Y175_D6 = 1'b1;
  assign CLBLL_L_X4Y110_SLICE_X5Y110_D2 = 1'b1;
  assign CLBLL_L_X4Y110_SLICE_X5Y110_D3 = 1'b1;
  assign CLBLL_L_X4Y110_SLICE_X5Y110_D4 = 1'b1;
  assign CLBLL_L_X4Y110_SLICE_X5Y110_D5 = 1'b1;
  assign CLBLL_L_X4Y110_SLICE_X5Y110_D6 = 1'b1;
  assign CLBLM_R_X5Y114_SLICE_X7Y114_A1 = LIOB33_X0Y119_IOB_X0Y119_I;
  assign CLBLM_R_X5Y114_SLICE_X7Y114_A2 = LIOB33_X0Y69_IOB_X0Y70_I;
  assign CLBLM_R_X5Y114_SLICE_X7Y114_A3 = RIOB33_X105Y159_IOB_X1Y159_I;
  assign CLBLM_R_X5Y114_SLICE_X7Y114_A4 = LIOB33_X0Y53_IOB_X0Y54_I;
  assign CLBLM_R_X5Y114_SLICE_X7Y114_A5 = LIOB33_X0Y67_IOB_X0Y68_I;
  assign CLBLM_R_X5Y114_SLICE_X7Y114_A6 = 1'b1;
  assign LIOI3_X0Y175_ILOGIC_X0Y176_D = LIOB33_X0Y175_IOB_X0Y176_I;
  assign CLBLM_R_X5Y114_SLICE_X7Y114_B1 = 1'b1;
  assign CLBLM_R_X5Y114_SLICE_X7Y114_B2 = 1'b1;
  assign CLBLM_R_X5Y114_SLICE_X7Y114_B3 = 1'b1;
  assign CLBLM_R_X5Y114_SLICE_X7Y114_B4 = 1'b1;
  assign CLBLM_R_X5Y114_SLICE_X7Y114_B5 = 1'b1;
  assign CLBLM_R_X5Y114_SLICE_X7Y114_B6 = 1'b1;
  assign CLBLM_R_X5Y114_SLICE_X7Y114_C1 = 1'b1;
  assign CLBLM_R_X5Y114_SLICE_X7Y114_C2 = 1'b1;
  assign CLBLM_R_X5Y114_SLICE_X7Y114_C3 = 1'b1;
  assign CLBLM_R_X5Y114_SLICE_X7Y114_C4 = 1'b1;
  assign CLBLM_R_X5Y114_SLICE_X7Y114_C5 = 1'b1;
  assign CLBLM_R_X5Y114_SLICE_X7Y114_C6 = 1'b1;
  assign LIOI3_X0Y175_ILOGIC_X0Y175_D = LIOB33_X0Y175_IOB_X0Y175_I;
  assign CLBLM_R_X5Y114_SLICE_X7Y114_D1 = 1'b1;
  assign CLBLM_R_X5Y114_SLICE_X7Y114_D2 = 1'b1;
  assign CLBLM_R_X5Y114_SLICE_X7Y114_D3 = 1'b1;
  assign CLBLM_R_X5Y114_SLICE_X7Y114_D4 = 1'b1;
  assign CLBLM_R_X5Y114_SLICE_X7Y114_D5 = 1'b1;
  assign CLBLM_R_X5Y114_SLICE_X7Y114_D6 = 1'b1;
  assign RIOB33_X105Y81_IOB_X1Y81_O = CLBLM_R_X103Y122_SLICE_X163Y122_CO6;
  assign RIOB33_X105Y81_IOB_X1Y82_O = CLBLM_R_X103Y107_SLICE_X163Y107_BO6;
  assign CLBLM_R_X5Y114_SLICE_X6Y114_A1 = CLBLM_R_X5Y114_SLICE_X7Y114_AO5;
  assign CLBLM_R_X5Y114_SLICE_X6Y114_A2 = LIOB33_X0Y57_IOB_X0Y58_I;
  assign CLBLM_R_X5Y114_SLICE_X6Y114_A3 = CLBLL_L_X4Y113_SLICE_X5Y113_AO6;
  assign CLBLM_R_X5Y114_SLICE_X6Y114_A4 = CLBLM_R_X5Y114_SLICE_X6Y114_BO6;
  assign CLBLM_R_X5Y114_SLICE_X6Y114_A5 = LIOB33_X0Y121_IOB_X0Y122_I;
  assign CLBLM_R_X5Y114_SLICE_X6Y114_A6 = CLBLM_R_X5Y111_SLICE_X7Y111_DO6;
  assign CLBLM_R_X5Y114_SLICE_X6Y114_B1 = LIOB33_X0Y71_IOB_X0Y72_I;
  assign CLBLM_R_X5Y114_SLICE_X6Y114_B2 = LIOB33_X0Y117_IOB_X0Y118_I;
  assign CLBLM_R_X5Y114_SLICE_X6Y114_B3 = LIOB33_SING_X0Y150_IOB_X0Y150_I;
  assign CLBLM_R_X5Y114_SLICE_X6Y114_B4 = LIOB33_X0Y151_IOB_X0Y151_I;
  assign CLBLM_R_X5Y114_SLICE_X6Y114_B5 = LIOB33_X0Y111_IOB_X0Y111_I;
  assign CLBLM_R_X5Y114_SLICE_X6Y114_B6 = LIOB33_X0Y63_IOB_X0Y63_I;
  assign CLBLM_R_X5Y114_SLICE_X6Y114_C1 = LIOB33_X0Y121_IOB_X0Y122_I;
  assign CLBLM_R_X5Y114_SLICE_X6Y114_C2 = CLBLL_L_X4Y113_SLICE_X5Y113_AO6;
  assign CLBLM_R_X5Y114_SLICE_X6Y114_C3 = LIOB33_X0Y57_IOB_X0Y58_I;
  assign CLBLM_R_X5Y114_SLICE_X6Y114_C4 = CLBLM_R_X7Y114_SLICE_X8Y114_AO6;
  assign CLBLM_R_X5Y114_SLICE_X6Y114_C5 = CLBLM_R_X5Y114_SLICE_X6Y114_DO6;
  assign CLBLM_R_X5Y114_SLICE_X6Y114_C6 = CLBLM_R_X5Y111_SLICE_X7Y111_DO6;
  assign RIOB33_X105Y141_IOB_X1Y142_O = CLBLM_R_X103Y123_SLICE_X162Y123_DO6;
  assign RIOB33_X105Y141_IOB_X1Y141_O = CLBLM_R_X101Y123_SLICE_X159Y123_BO6;
  assign CLBLM_R_X5Y114_SLICE_X6Y114_D1 = 1'b1;
  assign CLBLM_R_X5Y114_SLICE_X6Y114_D2 = CLBLM_R_X5Y114_SLICE_X7Y114_AO5;
  assign CLBLM_R_X5Y114_SLICE_X6Y114_D3 = LIOB33_X0Y111_IOB_X0Y111_I;
  assign CLBLM_R_X5Y114_SLICE_X6Y114_D4 = LIOB33_X0Y63_IOB_X0Y63_I;
  assign CLBLM_R_X5Y114_SLICE_X6Y114_D5 = LIOB33_X0Y71_IOB_X0Y72_I;
  assign CLBLM_R_X5Y114_SLICE_X6Y114_D6 = LIOB33_X0Y117_IOB_X0Y118_I;
  assign RIOB33_X105Y89_IOB_X1Y89_O = CLBLM_R_X49Y101_SLICE_X74Y101_AO5;
  assign RIOB33_X105Y89_IOB_X1Y90_O = CLBLM_L_X8Y113_SLICE_X10Y113_DO6;
  assign RIOI3_TBYTETERM_X105Y63_OLOGIC_X1Y64_T1 = 1'b1;
  assign RIOI3_X105Y173_OLOGIC_X1Y173_T1 = 1'b1;
  assign RIOI3_SING_X105Y50_OLOGIC_X1Y50_D1 = CLBLM_R_X49Y95_SLICE_X74Y95_AO6;
  assign CLBLL_L_X4Y111_SLICE_X4Y111_A1 = LIOB33_X0Y59_IOB_X0Y59_I;
  assign CLBLL_L_X4Y111_SLICE_X4Y111_A2 = LIOB33_X0Y57_IOB_X0Y58_I;
  assign CLBLL_L_X4Y111_SLICE_X4Y111_A3 = LIOB33_X0Y121_IOB_X0Y122_I;
  assign CLBLL_L_X4Y111_SLICE_X4Y111_A4 = CLBLM_R_X3Y111_SLICE_X2Y111_AO5;
  assign CLBLL_L_X4Y111_SLICE_X4Y111_A5 = LIOB33_X0Y95_IOB_X0Y96_I;
  assign CLBLL_L_X4Y111_SLICE_X4Y111_A6 = 1'b1;
  assign CLBLL_L_X4Y111_SLICE_X4Y111_B1 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLL_L_X4Y111_SLICE_X4Y111_B2 = LIOB33_X0Y59_IOB_X0Y60_I;
  assign CLBLL_L_X4Y111_SLICE_X4Y111_B3 = LIOB33_X0Y95_IOB_X0Y96_I;
  assign CLBLL_L_X4Y111_SLICE_X4Y111_B4 = CLBLL_L_X4Y111_SLICE_X5Y111_AO5;
  assign CLBLL_L_X4Y111_SLICE_X4Y111_B5 = CLBLL_L_X4Y111_SLICE_X4Y111_AO6;
  assign CLBLL_L_X4Y111_SLICE_X4Y111_B6 = LIOB33_X0Y115_IOB_X0Y116_I;
  assign CLBLL_L_X4Y111_SLICE_X4Y111_C1 = CLBLL_L_X4Y110_SLICE_X4Y110_BO6;
  assign CLBLL_L_X4Y111_SLICE_X4Y111_C2 = LIOB33_X0Y77_IOB_X0Y78_I;
  assign CLBLL_L_X4Y111_SLICE_X4Y111_C3 = LIOB33_X0Y79_IOB_X0Y79_I;
  assign CLBLL_L_X4Y111_SLICE_X4Y111_C4 = LIOB33_X0Y115_IOB_X0Y115_I;
  assign CLBLL_L_X4Y111_SLICE_X4Y111_C5 = LIOB33_X0Y95_IOB_X0Y96_I;
  assign CLBLL_L_X4Y111_SLICE_X4Y111_C6 = CLBLM_R_X3Y111_SLICE_X3Y111_AO6;
  assign CLBLL_L_X4Y111_SLICE_X4Y111_D1 = LIOB33_X0Y111_IOB_X0Y111_I;
  assign CLBLL_L_X4Y111_SLICE_X4Y111_D2 = CLBLL_L_X4Y110_SLICE_X4Y110_AO5;
  assign CLBLL_L_X4Y111_SLICE_X4Y111_D3 = CLBLL_L_X4Y111_SLICE_X4Y111_AO5;
  assign CLBLL_L_X4Y111_SLICE_X4Y111_D4 = LIOB33_X0Y115_IOB_X0Y116_I;
  assign CLBLL_L_X4Y111_SLICE_X4Y111_D5 = CLBLM_R_X3Y111_SLICE_X3Y111_AO5;
  assign CLBLL_L_X4Y111_SLICE_X4Y111_D6 = CLBLM_R_X3Y110_SLICE_X3Y110_AO6;
  assign RIOI3_SING_X105Y100_ILOGIC_X1Y100_D = RIOB33_SING_X105Y100_IOB_X1Y100_I;
  assign RIOI3_X105Y183_OLOGIC_X1Y184_D1 = RIOB33_SING_X105Y150_IOB_X1Y150_I;
  assign CLBLL_L_X4Y111_SLICE_X5Y111_A1 = LIOB33_X0Y53_IOB_X0Y54_I;
  assign CLBLL_L_X4Y111_SLICE_X5Y111_A2 = LIOB33_X0Y119_IOB_X0Y119_I;
  assign CLBLL_L_X4Y111_SLICE_X5Y111_A3 = CLBLM_R_X3Y111_SLICE_X3Y111_DO6;
  assign CLBLL_L_X4Y111_SLICE_X5Y111_A4 = LIOB33_X0Y55_IOB_X0Y55_I;
  assign CLBLL_L_X4Y111_SLICE_X5Y111_A5 = LIOB33_X0Y95_IOB_X0Y96_I;
  assign CLBLL_L_X4Y111_SLICE_X5Y111_A6 = 1'b1;
  assign RIOI3_X105Y183_OLOGIC_X1Y184_T1 = 1'b1;
  assign CLBLM_R_X3Y110_SLICE_X3Y110_B3 = 1'b1;
  assign CLBLL_L_X4Y111_SLICE_X5Y111_B1 = LIOB33_X0Y73_IOB_X0Y74_I;
  assign CLBLL_L_X4Y111_SLICE_X5Y111_B2 = CLBLL_L_X4Y112_SLICE_X5Y112_BO6;
  assign CLBLL_L_X4Y111_SLICE_X5Y111_B3 = LIOB33_X0Y71_IOB_X0Y72_I;
  assign CLBLL_L_X4Y111_SLICE_X5Y111_B4 = LIOB33_X0Y111_IOB_X0Y111_I;
  assign CLBLL_L_X4Y111_SLICE_X5Y111_B5 = LIOB33_X0Y95_IOB_X0Y96_I;
  assign CLBLL_L_X4Y111_SLICE_X5Y111_B6 = 1'b1;
  assign CLBLM_R_X3Y110_SLICE_X3Y110_B4 = 1'b1;
  assign RIOI3_X105Y91_OLOGIC_X1Y92_D1 = CLBLM_L_X10Y113_SLICE_X13Y113_AO6;
  assign CLBLM_R_X3Y110_SLICE_X3Y110_B5 = 1'b1;
  assign CLBLL_L_X4Y111_SLICE_X5Y111_C1 = CLBLL_L_X4Y111_SLICE_X5Y111_AO6;
  assign CLBLL_L_X4Y111_SLICE_X5Y111_C2 = CLBLM_R_X3Y111_SLICE_X3Y111_BO6;
  assign CLBLL_L_X4Y111_SLICE_X5Y111_C3 = CLBLL_L_X4Y111_SLICE_X4Y111_BO6;
  assign CLBLL_L_X4Y111_SLICE_X5Y111_C4 = CLBLL_L_X4Y112_SLICE_X4Y112_BO6;
  assign CLBLL_L_X4Y111_SLICE_X5Y111_C5 = CLBLL_L_X4Y111_SLICE_X5Y111_DO6;
  assign CLBLL_L_X4Y111_SLICE_X5Y111_C6 = LIOB33_X0Y117_IOB_X0Y118_I;
  assign CLBLM_R_X3Y110_SLICE_X3Y110_B6 = 1'b1;
  assign LIOI3_TBYTESRC_X0Y181_OLOGIC_X0Y182_D1 = LIOB33_X0Y97_IOB_X0Y97_I;
  assign RIOI3_X105Y61_OLOGIC_X1Y62_D1 = CLBLL_L_X100Y121_SLICE_X156Y121_BO6;
  assign RIOI3_X105Y91_OLOGIC_X1Y92_T1 = 1'b1;
  assign RIOI3_X105Y183_OLOGIC_X1Y183_T1 = 1'b1;
  assign LIOI3_TBYTESRC_X0Y181_OLOGIC_X0Y182_T1 = 1'b1;
  assign CLBLL_L_X4Y111_SLICE_X5Y111_D1 = LIOB33_X0Y55_IOB_X0Y55_I;
  assign CLBLL_L_X4Y111_SLICE_X5Y111_D2 = LIOB33_X0Y53_IOB_X0Y54_I;
  assign CLBLL_L_X4Y111_SLICE_X5Y111_D3 = LIOB33_X0Y95_IOB_X0Y96_I;
  assign CLBLL_L_X4Y111_SLICE_X5Y111_D4 = 1'b1;
  assign CLBLL_L_X4Y111_SLICE_X5Y111_D5 = LIOB33_X0Y119_IOB_X0Y119_I;
  assign CLBLL_L_X4Y111_SLICE_X5Y111_D6 = 1'b1;
  assign RIOI3_X105Y61_OLOGIC_X1Y62_T1 = 1'b1;
  assign RIOI3_X105Y91_OLOGIC_X1Y91_D1 = CLBLM_L_X10Y113_SLICE_X12Y113_CO6;
  assign RIOI3_X105Y61_OLOGIC_X1Y61_D1 = CLBLM_L_X8Y113_SLICE_X11Y113_BO6;
  assign LIOI3_TBYTESRC_X0Y181_OLOGIC_X0Y181_D1 = LIOB33_X0Y133_IOB_X0Y133_I;
  assign RIOI3_X105Y91_OLOGIC_X1Y91_T1 = 1'b1;
  assign CLBLM_R_X5Y115_SLICE_X7Y115_A1 = LIOB33_X0Y129_IOB_X0Y130_I;
  assign CLBLM_R_X5Y115_SLICE_X7Y115_A2 = CLBLM_R_X5Y115_SLICE_X6Y115_BO6;
  assign CLBLM_R_X5Y115_SLICE_X7Y115_A3 = CLBLM_L_X10Y123_SLICE_X12Y123_AO6;
  assign CLBLM_R_X5Y115_SLICE_X7Y115_A4 = CLBLM_R_X5Y115_SLICE_X6Y115_AO6;
  assign CLBLM_R_X5Y115_SLICE_X7Y115_A5 = CLBLM_R_X5Y111_SLICE_X6Y111_AO6;
  assign CLBLM_R_X5Y115_SLICE_X7Y115_A6 = CLBLM_R_X5Y111_SLICE_X7Y111_AO6;
  assign LIOI3_TBYTESRC_X0Y181_OLOGIC_X0Y181_T1 = 1'b1;
  assign RIOB33_X105Y83_IOB_X1Y83_O = CLBLM_R_X103Y102_SLICE_X163Y102_AO6;
  assign RIOB33_X105Y83_IOB_X1Y84_O = CLBLM_R_X103Y97_SLICE_X163Y97_BO6;
  assign CLBLM_R_X5Y115_SLICE_X7Y115_B1 = 1'b1;
  assign CLBLM_R_X5Y115_SLICE_X7Y115_B2 = 1'b1;
  assign CLBLM_R_X5Y115_SLICE_X7Y115_B3 = 1'b1;
  assign CLBLM_R_X5Y115_SLICE_X7Y115_B4 = 1'b1;
  assign CLBLM_R_X5Y115_SLICE_X7Y115_B5 = 1'b1;
  assign CLBLM_R_X5Y115_SLICE_X7Y115_B6 = 1'b1;
  assign CLBLM_R_X5Y115_SLICE_X7Y115_C1 = 1'b1;
  assign CLBLM_R_X5Y115_SLICE_X7Y115_C2 = 1'b1;
  assign CLBLM_R_X5Y115_SLICE_X7Y115_C3 = 1'b1;
  assign CLBLM_R_X5Y115_SLICE_X7Y115_C4 = 1'b1;
  assign CLBLM_R_X5Y115_SLICE_X7Y115_C5 = 1'b1;
  assign CLBLM_R_X5Y115_SLICE_X7Y115_C6 = 1'b1;
  assign CLBLM_R_X5Y115_SLICE_X7Y115_D1 = 1'b1;
  assign CLBLM_R_X5Y115_SLICE_X7Y115_D2 = 1'b1;
  assign CLBLM_R_X5Y115_SLICE_X7Y115_D3 = 1'b1;
  assign CLBLM_R_X5Y115_SLICE_X7Y115_D4 = 1'b1;
  assign CLBLM_R_X5Y115_SLICE_X7Y115_D5 = 1'b1;
  assign CLBLM_R_X5Y115_SLICE_X7Y115_D6 = 1'b1;
  assign CLBLM_R_X5Y115_SLICE_X6Y115_A1 = RIOB33_X105Y165_IOB_X1Y166_I;
  assign CLBLM_R_X5Y115_SLICE_X6Y115_A2 = LIOB33_X0Y63_IOB_X0Y63_I;
  assign CLBLM_R_X5Y115_SLICE_X6Y115_A3 = LIOB33_SING_X0Y150_IOB_X0Y150_I;
  assign CLBLM_R_X5Y115_SLICE_X6Y115_A4 = LIOB33_X0Y151_IOB_X0Y151_I;
  assign CLBLM_R_X5Y115_SLICE_X6Y115_A5 = LIOB33_X0Y117_IOB_X0Y118_I;
  assign CLBLM_R_X5Y115_SLICE_X6Y115_A6 = 1'b1;
  assign CLBLM_R_X103Y115_SLICE_X163Y115_B5 = 1'b1;
  assign RIOB33_X105Y143_IOB_X1Y143_O = CLBLM_L_X10Y123_SLICE_X12Y123_AO6;
  assign RIOB33_X105Y143_IOB_X1Y144_O = CLBLM_L_X10Y123_SLICE_X12Y123_AO6;
  assign CLBLM_R_X5Y115_SLICE_X6Y115_B1 = LIOB33_X0Y129_IOB_X0Y130_I;
  assign CLBLM_R_X5Y115_SLICE_X6Y115_B2 = LIOB33_X0Y57_IOB_X0Y58_I;
  assign CLBLM_R_X5Y115_SLICE_X6Y115_B3 = LIOB33_SING_X0Y150_IOB_X0Y150_I;
  assign CLBLM_R_X5Y115_SLICE_X6Y115_B4 = LIOB33_X0Y151_IOB_X0Y151_I;
  assign CLBLM_R_X5Y115_SLICE_X6Y115_B5 = LIOB33_X0Y121_IOB_X0Y122_I;
  assign CLBLM_R_X5Y115_SLICE_X6Y115_B6 = 1'b1;
  assign CLBLM_R_X5Y115_SLICE_X6Y115_C1 = 1'b1;
  assign CLBLM_R_X5Y115_SLICE_X6Y115_C2 = 1'b1;
  assign CLBLM_R_X5Y115_SLICE_X6Y115_C3 = 1'b1;
  assign CLBLM_R_X5Y115_SLICE_X6Y115_C4 = 1'b1;
  assign CLBLM_R_X5Y115_SLICE_X6Y115_C5 = 1'b1;
  assign CLBLM_R_X5Y115_SLICE_X6Y115_C6 = 1'b1;
  assign CLBLM_R_X5Y115_SLICE_X6Y115_D1 = 1'b1;
  assign CLBLM_R_X5Y115_SLICE_X6Y115_D2 = 1'b1;
  assign CLBLM_R_X5Y115_SLICE_X6Y115_D3 = 1'b1;
  assign CLBLM_R_X5Y115_SLICE_X6Y115_D4 = 1'b1;
  assign CLBLM_R_X5Y115_SLICE_X6Y115_D5 = 1'b1;
  assign CLBLM_R_X5Y115_SLICE_X6Y115_D6 = 1'b1;
  assign LIOB33_X0Y177_IOB_X0Y178_O = CLBLL_L_X2Y175_SLICE_X0Y175_AO6;
  assign LIOB33_SING_X0Y199_IOB_X0Y199_O = CLBLL_L_X4Y111_SLICE_X5Y111_CO6;
  assign CLBLL_L_X100Y113_SLICE_X156Y113_A1 = LIOB33_X0Y153_IOB_X0Y154_I;
  assign CLBLL_L_X100Y113_SLICE_X156Y113_A2 = CLBLM_R_X5Y111_SLICE_X7Y111_CO6;
  assign CLBLL_L_X100Y113_SLICE_X156Y113_A3 = LIOB33_X0Y165_IOB_X0Y165_I;
  assign CLBLL_L_X100Y113_SLICE_X156Y113_A4 = CLBLM_L_X8Y113_SLICE_X11Y113_BO6;
  assign CLBLL_L_X100Y113_SLICE_X156Y113_A5 = LIOB33_X0Y155_IOB_X0Y156_I;
  assign CLBLL_L_X100Y113_SLICE_X156Y113_A6 = RIOB33_X105Y117_IOB_X1Y117_I;
  assign LIOI3_X0Y171_ILOGIC_X0Y172_D = LIOB33_X0Y171_IOB_X0Y172_I;
  assign LIOI3_X0Y171_ILOGIC_X0Y171_D = LIOB33_X0Y171_IOB_X0Y171_I;
  assign CLBLL_L_X100Y113_SLICE_X156Y113_B1 = LIOB33_X0Y157_IOB_X0Y157_I;
  assign CLBLL_L_X100Y113_SLICE_X156Y113_B2 = CLBLM_R_X5Y111_SLICE_X7Y111_CO6;
  assign CLBLL_L_X100Y113_SLICE_X156Y113_B3 = LIOB33_X0Y165_IOB_X0Y165_I;
  assign CLBLL_L_X100Y113_SLICE_X156Y113_B4 = CLBLM_L_X8Y113_SLICE_X11Y113_BO6;
  assign CLBLL_L_X100Y113_SLICE_X156Y113_B5 = LIOB33_X0Y157_IOB_X0Y158_I;
  assign CLBLL_L_X100Y113_SLICE_X156Y113_B6 = RIOB33_X105Y117_IOB_X1Y117_I;
  assign LIOI3_X0Y139_ILOGIC_X0Y140_D = LIOB33_X0Y139_IOB_X0Y140_I;
  assign LIOI3_X0Y139_ILOGIC_X0Y139_D = LIOB33_X0Y139_IOB_X0Y139_I;
  assign LIOI3_X0Y109_ILOGIC_X0Y110_D = LIOB33_X0Y109_IOB_X0Y110_I;
  assign CLBLL_L_X100Y113_SLICE_X156Y113_C1 = 1'b1;
  assign CLBLL_L_X100Y113_SLICE_X156Y113_C2 = 1'b1;
  assign CLBLL_L_X100Y113_SLICE_X156Y113_C3 = 1'b1;
  assign CLBLL_L_X100Y113_SLICE_X156Y113_C4 = 1'b1;
  assign CLBLL_L_X100Y113_SLICE_X156Y113_C5 = 1'b1;
  assign CLBLL_L_X100Y113_SLICE_X156Y113_C6 = 1'b1;
  assign LIOI3_X0Y77_ILOGIC_X0Y78_D = LIOB33_X0Y77_IOB_X0Y78_I;
  assign LIOI3_X0Y109_ILOGIC_X0Y109_D = LIOB33_X0Y109_IOB_X0Y109_I;
  assign LIOI3_X0Y77_ILOGIC_X0Y77_D = LIOB33_X0Y77_IOB_X0Y77_I;
  assign RIOI3_X105Y153_ILOGIC_X1Y154_D = RIOB33_X105Y153_IOB_X1Y154_I;
  assign CLBLL_L_X100Y113_SLICE_X156Y113_D1 = 1'b1;
  assign CLBLM_R_X101Y117_SLICE_X158Y117_C6 = 1'b1;
  assign CLBLL_L_X100Y113_SLICE_X156Y113_D2 = 1'b1;
  assign CLBLL_L_X100Y113_SLICE_X156Y113_D3 = 1'b1;
  assign CLBLL_L_X100Y113_SLICE_X156Y113_D4 = 1'b1;
  assign CLBLL_L_X100Y113_SLICE_X156Y113_D5 = 1'b1;
  assign CLBLL_L_X100Y113_SLICE_X156Y113_D6 = 1'b1;
  assign RIOI3_X105Y123_ILOGIC_X1Y124_D = RIOB33_X105Y123_IOB_X1Y124_I;
  assign RIOI3_X105Y153_ILOGIC_X1Y153_D = RIOB33_X105Y153_IOB_X1Y153_I;
  assign RIOI3_X105Y123_ILOGIC_X1Y123_D = RIOB33_X105Y123_IOB_X1Y123_I;
  assign LIOI3_TBYTETERM_X0Y137_ILOGIC_X0Y138_D = LIOB33_X0Y137_IOB_X0Y138_I;
  assign LIOI3_TBYTETERM_X0Y137_ILOGIC_X0Y137_D = LIOB33_X0Y137_IOB_X0Y137_I;
  assign RIOI3_SING_X105Y149_OLOGIC_X1Y149_D1 = CLBLL_L_X4Y110_SLICE_X4Y110_CO6;
  assign CLBLL_L_X100Y113_SLICE_X157Y113_A1 = 1'b1;
  assign CLBLL_L_X100Y113_SLICE_X157Y113_A2 = 1'b1;
  assign CLBLL_L_X100Y113_SLICE_X157Y113_A3 = 1'b1;
  assign CLBLL_L_X100Y113_SLICE_X157Y113_A4 = 1'b1;
  assign CLBLL_L_X100Y113_SLICE_X157Y113_A5 = 1'b1;
  assign CLBLL_L_X100Y113_SLICE_X157Y113_A6 = 1'b1;
  assign CLBLL_L_X4Y112_SLICE_X4Y112_A1 = CLBLL_L_X4Y112_SLICE_X5Y112_AO5;
  assign CLBLL_L_X4Y112_SLICE_X4Y112_A2 = LIOB33_X0Y77_IOB_X0Y78_I;
  assign CLBLL_L_X4Y112_SLICE_X4Y112_A3 = LIOB33_X0Y79_IOB_X0Y79_I;
  assign CLBLL_L_X4Y112_SLICE_X4Y112_A4 = LIOB33_X0Y115_IOB_X0Y115_I;
  assign CLBLL_L_X100Y113_SLICE_X157Y113_B2 = 1'b1;
  assign CLBLL_L_X100Y113_SLICE_X157Y113_B3 = 1'b1;
  assign CLBLL_L_X4Y112_SLICE_X4Y112_B2 = LIOB33_X0Y113_IOB_X0Y114_I;
  assign CLBLL_L_X4Y112_SLICE_X4Y112_B3 = CLBLL_L_X4Y110_SLICE_X4Y110_AO6;
  assign CLBLL_L_X4Y112_SLICE_X4Y112_B4 = CLBLM_R_X3Y112_SLICE_X3Y112_AO6;
  assign CLBLL_L_X4Y112_SLICE_X4Y112_B5 = LIOB33_X0Y111_IOB_X0Y111_I;
  assign CLBLL_L_X4Y112_SLICE_X4Y112_B6 = CLBLL_L_X4Y110_SLICE_X4Y110_AO5;
  assign CLBLL_L_X100Y113_SLICE_X157Y113_B4 = 1'b1;
  assign CLBLL_L_X100Y113_SLICE_X157Y113_B5 = 1'b1;
  assign CLBLL_L_X100Y113_SLICE_X157Y113_B6 = 1'b1;
  assign CLBLL_L_X4Y112_SLICE_X4Y112_C1 = CLBLL_L_X4Y110_SLICE_X4Y110_AO6;
  assign CLBLL_L_X4Y112_SLICE_X4Y112_C2 = LIOB33_X0Y113_IOB_X0Y114_I;
  assign CLBLL_L_X4Y112_SLICE_X4Y112_C3 = CLBLL_L_X4Y112_SLICE_X5Y112_BO6;
  assign CLBLL_L_X4Y112_SLICE_X4Y112_C4 = CLBLL_L_X4Y112_SLICE_X4Y112_AO5;
  assign CLBLL_L_X4Y112_SLICE_X4Y112_C5 = LIOB33_X0Y111_IOB_X0Y112_I;
  assign CLBLL_L_X4Y112_SLICE_X4Y112_C6 = CLBLL_L_X4Y111_SLICE_X5Y111_BO5;
  assign CLBLL_L_X100Y113_SLICE_X157Y113_C3 = 1'b1;
  assign CLBLL_L_X100Y113_SLICE_X157Y113_C4 = 1'b1;
  assign CLBLL_L_X100Y113_SLICE_X157Y113_C5 = 1'b1;
  assign CLBLL_L_X100Y113_SLICE_X157Y113_C6 = 1'b1;
  assign RIOI3_TBYTESRC_X105Y107_ILOGIC_X1Y107_D = RIOB33_X105Y107_IOB_X1Y107_I;
  assign CLBLL_L_X100Y113_SLICE_X157Y113_D1 = 1'b1;
  assign CLBLL_L_X4Y112_SLICE_X4Y112_D1 = CLBLL_L_X4Y112_SLICE_X4Y112_AO6;
  assign CLBLL_L_X4Y112_SLICE_X4Y112_D2 = CLBLL_L_X4Y112_SLICE_X5Y112_AO5;
  assign CLBLL_L_X4Y112_SLICE_X4Y112_D3 = 1'b1;
  assign CLBLL_L_X4Y112_SLICE_X4Y112_D4 = CLBLL_L_X4Y111_SLICE_X5Y111_BO5;
  assign CLBLL_L_X4Y112_SLICE_X4Y112_D5 = 1'b1;
  assign CLBLL_L_X4Y112_SLICE_X4Y112_D6 = CLBLM_R_X3Y111_SLICE_X3Y111_AO6;
  assign CLBLL_L_X100Y113_SLICE_X157Y113_D2 = 1'b1;
  assign CLBLL_L_X100Y113_SLICE_X157Y113_D3 = 1'b1;
  assign CLBLL_L_X100Y113_SLICE_X157Y113_D4 = 1'b1;
  assign CLBLL_L_X100Y113_SLICE_X157Y113_D5 = 1'b1;
  assign CLBLL_L_X100Y113_SLICE_X157Y113_D6 = 1'b1;
  assign CLBLM_R_X103Y115_SLICE_X162Y115_A4 = 1'b1;
  assign LIOB33_SING_X0Y200_IOB_X0Y200_O = LIOB33_SING_X0Y100_IOB_X0Y100_I;
  assign CLBLL_L_X4Y112_SLICE_X5Y112_A1 = LIOB33_X0Y81_IOB_X0Y81_I;
  assign CLBLL_L_X4Y112_SLICE_X5Y112_A2 = 1'b1;
  assign CLBLL_L_X4Y112_SLICE_X5Y112_A3 = LIOB33_X0Y109_IOB_X0Y109_I;
  assign CLBLL_L_X4Y112_SLICE_X5Y112_A4 = LIOB33_X0Y79_IOB_X0Y80_I;
  assign CLBLL_L_X4Y112_SLICE_X5Y112_A5 = LIOB33_X0Y95_IOB_X0Y96_I;
  assign CLBLL_L_X4Y112_SLICE_X5Y112_A6 = 1'b1;
  assign CLBLL_L_X2Y98_SLICE_X0Y98_A1 = LIOB33_X0Y53_IOB_X0Y54_I;
  assign CLBLL_L_X2Y98_SLICE_X0Y98_A2 = 1'b1;
  assign CLBLL_L_X2Y98_SLICE_X0Y98_A3 = LIOB33_X0Y95_IOB_X0Y96_I;
  assign CLBLL_L_X2Y98_SLICE_X0Y98_A4 = LIOB33_X0Y81_IOB_X0Y82_I;
  assign CLBLL_L_X2Y98_SLICE_X0Y98_A5 = LIOB33_X0Y83_IOB_X0Y83_I;
  assign CLBLL_L_X2Y98_SLICE_X0Y98_A6 = LIOB33_X0Y55_IOB_X0Y55_I;
  assign CLBLL_L_X4Y112_SLICE_X5Y112_B1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLL_L_X4Y112_SLICE_X5Y112_B2 = LIOB33_X0Y75_IOB_X0Y75_I;
  assign CLBLL_L_X4Y112_SLICE_X5Y112_B3 = CLBLL_L_X4Y112_SLICE_X4Y112_AO6;
  assign CLBLL_L_X2Y98_SLICE_X0Y98_B1 = 1'b1;
  assign CLBLL_L_X2Y98_SLICE_X0Y98_B2 = 1'b1;
  assign CLBLL_L_X2Y98_SLICE_X0Y98_B3 = 1'b1;
  assign CLBLL_L_X2Y98_SLICE_X0Y98_B4 = 1'b1;
  assign CLBLL_L_X2Y98_SLICE_X0Y98_B5 = 1'b1;
  assign CLBLL_L_X2Y98_SLICE_X0Y98_B6 = 1'b1;
  assign CLBLL_L_X4Y112_SLICE_X5Y112_C1 = CLBLM_R_X3Y111_SLICE_X3Y111_DO6;
  assign CLBLL_L_X4Y112_SLICE_X5Y112_C2 = CLBLL_L_X4Y112_SLICE_X4Y112_AO5;
  assign CLBLL_L_X2Y98_SLICE_X0Y98_C1 = 1'b1;
  assign CLBLL_L_X2Y98_SLICE_X0Y98_C2 = 1'b1;
  assign CLBLL_L_X2Y98_SLICE_X0Y98_C3 = 1'b1;
  assign CLBLL_L_X2Y98_SLICE_X0Y98_C4 = 1'b1;
  assign CLBLL_L_X2Y98_SLICE_X0Y98_C5 = 1'b1;
  assign CLBLL_L_X2Y98_SLICE_X0Y98_C6 = 1'b1;
  assign CLBLL_L_X4Y112_SLICE_X5Y112_D1 = CLBLM_R_X3Y111_SLICE_X3Y111_BO5;
  assign CLBLL_L_X4Y112_SLICE_X5Y112_D2 = LIOB33_X0Y95_IOB_X0Y96_I;
  assign CLBLL_L_X4Y112_SLICE_X5Y112_D3 = CLBLL_L_X4Y112_SLICE_X5Y112_AO5;
  assign CLBLL_L_X4Y112_SLICE_X5Y112_D4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLL_L_X4Y112_SLICE_X5Y112_D5 = LIOB33_X0Y75_IOB_X0Y75_I;
  assign CLBLL_L_X4Y112_SLICE_X5Y112_D6 = LIOB33_X0Y113_IOB_X0Y114_I;
  assign CLBLL_L_X2Y98_SLICE_X0Y98_D1 = 1'b1;
  assign CLBLL_L_X2Y98_SLICE_X0Y98_D2 = 1'b1;
  assign CLBLL_L_X2Y98_SLICE_X0Y98_D3 = 1'b1;
  assign CLBLL_L_X2Y98_SLICE_X0Y98_D4 = 1'b1;
  assign CLBLL_L_X2Y98_SLICE_X0Y98_D5 = 1'b1;
  assign CLBLL_L_X2Y98_SLICE_X0Y98_D6 = 1'b1;
  assign CLBLM_R_X103Y115_SLICE_X162Y115_B6 = 1'b1;
  assign RIOB33_X105Y145_IOB_X1Y146_O = CLBLL_L_X100Y123_SLICE_X156Y123_AO5;
  assign RIOB33_X105Y145_IOB_X1Y145_O = CLBLL_L_X100Y123_SLICE_X156Y123_BO5;
  assign CLBLL_L_X2Y98_SLICE_X1Y98_A1 = 1'b1;
  assign CLBLL_L_X2Y98_SLICE_X1Y98_A2 = 1'b1;
  assign CLBLL_L_X2Y98_SLICE_X1Y98_A3 = 1'b1;
  assign CLBLL_L_X2Y98_SLICE_X1Y98_A4 = 1'b1;
  assign CLBLL_L_X2Y98_SLICE_X1Y98_A5 = 1'b1;
  assign CLBLL_L_X2Y98_SLICE_X1Y98_A6 = 1'b1;
  assign CLBLL_L_X2Y98_SLICE_X1Y98_B1 = 1'b1;
  assign CLBLL_L_X2Y98_SLICE_X1Y98_B2 = 1'b1;
  assign CLBLL_L_X2Y98_SLICE_X1Y98_B3 = 1'b1;
  assign CLBLL_L_X2Y98_SLICE_X1Y98_B4 = 1'b1;
  assign CLBLL_L_X2Y98_SLICE_X1Y98_B5 = 1'b1;
  assign CLBLL_L_X2Y98_SLICE_X1Y98_B6 = 1'b1;
  assign CLBLM_R_X103Y115_SLICE_X162Y115_C4 = 1'b1;
  assign CLBLM_R_X103Y115_SLICE_X162Y115_C5 = 1'b1;
  assign CLBLL_L_X2Y98_SLICE_X1Y98_C1 = 1'b1;
  assign CLBLL_L_X2Y98_SLICE_X1Y98_C2 = 1'b1;
  assign CLBLL_L_X2Y98_SLICE_X1Y98_C3 = 1'b1;
  assign CLBLL_L_X2Y98_SLICE_X1Y98_C4 = 1'b1;
  assign CLBLL_L_X2Y98_SLICE_X1Y98_C5 = 1'b1;
  assign CLBLL_L_X2Y98_SLICE_X1Y98_C6 = 1'b1;
  assign CLBLM_R_X103Y115_SLICE_X162Y115_C6 = 1'b1;
  assign CLBLL_L_X2Y98_SLICE_X1Y98_D1 = 1'b1;
  assign CLBLL_L_X2Y98_SLICE_X1Y98_D2 = 1'b1;
  assign CLBLL_L_X2Y98_SLICE_X1Y98_D3 = 1'b1;
  assign CLBLL_L_X2Y98_SLICE_X1Y98_D4 = 1'b1;
  assign CLBLL_L_X2Y98_SLICE_X1Y98_D5 = 1'b1;
  assign CLBLL_L_X2Y98_SLICE_X1Y98_D6 = 1'b1;
  assign LIOB33_X0Y179_IOB_X0Y180_O = LIOB33_X0Y133_IOB_X0Y133_I;
  assign LIOB33_X0Y179_IOB_X0Y179_O = LIOB33_X0Y133_IOB_X0Y134_I;
  assign CLBLM_R_X103Y115_SLICE_X162Y115_D1 = 1'b1;
  assign CLBLM_R_X103Y115_SLICE_X162Y115_D2 = 1'b1;
  assign CLBLM_R_X103Y115_SLICE_X162Y115_D3 = 1'b1;
  assign CLBLM_R_X103Y115_SLICE_X162Y115_D4 = 1'b1;
  assign CLBLM_R_X103Y115_SLICE_X162Y115_D5 = 1'b1;
  assign LIOI3_TBYTESRC_X0Y57_ILOGIC_X0Y58_D = LIOB33_X0Y57_IOB_X0Y58_I;
  assign CLBLM_R_X103Y115_SLICE_X162Y115_D6 = 1'b1;
  assign CLBLL_L_X4Y113_SLICE_X4Y113_A1 = 1'b1;
  assign CLBLL_L_X4Y113_SLICE_X4Y113_A2 = 1'b1;
  assign CLBLL_L_X4Y113_SLICE_X4Y113_A3 = 1'b1;
  assign CLBLL_L_X4Y113_SLICE_X4Y113_A4 = 1'b1;
  assign CLBLL_L_X4Y113_SLICE_X4Y113_A5 = 1'b1;
  assign CLBLL_L_X4Y113_SLICE_X4Y113_A6 = 1'b1;
  assign CLBLL_L_X4Y113_SLICE_X4Y113_B1 = 1'b1;
  assign CLBLL_L_X4Y113_SLICE_X4Y113_B2 = 1'b1;
  assign CLBLL_L_X4Y113_SLICE_X4Y113_B3 = 1'b1;
  assign CLBLL_L_X4Y113_SLICE_X4Y113_B4 = 1'b1;
  assign CLBLL_L_X4Y113_SLICE_X4Y113_B5 = 1'b1;
  assign CLBLL_L_X4Y113_SLICE_X4Y113_B6 = 1'b1;
  assign CLBLL_L_X4Y113_SLICE_X4Y113_C1 = 1'b1;
  assign CLBLL_L_X4Y113_SLICE_X4Y113_C2 = 1'b1;
  assign CLBLL_L_X4Y113_SLICE_X4Y113_C3 = 1'b1;
  assign CLBLL_L_X4Y113_SLICE_X4Y113_C4 = 1'b1;
  assign CLBLL_L_X4Y113_SLICE_X4Y113_C5 = 1'b1;
  assign CLBLL_L_X4Y113_SLICE_X4Y113_C6 = 1'b1;
  assign CLBLL_L_X4Y113_SLICE_X4Y113_D1 = 1'b1;
  assign CLBLL_L_X4Y113_SLICE_X4Y113_D2 = 1'b1;
  assign CLBLL_L_X4Y113_SLICE_X4Y113_D3 = 1'b1;
  assign CLBLL_L_X4Y113_SLICE_X4Y113_D4 = 1'b1;
  assign CLBLL_L_X4Y113_SLICE_X4Y113_D5 = 1'b1;
  assign CLBLL_L_X4Y113_SLICE_X4Y113_D6 = 1'b1;
  assign CLBLM_R_X25Y115_SLICE_X37Y115_A1 = 1'b1;
  assign CLBLM_R_X25Y115_SLICE_X37Y115_A2 = 1'b1;
  assign CLBLM_R_X25Y115_SLICE_X37Y115_A3 = 1'b1;
  assign CLBLM_R_X25Y115_SLICE_X37Y115_A4 = 1'b1;
  assign CLBLM_R_X25Y115_SLICE_X37Y115_A5 = 1'b1;
  assign CLBLM_R_X25Y115_SLICE_X37Y115_A6 = 1'b1;
  assign CLBLM_R_X25Y115_SLICE_X37Y115_B1 = 1'b1;
  assign CLBLM_R_X25Y115_SLICE_X37Y115_B2 = 1'b1;
  assign CLBLM_R_X25Y115_SLICE_X37Y115_B3 = 1'b1;
  assign CLBLM_R_X25Y115_SLICE_X37Y115_B4 = 1'b1;
  assign CLBLM_R_X25Y115_SLICE_X37Y115_B5 = 1'b1;
  assign CLBLM_R_X25Y115_SLICE_X37Y115_B6 = 1'b1;
  assign CLBLM_R_X25Y115_SLICE_X37Y115_C1 = 1'b1;
  assign CLBLM_R_X25Y115_SLICE_X37Y115_C2 = 1'b1;
  assign CLBLM_R_X25Y115_SLICE_X37Y115_C3 = 1'b1;
  assign CLBLM_R_X25Y115_SLICE_X37Y115_C4 = 1'b1;
  assign CLBLM_R_X25Y115_SLICE_X37Y115_C5 = 1'b1;
  assign CLBLM_R_X25Y115_SLICE_X37Y115_C6 = 1'b1;
  assign CLBLL_L_X4Y113_SLICE_X5Y113_A1 = LIOB33_X0Y119_IOB_X0Y120_I;
  assign CLBLL_L_X4Y113_SLICE_X5Y113_A2 = LIOB33_X0Y59_IOB_X0Y60_I;
  assign CLBLL_L_X4Y113_SLICE_X5Y113_A3 = LIOB33_X0Y115_IOB_X0Y116_I;
  assign CLBLL_L_X4Y113_SLICE_X5Y113_A4 = LIOB33_X0Y115_IOB_X0Y115_I;
  assign CLBLL_L_X4Y113_SLICE_X5Y113_A5 = LIOB33_X0Y77_IOB_X0Y78_I;
  assign CLBLL_L_X4Y113_SLICE_X5Y113_A6 = LIOB33_X0Y55_IOB_X0Y56_I;
  assign CLBLM_R_X25Y115_SLICE_X37Y115_D1 = 1'b1;
  assign CLBLM_R_X25Y115_SLICE_X37Y115_D2 = 1'b1;
  assign CLBLL_L_X4Y113_SLICE_X5Y113_B1 = LIOB33_X0Y111_IOB_X0Y111_I;
  assign CLBLL_L_X4Y113_SLICE_X5Y113_B2 = CLBLM_R_X3Y111_SLICE_X2Y111_AO5;
  assign CLBLL_L_X4Y113_SLICE_X5Y113_B3 = CLBLM_R_X3Y110_SLICE_X3Y110_AO5;
  assign CLBLL_L_X4Y113_SLICE_X5Y113_B4 = CLBLL_L_X4Y112_SLICE_X5Y112_AO6;
  assign CLBLL_L_X4Y113_SLICE_X5Y113_B5 = LIOB33_X0Y121_IOB_X0Y122_I;
  assign CLBLL_L_X4Y113_SLICE_X5Y113_B6 = CLBLL_L_X4Y110_SLICE_X4Y110_AO5;
  assign CLBLM_R_X25Y115_SLICE_X36Y115_A1 = LIOB33_X0Y59_IOB_X0Y60_I;
  assign CLBLM_R_X25Y115_SLICE_X36Y115_A2 = RIOB33_X105Y157_IOB_X1Y157_I;
  assign CLBLL_L_X4Y113_SLICE_X5Y113_C1 = 1'b1;
  assign CLBLL_L_X4Y113_SLICE_X5Y113_C2 = 1'b1;
  assign CLBLL_L_X4Y113_SLICE_X5Y113_C3 = 1'b1;
  assign CLBLL_L_X4Y113_SLICE_X5Y113_C4 = 1'b1;
  assign CLBLL_L_X4Y113_SLICE_X5Y113_C5 = 1'b1;
  assign CLBLL_L_X4Y113_SLICE_X5Y113_C6 = 1'b1;
  assign CLBLL_R_X57Y113_SLICE_X86Y113_A5 = CLBLM_R_X5Y113_SLICE_X6Y113_BO6;
  assign CLBLL_R_X57Y113_SLICE_X86Y113_A6 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLL_R_X57Y113_SLICE_X86Y113_A1 = LIOB33_X0Y153_IOB_X0Y154_I;
  assign CLBLL_R_X57Y113_SLICE_X86Y113_A2 = LIOB33_X0Y155_IOB_X0Y156_I;
  assign CLBLL_R_X57Y113_SLICE_X86Y113_A3 = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLL_R_X57Y113_SLICE_X86Y113_B3 = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLL_R_X57Y113_SLICE_X86Y113_B4 = CLBLM_R_X5Y113_SLICE_X6Y113_BO6;
  assign CLBLL_L_X4Y113_SLICE_X5Y113_D1 = 1'b1;
  assign CLBLL_L_X4Y113_SLICE_X5Y113_D2 = 1'b1;
  assign CLBLL_L_X4Y113_SLICE_X5Y113_D3 = 1'b1;
  assign CLBLL_L_X4Y113_SLICE_X5Y113_D4 = 1'b1;
  assign CLBLL_L_X4Y113_SLICE_X5Y113_D5 = 1'b1;
  assign CLBLL_L_X4Y113_SLICE_X5Y113_D6 = 1'b1;
  assign CLBLL_R_X57Y113_SLICE_X86Y113_B6 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLL_R_X57Y113_SLICE_X86Y113_C1 = 1'b1;
  assign CLBLL_R_X57Y113_SLICE_X86Y113_C2 = 1'b1;
  assign CLBLL_R_X57Y113_SLICE_X86Y113_C3 = 1'b1;
  assign CLBLL_R_X57Y113_SLICE_X86Y113_C4 = 1'b1;
  assign CLBLL_R_X57Y113_SLICE_X86Y113_C5 = 1'b1;
  assign CLBLL_R_X57Y113_SLICE_X86Y113_C6 = 1'b1;
  assign CLBLM_R_X25Y115_SLICE_X36Y115_C5 = 1'b1;
  assign CLBLM_R_X25Y115_SLICE_X36Y115_C6 = 1'b1;
  assign CLBLM_R_X25Y115_SLICE_X36Y115_D1 = 1'b1;
  assign CLBLL_R_X57Y113_SLICE_X86Y113_D1 = 1'b1;
  assign CLBLL_R_X57Y113_SLICE_X86Y113_D2 = 1'b1;
  assign CLBLL_R_X57Y113_SLICE_X86Y113_D3 = 1'b1;
  assign CLBLL_R_X57Y113_SLICE_X86Y113_D4 = 1'b1;
  assign CLBLL_R_X57Y113_SLICE_X86Y113_D5 = 1'b1;
  assign CLBLL_R_X57Y113_SLICE_X86Y113_D6 = 1'b1;
  assign CLBLM_R_X25Y115_SLICE_X36Y115_D2 = 1'b1;
  assign CLBLM_R_X25Y115_SLICE_X36Y115_D3 = 1'b1;
  assign CLBLM_R_X25Y115_SLICE_X36Y115_D4 = 1'b1;
  assign CLBLM_R_X25Y115_SLICE_X36Y115_D5 = 1'b1;
  assign CLBLM_R_X25Y115_SLICE_X36Y115_D6 = 1'b1;
  assign RIOI3_SING_X105Y150_ILOGIC_X1Y150_D = RIOB33_SING_X105Y150_IOB_X1Y150_I;
  assign CLBLL_R_X57Y113_SLICE_X87Y113_A1 = 1'b1;
  assign CLBLL_R_X57Y113_SLICE_X87Y113_A2 = 1'b1;
  assign CLBLL_R_X57Y113_SLICE_X87Y113_A3 = 1'b1;
  assign CLBLL_R_X57Y113_SLICE_X87Y113_A4 = 1'b1;
  assign CLBLL_R_X57Y113_SLICE_X87Y113_A5 = 1'b1;
  assign CLBLL_R_X57Y113_SLICE_X87Y113_A6 = 1'b1;
  assign CLBLL_R_X57Y113_SLICE_X87Y113_B1 = 1'b1;
  assign CLBLL_R_X57Y113_SLICE_X87Y113_B2 = 1'b1;
  assign CLBLL_R_X57Y113_SLICE_X87Y113_B3 = 1'b1;
  assign CLBLL_R_X57Y113_SLICE_X87Y113_B4 = 1'b1;
  assign CLBLL_R_X57Y113_SLICE_X87Y113_B5 = 1'b1;
  assign CLBLL_R_X57Y113_SLICE_X87Y113_B6 = 1'b1;
  assign LIOB33_X0Y181_IOB_X0Y181_O = LIOB33_X0Y133_IOB_X0Y133_I;
  assign LIOB33_X0Y181_IOB_X0Y182_O = LIOB33_X0Y97_IOB_X0Y97_I;
  assign CLBLL_R_X57Y113_SLICE_X87Y113_C1 = 1'b1;
  assign CLBLL_R_X57Y113_SLICE_X87Y113_C2 = 1'b1;
  assign CLBLL_R_X57Y113_SLICE_X87Y113_C3 = 1'b1;
  assign CLBLL_R_X57Y113_SLICE_X87Y113_C4 = 1'b1;
  assign CLBLL_R_X57Y113_SLICE_X87Y113_C5 = 1'b1;
  assign CLBLL_R_X57Y113_SLICE_X87Y113_C6 = 1'b1;
  assign RIOI3_X105Y185_OLOGIC_X1Y186_D1 = LIOB33_X0Y85_IOB_X0Y85_I;
  assign CLBLL_R_X57Y113_SLICE_X87Y113_D1 = 1'b1;
  assign CLBLL_R_X57Y113_SLICE_X87Y113_D2 = 1'b1;
  assign CLBLL_R_X57Y113_SLICE_X87Y113_D3 = 1'b1;
  assign CLBLL_R_X57Y113_SLICE_X87Y113_D4 = 1'b1;
  assign CLBLL_R_X57Y113_SLICE_X87Y113_D5 = 1'b1;
  assign CLBLL_R_X57Y113_SLICE_X87Y113_D6 = 1'b1;
  assign RIOI3_X105Y185_OLOGIC_X1Y186_T1 = 1'b1;
  assign RIOI3_X105Y95_OLOGIC_X1Y96_D1 = CLBLM_R_X25Y116_SLICE_X36Y116_BO6;
  assign RIOI3_X105Y185_OLOGIC_X1Y185_D1 = LIOB33_X0Y133_IOB_X0Y134_I;
  assign RIOI3_X105Y65_OLOGIC_X1Y66_D1 = CLBLM_R_X5Y112_SLICE_X6Y112_AO6;
  assign LIOI3_TBYTESRC_X0Y193_OLOGIC_X0Y194_D1 = 1'b0;
  assign RIOI3_X105Y95_OLOGIC_X1Y96_T1 = 1'b1;
  assign RIOI3_X105Y185_OLOGIC_X1Y185_T1 = 1'b1;
  assign CLBLM_L_X10Y114_SLICE_X12Y114_C1 = 1'b1;
  assign CLBLM_R_X103Y193_SLICE_X163Y193_A2 = 1'b1;
  assign RIOI3_X105Y65_OLOGIC_X1Y66_T1 = 1'b1;
  assign CLBLM_L_X10Y114_SLICE_X12Y114_C2 = 1'b1;
  assign LIOI3_TBYTESRC_X0Y193_OLOGIC_X0Y194_T1 = 1'b1;
  assign CLBLM_R_X103Y193_SLICE_X163Y193_A3 = 1'b1;
  assign RIOI3_X105Y95_OLOGIC_X1Y95_D1 = CLBLM_L_X10Y114_SLICE_X12Y114_BO6;
  assign CLBLM_L_X10Y114_SLICE_X12Y114_C3 = 1'b1;
  assign CLBLM_R_X103Y193_SLICE_X163Y193_A4 = LIOB33_X0Y85_IOB_X0Y85_I;
  assign CLBLM_L_X10Y114_SLICE_X12Y114_C4 = 1'b1;
  assign RIOI3_X105Y65_OLOGIC_X1Y65_D1 = CLBLM_R_X103Y107_SLICE_X163Y107_AO5;
  assign LIOI3_TBYTESRC_X0Y193_OLOGIC_X0Y193_D1 = CLBLM_R_X3Y112_SLICE_X3Y112_BO6;
  assign CLBLM_L_X10Y114_SLICE_X12Y114_C5 = 1'b1;
  assign RIOI3_X105Y95_OLOGIC_X1Y95_T1 = 1'b1;
  assign CLBLM_R_X103Y193_SLICE_X163Y193_A6 = 1'b1;
  assign CLBLM_L_X10Y114_SLICE_X12Y114_C6 = 1'b1;
  assign RIOI3_X105Y65_OLOGIC_X1Y65_T1 = 1'b1;
  assign LIOI3_TBYTESRC_X0Y193_OLOGIC_X0Y193_T1 = 1'b1;
  assign RIOI3_SING_X105Y199_OLOGIC_X1Y199_D1 = CLBLL_L_X2Y173_SLICE_X1Y173_BO5;
  assign CLBLM_R_X103Y193_SLICE_X163Y193_B1 = 1'b1;
  assign CLBLM_R_X103Y193_SLICE_X163Y193_B2 = 1'b1;
  assign CLBLM_R_X103Y193_SLICE_X163Y193_B3 = 1'b1;
  assign CLBLM_R_X103Y193_SLICE_X163Y193_B4 = 1'b1;
  assign CLBLM_R_X103Y193_SLICE_X163Y193_B5 = 1'b1;
  assign CLBLM_R_X103Y193_SLICE_X163Y193_B6 = 1'b1;
  assign RIOI3_SING_X105Y199_OLOGIC_X1Y199_T1 = 1'b1;
  assign CLBLM_R_X103Y193_SLICE_X163Y193_C1 = 1'b1;
  assign CLBLM_L_X10Y114_SLICE_X12Y114_D5 = 1'b1;
  assign CLBLM_R_X103Y193_SLICE_X163Y193_C2 = 1'b1;
  assign CLBLM_R_X103Y193_SLICE_X163Y193_C3 = 1'b1;
  assign CLBLM_R_X103Y193_SLICE_X163Y193_C4 = 1'b1;
  assign CLBLM_R_X103Y193_SLICE_X163Y193_C5 = 1'b1;
  assign CLBLM_R_X103Y193_SLICE_X163Y193_C6 = 1'b1;
  assign CLBLM_R_X25Y116_SLICE_X37Y116_A1 = 1'b1;
  assign CLBLM_R_X25Y116_SLICE_X37Y116_A2 = 1'b1;
  assign CLBLM_R_X25Y116_SLICE_X37Y116_A3 = 1'b1;
  assign CLBLM_R_X25Y116_SLICE_X37Y116_A4 = 1'b1;
  assign CLBLM_R_X25Y116_SLICE_X37Y116_A5 = 1'b1;
  assign CLBLM_R_X25Y116_SLICE_X37Y116_A6 = 1'b1;
  assign CLBLM_R_X103Y147_SLICE_X163Y147_A1 = RIOB33_X105Y103_IOB_X1Y103_I;
  assign CLBLL_L_X2Y146_SLICE_X0Y146_C2 = 1'b1;
  assign CLBLM_R_X103Y147_SLICE_X163Y147_A2 = 1'b1;
  assign CLBLM_R_X25Y116_SLICE_X37Y116_B1 = 1'b1;
  assign CLBLM_R_X25Y116_SLICE_X37Y116_B2 = 1'b1;
  assign CLBLM_R_X25Y116_SLICE_X37Y116_B3 = 1'b1;
  assign CLBLM_R_X25Y116_SLICE_X37Y116_B4 = 1'b1;
  assign CLBLM_R_X25Y116_SLICE_X37Y116_B5 = 1'b1;
  assign CLBLM_R_X25Y116_SLICE_X37Y116_B6 = 1'b1;
  assign CLBLM_R_X103Y147_SLICE_X163Y147_A3 = LIOB33_X0Y147_IOB_X0Y147_I;
  assign CLBLM_R_X103Y147_SLICE_X163Y147_A4 = 1'b1;
  assign CLBLM_R_X103Y147_SLICE_X163Y147_A6 = 1'b1;
  assign CLBLM_R_X25Y116_SLICE_X37Y116_C1 = 1'b1;
  assign CLBLM_R_X25Y116_SLICE_X37Y116_C2 = 1'b1;
  assign CLBLM_R_X25Y116_SLICE_X37Y116_C3 = 1'b1;
  assign CLBLM_R_X25Y116_SLICE_X37Y116_C4 = 1'b1;
  assign CLBLM_R_X25Y116_SLICE_X37Y116_C5 = 1'b1;
  assign CLBLM_R_X25Y116_SLICE_X37Y116_C6 = 1'b1;
  assign CLBLM_R_X103Y147_SLICE_X163Y147_B3 = 1'b1;
  assign CLBLL_L_X2Y146_SLICE_X0Y146_C6 = 1'b1;
  assign CLBLM_R_X103Y147_SLICE_X163Y147_B5 = 1'b1;
  assign CLBLM_R_X103Y147_SLICE_X163Y147_B6 = 1'b1;
  assign CLBLM_R_X103Y147_SLICE_X163Y147_C1 = 1'b1;
  assign CLBLM_R_X103Y147_SLICE_X163Y147_C2 = 1'b1;
  assign CLBLM_R_X103Y147_SLICE_X163Y147_C3 = 1'b1;
  assign CLBLM_R_X25Y116_SLICE_X37Y116_D1 = 1'b1;
  assign CLBLM_R_X25Y116_SLICE_X37Y116_D2 = 1'b1;
  assign CLBLM_R_X25Y116_SLICE_X37Y116_D3 = 1'b1;
  assign CLBLM_R_X25Y116_SLICE_X37Y116_D4 = 1'b1;
  assign CLBLM_R_X25Y116_SLICE_X37Y116_D5 = 1'b1;
  assign CLBLM_R_X25Y116_SLICE_X37Y116_D6 = 1'b1;
  assign CLBLM_R_X103Y147_SLICE_X163Y147_D1 = 1'b1;
  assign CLBLM_R_X103Y147_SLICE_X163Y147_D2 = 1'b1;
  assign CLBLM_R_X103Y147_SLICE_X163Y147_D3 = 1'b1;
  assign CLBLM_R_X103Y147_SLICE_X163Y147_D4 = 1'b1;
  assign CLBLM_R_X103Y147_SLICE_X163Y147_D5 = 1'b1;
  assign CLBLM_R_X25Y116_SLICE_X36Y116_A1 = LIOB33_SING_X0Y150_IOB_X0Y150_I;
  assign CLBLM_R_X25Y116_SLICE_X36Y116_A2 = LIOB33_X0Y151_IOB_X0Y151_I;
  assign CLBLM_R_X25Y116_SLICE_X36Y116_A3 = RIOB33_X105Y157_IOB_X1Y158_I;
  assign CLBLM_R_X25Y116_SLICE_X36Y116_A4 = LIOB33_X0Y55_IOB_X0Y56_I;
  assign CLBLM_R_X25Y116_SLICE_X36Y116_A5 = LIOB33_X0Y119_IOB_X0Y120_I;
  assign CLBLM_R_X25Y116_SLICE_X36Y116_A6 = 1'b1;
  assign CLBLM_R_X103Y147_SLICE_X162Y147_A1 = 1'b1;
  assign CLBLM_R_X103Y147_SLICE_X162Y147_A2 = 1'b1;
  assign CLBLM_R_X103Y147_SLICE_X162Y147_A3 = 1'b1;
  assign CLBLM_R_X103Y147_SLICE_X162Y147_A4 = 1'b1;
  assign CLBLM_R_X25Y116_SLICE_X36Y116_B1 = CLBLM_L_X10Y123_SLICE_X12Y123_AO6;
  assign CLBLM_R_X25Y116_SLICE_X36Y116_B2 = CLBLM_R_X5Y115_SLICE_X6Y115_AO6;
  assign CLBLM_R_X25Y116_SLICE_X36Y116_B3 = RIOB33_X105Y157_IOB_X1Y158_I;
  assign CLBLM_R_X25Y116_SLICE_X36Y116_B4 = CLBLM_R_X5Y111_SLICE_X6Y111_AO6;
  assign CLBLM_R_X25Y116_SLICE_X36Y116_B5 = CLBLM_R_X25Y116_SLICE_X36Y116_AO6;
  assign CLBLM_R_X25Y116_SLICE_X36Y116_B6 = CLBLM_R_X3Y111_SLICE_X2Y111_AO5;
  assign CLBLM_R_X103Y147_SLICE_X162Y147_A5 = 1'b1;
  assign CLBLM_R_X103Y147_SLICE_X162Y147_A6 = 1'b1;
  assign CLBLM_R_X103Y147_SLICE_X162Y147_B1 = 1'b1;
  assign CLBLM_R_X25Y116_SLICE_X36Y116_C1 = 1'b1;
  assign CLBLM_R_X25Y116_SLICE_X36Y116_C2 = 1'b1;
  assign CLBLM_R_X25Y116_SLICE_X36Y116_C3 = 1'b1;
  assign CLBLM_R_X25Y116_SLICE_X36Y116_C4 = 1'b1;
  assign CLBLM_R_X25Y116_SLICE_X36Y116_C5 = 1'b1;
  assign CLBLM_R_X25Y116_SLICE_X36Y116_C6 = 1'b1;
  assign CLBLM_R_X103Y147_SLICE_X162Y147_B4 = 1'b1;
  assign CLBLM_R_X103Y147_SLICE_X162Y147_B5 = 1'b1;
  assign CLBLM_R_X103Y147_SLICE_X162Y147_B6 = 1'b1;
  assign CLBLM_R_X103Y147_SLICE_X162Y147_C1 = 1'b1;
  assign CLBLM_R_X103Y147_SLICE_X162Y147_C2 = 1'b1;
  assign CLBLM_R_X103Y147_SLICE_X162Y147_C3 = 1'b1;
  assign CLBLM_R_X103Y147_SLICE_X162Y147_C4 = 1'b1;
  assign CLBLM_R_X103Y147_SLICE_X162Y147_C5 = 1'b1;
  assign CLBLM_R_X25Y116_SLICE_X36Y116_D1 = 1'b1;
  assign CLBLM_R_X25Y116_SLICE_X36Y116_D2 = 1'b1;
  assign CLBLM_R_X25Y116_SLICE_X36Y116_D3 = 1'b1;
  assign CLBLM_R_X25Y116_SLICE_X36Y116_D4 = 1'b1;
  assign CLBLM_R_X25Y116_SLICE_X36Y116_D5 = 1'b1;
  assign CLBLM_R_X25Y116_SLICE_X36Y116_D6 = 1'b1;
  assign CLBLM_R_X103Y147_SLICE_X162Y147_D1 = 1'b1;
  assign CLBLM_R_X103Y147_SLICE_X162Y147_D2 = 1'b1;
  assign CLBLM_R_X103Y147_SLICE_X162Y147_D3 = 1'b1;
  assign CLBLM_R_X103Y147_SLICE_X162Y147_D4 = 1'b1;
  assign CLBLM_R_X103Y147_SLICE_X162Y147_D5 = 1'b1;
  assign CLBLM_R_X103Y147_SLICE_X162Y147_D6 = 1'b1;
  assign RIOI3_TBYTESRC_X105Y119_ILOGIC_X1Y120_D = RIOB33_X105Y119_IOB_X1Y120_I;
  assign LIOB33_X0Y183_IOB_X0Y184_O = CLBLM_R_X103Y108_SLICE_X163Y108_AO5;
  assign LIOB33_X0Y183_IOB_X0Y183_O = LIOB33_X0Y101_IOB_X0Y102_I;
  assign RIOI3_TBYTESRC_X105Y119_ILOGIC_X1Y119_D = RIOB33_X105Y119_IOB_X1Y119_I;
  assign CLBLM_R_X103Y193_SLICE_X162Y193_A1 = 1'b1;
  assign CLBLM_R_X103Y193_SLICE_X162Y193_A2 = 1'b1;
  assign CLBLM_R_X103Y193_SLICE_X162Y193_A3 = 1'b1;
  assign CLBLM_R_X103Y193_SLICE_X162Y193_A4 = 1'b1;
  assign CLBLM_R_X103Y193_SLICE_X162Y193_A5 = 1'b1;
  assign LIOB33_X0Y193_IOB_X0Y194_O = 1'b0;
  assign CLBLM_R_X103Y193_SLICE_X162Y193_A6 = 1'b1;
  assign CLBLL_L_X4Y141_SLICE_X4Y141_A1 = 1'b1;
  assign CLBLL_L_X4Y141_SLICE_X4Y141_A2 = 1'b1;
  assign CLBLL_L_X4Y141_SLICE_X4Y141_A3 = LIOB33_X0Y159_IOB_X0Y160_I;
  assign CLBLL_L_X4Y141_SLICE_X4Y141_A4 = LIOB33_X0Y175_IOB_X0Y176_I;
  assign CLBLL_L_X4Y141_SLICE_X4Y141_A5 = 1'b1;
  assign CLBLL_L_X4Y141_SLICE_X4Y141_A6 = 1'b1;
  assign LIOB33_X0Y193_IOB_X0Y193_O = CLBLM_R_X3Y112_SLICE_X3Y112_BO6;
  assign RIOI3_TBYTESRC_X105Y93_OLOGIC_X1Y94_T1 = 1'b1;
  assign CLBLL_L_X4Y141_SLICE_X4Y141_B1 = 1'b1;
  assign CLBLL_L_X4Y141_SLICE_X4Y141_B2 = 1'b1;
  assign CLBLL_L_X4Y141_SLICE_X4Y141_B3 = 1'b1;
  assign CLBLL_L_X4Y141_SLICE_X4Y141_B4 = 1'b1;
  assign CLBLL_L_X4Y141_SLICE_X4Y141_B5 = 1'b1;
  assign CLBLL_L_X4Y141_SLICE_X4Y141_B6 = 1'b1;
  assign CLBLL_L_X4Y141_SLICE_X4Y141_C1 = 1'b1;
  assign CLBLL_L_X4Y141_SLICE_X4Y141_C2 = 1'b1;
  assign CLBLL_L_X4Y141_SLICE_X4Y141_C3 = 1'b1;
  assign CLBLL_L_X4Y141_SLICE_X4Y141_C4 = 1'b1;
  assign CLBLL_L_X4Y141_SLICE_X4Y141_C5 = 1'b1;
  assign CLBLL_L_X4Y141_SLICE_X4Y141_C6 = 1'b1;
  assign CLBLM_R_X103Y193_SLICE_X162Y193_B1 = 1'b1;
  assign CLBLM_R_X103Y193_SLICE_X162Y193_B2 = 1'b1;
  assign CLBLL_L_X4Y141_SLICE_X4Y141_D1 = 1'b1;
  assign CLBLL_L_X4Y141_SLICE_X4Y141_D2 = 1'b1;
  assign CLBLL_L_X4Y141_SLICE_X4Y141_D3 = 1'b1;
  assign CLBLL_L_X4Y141_SLICE_X4Y141_D4 = 1'b1;
  assign CLBLL_L_X4Y141_SLICE_X4Y141_D5 = 1'b1;
  assign CLBLL_L_X4Y141_SLICE_X4Y141_D6 = 1'b1;
  assign CLBLM_R_X103Y193_SLICE_X162Y193_B3 = 1'b1;
  assign CLBLM_R_X103Y193_SLICE_X162Y193_B4 = 1'b1;
  assign CLBLM_R_X103Y193_SLICE_X162Y193_B5 = 1'b1;
  assign CLBLM_R_X103Y193_SLICE_X162Y193_B6 = 1'b1;
  assign CLBLL_L_X4Y141_SLICE_X5Y141_A1 = 1'b1;
  assign CLBLL_L_X4Y141_SLICE_X5Y141_A2 = 1'b1;
  assign CLBLL_L_X4Y141_SLICE_X5Y141_A3 = 1'b1;
  assign CLBLL_L_X4Y141_SLICE_X5Y141_A4 = 1'b1;
  assign CLBLL_L_X4Y141_SLICE_X5Y141_A5 = 1'b1;
  assign CLBLL_L_X4Y141_SLICE_X5Y141_A6 = 1'b1;
  assign CLBLL_L_X4Y141_SLICE_X5Y141_B1 = 1'b1;
  assign CLBLL_L_X4Y141_SLICE_X5Y141_B2 = 1'b1;
  assign CLBLL_L_X4Y141_SLICE_X5Y141_B3 = 1'b1;
  assign CLBLL_L_X4Y141_SLICE_X5Y141_B4 = 1'b1;
  assign CLBLL_L_X4Y141_SLICE_X5Y141_B5 = 1'b1;
  assign CLBLL_L_X4Y141_SLICE_X5Y141_B6 = 1'b1;
  assign CLBLM_R_X103Y193_SLICE_X162Y193_C1 = 1'b1;
  assign CLBLL_L_X4Y141_SLICE_X5Y141_C1 = 1'b1;
  assign CLBLL_L_X4Y141_SLICE_X5Y141_C2 = 1'b1;
  assign CLBLL_L_X4Y141_SLICE_X5Y141_C3 = 1'b1;
  assign CLBLL_L_X4Y141_SLICE_X5Y141_C4 = 1'b1;
  assign CLBLL_L_X4Y141_SLICE_X5Y141_C5 = 1'b1;
  assign CLBLL_L_X4Y141_SLICE_X5Y141_C6 = 1'b1;
  assign CLBLM_R_X103Y193_SLICE_X162Y193_C2 = 1'b1;
  assign CLBLM_R_X103Y193_SLICE_X162Y193_C3 = 1'b1;
  assign CLBLM_R_X103Y193_SLICE_X162Y193_C4 = 1'b1;
  assign CLBLL_L_X4Y141_SLICE_X5Y141_D1 = 1'b1;
  assign CLBLL_L_X4Y141_SLICE_X5Y141_D2 = 1'b1;
  assign CLBLL_L_X4Y141_SLICE_X5Y141_D3 = 1'b1;
  assign CLBLL_L_X4Y141_SLICE_X5Y141_D4 = 1'b1;
  assign CLBLL_L_X4Y141_SLICE_X5Y141_D5 = 1'b1;
  assign CLBLL_L_X4Y141_SLICE_X5Y141_D6 = 1'b1;
  assign CLBLM_R_X103Y193_SLICE_X162Y193_C5 = 1'b1;
  assign CLBLM_R_X103Y193_SLICE_X162Y193_C6 = 1'b1;
  assign RIOB33_X105Y91_IOB_X1Y92_O = CLBLM_L_X10Y113_SLICE_X13Y113_AO6;
  assign RIOB33_X105Y91_IOB_X1Y91_O = CLBLM_L_X10Y113_SLICE_X12Y113_CO6;
  assign CLBLM_R_X103Y193_SLICE_X162Y193_D1 = 1'b1;
  assign CLBLM_R_X103Y193_SLICE_X162Y193_D2 = 1'b1;
  assign CLBLM_R_X103Y193_SLICE_X162Y193_D3 = 1'b1;
  assign CLBLM_R_X103Y193_SLICE_X162Y193_D4 = 1'b1;
  assign CLBLM_R_X103Y193_SLICE_X162Y193_D5 = 1'b1;
  assign CLBLM_R_X103Y122_SLICE_X163Y122_A1 = LIOB33_X0Y139_IOB_X0Y140_I;
  assign CLBLM_R_X103Y122_SLICE_X163Y122_A2 = 1'b1;
  assign CLBLM_R_X103Y122_SLICE_X163Y122_A3 = CLBLM_R_X103Y122_SLICE_X162Y122_AO6;
  assign CLBLM_R_X103Y122_SLICE_X163Y122_A4 = LIOB33_X0Y141_IOB_X0Y141_I;
  assign CLBLM_R_X103Y122_SLICE_X163Y122_A5 = RIOB33_X105Y103_IOB_X1Y104_I;
  assign CLBLM_R_X103Y122_SLICE_X163Y122_A6 = 1'b1;
  assign CLBLM_R_X103Y193_SLICE_X162Y193_D6 = 1'b1;
  assign CLBLM_R_X103Y122_SLICE_X163Y122_B1 = RIOB33_X105Y103_IOB_X1Y104_I;
  assign CLBLM_R_X103Y122_SLICE_X163Y122_B2 = LIOB33_X0Y141_IOB_X0Y142_I;
  assign CLBLM_R_X103Y122_SLICE_X163Y122_B3 = CLBLM_R_X103Y122_SLICE_X162Y122_AO6;
  assign CLBLM_R_X103Y122_SLICE_X163Y122_B4 = LIOB33_X0Y143_IOB_X0Y143_I;
  assign CLBLM_R_X103Y122_SLICE_X163Y122_B5 = 1'b1;
  assign CLBLM_R_X103Y122_SLICE_X163Y122_B6 = 1'b1;
  assign CLBLM_R_X103Y122_SLICE_X163Y122_C1 = CLBLM_R_X103Y115_SLICE_X163Y115_AO6;
  assign CLBLM_R_X103Y122_SLICE_X163Y122_C2 = LIOB33_X0Y141_IOB_X0Y141_I;
  assign CLBLM_R_X103Y122_SLICE_X163Y122_C3 = LIOB33_X0Y139_IOB_X0Y140_I;
  assign CLBLM_R_X103Y122_SLICE_X163Y122_C4 = CLBLM_R_X7Y121_SLICE_X8Y121_BO6;
  assign CLBLM_R_X103Y122_SLICE_X163Y122_C5 = RIOB33_X105Y103_IOB_X1Y104_I;
  assign CLBLM_R_X103Y122_SLICE_X163Y122_C6 = 1'b1;
  assign CLBLM_R_X103Y122_SLICE_X163Y122_D1 = CLBLM_R_X103Y115_SLICE_X163Y115_AO6;
  assign CLBLM_R_X103Y122_SLICE_X163Y122_D2 = CLBLM_R_X7Y121_SLICE_X8Y121_BO6;
  assign CLBLM_R_X103Y122_SLICE_X163Y122_D3 = LIOB33_X0Y141_IOB_X0Y142_I;
  assign CLBLM_R_X103Y122_SLICE_X163Y122_D4 = RIOB33_X105Y103_IOB_X1Y104_I;
  assign CLBLM_R_X103Y122_SLICE_X163Y122_D5 = LIOB33_X0Y143_IOB_X0Y143_I;
  assign CLBLM_R_X103Y122_SLICE_X163Y122_D6 = 1'b1;
  assign CLBLM_R_X103Y122_SLICE_X162Y122_A1 = RIOB33_X105Y123_IOB_X1Y123_I;
  assign CLBLM_R_X103Y122_SLICE_X162Y122_A2 = RIOB33_X105Y121_IOB_X1Y122_I;
  assign CLBLM_R_X103Y122_SLICE_X162Y122_A3 = CLBLM_L_X10Y113_SLICE_X12Y113_AO6;
  assign CLBLM_R_X103Y122_SLICE_X162Y122_A4 = 1'b1;
  assign CLBLM_R_X103Y122_SLICE_X162Y122_A5 = CLBLM_R_X5Y111_SLICE_X7Y111_BO6;
  assign CLBLM_R_X103Y122_SLICE_X162Y122_A6 = 1'b1;
  assign CLBLM_R_X103Y122_SLICE_X162Y122_B1 = 1'b1;
  assign CLBLM_R_X103Y122_SLICE_X162Y122_B2 = 1'b1;
  assign CLBLM_R_X103Y122_SLICE_X162Y122_B3 = 1'b1;
  assign CLBLM_R_X103Y122_SLICE_X162Y122_B4 = 1'b1;
  assign CLBLM_R_X103Y122_SLICE_X162Y122_B5 = 1'b1;
  assign CLBLM_R_X103Y122_SLICE_X162Y122_B6 = 1'b1;
  assign LIOB33_X0Y185_IOB_X0Y185_O = LIOB33_X0Y67_IOB_X0Y67_I;
  assign LIOB33_X0Y185_IOB_X0Y186_O = LIOB33_X0Y135_IOB_X0Y135_I;
  assign CLBLM_R_X103Y122_SLICE_X162Y122_C1 = 1'b1;
  assign CLBLM_R_X103Y122_SLICE_X162Y122_C2 = 1'b1;
  assign CLBLM_R_X103Y122_SLICE_X162Y122_C3 = 1'b1;
  assign CLBLM_R_X103Y122_SLICE_X162Y122_C4 = 1'b1;
  assign CLBLM_R_X103Y122_SLICE_X162Y122_C5 = 1'b1;
  assign CLBLM_R_X103Y122_SLICE_X162Y122_C6 = 1'b1;
  assign CLBLM_R_X103Y122_SLICE_X162Y122_D1 = 1'b1;
  assign CLBLM_R_X103Y122_SLICE_X162Y122_D2 = 1'b1;
  assign CLBLM_R_X103Y122_SLICE_X162Y122_D3 = 1'b1;
  assign CLBLM_R_X103Y122_SLICE_X162Y122_D4 = 1'b1;
  assign CLBLM_R_X103Y122_SLICE_X162Y122_D5 = 1'b1;
  assign CLBLM_R_X103Y122_SLICE_X162Y122_D6 = 1'b1;
  assign RIOI3_X105Y167_ILOGIC_X1Y167_D = RIOB33_X105Y167_IOB_X1Y167_I;
  assign CLBLM_R_X25Y115_SLICE_X37Y115_D3 = 1'b1;
  assign CLBLM_R_X25Y115_SLICE_X37Y115_D4 = 1'b1;
  assign CLBLM_R_X25Y115_SLICE_X37Y115_D5 = 1'b1;
  assign CLBLM_R_X25Y115_SLICE_X37Y115_D6 = 1'b1;
  assign RIOI3_TBYTESRC_X105Y93_OLOGIC_X1Y94_D1 = CLBLL_L_X4Y109_SLICE_X4Y109_AO5;
  assign RIOI3_X105Y189_OLOGIC_X1Y190_D1 = CLBLM_R_X103Y177_SLICE_X163Y177_AO5;
  assign RIOB33_X105Y93_IOB_X1Y94_O = CLBLL_L_X4Y109_SLICE_X4Y109_AO5;
  assign RIOB33_X105Y93_IOB_X1Y93_O = CLBLM_L_X10Y113_SLICE_X13Y113_BO6;
  assign RIOI3_X105Y189_OLOGIC_X1Y190_T1 = 1'b1;
  assign RIOI3_X105Y127_OLOGIC_X1Y128_D1 = CLBLM_R_X103Y123_SLICE_X162Y123_AO6;
  assign RIOI3_X105Y97_OLOGIC_X1Y98_D1 = CLBLM_R_X25Y115_SLICE_X36Y115_BO6;
  assign LIOI3_TBYTETERM_X0Y187_OLOGIC_X0Y188_D1 = CLBLL_L_X2Y173_SLICE_X1Y173_BO6;
  assign RIOI3_X105Y189_OLOGIC_X1Y189_D1 = CLBLL_L_X2Y173_SLICE_X1Y173_AO5;
  assign RIOI3_X105Y127_OLOGIC_X1Y128_T1 = 1'b1;
  assign RIOI3_X105Y67_OLOGIC_X1Y68_D1 = CLBLL_L_X4Y109_SLICE_X4Y109_AO6;
  assign RIOI3_X105Y97_OLOGIC_X1Y98_T1 = 1'b1;
  assign LIOI3_TBYTETERM_X0Y187_OLOGIC_X0Y188_T1 = 1'b1;
  assign RIOI3_X105Y189_OLOGIC_X1Y189_T1 = 1'b1;
  assign CLBLM_R_X25Y115_SLICE_X36Y115_A3 = LIOB33_SING_X0Y150_IOB_X0Y150_I;
  assign RIOI3_X105Y127_OLOGIC_X1Y127_D1 = CLBLL_R_X57Y113_SLICE_X86Y113_AO6;
  assign RIOI3_X105Y67_OLOGIC_X1Y68_T1 = 1'b1;
  assign CLBLM_R_X25Y115_SLICE_X36Y115_A4 = LIOB33_X0Y151_IOB_X0Y151_I;
  assign RIOI3_X105Y97_OLOGIC_X1Y97_D1 = CLBLM_R_X5Y115_SLICE_X7Y115_AO6;
  assign LIOI3_TBYTETERM_X0Y187_OLOGIC_X0Y187_D1 = CLBLL_L_X2Y173_SLICE_X1Y173_BO6;
  assign CLBLM_R_X25Y115_SLICE_X36Y115_A5 = LIOB33_X0Y115_IOB_X0Y116_I;
  assign RIOI3_X105Y127_OLOGIC_X1Y127_T1 = 1'b1;
  assign CLBLM_R_X25Y115_SLICE_X36Y115_A6 = 1'b1;
  assign RIOI3_X105Y67_OLOGIC_X1Y67_D1 = CLBLM_R_X5Y109_SLICE_X6Y109_AO6;
  assign RIOI3_X105Y97_OLOGIC_X1Y97_T1 = 1'b1;
  assign LIOI3_TBYTETERM_X0Y187_OLOGIC_X0Y187_T1 = 1'b1;
  assign CLBLM_R_X103Y123_SLICE_X163Y123_A1 = CLBLM_L_X8Y113_SLICE_X10Y113_DO6;
  assign CLBLM_R_X103Y123_SLICE_X163Y123_A2 = RIOB33_X105Y153_IOB_X1Y154_I;
  assign CLBLM_R_X103Y97_SLICE_X163Y97_A1 = 1'b1;
  assign CLBLM_R_X103Y97_SLICE_X163Y97_A2 = CLBLM_R_X5Y113_SLICE_X6Y113_BO6;
  assign CLBLM_R_X103Y97_SLICE_X163Y97_A3 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_R_X103Y97_SLICE_X163Y97_A4 = CLBLM_R_X5Y111_SLICE_X6Y111_BO6;
  assign CLBLM_R_X103Y97_SLICE_X163Y97_A5 = LIOB33_X0Y51_IOB_X0Y52_I;
  assign CLBLM_R_X103Y97_SLICE_X163Y97_A6 = CLBLM_R_X103Y122_SLICE_X163Y122_AO5;
  assign CLBLM_R_X103Y123_SLICE_X163Y123_A3 = RIOB33_X105Y113_IOB_X1Y114_I;
  assign CLBLM_R_X103Y123_SLICE_X163Y123_A4 = RIOB33_X105Y125_IOB_X1Y125_I;
  assign CLBLM_R_X103Y123_SLICE_X163Y123_A5 = RIOB33_X105Y153_IOB_X1Y153_I;
  assign CLBLM_R_X103Y97_SLICE_X163Y97_B1 = CLBLM_R_X103Y122_SLICE_X163Y122_BO5;
  assign CLBLM_R_X103Y97_SLICE_X163Y97_B2 = 1'b1;
  assign CLBLM_R_X103Y97_SLICE_X163Y97_B3 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_R_X103Y97_SLICE_X163Y97_B4 = CLBLM_R_X5Y113_SLICE_X6Y113_BO6;
  assign CLBLM_R_X103Y97_SLICE_X163Y97_B5 = CLBLM_R_X5Y111_SLICE_X6Y111_BO6;
  assign CLBLM_R_X103Y97_SLICE_X163Y97_B6 = LIOB33_X0Y51_IOB_X0Y52_I;
  assign CLBLM_R_X103Y123_SLICE_X163Y123_B1 = 1'b1;
  assign CLBLL_L_X2Y102_SLICE_X0Y102_A1 = LIOB33_X0Y63_IOB_X0Y63_I;
  assign CLBLL_L_X2Y102_SLICE_X0Y102_A2 = LIOB33_X0Y71_IOB_X0Y72_I;
  assign CLBLL_L_X2Y102_SLICE_X0Y102_A3 = LIOB33_X0Y75_IOB_X0Y75_I;
  assign CLBLL_L_X2Y102_SLICE_X0Y102_A4 = LIOB33_X0Y57_IOB_X0Y58_I;
  assign CLBLL_L_X2Y102_SLICE_X0Y102_A5 = LIOB33_X0Y53_IOB_X0Y54_I;
  assign CLBLL_L_X2Y102_SLICE_X0Y102_A6 = LIOB33_X0Y79_IOB_X0Y80_I;
  assign CLBLM_R_X25Y115_SLICE_X36Y115_B1 = CLBLM_L_X10Y123_SLICE_X12Y123_AO6;
  assign CLBLM_R_X103Y97_SLICE_X163Y97_C1 = 1'b1;
  assign CLBLM_R_X25Y115_SLICE_X36Y115_B2 = RIOB33_X105Y157_IOB_X1Y157_I;
  assign CLBLL_L_X2Y102_SLICE_X0Y102_B1 = 1'b1;
  assign CLBLL_L_X2Y102_SLICE_X0Y102_B2 = LIOB33_X0Y81_IOB_X0Y82_I;
  assign CLBLL_L_X2Y102_SLICE_X0Y102_B3 = LIOB33_X0Y77_IOB_X0Y78_I;
  assign CLBLL_L_X2Y102_SLICE_X0Y102_B4 = LIOB33_X0Y55_IOB_X0Y56_I;
  assign CLBLL_L_X2Y102_SLICE_X0Y102_B5 = CLBLL_L_X2Y102_SLICE_X0Y102_AO6;
  assign CLBLL_L_X2Y102_SLICE_X0Y102_B6 = LIOB33_X0Y59_IOB_X0Y60_I;
  assign CLBLM_R_X25Y115_SLICE_X36Y115_B3 = CLBLM_R_X5Y111_SLICE_X6Y111_AO6;
  assign CLBLM_R_X25Y115_SLICE_X36Y115_B4 = CLBLM_R_X5Y111_SLICE_X7Y111_AO5;
  assign CLBLL_L_X2Y102_SLICE_X0Y102_C1 = 1'b1;
  assign CLBLL_L_X2Y102_SLICE_X0Y102_C2 = 1'b1;
  assign CLBLL_L_X2Y102_SLICE_X0Y102_C3 = 1'b1;
  assign CLBLL_L_X2Y102_SLICE_X0Y102_C4 = 1'b1;
  assign CLBLL_L_X2Y102_SLICE_X0Y102_C5 = 1'b1;
  assign CLBLL_L_X2Y102_SLICE_X0Y102_C6 = 1'b1;
  assign CLBLM_R_X25Y115_SLICE_X36Y115_B5 = CLBLM_R_X25Y115_SLICE_X36Y115_AO6;
  assign CLBLM_R_X103Y97_SLICE_X163Y97_D3 = 1'b1;
  assign CLBLM_R_X25Y115_SLICE_X36Y115_B6 = CLBLM_R_X5Y115_SLICE_X6Y115_AO6;
  assign CLBLM_R_X103Y97_SLICE_X162Y97_A1 = 1'b1;
  assign CLBLM_R_X103Y97_SLICE_X162Y97_A2 = 1'b1;
  assign CLBLM_R_X103Y97_SLICE_X162Y97_A3 = 1'b1;
  assign CLBLM_R_X103Y97_SLICE_X162Y97_A4 = 1'b1;
  assign CLBLM_R_X103Y97_SLICE_X162Y97_A5 = 1'b1;
  assign CLBLL_L_X2Y102_SLICE_X0Y102_D1 = 1'b1;
  assign CLBLL_L_X2Y102_SLICE_X0Y102_D2 = 1'b1;
  assign CLBLL_L_X2Y102_SLICE_X0Y102_D3 = 1'b1;
  assign CLBLL_L_X2Y102_SLICE_X0Y102_D4 = 1'b1;
  assign CLBLL_L_X2Y102_SLICE_X0Y102_D5 = 1'b1;
  assign CLBLL_L_X2Y102_SLICE_X0Y102_D6 = 1'b1;
  assign CLBLM_R_X103Y97_SLICE_X162Y97_A6 = 1'b1;
  assign CLBLM_R_X103Y97_SLICE_X162Y97_B1 = 1'b1;
  assign CLBLM_R_X103Y97_SLICE_X162Y97_B2 = 1'b1;
  assign CLBLM_R_X103Y97_SLICE_X162Y97_B3 = 1'b1;
  assign CLBLM_R_X103Y97_SLICE_X162Y97_B4 = 1'b1;
  assign CLBLM_R_X103Y97_SLICE_X162Y97_B5 = 1'b1;
  assign CLBLM_R_X103Y97_SLICE_X162Y97_B6 = 1'b1;
  assign CLBLM_R_X103Y97_SLICE_X162Y97_C1 = 1'b1;
  assign CLBLM_R_X103Y97_SLICE_X162Y97_C2 = 1'b1;
  assign CLBLM_R_X103Y97_SLICE_X162Y97_C3 = 1'b1;
  assign CLBLM_R_X103Y97_SLICE_X162Y97_C4 = 1'b1;
  assign CLBLM_R_X103Y97_SLICE_X162Y97_C5 = 1'b1;
  assign CLBLM_R_X103Y97_SLICE_X162Y97_C6 = 1'b1;
  assign CLBLM_R_X25Y115_SLICE_X36Y115_C1 = 1'b1;
  assign CLBLM_R_X103Y123_SLICE_X162Y123_C2 = CLBLM_R_X103Y123_SLICE_X163Y123_AO5;
  assign CLBLM_R_X103Y123_SLICE_X162Y123_C3 = CLBLL_L_X4Y111_SLICE_X5Y111_AO5;
  assign CLBLM_R_X103Y123_SLICE_X162Y123_C4 = CLBLM_R_X103Y122_SLICE_X163Y122_AO5;
  assign CLBLM_R_X103Y123_SLICE_X162Y123_C5 = CLBLM_R_X5Y111_SLICE_X6Y111_AO6;
  assign CLBLM_R_X25Y115_SLICE_X36Y115_C2 = 1'b1;
  assign CLBLM_R_X103Y123_SLICE_X162Y123_D1 = CLBLM_R_X5Y114_SLICE_X7Y114_AO6;
  assign CLBLM_R_X103Y97_SLICE_X162Y97_D1 = 1'b1;
  assign CLBLM_R_X25Y115_SLICE_X36Y115_C3 = 1'b1;
  assign CLBLM_R_X103Y97_SLICE_X162Y97_D2 = 1'b1;
  assign CLBLL_L_X2Y102_SLICE_X1Y102_A1 = 1'b1;
  assign CLBLL_L_X2Y102_SLICE_X1Y102_A2 = 1'b1;
  assign CLBLL_L_X2Y102_SLICE_X1Y102_A3 = 1'b1;
  assign CLBLL_L_X2Y102_SLICE_X1Y102_A4 = 1'b1;
  assign CLBLL_L_X2Y102_SLICE_X1Y102_A5 = 1'b1;
  assign CLBLL_L_X2Y102_SLICE_X1Y102_A6 = 1'b1;
  assign CLBLM_R_X25Y115_SLICE_X36Y115_C4 = 1'b1;
  assign CLBLM_R_X103Y97_SLICE_X162Y97_D3 = 1'b1;
  assign CLBLM_R_X103Y97_SLICE_X162Y97_D4 = 1'b1;
  assign CLBLL_L_X2Y102_SLICE_X1Y102_B1 = 1'b1;
  assign CLBLL_L_X2Y102_SLICE_X1Y102_B2 = 1'b1;
  assign CLBLL_L_X2Y102_SLICE_X1Y102_B3 = 1'b1;
  assign CLBLL_L_X2Y102_SLICE_X1Y102_B4 = 1'b1;
  assign CLBLL_L_X2Y102_SLICE_X1Y102_B5 = 1'b1;
  assign CLBLL_L_X2Y102_SLICE_X1Y102_B6 = 1'b1;
  assign CLBLM_R_X103Y147_SLICE_X163Y147_B1 = 1'b1;
  assign CLBLM_R_X3Y110_SLICE_X3Y110_A1 = LIOB33_X0Y95_IOB_X0Y96_I;
  assign CLBLL_L_X2Y102_SLICE_X1Y102_C1 = 1'b1;
  assign CLBLL_L_X2Y102_SLICE_X1Y102_C2 = 1'b1;
  assign CLBLL_L_X2Y102_SLICE_X1Y102_C3 = 1'b1;
  assign CLBLL_L_X2Y102_SLICE_X1Y102_C4 = 1'b1;
  assign CLBLL_L_X2Y102_SLICE_X1Y102_C5 = 1'b1;
  assign CLBLL_L_X2Y102_SLICE_X1Y102_C6 = 1'b1;
  assign CLBLM_R_X3Y110_SLICE_X3Y110_A2 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X3Y110_SLICE_X3Y110_A3 = LIOB33_X0Y59_IOB_X0Y59_I;
  assign CLBLM_R_X3Y110_SLICE_X3Y110_A4 = LIOB33_X0Y57_IOB_X0Y58_I;
  assign CLBLM_R_X3Y110_SLICE_X3Y110_A5 = LIOB33_X0Y59_IOB_X0Y60_I;
  assign CLBLM_R_X3Y110_SLICE_X3Y110_A6 = 1'b1;
  assign CLBLM_R_X3Y110_SLICE_X3Y110_B1 = 1'b1;
  assign CLBLM_R_X3Y110_SLICE_X3Y110_B2 = 1'b1;
  assign CLBLL_L_X2Y102_SLICE_X1Y102_D1 = 1'b1;
  assign CLBLL_L_X2Y102_SLICE_X1Y102_D2 = 1'b1;
  assign CLBLL_L_X2Y102_SLICE_X1Y102_D3 = 1'b1;
  assign CLBLL_L_X2Y102_SLICE_X1Y102_D4 = 1'b1;
  assign CLBLL_L_X2Y102_SLICE_X1Y102_D5 = 1'b1;
  assign CLBLL_L_X2Y102_SLICE_X1Y102_D6 = 1'b1;
  assign CLBLM_R_X3Y110_SLICE_X3Y110_C1 = 1'b1;
  assign CLBLM_R_X3Y110_SLICE_X3Y110_C2 = 1'b1;
  assign CLBLM_R_X3Y110_SLICE_X3Y110_C3 = 1'b1;
  assign CLBLM_R_X3Y110_SLICE_X3Y110_C4 = 1'b1;
  assign CLBLM_R_X3Y110_SLICE_X3Y110_C5 = 1'b1;
  assign CLBLM_R_X3Y110_SLICE_X3Y110_C6 = 1'b1;
  assign LIOI3_X0Y115_ILOGIC_X0Y116_D = LIOB33_X0Y115_IOB_X0Y116_I;
  assign LIOI3_X0Y115_ILOGIC_X0Y115_D = LIOB33_X0Y115_IOB_X0Y115_I;
  assign RIOI3_X105Y101_ILOGIC_X1Y102_D = RIOB33_X105Y101_IOB_X1Y102_I;
  assign LIOI3_X0Y83_ILOGIC_X0Y84_D = LIOB33_X0Y83_IOB_X0Y84_I;
  assign CLBLM_R_X3Y110_SLICE_X3Y110_D1 = 1'b1;
  assign CLBLM_R_X3Y110_SLICE_X3Y110_D2 = 1'b1;
  assign CLBLM_R_X3Y110_SLICE_X3Y110_D3 = 1'b1;
  assign CLBLM_R_X3Y110_SLICE_X3Y110_D4 = 1'b1;
  assign CLBLM_R_X3Y110_SLICE_X3Y110_D5 = 1'b1;
  assign CLBLM_R_X3Y110_SLICE_X3Y110_D6 = 1'b1;
  assign LIOI3_X0Y83_ILOGIC_X0Y83_D = LIOB33_X0Y83_IOB_X0Y83_I;
  assign LIOI3_X0Y53_ILOGIC_X0Y54_D = LIOB33_X0Y53_IOB_X0Y54_I;
  assign RIOI3_X105Y159_ILOGIC_X1Y160_D = RIOB33_X105Y159_IOB_X1Y160_I;
  assign RIOI3_X105Y159_ILOGIC_X1Y159_D = RIOB33_X105Y159_IOB_X1Y159_I;
  assign LIOI3_X0Y53_ILOGIC_X0Y53_D = LIOB33_X0Y53_IOB_X0Y53_I;
  assign RIOI3_X105Y101_ILOGIC_X1Y101_D = RIOB33_X105Y101_IOB_X1Y101_I;
  assign CLBLM_R_X3Y110_SLICE_X2Y110_A1 = 1'b1;
  assign CLBLM_R_X3Y110_SLICE_X2Y110_A2 = 1'b1;
  assign CLBLM_R_X3Y110_SLICE_X2Y110_A3 = 1'b1;
  assign CLBLM_R_X3Y110_SLICE_X2Y110_A4 = 1'b1;
  assign CLBLM_R_X3Y110_SLICE_X2Y110_A5 = 1'b1;
  assign CLBLM_R_X3Y110_SLICE_X2Y110_A6 = 1'b1;
  assign CLBLM_R_X3Y110_SLICE_X2Y110_B1 = 1'b1;
  assign CLBLM_R_X3Y110_SLICE_X2Y110_B2 = 1'b1;
  assign CLBLM_R_X3Y110_SLICE_X2Y110_B3 = 1'b1;
  assign CLBLM_R_X3Y110_SLICE_X2Y110_B4 = 1'b1;
  assign CLBLM_R_X3Y110_SLICE_X2Y110_B5 = 1'b1;
  assign CLBLM_R_X3Y110_SLICE_X2Y110_B6 = 1'b1;
  assign CLBLM_R_X103Y147_SLICE_X163Y147_C4 = 1'b1;
  assign CLBLM_R_X103Y147_SLICE_X163Y147_C5 = 1'b1;
  assign CLBLM_R_X3Y110_SLICE_X2Y110_C1 = 1'b1;
  assign CLBLM_R_X3Y110_SLICE_X2Y110_C2 = 1'b1;
  assign CLBLM_R_X3Y110_SLICE_X2Y110_C3 = 1'b1;
  assign CLBLM_R_X3Y110_SLICE_X2Y110_C4 = 1'b1;
  assign CLBLM_R_X3Y110_SLICE_X2Y110_C5 = 1'b1;
  assign CLBLM_R_X3Y110_SLICE_X2Y110_C6 = 1'b1;
  assign CLBLM_R_X103Y147_SLICE_X163Y147_C6 = 1'b1;
  assign LIOI3_TBYTESRC_X0Y69_ILOGIC_X0Y70_D = LIOB33_X0Y69_IOB_X0Y70_I;
  assign CLBLM_R_X3Y110_SLICE_X2Y110_D1 = 1'b1;
  assign CLBLM_R_X3Y110_SLICE_X2Y110_D2 = 1'b1;
  assign CLBLM_R_X3Y110_SLICE_X2Y110_D3 = 1'b1;
  assign CLBLM_R_X3Y110_SLICE_X2Y110_D4 = 1'b1;
  assign CLBLM_R_X3Y110_SLICE_X2Y110_D5 = 1'b1;
  assign CLBLM_R_X3Y110_SLICE_X2Y110_D6 = 1'b1;
  assign LIOI3_TBYTESRC_X0Y81_ILOGIC_X0Y82_D = LIOB33_X0Y81_IOB_X0Y82_I;
  assign RIOB33_X105Y95_IOB_X1Y96_O = CLBLM_R_X25Y116_SLICE_X36Y116_BO6;
  assign RIOB33_X105Y95_IOB_X1Y95_O = CLBLM_L_X10Y114_SLICE_X12Y114_BO6;
  assign LIOI3_TBYTESRC_X0Y81_ILOGIC_X0Y81_D = LIOB33_X0Y81_IOB_X0Y81_I;
  assign CLBLM_R_X103Y147_SLICE_X163Y147_D6 = 1'b1;
  assign CLBLM_R_X101Y118_SLICE_X159Y118_A5 = 1'b1;
  assign CLBLM_R_X101Y118_SLICE_X159Y118_A6 = 1'b1;
  assign CLBLM_R_X101Y123_SLICE_X158Y123_B4 = CLBLM_R_X3Y111_SLICE_X2Y111_AO5;
  assign CLBLM_R_X101Y123_SLICE_X158Y123_B5 = CLBLM_R_X101Y123_SLICE_X158Y123_AO6;
  assign CLBLL_L_X4Y112_SLICE_X4Y112_A5 = LIOB33_X0Y95_IOB_X0Y96_I;
  assign CLBLM_R_X101Y123_SLICE_X158Y123_B6 = CLBLM_R_X25Y116_SLICE_X36Y116_AO5;
  assign CLBLL_L_X4Y112_SLICE_X4Y112_A6 = 1'b1;
  assign LIOB33_X0Y189_IOB_X0Y190_O = CLBLL_L_X2Y173_SLICE_X1Y173_BO6;
  assign LIOB33_X0Y189_IOB_X0Y189_O = CLBLL_L_X2Y173_SLICE_X1Y173_BO6;
  assign CLBLL_L_X4Y112_SLICE_X4Y112_B1 = CLBLL_L_X4Y112_SLICE_X4Y112_DO6;
  assign CLBLM_R_X101Y118_SLICE_X159Y118_C2 = 1'b1;
  assign CLBLM_R_X103Y147_SLICE_X162Y147_B2 = 1'b1;
  assign LIOI3_X0Y151_ILOGIC_X0Y151_D = LIOB33_X0Y151_IOB_X0Y151_I;
  assign CLBLM_R_X103Y147_SLICE_X162Y147_B3 = 1'b1;
  assign RIOI3_X105Y59_OLOGIC_X1Y60_T1 = 1'b1;
  assign CLBLM_R_X101Y118_SLICE_X159Y118_C6 = 1'b1;
  assign CLBLM_R_X3Y111_SLICE_X3Y111_A1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X3Y111_SLICE_X3Y111_A2 = LIOB33_X0Y95_IOB_X0Y96_I;
  assign CLBLM_R_X3Y111_SLICE_X3Y111_A3 = LIOB33_X0Y75_IOB_X0Y75_I;
  assign CLBLM_R_X3Y111_SLICE_X3Y111_A4 = 1'b1;
  assign CLBLM_R_X3Y111_SLICE_X3Y111_A5 = LIOB33_X0Y113_IOB_X0Y114_I;
  assign CLBLM_R_X3Y111_SLICE_X3Y111_A6 = 1'b1;
  assign CLBLM_R_X3Y111_SLICE_X3Y111_B1 = 1'b1;
  assign CLBLM_R_X3Y111_SLICE_X3Y111_B2 = LIOB33_X0Y95_IOB_X0Y96_I;
  assign CLBLM_R_X3Y111_SLICE_X3Y111_B3 = LIOB33_X0Y117_IOB_X0Y118_I;
  assign CLBLM_R_X3Y111_SLICE_X3Y111_B4 = LIOB33_X0Y63_IOB_X0Y63_I;
  assign CLBLM_R_X3Y111_SLICE_X3Y111_B5 = LIOB33_X0Y65_IOB_X0Y65_I;
  assign CLBLM_R_X3Y111_SLICE_X3Y111_B6 = 1'b1;
  assign CLBLM_R_X103Y147_SLICE_X162Y147_C6 = 1'b1;
  assign CLBLM_R_X3Y111_SLICE_X3Y111_C1 = LIOB33_X0Y117_IOB_X0Y118_I;
  assign CLBLM_R_X3Y111_SLICE_X3Y111_C2 = LIOB33_X0Y95_IOB_X0Y96_I;
  assign CLBLM_R_X3Y111_SLICE_X3Y111_C3 = CLBLL_L_X4Y111_SLICE_X4Y111_BO6;
  assign CLBLM_R_X3Y111_SLICE_X3Y111_C4 = LIOB33_X0Y65_IOB_X0Y65_I;
  assign CLBLM_R_X3Y111_SLICE_X3Y111_C5 = LIOB33_X0Y63_IOB_X0Y63_I;
  assign CLBLM_R_X3Y111_SLICE_X3Y111_C6 = 1'b1;
  assign CLBLM_R_X3Y111_SLICE_X3Y111_D1 = CLBLM_R_X3Y110_SLICE_X3Y110_AO6;
  assign CLBLM_R_X3Y111_SLICE_X3Y111_D2 = CLBLM_R_X3Y111_SLICE_X2Y111_AO6;
  assign CLBLM_R_X3Y111_SLICE_X3Y111_D3 = LIOB33_X0Y119_IOB_X0Y120_I;
  assign CLBLM_R_X3Y111_SLICE_X3Y111_D4 = LIOB33_X0Y115_IOB_X0Y116_I;
  assign CLBLM_R_X3Y111_SLICE_X3Y111_D5 = LIOB33_X0Y121_IOB_X0Y122_I;
  assign CLBLM_R_X3Y111_SLICE_X3Y111_D6 = CLBLM_R_X3Y110_SLICE_X3Y110_AO5;
  assign CLBLM_R_X3Y111_SLICE_X2Y111_A1 = LIOB33_X0Y55_IOB_X0Y56_I;
  assign CLBLM_R_X3Y111_SLICE_X2Y111_A2 = LIOB33_X0Y119_IOB_X0Y120_I;
  assign CLBLM_R_X3Y111_SLICE_X2Y111_A3 = LIOB33_X0Y57_IOB_X0Y57_I;
  assign CLBLM_R_X3Y111_SLICE_X2Y111_A4 = LIOB33_X0Y95_IOB_X0Y96_I;
  assign CLBLM_R_X3Y111_SLICE_X2Y111_A5 = 1'b1;
  assign CLBLM_R_X3Y111_SLICE_X2Y111_A6 = 1'b1;
  assign CLBLM_R_X3Y111_SLICE_X2Y111_B1 = 1'b1;
  assign CLBLM_R_X3Y111_SLICE_X2Y111_B2 = 1'b1;
  assign CLBLM_R_X3Y111_SLICE_X2Y111_B3 = 1'b1;
  assign CLBLM_R_X3Y111_SLICE_X2Y111_B4 = 1'b1;
  assign CLBLM_R_X3Y111_SLICE_X2Y111_B5 = 1'b1;
  assign CLBLM_R_X3Y111_SLICE_X2Y111_B6 = 1'b1;
  assign RIOI3_X105Y59_OLOGIC_X1Y59_T1 = 1'b1;
  assign CLBLM_R_X3Y111_SLICE_X2Y111_C1 = 1'b1;
  assign CLBLM_R_X3Y111_SLICE_X2Y111_C2 = 1'b1;
  assign CLBLM_R_X3Y111_SLICE_X2Y111_C3 = 1'b1;
  assign CLBLM_R_X3Y111_SLICE_X2Y111_C4 = 1'b1;
  assign CLBLM_R_X3Y111_SLICE_X2Y111_C5 = 1'b1;
  assign CLBLM_R_X3Y111_SLICE_X2Y111_C6 = 1'b1;
  assign RIOB33_X105Y97_IOB_X1Y97_O = CLBLM_R_X5Y115_SLICE_X7Y115_AO6;
  assign CLBLM_R_X3Y111_SLICE_X2Y111_D1 = 1'b1;
  assign CLBLM_R_X3Y111_SLICE_X2Y111_D2 = 1'b1;
  assign CLBLM_R_X3Y111_SLICE_X2Y111_D3 = 1'b1;
  assign CLBLM_R_X3Y111_SLICE_X2Y111_D4 = 1'b1;
  assign CLBLM_R_X3Y111_SLICE_X2Y111_D5 = 1'b1;
  assign CLBLM_R_X3Y111_SLICE_X2Y111_D6 = 1'b1;
  assign RIOB33_X105Y97_IOB_X1Y98_O = CLBLM_R_X25Y115_SLICE_X36Y115_BO6;
  assign CLBLM_R_X103Y193_SLICE_X163Y193_D1 = 1'b1;
  assign RIOI3_X105Y161_ILOGIC_X1Y161_D = RIOB33_X105Y161_IOB_X1Y161_I;
  assign CLBLM_R_X103Y193_SLICE_X163Y193_D2 = 1'b1;
  assign LIOB33_X0Y191_IOB_X0Y192_O = CLBLM_R_X5Y114_SLICE_X6Y114_AO6;
  assign LIOB33_X0Y191_IOB_X0Y191_O = CLBLM_R_X5Y113_SLICE_X7Y113_AO6;
  assign CLBLM_L_X56Y119_SLICE_X85Y119_C1 = 1'b1;
  assign CLBLM_L_X56Y119_SLICE_X85Y119_C2 = 1'b1;
  assign CLBLM_R_X103Y193_SLICE_X163Y193_D3 = 1'b1;
  assign CLBLM_R_X103Y177_SLICE_X163Y177_A1 = RIOB33_SING_X105Y150_IOB_X1Y150_I;
  assign CLBLM_R_X103Y177_SLICE_X163Y177_A2 = 1'b1;
  assign CLBLM_R_X103Y177_SLICE_X163Y177_A3 = LIOB33_X0Y107_IOB_X0Y108_I;
  assign CLBLM_R_X103Y177_SLICE_X163Y177_A4 = 1'b1;
  assign CLBLM_R_X103Y177_SLICE_X163Y177_A5 = 1'b1;
  assign CLBLM_R_X103Y177_SLICE_X163Y177_A6 = 1'b1;
  assign CLBLM_R_X103Y177_SLICE_X163Y177_B1 = 1'b1;
  assign CLBLM_L_X56Y119_SLICE_X85Y119_C5 = 1'b1;
  assign CLBLM_R_X103Y177_SLICE_X163Y177_B2 = 1'b1;
  assign CLBLM_R_X103Y177_SLICE_X163Y177_B3 = 1'b1;
  assign CLBLM_R_X103Y177_SLICE_X163Y177_B4 = 1'b1;
  assign CLBLM_R_X103Y177_SLICE_X163Y177_B6 = 1'b1;
  assign CLBLM_R_X103Y177_SLICE_X163Y177_B5 = 1'b1;
  assign RIOI3_X105Y89_OLOGIC_X1Y89_D1 = CLBLM_R_X49Y101_SLICE_X74Y101_AO5;
  assign CLBLM_R_X103Y177_SLICE_X163Y177_C1 = 1'b1;
  assign CLBLM_R_X103Y177_SLICE_X163Y177_C2 = 1'b1;
  assign CLBLM_R_X103Y177_SLICE_X163Y177_C3 = 1'b1;
  assign CLBLM_R_X103Y177_SLICE_X163Y177_C4 = 1'b1;
  assign CLBLM_R_X103Y177_SLICE_X163Y177_C5 = 1'b1;
  assign CLBLM_R_X103Y177_SLICE_X163Y177_C6 = 1'b1;
  assign CLBLM_R_X103Y193_SLICE_X163Y193_D4 = 1'b1;
  assign LIOI3_X0Y177_OLOGIC_X0Y178_D1 = CLBLL_L_X2Y175_SLICE_X0Y175_AO6;
  assign CLBLM_R_X103Y177_SLICE_X163Y177_D1 = 1'b1;
  assign CLBLM_R_X103Y177_SLICE_X163Y177_D2 = 1'b1;
  assign CLBLM_R_X103Y177_SLICE_X163Y177_D3 = 1'b1;
  assign CLBLM_R_X103Y177_SLICE_X163Y177_D4 = 1'b1;
  assign CLBLM_R_X103Y177_SLICE_X163Y177_D5 = 1'b1;
  assign CLBLM_R_X103Y177_SLICE_X163Y177_D6 = 1'b1;
  assign LIOI3_X0Y177_OLOGIC_X0Y178_T1 = 1'b1;
  assign CLBLM_R_X103Y177_SLICE_X162Y177_A1 = 1'b1;
  assign CLBLM_R_X103Y177_SLICE_X162Y177_A2 = 1'b1;
  assign CLBLM_R_X103Y177_SLICE_X162Y177_A3 = 1'b1;
  assign CLBLM_R_X103Y177_SLICE_X162Y177_A4 = 1'b1;
  assign CLBLM_R_X103Y177_SLICE_X162Y177_A5 = 1'b1;
  assign CLBLM_R_X103Y177_SLICE_X162Y177_A6 = 1'b1;
  assign CLBLM_R_X103Y193_SLICE_X163Y193_D5 = 1'b1;
  assign RIOI3_X105Y191_OLOGIC_X1Y192_D1 = CLBLM_R_X103Y177_SLICE_X163Y177_AO5;
  assign CLBLM_R_X103Y177_SLICE_X162Y177_B1 = 1'b1;
  assign CLBLM_R_X103Y177_SLICE_X162Y177_B2 = 1'b1;
  assign CLBLM_R_X103Y177_SLICE_X162Y177_B3 = 1'b1;
  assign CLBLM_R_X103Y177_SLICE_X162Y177_B4 = 1'b1;
  assign CLBLM_R_X103Y177_SLICE_X162Y177_B5 = 1'b1;
  assign CLBLM_R_X103Y177_SLICE_X162Y177_B6 = 1'b1;
  assign RIOI3_X105Y191_OLOGIC_X1Y192_T1 = 1'b1;
  assign CLBLM_R_X103Y177_SLICE_X162Y177_C1 = 1'b1;
  assign CLBLM_R_X103Y177_SLICE_X162Y177_C2 = 1'b1;
  assign CLBLM_R_X103Y177_SLICE_X162Y177_C3 = 1'b1;
  assign CLBLM_R_X103Y177_SLICE_X162Y177_C4 = 1'b1;
  assign CLBLM_R_X103Y177_SLICE_X162Y177_C5 = 1'b1;
  assign CLBLM_R_X103Y177_SLICE_X162Y177_C6 = 1'b1;
  assign CLBLL_L_X4Y112_SLICE_X5Y112_B4 = LIOB33_X0Y113_IOB_X0Y114_I;
  assign CLBLM_R_X103Y193_SLICE_X163Y193_D6 = 1'b1;
  assign RIOI3_X105Y129_OLOGIC_X1Y130_D1 = CLBLM_R_X101Y123_SLICE_X158Y123_BO6;
  assign RIOI3_X105Y191_OLOGIC_X1Y191_D1 = CLBLM_R_X103Y177_SLICE_X163Y177_AO5;
  assign CLBLL_L_X4Y112_SLICE_X5Y112_B5 = CLBLL_L_X4Y112_SLICE_X5Y112_AO6;
  assign RIOI3_X105Y129_OLOGIC_X1Y130_T1 = 1'b1;
  assign CLBLM_R_X103Y177_SLICE_X162Y177_D1 = 1'b1;
  assign CLBLL_L_X4Y112_SLICE_X5Y112_B6 = LIOB33_X0Y95_IOB_X0Y96_I;
  assign CLBLM_R_X103Y177_SLICE_X162Y177_D2 = 1'b1;
  assign CLBLM_R_X103Y177_SLICE_X162Y177_D3 = 1'b1;
  assign CLBLM_R_X103Y177_SLICE_X162Y177_D4 = 1'b1;
  assign CLBLM_R_X103Y177_SLICE_X162Y177_D5 = 1'b1;
  assign CLBLM_R_X103Y177_SLICE_X162Y177_D6 = 1'b1;
  assign RIOI3_X105Y71_OLOGIC_X1Y72_D1 = CLBLM_R_X103Y122_SLICE_X163Y122_BO6;
  assign RIOI3_X105Y191_OLOGIC_X1Y191_T1 = 1'b1;
  assign RIOI3_X105Y129_OLOGIC_X1Y129_D1 = CLBLM_R_X103Y123_SLICE_X162Y123_BO6;
  assign RIOI3_X105Y71_OLOGIC_X1Y72_T1 = 1'b1;
  assign RIOI3_X105Y129_OLOGIC_X1Y129_T1 = 1'b1;
  assign RIOI3_X105Y71_OLOGIC_X1Y71_D1 = CLBLM_R_X103Y122_SLICE_X163Y122_AO6;
  assign CLBLM_R_X3Y112_SLICE_X3Y112_A1 = 1'b1;
  assign CLBLM_R_X3Y112_SLICE_X3Y112_A2 = LIOB33_X0Y79_IOB_X0Y79_I;
  assign CLBLM_R_X3Y112_SLICE_X3Y112_A3 = LIOB33_X0Y115_IOB_X0Y115_I;
  assign CLBLM_R_X3Y112_SLICE_X3Y112_A4 = LIOB33_X0Y95_IOB_X0Y96_I;
  assign CLBLM_R_X3Y112_SLICE_X3Y112_A5 = LIOB33_X0Y77_IOB_X0Y78_I;
  assign CLBLM_R_X3Y112_SLICE_X3Y112_A6 = 1'b1;
  assign RIOI3_TBYTETERM_X105Y63_OLOGIC_X1Y64_D1 = CLBLM_R_X5Y113_SLICE_X6Y113_CO6;
  assign RIOI3_TBYTESRC_X105Y143_OLOGIC_X1Y144_D1 = CLBLM_L_X10Y123_SLICE_X12Y123_AO6;
  assign CLBLL_L_X4Y112_SLICE_X5Y112_C3 = CLBLL_L_X4Y111_SLICE_X4Y111_DO6;
  assign CLBLM_R_X3Y112_SLICE_X3Y112_B1 = LIOB33_X0Y111_IOB_X0Y111_I;
  assign CLBLM_R_X3Y112_SLICE_X3Y112_B2 = CLBLL_L_X4Y112_SLICE_X5Y112_BO6;
  assign CLBLM_R_X3Y112_SLICE_X3Y112_B3 = LIOB33_X0Y73_IOB_X0Y74_I;
  assign CLBLM_R_X3Y112_SLICE_X3Y112_B4 = LIOB33_X0Y95_IOB_X0Y96_I;
  assign CLBLL_L_X4Y112_SLICE_X5Y112_C4 = CLBLL_L_X4Y113_SLICE_X5Y113_BO6;
  assign CLBLM_R_X3Y112_SLICE_X3Y112_B5 = CLBLM_R_X3Y111_SLICE_X3Y111_CO5;
  assign CLBLM_R_X3Y112_SLICE_X3Y112_B6 = LIOB33_X0Y71_IOB_X0Y72_I;
  assign RIOI3_X105Y71_OLOGIC_X1Y71_T1 = 1'b1;
  assign CLBLL_L_X4Y112_SLICE_X5Y112_C5 = CLBLL_L_X4Y112_SLICE_X5Y112_DO6;
  assign CLBLM_R_X3Y112_SLICE_X3Y112_C1 = 1'b1;
  assign CLBLM_R_X3Y112_SLICE_X3Y112_C2 = 1'b1;
  assign CLBLM_R_X3Y112_SLICE_X3Y112_C3 = 1'b1;
  assign CLBLM_R_X3Y112_SLICE_X3Y112_C4 = 1'b1;
  assign CLBLL_L_X4Y112_SLICE_X5Y112_C6 = CLBLM_R_X5Y112_SLICE_X6Y112_CO6;
  assign CLBLM_R_X3Y112_SLICE_X3Y112_C5 = 1'b1;
  assign CLBLM_R_X3Y112_SLICE_X3Y112_C6 = 1'b1;
  assign RIOI3_TBYTESRC_X105Y143_OLOGIC_X1Y144_T1 = 1'b1;
  assign RIOI3_TBYTETERM_X105Y63_OLOGIC_X1Y63_D1 = CLBLM_R_X5Y111_SLICE_X6Y111_BO6;
  assign RIOI3_TBYTESRC_X105Y143_OLOGIC_X1Y143_D1 = CLBLM_L_X10Y123_SLICE_X12Y123_AO6;
  assign CLBLM_R_X3Y112_SLICE_X3Y112_D1 = 1'b1;
  assign CLBLM_R_X3Y112_SLICE_X3Y112_D2 = 1'b1;
  assign CLBLM_R_X3Y112_SLICE_X3Y112_D3 = 1'b1;
  assign CLBLM_R_X3Y112_SLICE_X3Y112_D4 = 1'b1;
  assign CLBLM_R_X3Y112_SLICE_X3Y112_D5 = 1'b1;
  assign CLBLM_R_X3Y112_SLICE_X3Y112_D6 = 1'b1;
  assign RIOI3_TBYTETERM_X105Y63_OLOGIC_X1Y63_T1 = 1'b1;
  assign RIOI3_TBYTESRC_X105Y143_OLOGIC_X1Y143_T1 = 1'b1;
  assign CLBLM_R_X3Y112_SLICE_X2Y112_A1 = 1'b1;
  assign CLBLM_R_X3Y112_SLICE_X2Y112_A2 = 1'b1;
  assign CLBLM_R_X3Y112_SLICE_X2Y112_A3 = 1'b1;
  assign CLBLM_R_X3Y112_SLICE_X2Y112_A4 = 1'b1;
  assign CLBLM_R_X3Y112_SLICE_X2Y112_A5 = 1'b1;
  assign CLBLM_R_X3Y112_SLICE_X2Y112_A6 = 1'b1;
  assign CLBLM_R_X3Y112_SLICE_X2Y112_B1 = 1'b1;
  assign CLBLM_R_X3Y112_SLICE_X2Y112_B2 = 1'b1;
  assign CLBLM_R_X3Y112_SLICE_X2Y112_B3 = 1'b1;
  assign CLBLM_R_X3Y112_SLICE_X2Y112_B4 = 1'b1;
  assign CLBLM_R_X3Y112_SLICE_X2Y112_B5 = 1'b1;
  assign CLBLM_R_X3Y112_SLICE_X2Y112_B6 = 1'b1;
  assign CLBLM_R_X3Y112_SLICE_X2Y112_C1 = 1'b1;
  assign CLBLM_R_X3Y112_SLICE_X2Y112_C2 = 1'b1;
  assign CLBLM_R_X3Y112_SLICE_X2Y112_C3 = 1'b1;
  assign CLBLM_R_X3Y112_SLICE_X2Y112_C4 = 1'b1;
  assign CLBLM_R_X3Y112_SLICE_X2Y112_C5 = 1'b1;
  assign CLBLM_R_X3Y112_SLICE_X2Y112_C6 = 1'b1;
  assign CLBLM_R_X3Y112_SLICE_X2Y112_D1 = 1'b1;
  assign CLBLM_R_X3Y112_SLICE_X2Y112_D2 = 1'b1;
  assign CLBLM_R_X3Y112_SLICE_X2Y112_D3 = 1'b1;
  assign CLBLM_R_X3Y112_SLICE_X2Y112_D4 = 1'b1;
  assign CLBLM_R_X3Y112_SLICE_X2Y112_D5 = 1'b1;
  assign CLBLM_R_X3Y112_SLICE_X2Y112_D6 = 1'b1;
  assign CLBLM_L_X10Y123_SLICE_X13Y123_A1 = 1'b1;
  assign CLBLM_L_X10Y123_SLICE_X13Y123_A2 = 1'b1;
  assign CLBLM_L_X10Y123_SLICE_X13Y123_A3 = 1'b1;
  assign CLBLM_L_X10Y123_SLICE_X13Y123_A4 = 1'b1;
  assign CLBLM_L_X10Y123_SLICE_X13Y123_A5 = 1'b1;
  assign CLBLM_L_X10Y123_SLICE_X13Y123_A6 = 1'b1;
  assign CLBLM_L_X10Y123_SLICE_X13Y123_B1 = 1'b1;
  assign CLBLM_L_X10Y123_SLICE_X13Y123_B2 = 1'b1;
  assign CLBLM_L_X10Y123_SLICE_X13Y123_B3 = 1'b1;
  assign CLBLM_L_X10Y123_SLICE_X13Y123_B4 = 1'b1;
  assign CLBLM_L_X10Y123_SLICE_X13Y123_B5 = 1'b1;
  assign CLBLM_L_X10Y123_SLICE_X13Y123_B6 = 1'b1;
  assign LIOI3_X0Y177_ILOGIC_X0Y177_D = LIOB33_X0Y177_IOB_X0Y177_I;
  assign CLBLM_L_X8Y113_SLICE_X11Y113_A1 = LIOB33_X0Y103_IOB_X0Y103_I;
  assign CLBLM_L_X8Y113_SLICE_X11Y113_A2 = LIOB33_X0Y95_IOB_X0Y95_I;
  assign CLBLM_L_X8Y113_SLICE_X11Y113_A3 = LIOB33_X0Y85_IOB_X0Y85_I;
  assign CLBLM_L_X8Y113_SLICE_X11Y113_A4 = LIOB33_X0Y103_IOB_X0Y104_I;
  assign CLBLM_L_X8Y113_SLICE_X11Y113_A5 = LIOB33_X0Y83_IOB_X0Y84_I;
  assign CLBLM_L_X8Y113_SLICE_X11Y113_A6 = 1'b1;
  assign CLBLM_L_X10Y123_SLICE_X13Y123_C1 = 1'b1;
  assign CLBLM_L_X10Y123_SLICE_X13Y123_C2 = 1'b1;
  assign CLBLM_L_X10Y123_SLICE_X13Y123_C3 = 1'b1;
  assign CLBLM_L_X8Y113_SLICE_X11Y113_B1 = LIOB33_SING_X0Y99_IOB_X0Y99_I;
  assign CLBLM_L_X8Y113_SLICE_X11Y113_B2 = CLBLM_R_X5Y115_SLICE_X6Y115_AO6;
  assign CLBLM_L_X8Y113_SLICE_X11Y113_B3 = LIOB33_X0Y129_IOB_X0Y129_I;
  assign CLBLM_L_X8Y113_SLICE_X11Y113_B4 = CLBLM_R_X7Y113_SLICE_X8Y113_AO5;
  assign CLBLM_L_X8Y113_SLICE_X11Y113_B5 = CLBLM_L_X10Y123_SLICE_X12Y123_AO6;
  assign CLBLM_L_X8Y113_SLICE_X11Y113_B6 = RIOB33_X105Y163_IOB_X1Y163_I;
  assign CLBLM_L_X10Y123_SLICE_X13Y123_D1 = 1'b1;
  assign CLBLM_L_X10Y123_SLICE_X13Y123_D2 = 1'b1;
  assign CLBLM_L_X8Y113_SLICE_X11Y113_C1 = CLBLM_R_X7Y113_SLICE_X8Y113_AO5;
  assign CLBLM_L_X8Y113_SLICE_X11Y113_C2 = CLBLM_R_X7Y113_SLICE_X8Y113_DO6;
  assign CLBLM_L_X8Y113_SLICE_X11Y113_C3 = CLBLM_R_X7Y113_SLICE_X8Y113_CO6;
  assign CLBLM_L_X8Y113_SLICE_X11Y113_C4 = CLBLM_L_X8Y113_SLICE_X10Y113_AO6;
  assign CLBLM_L_X8Y113_SLICE_X11Y113_C5 = CLBLM_L_X8Y113_SLICE_X11Y113_DO6;
  assign CLBLM_L_X8Y113_SLICE_X11Y113_C6 = CLBLM_R_X5Y113_SLICE_X6Y113_AO5;
  assign CLBLM_L_X10Y123_SLICE_X13Y123_D3 = 1'b1;
  assign CLBLM_L_X10Y123_SLICE_X13Y123_D4 = 1'b1;
  assign CLBLM_L_X10Y123_SLICE_X12Y123_A1 = 1'b1;
  assign CLBLM_L_X10Y123_SLICE_X12Y123_A2 = 1'b1;
  assign CLBLM_L_X10Y123_SLICE_X12Y123_A3 = LIOB33_X0Y159_IOB_X0Y160_I;
  assign CLBLM_L_X10Y123_SLICE_X12Y123_A4 = 1'b1;
  assign CLBLM_L_X10Y123_SLICE_X12Y123_A5 = LIOB33_X0Y159_IOB_X0Y159_I;
  assign CLBLM_L_X10Y123_SLICE_X12Y123_A6 = 1'b1;
  assign CLBLM_L_X8Y113_SLICE_X11Y113_D1 = CLBLM_L_X8Y113_SLICE_X11Y113_AO6;
  assign CLBLM_L_X8Y113_SLICE_X11Y113_D2 = LIOB33_X0Y125_IOB_X0Y125_I;
  assign CLBLM_L_X8Y113_SLICE_X11Y113_D3 = CLBLM_R_X7Y114_SLICE_X8Y114_BO5;
  assign CLBLM_L_X10Y123_SLICE_X12Y123_B1 = 1'b1;
  assign CLBLM_L_X10Y123_SLICE_X12Y123_B2 = 1'b1;
  assign CLBLM_L_X10Y123_SLICE_X12Y123_B3 = 1'b1;
  assign CLBLM_L_X10Y123_SLICE_X12Y123_B4 = 1'b1;
  assign CLBLM_L_X10Y123_SLICE_X12Y123_B5 = 1'b1;
  assign CLBLM_L_X10Y123_SLICE_X12Y123_B6 = 1'b1;
  assign CLBLM_L_X8Y113_SLICE_X11Y113_D4 = CLBLM_L_X8Y113_SLICE_X11Y113_AO5;
  assign CLBLM_L_X8Y113_SLICE_X11Y113_D5 = CLBLM_R_X5Y110_SLICE_X6Y110_AO6;
  assign CLBLM_L_X8Y113_SLICE_X11Y113_D6 = LIOB33_X0Y131_IOB_X0Y132_I;
  assign CLBLM_L_X8Y113_SLICE_X10Y113_A1 = 1'b1;
  assign CLBLM_L_X8Y113_SLICE_X10Y113_A2 = CLBLM_R_X5Y113_SLICE_X6Y113_AO6;
  assign CLBLM_L_X8Y113_SLICE_X10Y113_A3 = LIOB33_X0Y87_IOB_X0Y87_I;
  assign CLBLM_L_X8Y113_SLICE_X10Y113_A4 = LIOB33_X0Y95_IOB_X0Y95_I;
  assign CLBLM_L_X8Y113_SLICE_X10Y113_A5 = LIOB33_X0Y85_IOB_X0Y86_I;
  assign CLBLM_L_X8Y113_SLICE_X10Y113_A6 = 1'b1;
  assign CLBLM_L_X10Y123_SLICE_X12Y123_C1 = 1'b1;
  assign CLBLM_L_X10Y123_SLICE_X12Y123_C5 = 1'b1;
  assign CLBLM_L_X10Y123_SLICE_X12Y123_C6 = 1'b1;
  assign CLBLM_L_X8Y113_SLICE_X10Y113_B1 = LIOB33_X0Y153_IOB_X0Y153_I;
  assign CLBLM_L_X8Y113_SLICE_X10Y113_B2 = RIOB33_X105Y101_IOB_X1Y102_I;
  assign CLBLM_L_X8Y113_SLICE_X10Y113_B3 = CLBLM_R_X49Y101_SLICE_X74Y101_AO6;
  assign CLBLM_L_X8Y113_SLICE_X10Y113_B4 = LIOB33_X0Y151_IOB_X0Y152_I;
  assign CLBLM_L_X8Y113_SLICE_X10Y113_B5 = LIOB33_X0Y161_IOB_X0Y161_I;
  assign CLBLM_L_X8Y113_SLICE_X10Y113_B6 = CLBLM_L_X8Y113_SLICE_X10Y113_CO6;
  assign CLBLM_L_X10Y123_SLICE_X12Y123_D1 = 1'b1;
  assign CLBLM_L_X10Y123_SLICE_X12Y123_D2 = 1'b1;
  assign CLBLM_L_X10Y123_SLICE_X12Y123_D3 = 1'b1;
  assign CLBLM_L_X8Y113_SLICE_X10Y113_C1 = LIOB33_X0Y83_IOB_X0Y84_I;
  assign CLBLM_L_X8Y113_SLICE_X10Y113_C2 = CLBLM_L_X8Y113_SLICE_X11Y113_AO5;
  assign CLBLM_L_X8Y113_SLICE_X10Y113_C3 = LIOB33_X0Y65_IOB_X0Y66_I;
  assign CLBLM_L_X8Y113_SLICE_X10Y113_C4 = LIOB33_X0Y71_IOB_X0Y71_I;
  assign CLBLM_L_X8Y113_SLICE_X10Y113_C5 = RIOB33_X105Y167_IOB_X1Y167_I;
  assign CLBLM_L_X8Y113_SLICE_X10Y113_C6 = CLBLM_R_X5Y113_SLICE_X6Y113_AO6;
  assign CLBLM_L_X10Y123_SLICE_X12Y123_D4 = 1'b1;
  assign CLBLM_L_X10Y123_SLICE_X12Y123_D5 = 1'b1;
  assign CLBLM_L_X10Y123_SLICE_X12Y123_D6 = 1'b1;
  assign LIOI3_TBYTESRC_X0Y57_ILOGIC_X0Y57_D = LIOB33_X0Y57_IOB_X0Y57_I;
  assign CLBLM_L_X8Y113_SLICE_X10Y113_D1 = CLBLM_R_X5Y113_SLICE_X6Y113_AO6;
  assign CLBLM_L_X8Y113_SLICE_X10Y113_D2 = CLBLM_L_X8Y113_SLICE_X11Y113_AO5;
  assign CLBLM_L_X8Y113_SLICE_X10Y113_D3 = CLBLM_R_X7Y113_SLICE_X9Y113_CO6;
  assign CLBLM_L_X8Y113_SLICE_X10Y113_D4 = LIOB33_X0Y159_IOB_X0Y159_I;
  assign CLBLM_L_X8Y113_SLICE_X10Y113_D5 = RIOB33_X105Y167_IOB_X1Y167_I;
  assign CLBLM_L_X8Y113_SLICE_X10Y113_D6 = LIOB33_X0Y159_IOB_X0Y160_I;
  assign CLBLM_R_X101Y116_SLICE_X159Y116_A1 = 1'b1;
  assign CLBLM_R_X101Y116_SLICE_X159Y116_A2 = 1'b1;
  assign CLBLM_R_X101Y116_SLICE_X159Y116_A3 = 1'b1;
  assign CLBLM_R_X101Y116_SLICE_X159Y116_A4 = 1'b1;
  assign CLBLM_R_X101Y116_SLICE_X159Y116_A5 = 1'b1;
  assign CLBLM_R_X101Y116_SLICE_X159Y116_A6 = 1'b1;
  assign CLBLM_R_X101Y116_SLICE_X159Y116_B1 = 1'b1;
  assign CLBLM_R_X101Y116_SLICE_X159Y116_B2 = 1'b1;
  assign CLBLM_R_X101Y116_SLICE_X159Y116_B3 = 1'b1;
  assign CLBLM_R_X101Y116_SLICE_X159Y116_B4 = 1'b1;
  assign CLBLM_R_X101Y116_SLICE_X159Y116_B5 = 1'b1;
  assign CLBLM_R_X101Y116_SLICE_X159Y116_B6 = 1'b1;
  assign CLBLM_R_X101Y116_SLICE_X159Y116_C1 = 1'b1;
  assign CLBLM_R_X101Y116_SLICE_X159Y116_C2 = 1'b1;
  assign CLBLM_R_X101Y116_SLICE_X159Y116_C3 = 1'b1;
  assign CLBLM_R_X101Y116_SLICE_X159Y116_C4 = 1'b1;
  assign CLBLM_R_X101Y116_SLICE_X159Y116_C5 = 1'b1;
  assign CLBLM_R_X101Y116_SLICE_X159Y116_C6 = 1'b1;
  assign CLBLM_R_X101Y116_SLICE_X159Y116_D1 = 1'b1;
  assign CLBLM_R_X101Y116_SLICE_X159Y116_D2 = 1'b1;
  assign CLBLM_R_X101Y116_SLICE_X159Y116_D3 = 1'b1;
  assign CLBLM_R_X101Y116_SLICE_X159Y116_D4 = 1'b1;
  assign CLBLM_R_X101Y116_SLICE_X159Y116_D5 = 1'b1;
  assign CLBLM_R_X101Y116_SLICE_X159Y116_D6 = 1'b1;
  assign CLBLM_R_X101Y116_SLICE_X158Y116_A1 = CLBLM_R_X7Y113_SLICE_X8Y113_DO6;
  assign CLBLM_R_X101Y116_SLICE_X158Y116_A2 = CLBLM_R_X5Y110_SLICE_X6Y110_AO5;
  assign CLBLM_R_X101Y116_SLICE_X158Y116_A3 = RIOB33_X105Y115_IOB_X1Y116_I;
  assign CLBLM_R_X101Y116_SLICE_X158Y116_A4 = CLBLM_L_X10Y123_SLICE_X12Y123_AO6;
  assign CLBLM_R_X101Y116_SLICE_X158Y116_A5 = LIOB33_SING_X0Y50_IOB_X0Y50_I;
  assign CLBLM_R_X101Y116_SLICE_X158Y116_A6 = CLBLM_R_X7Y114_SLICE_X8Y114_AO5;
  assign CLBLM_R_X101Y116_SLICE_X158Y116_B1 = 1'b1;
  assign CLBLM_R_X101Y116_SLICE_X158Y116_B2 = 1'b1;
  assign CLBLM_R_X101Y116_SLICE_X158Y116_B3 = 1'b1;
  assign CLBLM_R_X101Y116_SLICE_X158Y116_B4 = 1'b1;
  assign CLBLM_R_X101Y116_SLICE_X158Y116_B5 = 1'b1;
  assign CLBLM_R_X101Y116_SLICE_X158Y116_B6 = 1'b1;
  assign CLBLM_R_X101Y116_SLICE_X158Y116_C1 = 1'b1;
  assign CLBLM_R_X101Y116_SLICE_X158Y116_C2 = 1'b1;
  assign CLBLM_R_X101Y116_SLICE_X158Y116_C3 = 1'b1;
  assign CLBLM_R_X101Y116_SLICE_X158Y116_C4 = 1'b1;
  assign CLBLM_R_X101Y116_SLICE_X158Y116_C5 = 1'b1;
  assign CLBLM_R_X101Y116_SLICE_X158Y116_C6 = 1'b1;
  assign CLBLM_R_X101Y116_SLICE_X158Y116_D1 = 1'b1;
  assign CLBLM_R_X101Y116_SLICE_X158Y116_D2 = 1'b1;
  assign CLBLM_R_X101Y116_SLICE_X158Y116_D3 = 1'b1;
  assign CLBLM_R_X101Y116_SLICE_X158Y116_D4 = 1'b1;
  assign CLBLM_R_X101Y116_SLICE_X158Y116_D5 = 1'b1;
  assign CLBLM_R_X101Y116_SLICE_X158Y116_D6 = 1'b1;
  assign RIOI3_X105Y125_ILOGIC_X1Y126_D = RIOB33_X105Y125_IOB_X1Y126_I;
  assign RIOI3_X105Y125_ILOGIC_X1Y125_D = RIOB33_X105Y125_IOB_X1Y125_I;
  assign LIOI3_X0Y55_ILOGIC_X0Y56_D = LIOB33_X0Y55_IOB_X0Y56_I;
  assign LIOI3_X0Y55_ILOGIC_X0Y55_D = LIOB33_X0Y55_IOB_X0Y55_I;
  assign CLBLL_L_X100Y121_SLICE_X156Y121_A1 = LIOB33_X0Y153_IOB_X0Y154_I;
  assign CLBLL_L_X100Y121_SLICE_X156Y121_A2 = CLBLM_R_X5Y111_SLICE_X7Y111_BO6;
  assign CLBLL_L_X100Y121_SLICE_X156Y121_A3 = CLBLM_L_X10Y113_SLICE_X12Y113_AO6;
  assign CLBLL_L_X100Y121_SLICE_X156Y121_A4 = RIOB33_X105Y155_IOB_X1Y155_I;
  assign CLBLL_L_X100Y121_SLICE_X156Y121_A5 = LIOB33_X0Y155_IOB_X0Y155_I;
  assign CLBLL_L_X100Y121_SLICE_X156Y121_A6 = LIOB33_X0Y155_IOB_X0Y156_I;
  assign CLBLL_L_X100Y121_SLICE_X156Y121_B1 = LIOB33_X0Y157_IOB_X0Y157_I;
  assign CLBLL_L_X100Y121_SLICE_X156Y121_B2 = CLBLM_R_X5Y111_SLICE_X7Y111_BO6;
  assign CLBLL_L_X100Y121_SLICE_X156Y121_B3 = LIOB33_X0Y157_IOB_X0Y158_I;
  assign CLBLL_L_X100Y121_SLICE_X156Y121_B4 = CLBLM_L_X10Y113_SLICE_X12Y113_AO6;
  assign CLBLL_L_X100Y121_SLICE_X156Y121_B5 = LIOB33_X0Y155_IOB_X0Y155_I;
  assign CLBLL_L_X100Y121_SLICE_X156Y121_B6 = RIOB33_X105Y155_IOB_X1Y155_I;
  assign LIOI3_TBYTETERM_X0Y163_ILOGIC_X0Y164_D = LIOB33_X0Y163_IOB_X0Y164_I;
  assign RIOI3_TBYTESRC_X105Y181_OLOGIC_X1Y182_T1 = 1'b1;
  assign CLBLL_L_X100Y121_SLICE_X156Y121_C1 = 1'b1;
  assign CLBLL_L_X100Y121_SLICE_X156Y121_C2 = 1'b1;
  assign CLBLL_L_X100Y121_SLICE_X156Y121_C3 = 1'b1;
  assign CLBLL_L_X100Y121_SLICE_X156Y121_C4 = 1'b1;
  assign CLBLL_L_X100Y121_SLICE_X156Y121_C5 = 1'b1;
  assign CLBLL_L_X100Y121_SLICE_X156Y121_C6 = 1'b1;
  assign CLBLL_L_X100Y121_SLICE_X156Y121_D1 = 1'b1;
  assign CLBLL_L_X100Y121_SLICE_X156Y121_D2 = 1'b1;
  assign CLBLL_L_X100Y121_SLICE_X156Y121_D3 = 1'b1;
  assign CLBLL_L_X100Y121_SLICE_X156Y121_D4 = 1'b1;
  assign CLBLL_L_X100Y121_SLICE_X156Y121_D5 = 1'b1;
  assign CLBLL_L_X100Y121_SLICE_X156Y121_D6 = 1'b1;
  assign CLBLL_L_X4Y107_SLICE_X5Y107_C6 = 1'b1;
  assign LIOB33_X0Y195_IOB_X0Y196_O = CLBLM_R_X3Y112_SLICE_X3Y112_BO6;
  assign LIOB33_X0Y195_IOB_X0Y195_O = 1'b0;
  assign CLBLL_L_X100Y121_SLICE_X157Y121_A1 = 1'b1;
  assign CLBLL_L_X100Y121_SLICE_X157Y121_A2 = 1'b1;
  assign CLBLL_L_X100Y121_SLICE_X157Y121_A3 = 1'b1;
  assign CLBLL_L_X100Y121_SLICE_X157Y121_A4 = 1'b1;
  assign CLBLL_L_X100Y121_SLICE_X157Y121_A5 = 1'b1;
  assign CLBLL_L_X100Y121_SLICE_X157Y121_A6 = 1'b1;
  assign CLBLL_L_X100Y121_SLICE_X157Y121_B1 = 1'b1;
  assign CLBLL_L_X100Y121_SLICE_X157Y121_B2 = 1'b1;
  assign CLBLL_L_X100Y121_SLICE_X157Y121_B3 = 1'b1;
  assign CLBLL_L_X100Y121_SLICE_X157Y121_B4 = 1'b1;
  assign CLBLL_L_X100Y121_SLICE_X157Y121_B5 = 1'b1;
  assign CLBLL_L_X100Y121_SLICE_X157Y121_B6 = 1'b1;
  assign CLBLL_L_X100Y121_SLICE_X157Y121_C1 = 1'b1;
  assign CLBLL_L_X100Y121_SLICE_X157Y121_C2 = 1'b1;
  assign CLBLL_L_X100Y121_SLICE_X157Y121_C3 = 1'b1;
  assign CLBLL_L_X100Y121_SLICE_X157Y121_C4 = 1'b1;
  assign CLBLL_L_X100Y121_SLICE_X157Y121_C5 = 1'b1;
  assign CLBLL_L_X100Y121_SLICE_X157Y121_C6 = 1'b1;
  assign CLBLL_L_X100Y121_SLICE_X157Y121_D1 = 1'b1;
  assign CLBLL_L_X100Y121_SLICE_X157Y121_D2 = 1'b1;
  assign CLBLL_L_X100Y121_SLICE_X157Y121_D3 = 1'b1;
  assign CLBLL_L_X100Y121_SLICE_X157Y121_D4 = 1'b1;
  assign CLBLL_L_X100Y121_SLICE_X157Y121_D5 = 1'b1;
  assign CLBLL_L_X100Y121_SLICE_X157Y121_D6 = 1'b1;
  assign CLBLL_L_X4Y107_SLICE_X5Y107_D3 = 1'b1;
  assign CLBLL_L_X4Y107_SLICE_X5Y107_D4 = 1'b1;
  assign CLBLL_L_X4Y107_SLICE_X5Y107_D5 = 1'b1;
  assign RIOI3_X105Y179_OLOGIC_X1Y180_T1 = 1'b1;
  assign RIOI3_X105Y155_ILOGIC_X1Y156_D = RIOB33_X105Y155_IOB_X1Y156_I;
  assign CLBLM_R_X101Y117_SLICE_X159Y117_A1 = 1'b1;
  assign CLBLM_R_X101Y117_SLICE_X159Y117_A2 = 1'b1;
  assign CLBLM_R_X101Y117_SLICE_X159Y117_A3 = 1'b1;
  assign CLBLM_R_X101Y117_SLICE_X159Y117_A4 = 1'b1;
  assign CLBLM_R_X101Y117_SLICE_X159Y117_A5 = 1'b1;
  assign CLBLM_R_X101Y117_SLICE_X159Y117_A6 = 1'b1;
  assign CLBLM_R_X101Y117_SLICE_X159Y117_B1 = 1'b1;
  assign CLBLM_R_X101Y117_SLICE_X159Y117_B2 = 1'b1;
  assign CLBLM_R_X101Y117_SLICE_X159Y117_B3 = 1'b1;
  assign CLBLM_R_X101Y117_SLICE_X159Y117_B4 = 1'b1;
  assign CLBLM_R_X101Y117_SLICE_X159Y117_B5 = 1'b1;
  assign CLBLM_R_X101Y117_SLICE_X159Y117_B6 = 1'b1;
  assign RIOI3_X105Y155_ILOGIC_X1Y155_D = RIOB33_X105Y155_IOB_X1Y155_I;
  assign LIOI3_X0Y85_ILOGIC_X0Y86_D = LIOB33_X0Y85_IOB_X0Y86_I;
  assign CLBLM_R_X101Y117_SLICE_X159Y117_C1 = 1'b1;
  assign CLBLM_R_X101Y117_SLICE_X159Y117_C2 = 1'b1;
  assign CLBLM_R_X101Y117_SLICE_X159Y117_C3 = 1'b1;
  assign CLBLM_R_X101Y117_SLICE_X159Y117_C4 = 1'b1;
  assign CLBLM_R_X101Y117_SLICE_X159Y117_C5 = 1'b1;
  assign CLBLM_R_X101Y117_SLICE_X159Y117_C6 = 1'b1;
  assign CLBLL_L_X4Y110_SLICE_X4Y110_C4 = CLBLL_L_X4Y109_SLICE_X4Y109_DO6;
  assign CLBLM_R_X101Y117_SLICE_X159Y117_D1 = 1'b1;
  assign CLBLM_R_X101Y117_SLICE_X159Y117_D2 = 1'b1;
  assign CLBLM_R_X101Y117_SLICE_X159Y117_D3 = 1'b1;
  assign CLBLM_R_X101Y117_SLICE_X159Y117_D4 = 1'b1;
  assign CLBLM_R_X101Y117_SLICE_X159Y117_D5 = 1'b1;
  assign CLBLM_R_X101Y117_SLICE_X159Y117_D6 = 1'b1;
  assign LIOI3_X0Y85_ILOGIC_X0Y85_D = LIOB33_X0Y85_IOB_X0Y85_I;
  assign CLBLM_R_X101Y117_SLICE_X158Y117_A1 = CLBLM_R_X7Y113_SLICE_X8Y113_DO6;
  assign CLBLM_R_X101Y117_SLICE_X158Y117_A2 = CLBLM_R_X5Y110_SLICE_X6Y110_AO5;
  assign CLBLM_R_X101Y117_SLICE_X158Y117_A3 = RIOB33_X105Y151_IOB_X1Y151_I;
  assign CLBLM_R_X101Y117_SLICE_X158Y117_A4 = CLBLM_L_X10Y123_SLICE_X12Y123_AO6;
  assign CLBLM_R_X101Y117_SLICE_X158Y117_A5 = RIOB33_X105Y151_IOB_X1Y152_I;
  assign CLBLM_R_X101Y117_SLICE_X158Y117_A6 = CLBLM_R_X7Y114_SLICE_X8Y114_AO5;
  assign CLBLM_R_X101Y117_SLICE_X158Y117_B1 = 1'b1;
  assign CLBLM_R_X101Y117_SLICE_X158Y117_B2 = 1'b1;
  assign CLBLM_R_X101Y117_SLICE_X158Y117_B3 = 1'b1;
  assign CLBLM_R_X101Y117_SLICE_X158Y117_B4 = 1'b1;
  assign CLBLM_R_X101Y117_SLICE_X158Y117_B5 = 1'b1;
  assign CLBLM_R_X101Y117_SLICE_X158Y117_B6 = 1'b1;
  assign CLBLM_L_X56Y119_SLICE_X85Y119_A1 = 1'b1;
  assign CLBLM_L_X56Y119_SLICE_X85Y119_A2 = 1'b1;
  assign CLBLM_L_X56Y119_SLICE_X85Y119_A3 = 1'b1;
  assign CLBLM_L_X56Y119_SLICE_X85Y119_A4 = 1'b1;
  assign CLBLM_R_X101Y117_SLICE_X158Y117_C1 = 1'b1;
  assign CLBLM_R_X101Y117_SLICE_X158Y117_C2 = 1'b1;
  assign CLBLM_R_X101Y117_SLICE_X158Y117_C3 = 1'b1;
  assign CLBLM_R_X101Y117_SLICE_X158Y117_C4 = 1'b1;
  assign CLBLM_R_X101Y117_SLICE_X158Y117_C5 = 1'b1;
  assign CLBLM_L_X56Y119_SLICE_X85Y119_A5 = 1'b1;
  assign CLBLM_L_X56Y119_SLICE_X85Y119_A6 = 1'b1;
  assign CLBLM_L_X56Y119_SLICE_X85Y119_B1 = 1'b1;
  assign CLBLM_L_X56Y119_SLICE_X85Y119_B2 = 1'b1;
  assign CLBLM_L_X56Y119_SLICE_X85Y119_B3 = 1'b1;
  assign CLBLM_L_X56Y119_SLICE_X85Y119_B4 = 1'b1;
  assign CLBLM_L_X56Y119_SLICE_X85Y119_B5 = 1'b1;
  assign CLBLM_L_X56Y119_SLICE_X85Y119_B6 = 1'b1;
  assign CLBLM_R_X101Y117_SLICE_X158Y117_D1 = 1'b1;
  assign CLBLM_R_X101Y117_SLICE_X158Y117_D2 = 1'b1;
  assign CLBLM_R_X101Y117_SLICE_X158Y117_D3 = 1'b1;
  assign CLBLM_R_X101Y117_SLICE_X158Y117_D4 = 1'b1;
  assign CLBLM_R_X101Y117_SLICE_X158Y117_D5 = 1'b1;
  assign CLBLM_L_X56Y119_SLICE_X85Y119_C6 = 1'b1;
  assign CLBLM_R_X101Y117_SLICE_X158Y117_D6 = 1'b1;
  assign CLBLM_L_X56Y119_SLICE_X85Y119_C3 = 1'b1;
  assign CLBLM_L_X56Y119_SLICE_X85Y119_C4 = 1'b1;
  assign CLBLM_L_X56Y119_SLICE_X85Y119_D1 = 1'b1;
  assign CLBLM_L_X56Y119_SLICE_X85Y119_D2 = 1'b1;
  assign CLBLM_L_X56Y119_SLICE_X85Y119_D3 = 1'b1;
  assign CLBLM_L_X56Y119_SLICE_X85Y119_D4 = 1'b1;
  assign CLBLM_L_X56Y119_SLICE_X85Y119_D5 = 1'b1;
  assign CLBLM_L_X56Y119_SLICE_X85Y119_D6 = 1'b1;
  assign LIOI3_TBYTETERM_X0Y163_ILOGIC_X0Y163_D = LIOB33_X0Y163_IOB_X0Y163_I;
  assign CLBLM_L_X56Y119_SLICE_X84Y119_A1 = LIOB33_X0Y175_IOB_X0Y175_I;
  assign CLBLM_L_X56Y119_SLICE_X84Y119_A2 = RIOB33_X105Y119_IOB_X1Y119_I;
  assign CLBLM_L_X56Y119_SLICE_X84Y119_A3 = LIOB33_X0Y113_IOB_X0Y113_I;
  assign CLBLM_L_X56Y119_SLICE_X84Y119_A4 = CLBLM_L_X10Y113_SLICE_X13Y113_BO6;
  assign CLBLM_L_X56Y119_SLICE_X84Y119_A5 = LIOB33_X0Y53_IOB_X0Y53_I;
  assign CLBLM_L_X56Y119_SLICE_X84Y119_A6 = 1'b1;
  assign CLBLM_L_X56Y119_SLICE_X84Y119_B1 = 1'b1;
  assign CLBLM_L_X56Y119_SLICE_X84Y119_B2 = 1'b1;
  assign CLBLM_L_X56Y119_SLICE_X84Y119_B3 = 1'b1;
  assign CLBLM_L_X56Y119_SLICE_X84Y119_B4 = 1'b1;
  assign CLBLM_L_X56Y119_SLICE_X84Y119_B5 = 1'b1;
  assign CLBLM_L_X56Y119_SLICE_X84Y119_B6 = 1'b1;
  assign LIOI3_X0Y179_OLOGIC_X0Y180_D1 = LIOB33_X0Y133_IOB_X0Y133_I;
  assign LIOI3_SING_X0Y50_ILOGIC_X0Y50_D = LIOB33_SING_X0Y50_IOB_X0Y50_I;
  assign CLBLM_L_X56Y119_SLICE_X84Y119_C1 = 1'b1;
  assign CLBLM_L_X56Y119_SLICE_X84Y119_C2 = 1'b1;
  assign CLBLM_L_X56Y119_SLICE_X84Y119_C3 = 1'b1;
  assign CLBLM_L_X56Y119_SLICE_X84Y119_C4 = 1'b1;
  assign CLBLM_L_X56Y119_SLICE_X84Y119_C5 = 1'b1;
  assign CLBLM_L_X56Y119_SLICE_X84Y119_C6 = 1'b1;
  assign LIOI3_X0Y179_OLOGIC_X0Y180_T1 = 1'b1;
  assign LIOI3_X0Y179_OLOGIC_X0Y179_D1 = LIOB33_X0Y133_IOB_X0Y134_I;
  assign CLBLM_L_X56Y119_SLICE_X84Y119_D1 = 1'b1;
  assign CLBLM_L_X56Y119_SLICE_X84Y119_D2 = 1'b1;
  assign CLBLM_L_X56Y119_SLICE_X84Y119_D3 = 1'b1;
  assign CLBLM_L_X56Y119_SLICE_X84Y119_D4 = 1'b1;
  assign CLBLM_L_X56Y119_SLICE_X84Y119_D5 = 1'b1;
  assign CLBLM_L_X56Y119_SLICE_X84Y119_D6 = 1'b1;
  assign RIOB33_X105Y59_IOB_X1Y60_O = CLBLM_L_X10Y113_SLICE_X12Y113_BO6;
  assign RIOI3_X105Y195_OLOGIC_X1Y196_D1 = CLBLL_L_X2Y173_SLICE_X0Y173_AO6;
  assign RIOI3_X105Y195_OLOGIC_X1Y196_T1 = 1'b1;
  assign LIOI3_X0Y179_OLOGIC_X0Y179_T1 = 1'b1;
  assign RIOI3_X105Y133_OLOGIC_X1Y134_D1 = CLBLM_R_X101Y118_SLICE_X158Y118_BO6;
  assign RIOI3_X105Y195_OLOGIC_X1Y195_D1 = LIOB33_X0Y85_IOB_X0Y85_I;
  assign LIOB33_X0Y197_IOB_X0Y198_O = CLBLL_L_X2Y102_SLICE_X0Y102_BO6;
  assign LIOB33_X0Y197_IOB_X0Y197_O = CLBLL_L_X4Y110_SLICE_X4Y110_CO5;
  assign RIOI3_X105Y133_OLOGIC_X1Y134_T1 = 1'b1;
  assign RIOI3_X105Y73_OLOGIC_X1Y74_D1 = CLBLL_L_X100Y113_SLICE_X156Y113_AO6;
  assign RIOI3_X105Y195_OLOGIC_X1Y195_T1 = 1'b1;
  assign RIOI3_X105Y133_OLOGIC_X1Y133_D1 = CLBLM_R_X101Y123_SLICE_X158Y123_CO6;
  assign RIOI3_X105Y73_OLOGIC_X1Y74_T1 = 1'b1;
  assign RIOI3_X105Y133_OLOGIC_X1Y133_T1 = 1'b1;
  assign RIOI3_X105Y73_OLOGIC_X1Y73_D1 = CLBLL_L_X36Y113_SLICE_X54Y113_AO6;
  assign RIOI3_TBYTETERM_X105Y87_OLOGIC_X1Y88_D1 = CLBLM_L_X8Y113_SLICE_X10Y113_BO6;
  assign RIOI3_X105Y73_OLOGIC_X1Y73_T1 = 1'b1;
  assign RIOI3_TBYTETERM_X105Y87_OLOGIC_X1Y88_T1 = 1'b1;
  assign RIOI3_TBYTETERM_X105Y87_OLOGIC_X1Y87_D1 = CLBLM_R_X103Y102_SLICE_X163Y102_BO6;
  assign LIOI3_X0Y117_ILOGIC_X0Y118_D = LIOB33_X0Y117_IOB_X0Y118_I;
  assign RIOI3_TBYTETERM_X105Y87_OLOGIC_X1Y87_T1 = 1'b1;
  assign CLBLM_R_X29Y115_SLICE_X43Y115_A1 = 1'b1;
  assign CLBLM_R_X29Y115_SLICE_X43Y115_A2 = 1'b1;
  assign CLBLM_R_X29Y115_SLICE_X43Y115_A3 = 1'b1;
  assign CLBLM_R_X29Y115_SLICE_X43Y115_A4 = 1'b1;
  assign CLBLM_R_X29Y115_SLICE_X43Y115_A5 = 1'b1;
  assign CLBLM_R_X29Y115_SLICE_X43Y115_A6 = 1'b1;
  assign LIOI3_X0Y117_ILOGIC_X0Y117_D = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLM_R_X29Y115_SLICE_X43Y115_B1 = 1'b1;
  assign CLBLM_R_X29Y115_SLICE_X43Y115_B2 = 1'b1;
  assign CLBLM_R_X29Y115_SLICE_X43Y115_B3 = 1'b1;
  assign CLBLM_R_X29Y115_SLICE_X43Y115_B4 = 1'b1;
  assign CLBLM_R_X29Y115_SLICE_X43Y115_B5 = 1'b1;
  assign CLBLM_R_X29Y115_SLICE_X43Y115_B6 = 1'b1;
  assign CLBLM_R_X29Y115_SLICE_X43Y115_C1 = 1'b1;
  assign CLBLM_R_X29Y115_SLICE_X43Y115_C2 = 1'b1;
  assign CLBLM_R_X29Y115_SLICE_X43Y115_C3 = 1'b1;
  assign CLBLM_R_X29Y115_SLICE_X43Y115_C4 = 1'b1;
  assign CLBLM_R_X29Y115_SLICE_X43Y115_C5 = 1'b1;
  assign CLBLM_R_X29Y115_SLICE_X43Y115_C6 = 1'b1;
  assign CLBLM_R_X29Y115_SLICE_X43Y115_D1 = 1'b1;
  assign CLBLM_R_X29Y115_SLICE_X43Y115_D2 = 1'b1;
  assign CLBLM_R_X29Y115_SLICE_X43Y115_D3 = 1'b1;
  assign CLBLM_R_X29Y115_SLICE_X43Y115_D4 = 1'b1;
  assign CLBLM_R_X29Y115_SLICE_X43Y115_D5 = 1'b1;
  assign CLBLM_R_X29Y115_SLICE_X43Y115_D6 = 1'b1;
  assign CLBLM_R_X103Y102_SLICE_X163Y102_A1 = CLBLM_R_X5Y113_SLICE_X6Y113_CO6;
  assign CLBLM_R_X103Y102_SLICE_X163Y102_A2 = CLBLM_L_X10Y113_SLICE_X12Y113_BO6;
  assign CLBLM_R_X103Y102_SLICE_X163Y102_A3 = CLBLM_R_X103Y122_SLICE_X163Y122_AO5;
  assign CLBLM_R_X103Y102_SLICE_X163Y102_A4 = RIOB33_X105Y109_IOB_X1Y110_I;
  assign CLBLM_R_X29Y115_SLICE_X42Y115_A1 = LIOB33_X0Y155_IOB_X0Y156_I;
  assign CLBLM_R_X29Y115_SLICE_X42Y115_A2 = LIOB33_X0Y163_IOB_X0Y164_I;
  assign CLBLM_R_X29Y115_SLICE_X42Y115_A3 = CLBLM_L_X10Y114_SLICE_X12Y114_AO6;
  assign CLBLM_R_X29Y115_SLICE_X42Y115_A4 = LIOB33_X0Y163_IOB_X0Y163_I;
  assign CLBLM_R_X29Y115_SLICE_X42Y115_A5 = LIOB33_X0Y153_IOB_X0Y154_I;
  assign CLBLM_R_X29Y115_SLICE_X42Y115_A6 = CLBLM_R_X5Y112_SLICE_X6Y112_AO6;
  assign CLBLM_R_X103Y102_SLICE_X163Y102_A5 = 1'b1;
  assign CLBLM_R_X103Y102_SLICE_X163Y102_A6 = RIOB33_X105Y109_IOB_X1Y109_I;
  assign CLBLM_R_X103Y102_SLICE_X163Y102_B1 = CLBLM_R_X5Y113_SLICE_X6Y113_CO6;
  assign CLBLM_R_X29Y115_SLICE_X42Y115_B1 = LIOB33_X0Y157_IOB_X0Y158_I;
  assign CLBLM_R_X29Y115_SLICE_X42Y115_B2 = LIOB33_X0Y163_IOB_X0Y164_I;
  assign CLBLM_R_X29Y115_SLICE_X42Y115_B3 = CLBLM_L_X10Y114_SLICE_X12Y114_AO6;
  assign CLBLM_R_X29Y115_SLICE_X42Y115_B4 = CLBLM_R_X5Y112_SLICE_X6Y112_AO6;
  assign CLBLM_R_X29Y115_SLICE_X42Y115_B5 = LIOB33_X0Y157_IOB_X0Y157_I;
  assign CLBLM_R_X29Y115_SLICE_X42Y115_B6 = LIOB33_X0Y163_IOB_X0Y163_I;
  assign CLBLM_R_X101Y118_SLICE_X159Y118_A1 = 1'b1;
  assign CLBLM_R_X101Y118_SLICE_X159Y118_A2 = 1'b1;
  assign CLBLM_R_X101Y118_SLICE_X159Y118_A3 = 1'b1;
  assign CLBLM_R_X101Y118_SLICE_X159Y118_A4 = 1'b1;
  assign CLBLM_R_X29Y115_SLICE_X42Y115_C1 = 1'b1;
  assign CLBLM_R_X29Y115_SLICE_X42Y115_C2 = 1'b1;
  assign CLBLM_R_X29Y115_SLICE_X42Y115_C3 = 1'b1;
  assign CLBLM_R_X29Y115_SLICE_X42Y115_C4 = 1'b1;
  assign CLBLM_R_X29Y115_SLICE_X42Y115_C5 = 1'b1;
  assign CLBLM_R_X29Y115_SLICE_X42Y115_C6 = 1'b1;
  assign CLBLM_R_X101Y118_SLICE_X159Y118_B1 = 1'b1;
  assign CLBLM_R_X101Y118_SLICE_X159Y118_B2 = 1'b1;
  assign CLBLM_R_X101Y118_SLICE_X159Y118_B3 = 1'b1;
  assign CLBLM_R_X101Y118_SLICE_X159Y118_B4 = 1'b1;
  assign CLBLM_R_X101Y118_SLICE_X159Y118_B5 = 1'b1;
  assign CLBLM_R_X101Y118_SLICE_X159Y118_B6 = 1'b1;
  assign CLBLM_R_X101Y118_SLICE_X159Y118_C1 = 1'b1;
  assign CLBLM_R_X29Y115_SLICE_X42Y115_D1 = 1'b1;
  assign CLBLM_R_X29Y115_SLICE_X42Y115_D2 = 1'b1;
  assign CLBLM_R_X29Y115_SLICE_X42Y115_D3 = 1'b1;
  assign CLBLM_R_X29Y115_SLICE_X42Y115_D4 = 1'b1;
  assign CLBLM_R_X29Y115_SLICE_X42Y115_D5 = 1'b1;
  assign CLBLM_R_X29Y115_SLICE_X42Y115_D6 = 1'b1;
  assign CLBLM_R_X101Y118_SLICE_X159Y118_C3 = 1'b1;
  assign CLBLM_R_X101Y118_SLICE_X159Y118_C4 = 1'b1;
  assign CLBLM_R_X101Y118_SLICE_X159Y118_C5 = 1'b1;
  assign CLBLM_R_X101Y118_SLICE_X159Y118_D1 = 1'b1;
  assign CLBLM_R_X101Y118_SLICE_X159Y118_D2 = 1'b1;
  assign CLBLM_R_X101Y118_SLICE_X159Y118_D3 = 1'b1;
  assign CLBLM_R_X101Y118_SLICE_X159Y118_D4 = 1'b1;
  assign CLBLM_R_X101Y118_SLICE_X159Y118_D5 = 1'b1;
  assign CLBLM_R_X101Y118_SLICE_X159Y118_D6 = 1'b1;
  assign CLBLM_R_X103Y102_SLICE_X162Y102_A4 = 1'b1;
  assign CLBLM_R_X103Y102_SLICE_X162Y102_A6 = 1'b1;
  assign CLBLM_R_X103Y102_SLICE_X162Y102_B1 = 1'b1;
  assign CLBLM_R_X103Y102_SLICE_X162Y102_B2 = 1'b1;
  assign CLBLM_R_X101Y118_SLICE_X158Y118_A1 = CLBLM_R_X5Y115_SLICE_X6Y115_BO5;
  assign CLBLM_R_X101Y118_SLICE_X158Y118_A2 = CLBLM_L_X10Y123_SLICE_X12Y123_AO6;
  assign CLBLM_R_X101Y118_SLICE_X158Y118_A3 = CLBLM_R_X101Y117_SLICE_X158Y117_AO6;
  assign CLBLM_R_X101Y118_SLICE_X158Y118_A4 = CLBLL_L_X100Y123_SLICE_X156Y123_BO6;
  assign CLBLM_R_X101Y118_SLICE_X158Y118_A5 = CLBLM_R_X5Y111_SLICE_X6Y111_AO6;
  assign CLBLM_R_X101Y118_SLICE_X158Y118_A6 = CLBLM_R_X5Y111_SLICE_X7Y111_AO6;
  assign CLBLM_R_X103Y102_SLICE_X162Y102_B5 = 1'b1;
  assign CLBLM_R_X103Y102_SLICE_X162Y102_B6 = 1'b1;
  assign CLBLM_R_X103Y102_SLICE_X162Y102_C1 = 1'b1;
  assign CLBLM_R_X101Y118_SLICE_X158Y118_B1 = CLBLM_R_X5Y115_SLICE_X6Y115_BO5;
  assign CLBLM_R_X101Y118_SLICE_X158Y118_B2 = CLBLM_L_X10Y123_SLICE_X12Y123_AO6;
  assign CLBLM_R_X101Y118_SLICE_X158Y118_B3 = CLBLM_R_X101Y117_SLICE_X158Y117_AO6;
  assign CLBLM_R_X101Y118_SLICE_X158Y118_B4 = CLBLL_L_X100Y123_SLICE_X156Y123_AO6;
  assign CLBLM_R_X101Y118_SLICE_X158Y118_B5 = CLBLM_R_X5Y111_SLICE_X6Y111_AO6;
  assign CLBLM_R_X101Y118_SLICE_X158Y118_B6 = CLBLM_R_X5Y111_SLICE_X7Y111_AO6;
  assign CLBLM_R_X103Y102_SLICE_X162Y102_C5 = 1'b1;
  assign CLBLM_R_X103Y102_SLICE_X162Y102_C6 = 1'b1;
  assign CLBLM_R_X103Y102_SLICE_X162Y102_D1 = 1'b1;
  assign CLBLM_R_X101Y118_SLICE_X158Y118_C1 = CLBLM_R_X5Y111_SLICE_X6Y111_AO6;
  assign CLBLM_R_X101Y118_SLICE_X158Y118_C2 = CLBLM_R_X101Y116_SLICE_X158Y116_AO6;
  assign CLBLM_R_X101Y118_SLICE_X158Y118_C3 = CLBLM_R_X5Y115_SLICE_X6Y115_BO5;
  assign CLBLM_R_X101Y118_SLICE_X158Y118_C4 = CLBLM_R_X5Y111_SLICE_X7Y111_AO6;
  assign CLBLM_R_X101Y118_SLICE_X158Y118_C5 = CLBLM_R_X103Y122_SLICE_X163Y122_AO5;
  assign CLBLM_R_X101Y118_SLICE_X158Y118_C6 = CLBLM_L_X10Y123_SLICE_X12Y123_AO6;
  assign CLBLM_R_X103Y102_SLICE_X162Y102_D3 = 1'b1;
  assign CLBLM_R_X103Y102_SLICE_X162Y102_D4 = 1'b1;
  assign CLBLM_R_X103Y102_SLICE_X162Y102_D5 = 1'b1;
  assign CLBLM_R_X103Y102_SLICE_X162Y102_D6 = 1'b1;
  assign LIOI3_TBYTESRC_X0Y93_ILOGIC_X0Y94_D = LIOB33_X0Y93_IOB_X0Y94_I;
  assign LIOI3_TBYTESRC_X0Y93_ILOGIC_X0Y93_D = LIOB33_X0Y93_IOB_X0Y93_I;
  assign CLBLM_R_X101Y118_SLICE_X158Y118_D1 = CLBLM_R_X5Y111_SLICE_X6Y111_AO6;
  assign CLBLM_R_X101Y118_SLICE_X158Y118_D2 = CLBLM_R_X101Y116_SLICE_X158Y116_AO6;
  assign CLBLM_R_X101Y118_SLICE_X158Y118_D3 = CLBLM_R_X5Y115_SLICE_X6Y115_BO5;
  assign CLBLM_R_X101Y118_SLICE_X158Y118_D4 = CLBLM_R_X5Y111_SLICE_X7Y111_AO6;
  assign CLBLM_R_X101Y118_SLICE_X158Y118_D5 = CLBLM_R_X103Y122_SLICE_X163Y122_BO5;
  assign CLBLM_R_X101Y118_SLICE_X158Y118_D6 = CLBLM_L_X10Y123_SLICE_X12Y123_AO6;
  assign RIOI3_TBYTESRC_X105Y157_ILOGIC_X1Y158_D = RIOB33_X105Y157_IOB_X1Y158_I;
  assign RIOI3_TBYTESRC_X105Y157_ILOGIC_X1Y157_D = RIOB33_X105Y157_IOB_X1Y157_I;
  assign CLBLL_L_X100Y123_SLICE_X156Y123_A1 = 1'b1;
  assign CLBLL_L_X100Y123_SLICE_X156Y123_A2 = LIOB33_X0Y157_IOB_X0Y157_I;
  assign CLBLL_L_X100Y123_SLICE_X156Y123_A3 = 1'b1;
  assign CLBLL_L_X100Y123_SLICE_X156Y123_A4 = CLBLM_R_X7Y121_SLICE_X8Y121_AO6;
  assign CLBLL_L_X100Y123_SLICE_X156Y123_A5 = LIOB33_X0Y157_IOB_X0Y158_I;
  assign CLBLL_L_X100Y123_SLICE_X156Y123_A6 = 1'b1;
  assign CLBLL_L_X100Y123_SLICE_X156Y123_B1 = LIOB33_X0Y153_IOB_X0Y154_I;
  assign CLBLL_L_X100Y123_SLICE_X156Y123_B2 = CLBLM_R_X7Y121_SLICE_X8Y121_AO6;
  assign CLBLL_L_X100Y123_SLICE_X156Y123_B3 = 1'b1;
  assign CLBLL_L_X100Y123_SLICE_X156Y123_B4 = 1'b1;
  assign CLBLL_L_X100Y123_SLICE_X156Y123_B5 = LIOB33_X0Y155_IOB_X0Y156_I;
  assign CLBLL_L_X100Y123_SLICE_X156Y123_B6 = 1'b1;
  assign CLBLL_L_X100Y123_SLICE_X156Y123_C1 = 1'b1;
  assign CLBLL_L_X100Y123_SLICE_X156Y123_C2 = 1'b1;
  assign CLBLL_L_X100Y123_SLICE_X156Y123_C3 = 1'b1;
  assign CLBLL_L_X100Y123_SLICE_X156Y123_C4 = 1'b1;
  assign CLBLL_L_X100Y123_SLICE_X156Y123_C5 = 1'b1;
  assign CLBLL_L_X100Y123_SLICE_X156Y123_C6 = 1'b1;
  assign LIOI3_X0Y147_ILOGIC_X0Y147_D = LIOB33_X0Y147_IOB_X0Y147_I;
  assign CLBLL_L_X100Y123_SLICE_X156Y123_D1 = 1'b1;
  assign CLBLL_L_X100Y123_SLICE_X156Y123_D2 = 1'b1;
  assign CLBLL_L_X100Y123_SLICE_X156Y123_D3 = 1'b1;
  assign CLBLL_L_X100Y123_SLICE_X156Y123_D4 = 1'b1;
  assign CLBLL_L_X100Y123_SLICE_X156Y123_D5 = 1'b1;
  assign CLBLL_L_X100Y123_SLICE_X156Y123_D6 = 1'b1;
  assign LIOI3_SING_X0Y99_ILOGIC_X0Y99_D = LIOB33_SING_X0Y99_IOB_X0Y99_I;
  assign LIOI3_X0Y51_ILOGIC_X0Y52_D = LIOB33_X0Y51_IOB_X0Y52_I;
  assign CLBLL_L_X100Y123_SLICE_X157Y123_A1 = 1'b1;
  assign CLBLL_L_X100Y123_SLICE_X157Y123_A2 = 1'b1;
  assign CLBLL_L_X100Y123_SLICE_X157Y123_A3 = 1'b1;
  assign CLBLL_L_X100Y123_SLICE_X157Y123_A4 = 1'b1;
  assign CLBLL_L_X100Y123_SLICE_X157Y123_A5 = 1'b1;
  assign CLBLL_L_X100Y123_SLICE_X157Y123_A6 = 1'b1;
  assign CLBLL_L_X100Y123_SLICE_X157Y123_B1 = 1'b1;
  assign CLBLL_L_X100Y123_SLICE_X157Y123_B2 = 1'b1;
  assign CLBLL_L_X100Y123_SLICE_X157Y123_B3 = 1'b1;
  assign CLBLL_L_X100Y123_SLICE_X157Y123_B4 = 1'b1;
  assign CLBLL_L_X100Y123_SLICE_X157Y123_B5 = 1'b1;
  assign CLBLL_L_X100Y123_SLICE_X157Y123_B6 = 1'b1;
  assign LIOI3_X0Y51_ILOGIC_X0Y51_D = LIOB33_X0Y51_IOB_X0Y51_I;
  assign CLBLL_L_X100Y123_SLICE_X157Y123_C1 = 1'b1;
  assign CLBLL_L_X100Y123_SLICE_X157Y123_C2 = 1'b1;
  assign CLBLL_L_X100Y123_SLICE_X157Y123_C3 = 1'b1;
  assign CLBLL_L_X100Y123_SLICE_X157Y123_C4 = 1'b1;
  assign CLBLL_L_X100Y123_SLICE_X157Y123_C5 = 1'b1;
  assign CLBLL_L_X100Y123_SLICE_X157Y123_C6 = 1'b1;
  assign CLBLL_L_X100Y123_SLICE_X157Y123_D1 = 1'b1;
  assign CLBLL_L_X100Y123_SLICE_X157Y123_D2 = 1'b1;
  assign CLBLL_L_X100Y123_SLICE_X157Y123_D3 = 1'b1;
  assign CLBLL_L_X100Y123_SLICE_X157Y123_D4 = 1'b1;
  assign CLBLL_L_X100Y123_SLICE_X157Y123_D5 = 1'b1;
  assign CLBLL_L_X100Y123_SLICE_X157Y123_D6 = 1'b1;
  assign CLBLM_R_X101Y119_SLICE_X159Y119_A1 = 1'b1;
  assign CLBLM_R_X101Y119_SLICE_X159Y119_A2 = 1'b1;
  assign CLBLM_R_X101Y119_SLICE_X159Y119_A3 = 1'b1;
  assign CLBLM_R_X101Y119_SLICE_X159Y119_A4 = 1'b1;
  assign CLBLM_R_X101Y119_SLICE_X159Y119_A5 = 1'b1;
  assign CLBLM_R_X101Y119_SLICE_X159Y119_A6 = 1'b1;
  assign CLBLM_R_X101Y119_SLICE_X159Y119_B1 = 1'b1;
  assign CLBLM_R_X101Y119_SLICE_X159Y119_B2 = 1'b1;
  assign CLBLM_R_X101Y119_SLICE_X159Y119_B3 = 1'b1;
  assign CLBLM_R_X101Y119_SLICE_X159Y119_B4 = 1'b1;
  assign CLBLM_R_X101Y119_SLICE_X159Y119_B5 = 1'b1;
  assign CLBLM_R_X101Y119_SLICE_X159Y119_B6 = 1'b1;
  assign CLBLM_R_X101Y119_SLICE_X159Y119_C1 = 1'b1;
  assign CLBLM_R_X101Y119_SLICE_X159Y119_C2 = 1'b1;
  assign CLBLM_R_X101Y119_SLICE_X159Y119_C3 = 1'b1;
  assign CLBLM_R_X101Y119_SLICE_X159Y119_C4 = 1'b1;
  assign CLBLM_R_X101Y119_SLICE_X159Y119_C5 = 1'b1;
  assign CLBLM_R_X101Y119_SLICE_X159Y119_C6 = 1'b1;
  assign CLBLM_R_X101Y119_SLICE_X159Y119_D1 = 1'b1;
  assign CLBLM_R_X101Y119_SLICE_X159Y119_D2 = 1'b1;
  assign CLBLM_R_X101Y119_SLICE_X159Y119_D3 = 1'b1;
  assign CLBLM_R_X101Y119_SLICE_X159Y119_D4 = 1'b1;
  assign CLBLM_R_X101Y119_SLICE_X159Y119_D5 = 1'b1;
  assign CLBLM_R_X101Y119_SLICE_X159Y119_D6 = 1'b1;
  assign CLBLM_R_X101Y119_SLICE_X158Y119_A1 = CLBLM_L_X10Y123_SLICE_X12Y123_AO6;
  assign CLBLM_R_X101Y119_SLICE_X158Y119_A2 = CLBLL_L_X100Y123_SLICE_X156Y123_BO6;
  assign CLBLM_R_X101Y119_SLICE_X158Y119_A3 = CLBLM_R_X5Y111_SLICE_X7Y111_AO5;
  assign CLBLM_R_X101Y119_SLICE_X158Y119_A4 = CLBLM_L_X56Y119_SLICE_X84Y119_AO6;
  assign CLBLM_R_X101Y119_SLICE_X158Y119_A5 = CLBLM_R_X5Y111_SLICE_X6Y111_AO6;
  assign CLBLM_R_X101Y119_SLICE_X158Y119_A6 = CLBLM_R_X25Y115_SLICE_X36Y115_AO5;
  assign CLBLM_R_X101Y119_SLICE_X158Y119_B1 = CLBLM_L_X56Y119_SLICE_X84Y119_AO6;
  assign CLBLM_R_X101Y119_SLICE_X158Y119_B2 = CLBLM_L_X10Y123_SLICE_X12Y123_AO6;
  assign CLBLM_R_X101Y119_SLICE_X158Y119_B3 = CLBLM_R_X5Y111_SLICE_X7Y111_AO5;
  assign CLBLM_R_X101Y119_SLICE_X158Y119_B4 = CLBLL_L_X100Y123_SLICE_X156Y123_AO6;
  assign CLBLM_R_X101Y119_SLICE_X158Y119_B5 = CLBLM_R_X5Y111_SLICE_X6Y111_AO6;
  assign CLBLM_R_X101Y119_SLICE_X158Y119_B6 = CLBLM_R_X25Y115_SLICE_X36Y115_AO5;
  assign CLBLM_R_X101Y119_SLICE_X158Y119_C1 = CLBLM_R_X5Y111_SLICE_X6Y111_AO6;
  assign CLBLM_R_X101Y119_SLICE_X158Y119_C2 = CLBLM_R_X25Y115_SLICE_X36Y115_AO5;
  assign CLBLM_R_X101Y119_SLICE_X158Y119_C3 = CLBLM_R_X5Y111_SLICE_X7Y111_AO5;
  assign CLBLM_R_X101Y119_SLICE_X158Y119_C4 = CLBLM_R_X103Y122_SLICE_X163Y122_AO5;
  assign CLBLM_R_X101Y119_SLICE_X158Y119_C5 = CLBLM_L_X56Y119_SLICE_X84Y119_AO5;
  assign CLBLM_R_X101Y119_SLICE_X158Y119_C6 = CLBLM_L_X10Y123_SLICE_X12Y123_AO6;
  assign CLBLM_R_X101Y119_SLICE_X158Y119_D1 = CLBLM_R_X5Y111_SLICE_X7Y111_AO5;
  assign CLBLM_R_X101Y119_SLICE_X158Y119_D2 = CLBLM_R_X103Y122_SLICE_X163Y122_BO5;
  assign CLBLM_R_X101Y119_SLICE_X158Y119_D3 = CLBLM_L_X56Y119_SLICE_X84Y119_AO5;
  assign CLBLM_R_X101Y119_SLICE_X158Y119_D4 = CLBLM_R_X25Y115_SLICE_X36Y115_AO5;
  assign CLBLM_R_X101Y119_SLICE_X158Y119_D5 = CLBLM_L_X10Y123_SLICE_X12Y123_AO6;
  assign CLBLM_R_X101Y119_SLICE_X158Y119_D6 = CLBLM_R_X5Y111_SLICE_X6Y111_AO6;
  assign LIOI3_X0Y79_ILOGIC_X0Y80_D = LIOB33_X0Y79_IOB_X0Y80_I;
  assign LIOI3_X0Y79_ILOGIC_X0Y79_D = LIOB33_X0Y79_IOB_X0Y79_I;
  assign CLBLL_L_X100Y113_SLICE_X157Y113_B1 = 1'b1;
  assign LIOI3_SING_X0Y100_ILOGIC_X0Y100_D = LIOB33_SING_X0Y100_IOB_X0Y100_I;
  assign LIOI3_X0Y183_OLOGIC_X0Y184_D1 = CLBLM_R_X103Y108_SLICE_X163Y108_AO5;
  assign LIOI3_X0Y183_OLOGIC_X0Y184_T1 = 1'b1;
  assign CLBLL_L_X100Y113_SLICE_X157Y113_C1 = 1'b1;
  assign RIOB33_X105Y51_IOB_X1Y52_O = CLBLM_R_X49Y95_SLICE_X74Y95_AO6;
  assign RIOB33_X105Y51_IOB_X1Y51_O = CLBLL_L_X4Y111_SLICE_X5Y111_CO6;
  assign RIOI3_X105Y197_OLOGIC_X1Y198_D1 = CLBLL_L_X2Y173_SLICE_X1Y173_AO6;
  assign LIOI3_X0Y183_OLOGIC_X0Y183_D1 = LIOB33_X0Y101_IOB_X0Y102_I;
  assign CLBLL_L_X100Y113_SLICE_X157Y113_C2 = 1'b1;
  assign RIOI3_X105Y197_OLOGIC_X1Y198_T1 = 1'b1;
  assign LIOI3_X0Y183_OLOGIC_X0Y183_T1 = 1'b1;
  assign RIOI3_X105Y135_OLOGIC_X1Y136_D1 = CLBLM_R_X101Y118_SLICE_X158Y118_CO6;
  assign RIOI3_X105Y197_OLOGIC_X1Y197_D1 = CLBLL_L_X2Y173_SLICE_X1Y173_AO6;
  assign RIOI3_X105Y135_OLOGIC_X1Y136_T1 = 1'b1;
  assign RIOI3_X105Y75_OLOGIC_X1Y76_D1 = CLBLL_R_X57Y113_SLICE_X86Y113_BO6;
  assign RIOI3_X105Y197_OLOGIC_X1Y197_T1 = 1'b1;
  assign RIOI3_X105Y135_OLOGIC_X1Y135_D1 = CLBLM_R_X101Y119_SLICE_X158Y119_CO6;
  assign RIOI3_X105Y75_OLOGIC_X1Y76_T1 = 1'b1;
  assign LIOI3_X0Y111_ILOGIC_X0Y112_D = LIOB33_X0Y111_IOB_X0Y112_I;
  assign RIOI3_X105Y135_OLOGIC_X1Y135_T1 = 1'b1;
  assign RIOI3_X105Y75_OLOGIC_X1Y75_D1 = CLBLM_R_X29Y115_SLICE_X42Y115_AO6;
  assign RIOI3_X105Y75_OLOGIC_X1Y75_T1 = 1'b1;
  assign LIOI3_X0Y111_ILOGIC_X0Y111_D = LIOB33_X0Y111_IOB_X0Y111_I;
  assign CLBLM_R_X103Y107_SLICE_X163Y107_C3 = 1'b1;
  assign CLBLM_R_X103Y107_SLICE_X163Y107_C4 = 1'b1;
  assign CLBLM_R_X103Y107_SLICE_X163Y107_C5 = 1'b1;
  assign RIOI3_X105Y109_ILOGIC_X1Y109_D = RIOB33_X105Y109_IOB_X1Y109_I;
  assign LIOI3_X0Y153_ILOGIC_X0Y154_D = LIOB33_X0Y153_IOB_X0Y154_I;
  assign LIOI3_X0Y153_ILOGIC_X0Y153_D = LIOB33_X0Y153_IOB_X0Y153_I;
  assign LIOI3_X0Y123_ILOGIC_X0Y124_D = LIOB33_X0Y123_IOB_X0Y124_I;
  assign CLBLL_L_X2Y136_SLICE_X0Y136_A1 = LIOB33_X0Y137_IOB_X0Y138_I;
  assign CLBLL_L_X2Y136_SLICE_X0Y136_A2 = LIOB33_X0Y109_IOB_X0Y110_I;
  assign CLBLL_L_X2Y136_SLICE_X0Y136_A3 = LIOB33_X0Y135_IOB_X0Y136_I;
  assign CLBLL_L_X2Y136_SLICE_X0Y136_A4 = LIOB33_X0Y135_IOB_X0Y135_I;
  assign CLBLL_L_X2Y136_SLICE_X0Y136_A5 = LIOB33_X0Y67_IOB_X0Y67_I;
  assign CLBLL_L_X2Y136_SLICE_X0Y136_A6 = LIOB33_X0Y137_IOB_X0Y137_I;
  assign CLBLM_R_X103Y107_SLICE_X163Y107_D1 = 1'b1;
  assign LIOI3_X0Y91_ILOGIC_X0Y92_D = LIOB33_X0Y91_IOB_X0Y92_I;
  assign LIOI3_X0Y123_ILOGIC_X0Y123_D = LIOB33_X0Y123_IOB_X0Y123_I;
  assign CLBLL_L_X2Y136_SLICE_X0Y136_B1 = 1'b1;
  assign CLBLL_L_X2Y136_SLICE_X0Y136_B2 = 1'b1;
  assign CLBLL_L_X2Y136_SLICE_X0Y136_B3 = LIOB33_X0Y109_IOB_X0Y110_I;
  assign CLBLL_L_X2Y136_SLICE_X0Y136_B4 = 1'b1;
  assign CLBLL_L_X2Y136_SLICE_X0Y136_B5 = LIOB33_X0Y135_IOB_X0Y136_I;
  assign CLBLL_L_X2Y136_SLICE_X0Y136_B6 = 1'b1;
  assign LIOI3_X0Y61_ILOGIC_X0Y62_D = LIOB33_X0Y61_IOB_X0Y62_I;
  assign LIOI3_X0Y91_ILOGIC_X0Y91_D = LIOB33_X0Y91_IOB_X0Y91_I;
  assign RIOI3_X105Y167_ILOGIC_X1Y168_D = RIOB33_X105Y167_IOB_X1Y168_I;
  assign CLBLL_L_X2Y136_SLICE_X0Y136_C1 = 1'b1;
  assign CLBLL_L_X2Y136_SLICE_X0Y136_C2 = 1'b1;
  assign CLBLL_L_X2Y136_SLICE_X0Y136_C3 = 1'b1;
  assign CLBLL_L_X2Y136_SLICE_X0Y136_C4 = 1'b1;
  assign CLBLL_L_X2Y136_SLICE_X0Y136_C5 = 1'b1;
  assign CLBLL_L_X2Y136_SLICE_X0Y136_C6 = 1'b1;
  assign CLBLM_R_X103Y107_SLICE_X163Y107_D5 = 1'b1;
  assign RIOI3_X105Y105_ILOGIC_X1Y106_D = RIOB33_X105Y105_IOB_X1Y106_I;
  assign CLBLM_R_X103Y107_SLICE_X163Y107_D6 = 1'b1;
  assign RIOI3_X105Y105_ILOGIC_X1Y105_D = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLL_L_X2Y136_SLICE_X0Y136_D1 = 1'b1;
  assign CLBLL_L_X2Y136_SLICE_X0Y136_D2 = 1'b1;
  assign CLBLL_L_X2Y136_SLICE_X0Y136_D3 = 1'b1;
  assign CLBLL_L_X2Y136_SLICE_X0Y136_D4 = 1'b1;
  assign CLBLL_L_X2Y136_SLICE_X0Y136_D5 = 1'b1;
  assign CLBLL_L_X2Y136_SLICE_X0Y136_D6 = 1'b1;
  assign RIOB33_SING_X105Y50_IOB_X1Y50_O = CLBLM_R_X49Y95_SLICE_X74Y95_AO6;
  assign LIOI3_TBYTESRC_X0Y107_ILOGIC_X0Y108_D = LIOB33_X0Y107_IOB_X0Y108_I;
  assign LIOI3_TBYTESRC_X0Y107_ILOGIC_X0Y107_D = LIOB33_X0Y107_IOB_X0Y107_I;
  assign LIOI3_TBYTESRC_X0Y119_ILOGIC_X0Y120_D = LIOB33_X0Y119_IOB_X0Y120_I;
  assign RIOI3_TBYTETERM_X105Y113_ILOGIC_X1Y114_D = RIOB33_X105Y113_IOB_X1Y114_I;
  assign RIOI3_TBYTETERM_X105Y113_ILOGIC_X1Y113_D = RIOB33_X105Y113_IOB_X1Y113_I;
  assign LIOI3_X0Y141_ILOGIC_X0Y142_D = LIOB33_X0Y141_IOB_X0Y142_I;
  assign RIOI3_TBYTESRC_X105Y169_ILOGIC_X1Y170_D = RIOB33_X105Y169_IOB_X1Y170_I;
  assign CLBLL_L_X2Y136_SLICE_X1Y136_A1 = 1'b1;
  assign CLBLL_L_X2Y136_SLICE_X1Y136_A2 = 1'b1;
  assign CLBLL_L_X2Y136_SLICE_X1Y136_A3 = 1'b1;
  assign CLBLL_L_X2Y136_SLICE_X1Y136_A4 = 1'b1;
  assign CLBLL_L_X2Y136_SLICE_X1Y136_A5 = 1'b1;
  assign CLBLL_L_X2Y136_SLICE_X1Y136_A6 = 1'b1;
  assign RIOI3_TBYTESRC_X105Y169_ILOGIC_X1Y169_D = RIOB33_X105Y169_IOB_X1Y169_I;
  assign CLBLL_L_X2Y136_SLICE_X1Y136_B1 = 1'b1;
  assign CLBLL_L_X2Y136_SLICE_X1Y136_B2 = 1'b1;
  assign CLBLL_L_X2Y136_SLICE_X1Y136_B3 = 1'b1;
  assign CLBLL_L_X2Y136_SLICE_X1Y136_B4 = 1'b1;
  assign CLBLL_L_X2Y136_SLICE_X1Y136_B5 = 1'b1;
  assign CLBLL_L_X2Y136_SLICE_X1Y136_B6 = 1'b1;
  assign RIOB33_X105Y53_IOB_X1Y53_O = CLBLM_L_X10Y113_SLICE_X12Y113_AO6;
  assign LIOI3_X0Y141_ILOGIC_X0Y141_D = LIOB33_X0Y141_IOB_X0Y141_I;
  assign RIOB33_X105Y53_IOB_X1Y54_O = CLBLM_R_X103Y108_SLICE_X163Y108_AO6;
  assign CLBLL_L_X2Y136_SLICE_X1Y136_C1 = 1'b1;
  assign CLBLL_L_X2Y136_SLICE_X1Y136_C2 = 1'b1;
  assign CLBLL_L_X2Y136_SLICE_X1Y136_C3 = 1'b1;
  assign CLBLL_L_X2Y136_SLICE_X1Y136_C4 = 1'b1;
  assign CLBLL_L_X2Y136_SLICE_X1Y136_C5 = 1'b1;
  assign CLBLL_L_X2Y136_SLICE_X1Y136_C6 = 1'b1;
  assign CLBLM_R_X103Y107_SLICE_X162Y107_A6 = 1'b1;
  assign CLBLL_L_X2Y136_SLICE_X1Y136_D1 = 1'b1;
  assign CLBLL_L_X2Y136_SLICE_X1Y136_D2 = 1'b1;
  assign CLBLL_L_X2Y136_SLICE_X1Y136_D3 = 1'b1;
  assign CLBLL_L_X2Y136_SLICE_X1Y136_D4 = 1'b1;
  assign CLBLL_L_X2Y136_SLICE_X1Y136_D5 = 1'b1;
  assign CLBLL_L_X2Y136_SLICE_X1Y136_D6 = 1'b1;
  assign RIOI3_TBYTESRC_X105Y131_OLOGIC_X1Y132_D1 = CLBLM_R_X101Y119_SLICE_X158Y119_AO6;
  assign CLBLM_R_X103Y107_SLICE_X162Y107_B3 = 1'b1;
  assign CLBLM_R_X103Y107_SLICE_X162Y107_B4 = 1'b1;
  assign CLBLM_R_X103Y107_SLICE_X162Y107_B5 = 1'b1;
  assign CLBLM_R_X103Y107_SLICE_X162Y107_B6 = 1'b1;
  assign CLBLM_R_X103Y102_SLICE_X163Y102_B2 = CLBLM_L_X10Y113_SLICE_X12Y113_BO6;
  assign LIOI3_TBYTESRC_X0Y119_ILOGIC_X0Y119_D = LIOB33_X0Y119_IOB_X0Y119_I;
  assign CLBLM_R_X103Y102_SLICE_X163Y102_B3 = 1'b1;
  assign CLBLM_R_X103Y102_SLICE_X163Y102_B4 = RIOB33_X105Y109_IOB_X1Y110_I;
  assign CLBLM_R_X103Y102_SLICE_X163Y102_B5 = CLBLM_R_X103Y122_SLICE_X163Y122_BO5;
  assign RIOI3_TBYTESRC_X105Y131_OLOGIC_X1Y132_T1 = 1'b1;
  assign RIOB33_X105Y173_IOB_X1Y174_O = LIOB33_X0Y133_IOB_X0Y133_I;
  assign CLBLM_R_X103Y102_SLICE_X163Y102_B6 = RIOB33_X105Y109_IOB_X1Y109_I;
  assign RIOB33_X105Y173_IOB_X1Y173_O = CLBLM_R_X103Y147_SLICE_X163Y147_AO5;
  assign RIOB33_SING_X105Y99_IOB_X1Y99_O = CLBLM_R_X101Y119_SLICE_X158Y119_BO6;
  assign CLBLM_R_X103Y107_SLICE_X162Y107_C1 = 1'b1;
  assign CLBLM_R_X103Y107_SLICE_X162Y107_C2 = 1'b1;
  assign CLBLM_R_X103Y107_SLICE_X162Y107_C3 = 1'b1;
  assign CLBLM_R_X103Y107_SLICE_X162Y107_C4 = 1'b1;
  assign CLBLM_R_X103Y102_SLICE_X163Y102_C1 = 1'b1;
  assign CLBLM_R_X103Y107_SLICE_X162Y107_C5 = 1'b1;
  assign CLBLM_R_X103Y102_SLICE_X163Y102_C2 = 1'b1;
  assign CLBLM_R_X103Y107_SLICE_X162Y107_C6 = 1'b1;
  assign CLBLM_R_X103Y102_SLICE_X163Y102_C3 = 1'b1;
  assign CLBLM_R_X103Y102_SLICE_X163Y102_C4 = 1'b1;
  assign CLBLM_R_X103Y102_SLICE_X163Y102_C5 = 1'b1;
  assign CLBLM_R_X103Y102_SLICE_X163Y102_C6 = 1'b1;
  assign RIOI3_TBYTESRC_X105Y131_OLOGIC_X1Y131_D1 = CLBLM_R_X101Y118_SLICE_X158Y118_AO6;
  assign CLBLM_R_X103Y107_SLICE_X162Y107_D1 = 1'b1;
  assign CLBLM_R_X103Y107_SLICE_X162Y107_D2 = 1'b1;
  assign CLBLM_R_X103Y107_SLICE_X162Y107_D3 = 1'b1;
  assign CLBLM_R_X103Y102_SLICE_X163Y102_D1 = 1'b1;
  assign CLBLM_R_X103Y107_SLICE_X162Y107_D4 = 1'b1;
  assign CLBLM_R_X103Y102_SLICE_X163Y102_D2 = 1'b1;
  assign CLBLM_R_X103Y107_SLICE_X162Y107_D5 = 1'b1;
  assign CLBLM_R_X103Y102_SLICE_X163Y102_D3 = 1'b1;
  assign LIOI3_X0Y173_ILOGIC_X0Y174_D = LIOB33_X0Y173_IOB_X0Y174_I;
  assign CLBLM_R_X103Y107_SLICE_X162Y107_D6 = 1'b1;
  assign CLBLM_R_X103Y102_SLICE_X163Y102_D4 = 1'b1;
  assign RIOI3_TBYTESRC_X105Y131_OLOGIC_X1Y131_T1 = 1'b1;
  assign CLBLM_R_X103Y102_SLICE_X163Y102_D5 = 1'b1;
  assign CLBLM_R_X103Y102_SLICE_X163Y102_D6 = 1'b1;
  assign LIOI3_X0Y173_ILOGIC_X0Y173_D = LIOB33_X0Y173_IOB_X0Y173_I;
  assign CLBLM_R_X49Y95_SLICE_X75Y95_A1 = 1'b1;
  assign CLBLM_R_X49Y95_SLICE_X75Y95_A2 = 1'b1;
  assign CLBLM_R_X49Y95_SLICE_X75Y95_A3 = 1'b1;
  assign CLBLM_R_X49Y95_SLICE_X75Y95_A4 = 1'b1;
  assign CLBLM_R_X49Y95_SLICE_X75Y95_A5 = 1'b1;
  assign CLBLM_R_X49Y95_SLICE_X75Y95_A6 = 1'b1;
  assign CLBLM_R_X49Y95_SLICE_X75Y95_B1 = 1'b1;
  assign CLBLM_R_X49Y95_SLICE_X75Y95_B2 = 1'b1;
  assign CLBLM_R_X49Y95_SLICE_X75Y95_B3 = 1'b1;
  assign CLBLM_R_X49Y95_SLICE_X75Y95_B4 = 1'b1;
  assign CLBLM_R_X49Y95_SLICE_X75Y95_B5 = 1'b1;
  assign CLBLM_R_X49Y95_SLICE_X75Y95_B6 = 1'b1;
  assign CLBLM_R_X103Y102_SLICE_X162Y102_A1 = 1'b1;
  assign CLBLM_R_X49Y95_SLICE_X75Y95_C1 = 1'b1;
  assign CLBLM_R_X49Y95_SLICE_X75Y95_C2 = 1'b1;
  assign CLBLM_R_X49Y95_SLICE_X75Y95_C3 = 1'b1;
  assign CLBLM_R_X49Y95_SLICE_X75Y95_C4 = 1'b1;
  assign CLBLM_R_X49Y95_SLICE_X75Y95_C5 = 1'b1;
  assign CLBLM_R_X49Y95_SLICE_X75Y95_C6 = 1'b1;
  assign CLBLM_R_X103Y102_SLICE_X162Y102_A2 = 1'b1;
  assign CLBLM_R_X103Y102_SLICE_X162Y102_A3 = 1'b1;
  assign CLBLM_R_X49Y95_SLICE_X75Y95_D1 = 1'b1;
  assign CLBLM_R_X49Y95_SLICE_X75Y95_D2 = 1'b1;
  assign CLBLM_R_X49Y95_SLICE_X75Y95_D3 = 1'b1;
  assign CLBLM_R_X49Y95_SLICE_X75Y95_D4 = 1'b1;
  assign CLBLM_R_X49Y95_SLICE_X75Y95_D5 = 1'b1;
  assign CLBLM_R_X49Y95_SLICE_X75Y95_D6 = 1'b1;
  assign CLBLM_R_X103Y102_SLICE_X162Y102_A5 = 1'b1;
  assign RIOB33_X105Y55_IOB_X1Y56_O = CLBLM_R_X5Y111_SLICE_X7Y111_BO6;
  assign RIOB33_X105Y55_IOB_X1Y55_O = CLBLM_L_X10Y114_SLICE_X12Y114_AO6;
  assign CLBLM_R_X49Y95_SLICE_X74Y95_A1 = 1'b1;
  assign CLBLM_R_X49Y95_SLICE_X74Y95_A2 = CLBLM_R_X5Y113_SLICE_X6Y113_AO6;
  assign CLBLM_R_X49Y95_SLICE_X74Y95_A3 = LIOB33_X0Y83_IOB_X0Y84_I;
  assign CLBLM_R_X49Y95_SLICE_X74Y95_A4 = LIOB33_X0Y85_IOB_X0Y85_I;
  assign CLBLM_R_X49Y95_SLICE_X74Y95_A5 = LIOB33_X0Y95_IOB_X0Y95_I;
  assign CLBLM_R_X49Y95_SLICE_X74Y95_A6 = 1'b1;
  assign CLBLM_R_X49Y95_SLICE_X74Y95_B1 = 1'b1;
  assign CLBLM_R_X49Y95_SLICE_X74Y95_B2 = 1'b1;
  assign CLBLM_R_X49Y95_SLICE_X74Y95_B3 = 1'b1;
  assign CLBLM_R_X49Y95_SLICE_X74Y95_B4 = 1'b1;
  assign CLBLM_R_X49Y95_SLICE_X74Y95_B5 = 1'b1;
  assign CLBLM_R_X49Y95_SLICE_X74Y95_B6 = 1'b1;
  assign CLBLM_R_X49Y95_SLICE_X74Y95_C1 = 1'b1;
  assign CLBLM_R_X49Y95_SLICE_X74Y95_C2 = 1'b1;
  assign CLBLM_R_X49Y95_SLICE_X74Y95_C3 = 1'b1;
  assign CLBLM_R_X49Y95_SLICE_X74Y95_C4 = 1'b1;
  assign CLBLM_R_X49Y95_SLICE_X74Y95_C5 = 1'b1;
  assign CLBLM_R_X49Y95_SLICE_X74Y95_C6 = 1'b1;
  assign CLBLM_R_X103Y102_SLICE_X162Y102_B3 = 1'b1;
  assign CLBLM_R_X49Y95_SLICE_X74Y95_D1 = 1'b1;
  assign CLBLM_R_X49Y95_SLICE_X74Y95_D2 = 1'b1;
  assign CLBLM_R_X49Y95_SLICE_X74Y95_D3 = 1'b1;
  assign CLBLM_R_X49Y95_SLICE_X74Y95_D4 = 1'b1;
  assign CLBLM_R_X49Y95_SLICE_X74Y95_D5 = 1'b1;
  assign CLBLM_R_X49Y95_SLICE_X74Y95_D6 = 1'b1;
  assign CLBLM_R_X103Y102_SLICE_X162Y102_B4 = 1'b1;
endmodule
