module top(
  input LIOB33_SING_X0Y100_IOB_X0Y100_IPAD,
  input LIOB33_X0Y101_IOB_X0Y101_IPAD,
  input LIOB33_X0Y101_IOB_X0Y102_IPAD,
  input LIOB33_X0Y103_IOB_X0Y103_IPAD,
  input LIOB33_X0Y103_IOB_X0Y104_IPAD,
  input LIOB33_X0Y105_IOB_X0Y105_IPAD,
  input LIOB33_X0Y105_IOB_X0Y106_IPAD,
  input LIOB33_X0Y107_IOB_X0Y107_IPAD,
  input LIOB33_X0Y107_IOB_X0Y108_IPAD,
  input LIOB33_X0Y109_IOB_X0Y109_IPAD,
  input LIOB33_X0Y109_IOB_X0Y110_IPAD,
  input LIOB33_X0Y111_IOB_X0Y111_IPAD,
  input LIOB33_X0Y111_IOB_X0Y112_IPAD,
  input LIOB33_X0Y113_IOB_X0Y113_IPAD,
  input LIOB33_X0Y113_IOB_X0Y114_IPAD,
  input LIOB33_X0Y115_IOB_X0Y115_IPAD,
  input LIOB33_X0Y115_IOB_X0Y116_IPAD,
  input LIOB33_X0Y117_IOB_X0Y117_IPAD,
  input RIOB33_SING_X105Y100_IOB_X1Y100_IPAD,
  input RIOB33_X105Y101_IOB_X1Y101_IPAD,
  input RIOB33_X105Y101_IOB_X1Y102_IPAD,
  input RIOB33_X105Y103_IOB_X1Y103_IPAD,
  input RIOB33_X105Y103_IOB_X1Y104_IPAD,
  input RIOB33_X105Y105_IOB_X1Y105_IPAD,
  input RIOB33_X105Y105_IOB_X1Y106_IPAD,
  input RIOB33_X105Y107_IOB_X1Y107_IPAD,
  input RIOB33_X105Y107_IOB_X1Y108_IPAD,
  input RIOB33_X105Y109_IOB_X1Y109_IPAD,
  input RIOB33_X105Y109_IOB_X1Y110_IPAD,
  input RIOB33_X105Y111_IOB_X1Y111_IPAD,
  input RIOB33_X105Y111_IOB_X1Y112_IPAD,
  input RIOB33_X105Y113_IOB_X1Y113_IPAD,
  output LIOB33_SING_X0Y149_IOB_X0Y149_OPAD,
  output LIOB33_X0Y117_IOB_X0Y118_OPAD,
  output LIOB33_X0Y119_IOB_X0Y119_OPAD,
  output LIOB33_X0Y119_IOB_X0Y120_OPAD,
  output LIOB33_X0Y121_IOB_X0Y121_OPAD,
  output LIOB33_X0Y121_IOB_X0Y122_OPAD,
  output LIOB33_X0Y123_IOB_X0Y123_OPAD,
  output LIOB33_X0Y123_IOB_X0Y124_OPAD,
  output LIOB33_X0Y125_IOB_X0Y125_OPAD,
  output LIOB33_X0Y125_IOB_X0Y126_OPAD,
  output LIOB33_X0Y127_IOB_X0Y127_OPAD,
  output LIOB33_X0Y127_IOB_X0Y128_OPAD,
  output LIOB33_X0Y129_IOB_X0Y129_OPAD,
  output LIOB33_X0Y129_IOB_X0Y130_OPAD,
  output LIOB33_X0Y131_IOB_X0Y131_OPAD,
  output LIOB33_X0Y131_IOB_X0Y132_OPAD,
  output LIOB33_X0Y133_IOB_X0Y133_OPAD,
  output LIOB33_X0Y133_IOB_X0Y134_OPAD,
  output LIOB33_X0Y135_IOB_X0Y135_OPAD,
  output LIOB33_X0Y135_IOB_X0Y136_OPAD,
  output LIOB33_X0Y137_IOB_X0Y137_OPAD,
  output LIOB33_X0Y137_IOB_X0Y138_OPAD,
  output LIOB33_X0Y139_IOB_X0Y139_OPAD,
  output LIOB33_X0Y139_IOB_X0Y140_OPAD,
  output LIOB33_X0Y141_IOB_X0Y141_OPAD,
  output LIOB33_X0Y141_IOB_X0Y142_OPAD,
  output LIOB33_X0Y143_IOB_X0Y143_OPAD,
  output LIOB33_X0Y145_IOB_X0Y145_OPAD,
  output LIOB33_X0Y145_IOB_X0Y146_OPAD,
  output LIOB33_X0Y147_IOB_X0Y147_OPAD,
  output LIOB33_X0Y147_IOB_X0Y148_OPAD
  );
  wire [0:0] CLBLL_L_X2Y104_SLICE_X0Y104_A;
  wire [0:0] CLBLL_L_X2Y104_SLICE_X0Y104_A1;
  wire [0:0] CLBLL_L_X2Y104_SLICE_X0Y104_A2;
  wire [0:0] CLBLL_L_X2Y104_SLICE_X0Y104_A3;
  wire [0:0] CLBLL_L_X2Y104_SLICE_X0Y104_A4;
  wire [0:0] CLBLL_L_X2Y104_SLICE_X0Y104_A5;
  wire [0:0] CLBLL_L_X2Y104_SLICE_X0Y104_A6;
  wire [0:0] CLBLL_L_X2Y104_SLICE_X0Y104_AMUX;
  wire [0:0] CLBLL_L_X2Y104_SLICE_X0Y104_AO5;
  wire [0:0] CLBLL_L_X2Y104_SLICE_X0Y104_AO6;
  wire [0:0] CLBLL_L_X2Y104_SLICE_X0Y104_A_CY;
  wire [0:0] CLBLL_L_X2Y104_SLICE_X0Y104_A_XOR;
  wire [0:0] CLBLL_L_X2Y104_SLICE_X0Y104_B;
  wire [0:0] CLBLL_L_X2Y104_SLICE_X0Y104_B1;
  wire [0:0] CLBLL_L_X2Y104_SLICE_X0Y104_B2;
  wire [0:0] CLBLL_L_X2Y104_SLICE_X0Y104_B3;
  wire [0:0] CLBLL_L_X2Y104_SLICE_X0Y104_B4;
  wire [0:0] CLBLL_L_X2Y104_SLICE_X0Y104_B5;
  wire [0:0] CLBLL_L_X2Y104_SLICE_X0Y104_B6;
  wire [0:0] CLBLL_L_X2Y104_SLICE_X0Y104_BMUX;
  wire [0:0] CLBLL_L_X2Y104_SLICE_X0Y104_BO5;
  wire [0:0] CLBLL_L_X2Y104_SLICE_X0Y104_BO6;
  wire [0:0] CLBLL_L_X2Y104_SLICE_X0Y104_B_CY;
  wire [0:0] CLBLL_L_X2Y104_SLICE_X0Y104_B_XOR;
  wire [0:0] CLBLL_L_X2Y104_SLICE_X0Y104_C;
  wire [0:0] CLBLL_L_X2Y104_SLICE_X0Y104_C1;
  wire [0:0] CLBLL_L_X2Y104_SLICE_X0Y104_C2;
  wire [0:0] CLBLL_L_X2Y104_SLICE_X0Y104_C3;
  wire [0:0] CLBLL_L_X2Y104_SLICE_X0Y104_C4;
  wire [0:0] CLBLL_L_X2Y104_SLICE_X0Y104_C5;
  wire [0:0] CLBLL_L_X2Y104_SLICE_X0Y104_C6;
  wire [0:0] CLBLL_L_X2Y104_SLICE_X0Y104_CMUX;
  wire [0:0] CLBLL_L_X2Y104_SLICE_X0Y104_CO5;
  wire [0:0] CLBLL_L_X2Y104_SLICE_X0Y104_CO6;
  wire [0:0] CLBLL_L_X2Y104_SLICE_X0Y104_C_CY;
  wire [0:0] CLBLL_L_X2Y104_SLICE_X0Y104_C_XOR;
  wire [0:0] CLBLL_L_X2Y104_SLICE_X0Y104_D;
  wire [0:0] CLBLL_L_X2Y104_SLICE_X0Y104_D1;
  wire [0:0] CLBLL_L_X2Y104_SLICE_X0Y104_D2;
  wire [0:0] CLBLL_L_X2Y104_SLICE_X0Y104_D3;
  wire [0:0] CLBLL_L_X2Y104_SLICE_X0Y104_D4;
  wire [0:0] CLBLL_L_X2Y104_SLICE_X0Y104_D5;
  wire [0:0] CLBLL_L_X2Y104_SLICE_X0Y104_D6;
  wire [0:0] CLBLL_L_X2Y104_SLICE_X0Y104_DO5;
  wire [0:0] CLBLL_L_X2Y104_SLICE_X0Y104_DO6;
  wire [0:0] CLBLL_L_X2Y104_SLICE_X0Y104_D_CY;
  wire [0:0] CLBLL_L_X2Y104_SLICE_X0Y104_D_XOR;
  wire [0:0] CLBLL_L_X2Y104_SLICE_X1Y104_A;
  wire [0:0] CLBLL_L_X2Y104_SLICE_X1Y104_A1;
  wire [0:0] CLBLL_L_X2Y104_SLICE_X1Y104_A2;
  wire [0:0] CLBLL_L_X2Y104_SLICE_X1Y104_A3;
  wire [0:0] CLBLL_L_X2Y104_SLICE_X1Y104_A4;
  wire [0:0] CLBLL_L_X2Y104_SLICE_X1Y104_A5;
  wire [0:0] CLBLL_L_X2Y104_SLICE_X1Y104_A6;
  wire [0:0] CLBLL_L_X2Y104_SLICE_X1Y104_AMUX;
  wire [0:0] CLBLL_L_X2Y104_SLICE_X1Y104_AO5;
  wire [0:0] CLBLL_L_X2Y104_SLICE_X1Y104_AO6;
  wire [0:0] CLBLL_L_X2Y104_SLICE_X1Y104_A_CY;
  wire [0:0] CLBLL_L_X2Y104_SLICE_X1Y104_A_XOR;
  wire [0:0] CLBLL_L_X2Y104_SLICE_X1Y104_B;
  wire [0:0] CLBLL_L_X2Y104_SLICE_X1Y104_B1;
  wire [0:0] CLBLL_L_X2Y104_SLICE_X1Y104_B2;
  wire [0:0] CLBLL_L_X2Y104_SLICE_X1Y104_B3;
  wire [0:0] CLBLL_L_X2Y104_SLICE_X1Y104_B4;
  wire [0:0] CLBLL_L_X2Y104_SLICE_X1Y104_B5;
  wire [0:0] CLBLL_L_X2Y104_SLICE_X1Y104_B6;
  wire [0:0] CLBLL_L_X2Y104_SLICE_X1Y104_BO5;
  wire [0:0] CLBLL_L_X2Y104_SLICE_X1Y104_BO6;
  wire [0:0] CLBLL_L_X2Y104_SLICE_X1Y104_B_CY;
  wire [0:0] CLBLL_L_X2Y104_SLICE_X1Y104_B_XOR;
  wire [0:0] CLBLL_L_X2Y104_SLICE_X1Y104_C;
  wire [0:0] CLBLL_L_X2Y104_SLICE_X1Y104_C1;
  wire [0:0] CLBLL_L_X2Y104_SLICE_X1Y104_C2;
  wire [0:0] CLBLL_L_X2Y104_SLICE_X1Y104_C3;
  wire [0:0] CLBLL_L_X2Y104_SLICE_X1Y104_C4;
  wire [0:0] CLBLL_L_X2Y104_SLICE_X1Y104_C5;
  wire [0:0] CLBLL_L_X2Y104_SLICE_X1Y104_C6;
  wire [0:0] CLBLL_L_X2Y104_SLICE_X1Y104_CO5;
  wire [0:0] CLBLL_L_X2Y104_SLICE_X1Y104_CO6;
  wire [0:0] CLBLL_L_X2Y104_SLICE_X1Y104_C_CY;
  wire [0:0] CLBLL_L_X2Y104_SLICE_X1Y104_C_XOR;
  wire [0:0] CLBLL_L_X2Y104_SLICE_X1Y104_D;
  wire [0:0] CLBLL_L_X2Y104_SLICE_X1Y104_D1;
  wire [0:0] CLBLL_L_X2Y104_SLICE_X1Y104_D2;
  wire [0:0] CLBLL_L_X2Y104_SLICE_X1Y104_D3;
  wire [0:0] CLBLL_L_X2Y104_SLICE_X1Y104_D4;
  wire [0:0] CLBLL_L_X2Y104_SLICE_X1Y104_D5;
  wire [0:0] CLBLL_L_X2Y104_SLICE_X1Y104_D6;
  wire [0:0] CLBLL_L_X2Y104_SLICE_X1Y104_DO5;
  wire [0:0] CLBLL_L_X2Y104_SLICE_X1Y104_DO6;
  wire [0:0] CLBLL_L_X2Y104_SLICE_X1Y104_D_CY;
  wire [0:0] CLBLL_L_X2Y104_SLICE_X1Y104_D_XOR;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X0Y106_A;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X0Y106_A1;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X0Y106_A2;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X0Y106_A3;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X0Y106_A4;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X0Y106_A5;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X0Y106_A6;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X0Y106_AMUX;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X0Y106_AO5;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X0Y106_AO6;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X0Y106_A_CY;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X0Y106_A_XOR;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X0Y106_B;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X0Y106_B1;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X0Y106_B2;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X0Y106_B3;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X0Y106_B4;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X0Y106_B5;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X0Y106_B6;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X0Y106_BO5;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X0Y106_BO6;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X0Y106_B_CY;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X0Y106_B_XOR;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X0Y106_C;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X0Y106_C1;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X0Y106_C2;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X0Y106_C3;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X0Y106_C4;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X0Y106_C5;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X0Y106_C6;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X0Y106_CO5;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X0Y106_CO6;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X0Y106_C_CY;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X0Y106_C_XOR;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X0Y106_D;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X0Y106_D1;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X0Y106_D2;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X0Y106_D3;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X0Y106_D4;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X0Y106_D5;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X0Y106_D6;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X0Y106_DO5;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X0Y106_DO6;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X0Y106_D_CY;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X0Y106_D_XOR;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X1Y106_A;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X1Y106_A1;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X1Y106_A2;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X1Y106_A3;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X1Y106_A4;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X1Y106_A5;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X1Y106_A6;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X1Y106_AMUX;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X1Y106_AO5;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X1Y106_AO6;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X1Y106_A_CY;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X1Y106_A_XOR;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X1Y106_B;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X1Y106_B1;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X1Y106_B2;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X1Y106_B3;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X1Y106_B4;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X1Y106_B5;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X1Y106_B6;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X1Y106_BO5;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X1Y106_BO6;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X1Y106_B_CY;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X1Y106_B_XOR;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X1Y106_C;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X1Y106_C1;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X1Y106_C2;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X1Y106_C3;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X1Y106_C4;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X1Y106_C5;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X1Y106_C6;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X1Y106_CMUX;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X1Y106_CO5;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X1Y106_CO6;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X1Y106_C_CY;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X1Y106_C_XOR;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X1Y106_D;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X1Y106_D1;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X1Y106_D2;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X1Y106_D3;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X1Y106_D4;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X1Y106_D5;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X1Y106_D6;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X1Y106_DO5;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X1Y106_DO6;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X1Y106_D_CY;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X1Y106_D_XOR;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X0Y107_A;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X0Y107_A1;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X0Y107_A2;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X0Y107_A3;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X0Y107_A4;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X0Y107_A5;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X0Y107_A6;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X0Y107_AO5;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X0Y107_AO6;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X0Y107_A_CY;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X0Y107_A_XOR;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X0Y107_B;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X0Y107_B1;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X0Y107_B2;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X0Y107_B3;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X0Y107_B4;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X0Y107_B5;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X0Y107_B6;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X0Y107_BO5;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X0Y107_BO6;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X0Y107_B_CY;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X0Y107_B_XOR;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X0Y107_C;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X0Y107_C1;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X0Y107_C2;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X0Y107_C3;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X0Y107_C4;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X0Y107_C5;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X0Y107_C6;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X0Y107_CO5;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X0Y107_CO6;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X0Y107_C_CY;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X0Y107_C_XOR;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X0Y107_D;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X0Y107_D1;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X0Y107_D2;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X0Y107_D3;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X0Y107_D4;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X0Y107_D5;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X0Y107_D6;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X0Y107_DO5;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X0Y107_DO6;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X0Y107_D_CY;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X0Y107_D_XOR;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X1Y107_A;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X1Y107_A1;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X1Y107_A2;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X1Y107_A3;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X1Y107_A4;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X1Y107_A5;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X1Y107_A6;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X1Y107_AO5;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X1Y107_AO6;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X1Y107_A_CY;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X1Y107_A_XOR;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X1Y107_B;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X1Y107_B1;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X1Y107_B2;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X1Y107_B3;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X1Y107_B4;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X1Y107_B5;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X1Y107_B6;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X1Y107_BO5;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X1Y107_BO6;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X1Y107_B_CY;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X1Y107_B_XOR;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X1Y107_C;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X1Y107_C1;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X1Y107_C2;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X1Y107_C3;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X1Y107_C4;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X1Y107_C5;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X1Y107_C6;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X1Y107_CO5;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X1Y107_CO6;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X1Y107_C_CY;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X1Y107_C_XOR;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X1Y107_D;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X1Y107_D1;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X1Y107_D2;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X1Y107_D3;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X1Y107_D4;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X1Y107_D5;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X1Y107_D6;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X1Y107_DO5;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X1Y107_DO6;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X1Y107_D_CY;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X1Y107_D_XOR;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X0Y109_A;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X0Y109_A1;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X0Y109_A2;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X0Y109_A3;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X0Y109_A4;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X0Y109_A5;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X0Y109_A6;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X0Y109_AMUX;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X0Y109_AO5;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X0Y109_AO6;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X0Y109_A_CY;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X0Y109_A_XOR;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X0Y109_B;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X0Y109_B1;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X0Y109_B2;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X0Y109_B3;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X0Y109_B4;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X0Y109_B5;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X0Y109_B6;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X0Y109_BO5;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X0Y109_BO6;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X0Y109_B_CY;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X0Y109_B_XOR;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X0Y109_C;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X0Y109_C1;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X0Y109_C2;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X0Y109_C3;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X0Y109_C4;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X0Y109_C5;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X0Y109_C6;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X0Y109_CO5;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X0Y109_CO6;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X0Y109_C_CY;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X0Y109_C_XOR;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X0Y109_D;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X0Y109_D1;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X0Y109_D2;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X0Y109_D3;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X0Y109_D4;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X0Y109_D5;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X0Y109_D6;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X0Y109_DO5;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X0Y109_DO6;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X0Y109_D_CY;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X0Y109_D_XOR;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X1Y109_A;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X1Y109_A1;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X1Y109_A2;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X1Y109_A3;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X1Y109_A4;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X1Y109_A5;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X1Y109_A6;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X1Y109_AO5;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X1Y109_AO6;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X1Y109_A_CY;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X1Y109_A_XOR;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X1Y109_B;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X1Y109_B1;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X1Y109_B2;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X1Y109_B3;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X1Y109_B4;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X1Y109_B5;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X1Y109_B6;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X1Y109_BO5;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X1Y109_BO6;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X1Y109_B_CY;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X1Y109_B_XOR;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X1Y109_C;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X1Y109_C1;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X1Y109_C2;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X1Y109_C3;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X1Y109_C4;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X1Y109_C5;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X1Y109_C6;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X1Y109_CO5;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X1Y109_CO6;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X1Y109_C_CY;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X1Y109_C_XOR;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X1Y109_D;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X1Y109_D1;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X1Y109_D2;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X1Y109_D3;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X1Y109_D4;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X1Y109_D5;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X1Y109_D6;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X1Y109_DO5;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X1Y109_DO6;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X1Y109_D_CY;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X1Y109_D_XOR;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X0Y110_A;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X0Y110_A1;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X0Y110_A2;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X0Y110_A3;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X0Y110_A4;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X0Y110_A5;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X0Y110_A6;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X0Y110_AMUX;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X0Y110_AO5;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X0Y110_AO6;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X0Y110_A_CY;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X0Y110_A_XOR;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X0Y110_B;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X0Y110_B1;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X0Y110_B2;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X0Y110_B3;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X0Y110_B4;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X0Y110_B5;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X0Y110_B6;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X0Y110_BO5;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X0Y110_BO6;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X0Y110_B_CY;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X0Y110_B_XOR;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X0Y110_C;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X0Y110_C1;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X0Y110_C2;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X0Y110_C3;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X0Y110_C4;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X0Y110_C5;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X0Y110_C6;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X0Y110_CO5;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X0Y110_CO6;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X0Y110_C_CY;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X0Y110_C_XOR;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X0Y110_D;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X0Y110_D1;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X0Y110_D2;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X0Y110_D3;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X0Y110_D4;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X0Y110_D5;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X0Y110_D6;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X0Y110_DO5;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X0Y110_DO6;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X0Y110_D_CY;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X0Y110_D_XOR;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X1Y110_A;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X1Y110_A1;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X1Y110_A2;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X1Y110_A3;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X1Y110_A4;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X1Y110_A5;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X1Y110_A6;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X1Y110_AO5;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X1Y110_AO6;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X1Y110_A_CY;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X1Y110_A_XOR;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X1Y110_B;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X1Y110_B1;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X1Y110_B2;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X1Y110_B3;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X1Y110_B4;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X1Y110_B5;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X1Y110_B6;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X1Y110_BO5;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X1Y110_BO6;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X1Y110_B_CY;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X1Y110_B_XOR;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X1Y110_C;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X1Y110_C1;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X1Y110_C2;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X1Y110_C3;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X1Y110_C4;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X1Y110_C5;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X1Y110_C6;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X1Y110_CO5;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X1Y110_CO6;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X1Y110_C_CY;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X1Y110_C_XOR;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X1Y110_D;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X1Y110_D1;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X1Y110_D2;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X1Y110_D3;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X1Y110_D4;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X1Y110_D5;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X1Y110_D6;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X1Y110_DO5;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X1Y110_DO6;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X1Y110_D_CY;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X1Y110_D_XOR;
  wire [0:0] CLBLL_L_X4Y103_SLICE_X4Y103_A;
  wire [0:0] CLBLL_L_X4Y103_SLICE_X4Y103_A1;
  wire [0:0] CLBLL_L_X4Y103_SLICE_X4Y103_A2;
  wire [0:0] CLBLL_L_X4Y103_SLICE_X4Y103_A3;
  wire [0:0] CLBLL_L_X4Y103_SLICE_X4Y103_A4;
  wire [0:0] CLBLL_L_X4Y103_SLICE_X4Y103_A5;
  wire [0:0] CLBLL_L_X4Y103_SLICE_X4Y103_A6;
  wire [0:0] CLBLL_L_X4Y103_SLICE_X4Y103_AMUX;
  wire [0:0] CLBLL_L_X4Y103_SLICE_X4Y103_AO5;
  wire [0:0] CLBLL_L_X4Y103_SLICE_X4Y103_AO6;
  wire [0:0] CLBLL_L_X4Y103_SLICE_X4Y103_A_CY;
  wire [0:0] CLBLL_L_X4Y103_SLICE_X4Y103_A_XOR;
  wire [0:0] CLBLL_L_X4Y103_SLICE_X4Y103_B;
  wire [0:0] CLBLL_L_X4Y103_SLICE_X4Y103_B1;
  wire [0:0] CLBLL_L_X4Y103_SLICE_X4Y103_B2;
  wire [0:0] CLBLL_L_X4Y103_SLICE_X4Y103_B3;
  wire [0:0] CLBLL_L_X4Y103_SLICE_X4Y103_B4;
  wire [0:0] CLBLL_L_X4Y103_SLICE_X4Y103_B5;
  wire [0:0] CLBLL_L_X4Y103_SLICE_X4Y103_B6;
  wire [0:0] CLBLL_L_X4Y103_SLICE_X4Y103_BO5;
  wire [0:0] CLBLL_L_X4Y103_SLICE_X4Y103_BO6;
  wire [0:0] CLBLL_L_X4Y103_SLICE_X4Y103_B_CY;
  wire [0:0] CLBLL_L_X4Y103_SLICE_X4Y103_B_XOR;
  wire [0:0] CLBLL_L_X4Y103_SLICE_X4Y103_C;
  wire [0:0] CLBLL_L_X4Y103_SLICE_X4Y103_C1;
  wire [0:0] CLBLL_L_X4Y103_SLICE_X4Y103_C2;
  wire [0:0] CLBLL_L_X4Y103_SLICE_X4Y103_C3;
  wire [0:0] CLBLL_L_X4Y103_SLICE_X4Y103_C4;
  wire [0:0] CLBLL_L_X4Y103_SLICE_X4Y103_C5;
  wire [0:0] CLBLL_L_X4Y103_SLICE_X4Y103_C6;
  wire [0:0] CLBLL_L_X4Y103_SLICE_X4Y103_CO5;
  wire [0:0] CLBLL_L_X4Y103_SLICE_X4Y103_CO6;
  wire [0:0] CLBLL_L_X4Y103_SLICE_X4Y103_C_CY;
  wire [0:0] CLBLL_L_X4Y103_SLICE_X4Y103_C_XOR;
  wire [0:0] CLBLL_L_X4Y103_SLICE_X4Y103_D;
  wire [0:0] CLBLL_L_X4Y103_SLICE_X4Y103_D1;
  wire [0:0] CLBLL_L_X4Y103_SLICE_X4Y103_D2;
  wire [0:0] CLBLL_L_X4Y103_SLICE_X4Y103_D3;
  wire [0:0] CLBLL_L_X4Y103_SLICE_X4Y103_D4;
  wire [0:0] CLBLL_L_X4Y103_SLICE_X4Y103_D5;
  wire [0:0] CLBLL_L_X4Y103_SLICE_X4Y103_D6;
  wire [0:0] CLBLL_L_X4Y103_SLICE_X4Y103_DO5;
  wire [0:0] CLBLL_L_X4Y103_SLICE_X4Y103_DO6;
  wire [0:0] CLBLL_L_X4Y103_SLICE_X4Y103_D_CY;
  wire [0:0] CLBLL_L_X4Y103_SLICE_X4Y103_D_XOR;
  wire [0:0] CLBLL_L_X4Y103_SLICE_X5Y103_A;
  wire [0:0] CLBLL_L_X4Y103_SLICE_X5Y103_A1;
  wire [0:0] CLBLL_L_X4Y103_SLICE_X5Y103_A2;
  wire [0:0] CLBLL_L_X4Y103_SLICE_X5Y103_A3;
  wire [0:0] CLBLL_L_X4Y103_SLICE_X5Y103_A4;
  wire [0:0] CLBLL_L_X4Y103_SLICE_X5Y103_A5;
  wire [0:0] CLBLL_L_X4Y103_SLICE_X5Y103_A6;
  wire [0:0] CLBLL_L_X4Y103_SLICE_X5Y103_AMUX;
  wire [0:0] CLBLL_L_X4Y103_SLICE_X5Y103_AO5;
  wire [0:0] CLBLL_L_X4Y103_SLICE_X5Y103_AO6;
  wire [0:0] CLBLL_L_X4Y103_SLICE_X5Y103_A_CY;
  wire [0:0] CLBLL_L_X4Y103_SLICE_X5Y103_A_XOR;
  wire [0:0] CLBLL_L_X4Y103_SLICE_X5Y103_B;
  wire [0:0] CLBLL_L_X4Y103_SLICE_X5Y103_B1;
  wire [0:0] CLBLL_L_X4Y103_SLICE_X5Y103_B2;
  wire [0:0] CLBLL_L_X4Y103_SLICE_X5Y103_B3;
  wire [0:0] CLBLL_L_X4Y103_SLICE_X5Y103_B4;
  wire [0:0] CLBLL_L_X4Y103_SLICE_X5Y103_B5;
  wire [0:0] CLBLL_L_X4Y103_SLICE_X5Y103_B6;
  wire [0:0] CLBLL_L_X4Y103_SLICE_X5Y103_BO5;
  wire [0:0] CLBLL_L_X4Y103_SLICE_X5Y103_BO6;
  wire [0:0] CLBLL_L_X4Y103_SLICE_X5Y103_B_CY;
  wire [0:0] CLBLL_L_X4Y103_SLICE_X5Y103_B_XOR;
  wire [0:0] CLBLL_L_X4Y103_SLICE_X5Y103_C;
  wire [0:0] CLBLL_L_X4Y103_SLICE_X5Y103_C1;
  wire [0:0] CLBLL_L_X4Y103_SLICE_X5Y103_C2;
  wire [0:0] CLBLL_L_X4Y103_SLICE_X5Y103_C3;
  wire [0:0] CLBLL_L_X4Y103_SLICE_X5Y103_C4;
  wire [0:0] CLBLL_L_X4Y103_SLICE_X5Y103_C5;
  wire [0:0] CLBLL_L_X4Y103_SLICE_X5Y103_C6;
  wire [0:0] CLBLL_L_X4Y103_SLICE_X5Y103_CO5;
  wire [0:0] CLBLL_L_X4Y103_SLICE_X5Y103_CO6;
  wire [0:0] CLBLL_L_X4Y103_SLICE_X5Y103_C_CY;
  wire [0:0] CLBLL_L_X4Y103_SLICE_X5Y103_C_XOR;
  wire [0:0] CLBLL_L_X4Y103_SLICE_X5Y103_D;
  wire [0:0] CLBLL_L_X4Y103_SLICE_X5Y103_D1;
  wire [0:0] CLBLL_L_X4Y103_SLICE_X5Y103_D2;
  wire [0:0] CLBLL_L_X4Y103_SLICE_X5Y103_D3;
  wire [0:0] CLBLL_L_X4Y103_SLICE_X5Y103_D4;
  wire [0:0] CLBLL_L_X4Y103_SLICE_X5Y103_D5;
  wire [0:0] CLBLL_L_X4Y103_SLICE_X5Y103_D6;
  wire [0:0] CLBLL_L_X4Y103_SLICE_X5Y103_DO5;
  wire [0:0] CLBLL_L_X4Y103_SLICE_X5Y103_DO6;
  wire [0:0] CLBLL_L_X4Y103_SLICE_X5Y103_D_CY;
  wire [0:0] CLBLL_L_X4Y103_SLICE_X5Y103_D_XOR;
  wire [0:0] CLBLL_L_X4Y104_SLICE_X4Y104_A;
  wire [0:0] CLBLL_L_X4Y104_SLICE_X4Y104_A1;
  wire [0:0] CLBLL_L_X4Y104_SLICE_X4Y104_A2;
  wire [0:0] CLBLL_L_X4Y104_SLICE_X4Y104_A3;
  wire [0:0] CLBLL_L_X4Y104_SLICE_X4Y104_A4;
  wire [0:0] CLBLL_L_X4Y104_SLICE_X4Y104_A5;
  wire [0:0] CLBLL_L_X4Y104_SLICE_X4Y104_A6;
  wire [0:0] CLBLL_L_X4Y104_SLICE_X4Y104_AO5;
  wire [0:0] CLBLL_L_X4Y104_SLICE_X4Y104_AO6;
  wire [0:0] CLBLL_L_X4Y104_SLICE_X4Y104_A_CY;
  wire [0:0] CLBLL_L_X4Y104_SLICE_X4Y104_A_XOR;
  wire [0:0] CLBLL_L_X4Y104_SLICE_X4Y104_B;
  wire [0:0] CLBLL_L_X4Y104_SLICE_X4Y104_B1;
  wire [0:0] CLBLL_L_X4Y104_SLICE_X4Y104_B2;
  wire [0:0] CLBLL_L_X4Y104_SLICE_X4Y104_B3;
  wire [0:0] CLBLL_L_X4Y104_SLICE_X4Y104_B4;
  wire [0:0] CLBLL_L_X4Y104_SLICE_X4Y104_B5;
  wire [0:0] CLBLL_L_X4Y104_SLICE_X4Y104_B6;
  wire [0:0] CLBLL_L_X4Y104_SLICE_X4Y104_BO5;
  wire [0:0] CLBLL_L_X4Y104_SLICE_X4Y104_BO6;
  wire [0:0] CLBLL_L_X4Y104_SLICE_X4Y104_B_CY;
  wire [0:0] CLBLL_L_X4Y104_SLICE_X4Y104_B_XOR;
  wire [0:0] CLBLL_L_X4Y104_SLICE_X4Y104_C;
  wire [0:0] CLBLL_L_X4Y104_SLICE_X4Y104_C1;
  wire [0:0] CLBLL_L_X4Y104_SLICE_X4Y104_C2;
  wire [0:0] CLBLL_L_X4Y104_SLICE_X4Y104_C3;
  wire [0:0] CLBLL_L_X4Y104_SLICE_X4Y104_C4;
  wire [0:0] CLBLL_L_X4Y104_SLICE_X4Y104_C5;
  wire [0:0] CLBLL_L_X4Y104_SLICE_X4Y104_C6;
  wire [0:0] CLBLL_L_X4Y104_SLICE_X4Y104_CO5;
  wire [0:0] CLBLL_L_X4Y104_SLICE_X4Y104_CO6;
  wire [0:0] CLBLL_L_X4Y104_SLICE_X4Y104_C_CY;
  wire [0:0] CLBLL_L_X4Y104_SLICE_X4Y104_C_XOR;
  wire [0:0] CLBLL_L_X4Y104_SLICE_X4Y104_D;
  wire [0:0] CLBLL_L_X4Y104_SLICE_X4Y104_D1;
  wire [0:0] CLBLL_L_X4Y104_SLICE_X4Y104_D2;
  wire [0:0] CLBLL_L_X4Y104_SLICE_X4Y104_D3;
  wire [0:0] CLBLL_L_X4Y104_SLICE_X4Y104_D4;
  wire [0:0] CLBLL_L_X4Y104_SLICE_X4Y104_D5;
  wire [0:0] CLBLL_L_X4Y104_SLICE_X4Y104_D6;
  wire [0:0] CLBLL_L_X4Y104_SLICE_X4Y104_DO5;
  wire [0:0] CLBLL_L_X4Y104_SLICE_X4Y104_DO6;
  wire [0:0] CLBLL_L_X4Y104_SLICE_X4Y104_D_CY;
  wire [0:0] CLBLL_L_X4Y104_SLICE_X4Y104_D_XOR;
  wire [0:0] CLBLL_L_X4Y104_SLICE_X5Y104_A;
  wire [0:0] CLBLL_L_X4Y104_SLICE_X5Y104_A1;
  wire [0:0] CLBLL_L_X4Y104_SLICE_X5Y104_A2;
  wire [0:0] CLBLL_L_X4Y104_SLICE_X5Y104_A3;
  wire [0:0] CLBLL_L_X4Y104_SLICE_X5Y104_A4;
  wire [0:0] CLBLL_L_X4Y104_SLICE_X5Y104_A5;
  wire [0:0] CLBLL_L_X4Y104_SLICE_X5Y104_A6;
  wire [0:0] CLBLL_L_X4Y104_SLICE_X5Y104_AMUX;
  wire [0:0] CLBLL_L_X4Y104_SLICE_X5Y104_AO5;
  wire [0:0] CLBLL_L_X4Y104_SLICE_X5Y104_AO6;
  wire [0:0] CLBLL_L_X4Y104_SLICE_X5Y104_A_CY;
  wire [0:0] CLBLL_L_X4Y104_SLICE_X5Y104_A_XOR;
  wire [0:0] CLBLL_L_X4Y104_SLICE_X5Y104_B;
  wire [0:0] CLBLL_L_X4Y104_SLICE_X5Y104_B1;
  wire [0:0] CLBLL_L_X4Y104_SLICE_X5Y104_B2;
  wire [0:0] CLBLL_L_X4Y104_SLICE_X5Y104_B3;
  wire [0:0] CLBLL_L_X4Y104_SLICE_X5Y104_B4;
  wire [0:0] CLBLL_L_X4Y104_SLICE_X5Y104_B5;
  wire [0:0] CLBLL_L_X4Y104_SLICE_X5Y104_B6;
  wire [0:0] CLBLL_L_X4Y104_SLICE_X5Y104_BO5;
  wire [0:0] CLBLL_L_X4Y104_SLICE_X5Y104_BO6;
  wire [0:0] CLBLL_L_X4Y104_SLICE_X5Y104_B_CY;
  wire [0:0] CLBLL_L_X4Y104_SLICE_X5Y104_B_XOR;
  wire [0:0] CLBLL_L_X4Y104_SLICE_X5Y104_C;
  wire [0:0] CLBLL_L_X4Y104_SLICE_X5Y104_C1;
  wire [0:0] CLBLL_L_X4Y104_SLICE_X5Y104_C2;
  wire [0:0] CLBLL_L_X4Y104_SLICE_X5Y104_C3;
  wire [0:0] CLBLL_L_X4Y104_SLICE_X5Y104_C4;
  wire [0:0] CLBLL_L_X4Y104_SLICE_X5Y104_C5;
  wire [0:0] CLBLL_L_X4Y104_SLICE_X5Y104_C6;
  wire [0:0] CLBLL_L_X4Y104_SLICE_X5Y104_CO5;
  wire [0:0] CLBLL_L_X4Y104_SLICE_X5Y104_CO6;
  wire [0:0] CLBLL_L_X4Y104_SLICE_X5Y104_C_CY;
  wire [0:0] CLBLL_L_X4Y104_SLICE_X5Y104_C_XOR;
  wire [0:0] CLBLL_L_X4Y104_SLICE_X5Y104_D;
  wire [0:0] CLBLL_L_X4Y104_SLICE_X5Y104_D1;
  wire [0:0] CLBLL_L_X4Y104_SLICE_X5Y104_D2;
  wire [0:0] CLBLL_L_X4Y104_SLICE_X5Y104_D3;
  wire [0:0] CLBLL_L_X4Y104_SLICE_X5Y104_D4;
  wire [0:0] CLBLL_L_X4Y104_SLICE_X5Y104_D5;
  wire [0:0] CLBLL_L_X4Y104_SLICE_X5Y104_D6;
  wire [0:0] CLBLL_L_X4Y104_SLICE_X5Y104_DO5;
  wire [0:0] CLBLL_L_X4Y104_SLICE_X5Y104_DO6;
  wire [0:0] CLBLL_L_X4Y104_SLICE_X5Y104_D_CY;
  wire [0:0] CLBLL_L_X4Y104_SLICE_X5Y104_D_XOR;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X4Y105_A;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X4Y105_A1;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X4Y105_A2;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X4Y105_A3;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X4Y105_A4;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X4Y105_A5;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X4Y105_A6;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X4Y105_AMUX;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X4Y105_AO5;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X4Y105_AO6;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X4Y105_A_CY;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X4Y105_A_XOR;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X4Y105_B;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X4Y105_B1;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X4Y105_B2;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X4Y105_B3;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X4Y105_B4;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X4Y105_B5;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X4Y105_B6;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X4Y105_BO5;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X4Y105_BO6;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X4Y105_B_CY;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X4Y105_B_XOR;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X4Y105_C;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X4Y105_C1;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X4Y105_C2;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X4Y105_C3;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X4Y105_C4;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X4Y105_C5;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X4Y105_C6;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X4Y105_CO5;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X4Y105_CO6;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X4Y105_C_CY;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X4Y105_C_XOR;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X4Y105_D;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X4Y105_D1;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X4Y105_D2;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X4Y105_D3;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X4Y105_D4;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X4Y105_D5;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X4Y105_D6;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X4Y105_DO5;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X4Y105_DO6;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X4Y105_D_CY;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X4Y105_D_XOR;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X5Y105_A;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X5Y105_A1;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X5Y105_A2;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X5Y105_A3;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X5Y105_A4;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X5Y105_A5;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X5Y105_A6;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X5Y105_AO5;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X5Y105_AO6;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X5Y105_A_CY;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X5Y105_A_XOR;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X5Y105_B;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X5Y105_B1;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X5Y105_B2;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X5Y105_B3;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X5Y105_B4;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X5Y105_B5;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X5Y105_B6;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X5Y105_BO5;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X5Y105_BO6;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X5Y105_B_CY;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X5Y105_B_XOR;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X5Y105_C;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X5Y105_C1;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X5Y105_C2;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X5Y105_C3;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X5Y105_C4;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X5Y105_C5;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X5Y105_C6;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X5Y105_CO5;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X5Y105_CO6;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X5Y105_C_CY;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X5Y105_C_XOR;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X5Y105_D;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X5Y105_D1;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X5Y105_D2;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X5Y105_D3;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X5Y105_D4;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X5Y105_D5;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X5Y105_D6;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X5Y105_DO5;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X5Y105_DO6;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X5Y105_D_CY;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X5Y105_D_XOR;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X4Y106_A;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X4Y106_A1;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X4Y106_A2;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X4Y106_A3;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X4Y106_A4;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X4Y106_A5;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X4Y106_A6;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X4Y106_AO5;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X4Y106_AO6;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X4Y106_A_CY;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X4Y106_A_XOR;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X4Y106_B;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X4Y106_B1;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X4Y106_B2;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X4Y106_B3;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X4Y106_B4;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X4Y106_B5;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X4Y106_B6;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X4Y106_BO5;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X4Y106_BO6;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X4Y106_B_CY;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X4Y106_B_XOR;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X4Y106_C;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X4Y106_C1;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X4Y106_C2;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X4Y106_C3;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X4Y106_C4;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X4Y106_C5;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X4Y106_C6;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X4Y106_CO5;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X4Y106_CO6;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X4Y106_C_CY;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X4Y106_C_XOR;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X4Y106_D;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X4Y106_D1;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X4Y106_D2;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X4Y106_D3;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X4Y106_D4;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X4Y106_D5;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X4Y106_D6;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X4Y106_DO5;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X4Y106_DO6;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X4Y106_D_CY;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X4Y106_D_XOR;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X5Y106_A;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X5Y106_A1;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X5Y106_A2;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X5Y106_A3;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X5Y106_A4;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X5Y106_A5;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X5Y106_A6;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X5Y106_AO5;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X5Y106_AO6;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X5Y106_A_CY;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X5Y106_A_XOR;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X5Y106_B;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X5Y106_B1;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X5Y106_B2;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X5Y106_B3;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X5Y106_B4;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X5Y106_B5;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X5Y106_B6;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X5Y106_BO5;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X5Y106_BO6;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X5Y106_B_CY;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X5Y106_B_XOR;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X5Y106_C;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X5Y106_C1;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X5Y106_C2;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X5Y106_C3;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X5Y106_C4;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X5Y106_C5;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X5Y106_C6;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X5Y106_CO5;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X5Y106_CO6;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X5Y106_C_CY;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X5Y106_C_XOR;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X5Y106_D;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X5Y106_D1;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X5Y106_D2;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X5Y106_D3;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X5Y106_D4;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X5Y106_D5;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X5Y106_D6;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X5Y106_DO5;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X5Y106_DO6;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X5Y106_D_CY;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X5Y106_D_XOR;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X4Y107_A;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X4Y107_A1;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X4Y107_A2;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X4Y107_A3;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X4Y107_A4;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X4Y107_A5;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X4Y107_A6;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X4Y107_AO5;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X4Y107_AO6;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X4Y107_A_CY;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X4Y107_A_XOR;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X4Y107_B;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X4Y107_B1;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X4Y107_B2;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X4Y107_B3;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X4Y107_B4;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X4Y107_B5;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X4Y107_B6;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X4Y107_BO5;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X4Y107_BO6;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X4Y107_B_CY;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X4Y107_B_XOR;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X4Y107_C;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X4Y107_C1;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X4Y107_C2;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X4Y107_C3;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X4Y107_C4;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X4Y107_C5;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X4Y107_C6;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X4Y107_CO5;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X4Y107_CO6;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X4Y107_C_CY;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X4Y107_C_XOR;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X4Y107_D;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X4Y107_D1;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X4Y107_D2;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X4Y107_D3;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X4Y107_D4;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X4Y107_D5;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X4Y107_D6;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X4Y107_DO5;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X4Y107_DO6;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X4Y107_D_CY;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X4Y107_D_XOR;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X5Y107_A;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X5Y107_A1;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X5Y107_A2;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X5Y107_A3;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X5Y107_A4;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X5Y107_A5;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X5Y107_A6;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X5Y107_AMUX;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X5Y107_AO5;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X5Y107_AO6;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X5Y107_A_CY;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X5Y107_A_XOR;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X5Y107_B;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X5Y107_B1;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X5Y107_B2;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X5Y107_B3;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X5Y107_B4;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X5Y107_B5;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X5Y107_B6;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X5Y107_BO5;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X5Y107_BO6;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X5Y107_B_CY;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X5Y107_B_XOR;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X5Y107_C;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X5Y107_C1;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X5Y107_C2;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X5Y107_C3;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X5Y107_C4;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X5Y107_C5;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X5Y107_C6;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X5Y107_CMUX;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X5Y107_CO5;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X5Y107_CO6;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X5Y107_C_CY;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X5Y107_C_XOR;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X5Y107_D;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X5Y107_D1;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X5Y107_D2;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X5Y107_D3;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X5Y107_D4;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X5Y107_D5;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X5Y107_D6;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X5Y107_DO5;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X5Y107_DO6;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X5Y107_D_CY;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X5Y107_D_XOR;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X4Y108_A;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X4Y108_A1;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X4Y108_A2;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X4Y108_A3;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X4Y108_A4;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X4Y108_A5;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X4Y108_A6;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X4Y108_AMUX;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X4Y108_AO5;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X4Y108_AO6;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X4Y108_A_CY;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X4Y108_A_XOR;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X4Y108_B;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X4Y108_B1;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X4Y108_B2;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X4Y108_B3;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X4Y108_B4;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X4Y108_B5;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X4Y108_B6;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X4Y108_BO5;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X4Y108_BO6;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X4Y108_B_CY;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X4Y108_B_XOR;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X4Y108_C;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X4Y108_C1;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X4Y108_C2;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X4Y108_C3;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X4Y108_C4;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X4Y108_C5;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X4Y108_C6;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X4Y108_CO5;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X4Y108_CO6;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X4Y108_C_CY;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X4Y108_C_XOR;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X4Y108_D;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X4Y108_D1;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X4Y108_D2;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X4Y108_D3;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X4Y108_D4;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X4Y108_D5;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X4Y108_D6;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X4Y108_DO5;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X4Y108_DO6;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X4Y108_D_CY;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X4Y108_D_XOR;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X5Y108_A;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X5Y108_A1;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X5Y108_A2;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X5Y108_A3;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X5Y108_A4;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X5Y108_A5;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X5Y108_A6;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X5Y108_AO5;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X5Y108_AO6;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X5Y108_A_CY;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X5Y108_A_XOR;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X5Y108_B;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X5Y108_B1;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X5Y108_B2;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X5Y108_B3;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X5Y108_B4;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X5Y108_B5;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X5Y108_B6;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X5Y108_BO5;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X5Y108_BO6;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X5Y108_B_CY;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X5Y108_B_XOR;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X5Y108_C;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X5Y108_C1;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X5Y108_C2;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X5Y108_C3;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X5Y108_C4;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X5Y108_C5;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X5Y108_C6;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X5Y108_CO5;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X5Y108_CO6;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X5Y108_C_CY;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X5Y108_C_XOR;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X5Y108_D;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X5Y108_D1;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X5Y108_D2;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X5Y108_D3;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X5Y108_D4;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X5Y108_D5;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X5Y108_D6;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X5Y108_DO5;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X5Y108_DO6;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X5Y108_D_CY;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X5Y108_D_XOR;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X4Y109_A;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X4Y109_A1;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X4Y109_A2;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X4Y109_A3;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X4Y109_A4;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X4Y109_A5;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X4Y109_A6;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X4Y109_AMUX;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X4Y109_AO5;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X4Y109_AO6;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X4Y109_A_CY;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X4Y109_A_XOR;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X4Y109_B;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X4Y109_B1;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X4Y109_B2;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X4Y109_B3;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X4Y109_B4;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X4Y109_B5;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X4Y109_B6;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X4Y109_BO5;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X4Y109_BO6;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X4Y109_B_CY;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X4Y109_B_XOR;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X4Y109_C;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X4Y109_C1;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X4Y109_C2;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X4Y109_C3;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X4Y109_C4;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X4Y109_C5;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X4Y109_C6;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X4Y109_CO5;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X4Y109_CO6;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X4Y109_C_CY;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X4Y109_C_XOR;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X4Y109_D;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X4Y109_D1;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X4Y109_D2;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X4Y109_D3;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X4Y109_D4;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X4Y109_D5;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X4Y109_D6;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X4Y109_DO5;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X4Y109_DO6;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X4Y109_D_CY;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X4Y109_D_XOR;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X5Y109_A;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X5Y109_A1;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X5Y109_A2;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X5Y109_A3;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X5Y109_A4;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X5Y109_A5;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X5Y109_A6;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X5Y109_AMUX;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X5Y109_AO5;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X5Y109_AO6;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X5Y109_A_CY;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X5Y109_A_XOR;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X5Y109_B;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X5Y109_B1;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X5Y109_B2;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X5Y109_B3;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X5Y109_B4;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X5Y109_B5;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X5Y109_B6;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X5Y109_BO5;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X5Y109_BO6;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X5Y109_B_CY;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X5Y109_B_XOR;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X5Y109_C;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X5Y109_C1;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X5Y109_C2;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X5Y109_C3;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X5Y109_C4;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X5Y109_C5;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X5Y109_C6;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X5Y109_CO5;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X5Y109_CO6;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X5Y109_C_CY;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X5Y109_C_XOR;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X5Y109_D;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X5Y109_D1;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X5Y109_D2;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X5Y109_D3;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X5Y109_D4;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X5Y109_D5;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X5Y109_D6;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X5Y109_DO5;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X5Y109_DO6;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X5Y109_D_CY;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X5Y109_D_XOR;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X4Y110_A;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X4Y110_A1;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X4Y110_A2;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X4Y110_A3;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X4Y110_A4;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X4Y110_A5;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X4Y110_A6;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X4Y110_AO5;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X4Y110_AO6;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X4Y110_A_CY;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X4Y110_A_XOR;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X4Y110_B;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X4Y110_B1;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X4Y110_B2;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X4Y110_B3;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X4Y110_B4;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X4Y110_B5;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X4Y110_B6;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X4Y110_BO5;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X4Y110_BO6;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X4Y110_B_CY;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X4Y110_B_XOR;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X4Y110_C;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X4Y110_C1;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X4Y110_C2;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X4Y110_C3;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X4Y110_C4;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X4Y110_C5;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X4Y110_C6;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X4Y110_CO5;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X4Y110_CO6;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X4Y110_C_CY;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X4Y110_C_XOR;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X4Y110_D;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X4Y110_D1;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X4Y110_D2;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X4Y110_D3;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X4Y110_D4;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X4Y110_D5;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X4Y110_D6;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X4Y110_DO5;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X4Y110_DO6;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X4Y110_D_CY;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X4Y110_D_XOR;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X5Y110_A;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X5Y110_A1;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X5Y110_A2;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X5Y110_A3;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X5Y110_A4;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X5Y110_A5;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X5Y110_A6;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X5Y110_AMUX;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X5Y110_AO5;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X5Y110_AO6;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X5Y110_A_CY;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X5Y110_A_XOR;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X5Y110_B;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X5Y110_B1;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X5Y110_B2;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X5Y110_B3;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X5Y110_B4;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X5Y110_B5;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X5Y110_B6;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X5Y110_BMUX;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X5Y110_BO5;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X5Y110_BO6;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X5Y110_B_CY;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X5Y110_B_XOR;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X5Y110_C;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X5Y110_C1;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X5Y110_C2;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X5Y110_C3;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X5Y110_C4;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X5Y110_C5;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X5Y110_C6;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X5Y110_CO5;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X5Y110_CO6;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X5Y110_C_CY;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X5Y110_C_XOR;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X5Y110_D;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X5Y110_D1;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X5Y110_D2;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X5Y110_D3;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X5Y110_D4;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X5Y110_D5;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X5Y110_D6;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X5Y110_DO5;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X5Y110_DO6;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X5Y110_D_CY;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X5Y110_D_XOR;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X4Y111_A;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X4Y111_A1;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X4Y111_A2;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X4Y111_A3;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X4Y111_A4;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X4Y111_A5;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X4Y111_A6;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X4Y111_AMUX;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X4Y111_AO5;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X4Y111_AO6;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X4Y111_A_CY;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X4Y111_A_XOR;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X4Y111_B;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X4Y111_B1;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X4Y111_B2;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X4Y111_B3;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X4Y111_B4;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X4Y111_B5;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X4Y111_B6;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X4Y111_BMUX;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X4Y111_BO5;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X4Y111_BO6;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X4Y111_B_CY;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X4Y111_B_XOR;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X4Y111_C;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X4Y111_C1;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X4Y111_C2;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X4Y111_C3;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X4Y111_C4;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X4Y111_C5;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X4Y111_C6;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X4Y111_CMUX;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X4Y111_CO5;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X4Y111_CO6;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X4Y111_C_CY;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X4Y111_C_XOR;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X4Y111_D;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X4Y111_D1;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X4Y111_D2;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X4Y111_D3;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X4Y111_D4;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X4Y111_D5;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X4Y111_D6;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X4Y111_DMUX;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X4Y111_DO5;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X4Y111_DO6;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X4Y111_D_CY;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X4Y111_D_XOR;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X5Y111_A;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X5Y111_A1;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X5Y111_A2;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X5Y111_A3;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X5Y111_A4;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X5Y111_A5;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X5Y111_A6;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X5Y111_AMUX;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X5Y111_AO5;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X5Y111_AO6;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X5Y111_A_CY;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X5Y111_A_XOR;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X5Y111_B;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X5Y111_B1;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X5Y111_B2;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X5Y111_B3;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X5Y111_B4;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X5Y111_B5;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X5Y111_B6;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X5Y111_BO5;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X5Y111_BO6;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X5Y111_B_CY;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X5Y111_B_XOR;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X5Y111_C;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X5Y111_C1;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X5Y111_C2;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X5Y111_C3;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X5Y111_C4;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X5Y111_C5;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X5Y111_C6;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X5Y111_CO5;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X5Y111_CO6;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X5Y111_C_CY;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X5Y111_C_XOR;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X5Y111_D;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X5Y111_D1;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X5Y111_D2;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X5Y111_D3;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X5Y111_D4;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X5Y111_D5;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X5Y111_D6;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X5Y111_DO5;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X5Y111_DO6;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X5Y111_D_CY;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X5Y111_D_XOR;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X4Y112_A;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X4Y112_A1;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X4Y112_A2;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X4Y112_A3;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X4Y112_A4;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X4Y112_A5;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X4Y112_A6;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X4Y112_AMUX;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X4Y112_AO5;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X4Y112_AO6;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X4Y112_A_CY;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X4Y112_A_XOR;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X4Y112_B;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X4Y112_B1;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X4Y112_B2;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X4Y112_B3;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X4Y112_B4;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X4Y112_B5;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X4Y112_B6;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X4Y112_BO5;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X4Y112_BO6;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X4Y112_B_CY;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X4Y112_B_XOR;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X4Y112_C;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X4Y112_C1;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X4Y112_C2;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X4Y112_C3;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X4Y112_C4;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X4Y112_C5;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X4Y112_C6;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X4Y112_CO5;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X4Y112_CO6;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X4Y112_C_CY;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X4Y112_C_XOR;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X4Y112_D;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X4Y112_D1;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X4Y112_D2;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X4Y112_D3;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X4Y112_D4;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X4Y112_D5;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X4Y112_D6;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X4Y112_DO5;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X4Y112_DO6;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X4Y112_D_CY;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X4Y112_D_XOR;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X5Y112_A;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X5Y112_A1;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X5Y112_A2;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X5Y112_A3;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X5Y112_A4;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X5Y112_A5;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X5Y112_A6;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X5Y112_AO5;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X5Y112_AO6;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X5Y112_A_CY;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X5Y112_A_XOR;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X5Y112_B;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X5Y112_B1;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X5Y112_B2;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X5Y112_B3;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X5Y112_B4;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X5Y112_B5;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X5Y112_B6;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X5Y112_BO5;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X5Y112_BO6;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X5Y112_B_CY;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X5Y112_B_XOR;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X5Y112_C;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X5Y112_C1;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X5Y112_C2;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X5Y112_C3;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X5Y112_C4;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X5Y112_C5;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X5Y112_C6;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X5Y112_CMUX;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X5Y112_CO5;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X5Y112_CO6;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X5Y112_C_CY;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X5Y112_C_XOR;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X5Y112_D;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X5Y112_D1;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X5Y112_D2;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X5Y112_D3;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X5Y112_D4;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X5Y112_D5;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X5Y112_D6;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X5Y112_DO5;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X5Y112_DO6;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X5Y112_D_CY;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X5Y112_D_XOR;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_A;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_A1;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_A2;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_A3;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_A4;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_A5;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_A6;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_AMUX;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_AO5;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_AO6;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_A_CY;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_A_XOR;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_B;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_B1;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_B2;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_B3;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_B4;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_B5;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_B6;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_BO5;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_BO6;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_B_CY;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_B_XOR;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_C;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_C1;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_C2;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_C3;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_C4;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_C5;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_C6;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_CO5;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_CO6;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_C_CY;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_C_XOR;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_D;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_D1;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_D2;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_D3;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_D4;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_D5;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_D6;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_DO5;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_DO6;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_D_CY;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_D_XOR;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_A;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_A1;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_A2;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_A3;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_A4;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_A5;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_A6;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_AMUX;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_AO5;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_AO6;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_A_CY;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_A_XOR;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_B;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_B1;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_B2;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_B3;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_B4;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_B5;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_B6;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_BO5;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_BO6;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_B_CY;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_B_XOR;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_C;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_C1;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_C2;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_C3;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_C4;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_C5;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_C6;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_CO5;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_CO6;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_C_CY;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_C_XOR;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_D;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_D1;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_D2;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_D3;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_D4;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_D5;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_D6;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_DO5;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_DO6;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_D_CY;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_D_XOR;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X4Y114_A;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X4Y114_A1;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X4Y114_A2;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X4Y114_A3;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X4Y114_A4;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X4Y114_A5;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X4Y114_A6;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X4Y114_AMUX;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X4Y114_AO5;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X4Y114_AO6;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X4Y114_A_CY;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X4Y114_A_XOR;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X4Y114_B;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X4Y114_B1;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X4Y114_B2;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X4Y114_B3;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X4Y114_B4;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X4Y114_B5;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X4Y114_B6;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X4Y114_BMUX;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X4Y114_BO5;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X4Y114_BO6;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X4Y114_B_CY;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X4Y114_B_XOR;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X4Y114_C;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X4Y114_C1;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X4Y114_C2;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X4Y114_C3;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X4Y114_C4;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X4Y114_C5;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X4Y114_C6;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X4Y114_CO5;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X4Y114_CO6;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X4Y114_C_CY;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X4Y114_C_XOR;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X4Y114_D;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X4Y114_D1;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X4Y114_D2;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X4Y114_D3;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X4Y114_D4;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X4Y114_D5;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X4Y114_D6;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X4Y114_DO5;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X4Y114_DO6;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X4Y114_D_CY;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X4Y114_D_XOR;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X5Y114_A;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X5Y114_A1;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X5Y114_A2;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X5Y114_A3;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X5Y114_A4;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X5Y114_A5;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X5Y114_A6;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X5Y114_AO5;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X5Y114_AO6;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X5Y114_A_CY;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X5Y114_A_XOR;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X5Y114_B;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X5Y114_B1;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X5Y114_B2;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X5Y114_B3;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X5Y114_B4;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X5Y114_B5;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X5Y114_B6;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X5Y114_BO5;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X5Y114_BO6;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X5Y114_B_CY;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X5Y114_B_XOR;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X5Y114_C;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X5Y114_C1;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X5Y114_C2;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X5Y114_C3;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X5Y114_C4;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X5Y114_C5;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X5Y114_C6;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X5Y114_CO5;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X5Y114_CO6;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X5Y114_C_CY;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X5Y114_C_XOR;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X5Y114_D;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X5Y114_D1;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X5Y114_D2;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X5Y114_D3;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X5Y114_D4;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X5Y114_D5;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X5Y114_D6;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X5Y114_DO5;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X5Y114_DO6;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X5Y114_D_CY;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X5Y114_D_XOR;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X4Y115_A;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X4Y115_A1;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X4Y115_A2;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X4Y115_A3;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X4Y115_A4;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X4Y115_A5;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X4Y115_A6;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X4Y115_AMUX;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X4Y115_AO5;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X4Y115_AO6;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X4Y115_A_CY;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X4Y115_A_XOR;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X4Y115_B;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X4Y115_B1;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X4Y115_B2;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X4Y115_B3;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X4Y115_B4;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X4Y115_B5;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X4Y115_B6;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X4Y115_BO5;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X4Y115_BO6;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X4Y115_B_CY;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X4Y115_B_XOR;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X4Y115_C;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X4Y115_C1;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X4Y115_C2;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X4Y115_C3;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X4Y115_C4;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X4Y115_C5;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X4Y115_C6;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X4Y115_CO5;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X4Y115_CO6;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X4Y115_C_CY;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X4Y115_C_XOR;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X4Y115_D;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X4Y115_D1;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X4Y115_D2;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X4Y115_D3;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X4Y115_D4;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X4Y115_D5;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X4Y115_D6;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X4Y115_DO5;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X4Y115_DO6;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X4Y115_D_CY;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X4Y115_D_XOR;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X5Y115_A;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X5Y115_A1;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X5Y115_A2;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X5Y115_A3;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X5Y115_A4;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X5Y115_A5;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X5Y115_A6;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X5Y115_AO5;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X5Y115_AO6;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X5Y115_A_CY;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X5Y115_A_XOR;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X5Y115_B;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X5Y115_B1;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X5Y115_B2;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X5Y115_B3;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X5Y115_B4;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X5Y115_B5;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X5Y115_B6;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X5Y115_BO5;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X5Y115_BO6;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X5Y115_B_CY;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X5Y115_B_XOR;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X5Y115_C;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X5Y115_C1;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X5Y115_C2;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X5Y115_C3;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X5Y115_C4;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X5Y115_C5;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X5Y115_C6;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X5Y115_CO5;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X5Y115_CO6;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X5Y115_C_CY;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X5Y115_C_XOR;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X5Y115_D;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X5Y115_D1;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X5Y115_D2;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X5Y115_D3;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X5Y115_D4;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X5Y115_D5;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X5Y115_D6;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X5Y115_DO5;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X5Y115_DO6;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X5Y115_D_CY;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X5Y115_D_XOR;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X4Y116_A;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X4Y116_A1;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X4Y116_A2;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X4Y116_A3;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X4Y116_A4;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X4Y116_A5;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X4Y116_A6;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X4Y116_AO5;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X4Y116_AO6;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X4Y116_A_CY;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X4Y116_A_XOR;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X4Y116_B;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X4Y116_B1;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X4Y116_B2;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X4Y116_B3;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X4Y116_B4;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X4Y116_B5;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X4Y116_B6;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X4Y116_BO5;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X4Y116_BO6;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X4Y116_B_CY;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X4Y116_B_XOR;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X4Y116_C;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X4Y116_C1;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X4Y116_C2;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X4Y116_C3;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X4Y116_C4;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X4Y116_C5;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X4Y116_C6;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X4Y116_CO5;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X4Y116_CO6;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X4Y116_C_CY;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X4Y116_C_XOR;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X4Y116_D;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X4Y116_D1;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X4Y116_D2;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X4Y116_D3;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X4Y116_D4;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X4Y116_D5;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X4Y116_D6;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X4Y116_DO5;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X4Y116_DO6;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X4Y116_D_CY;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X4Y116_D_XOR;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X5Y116_A;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X5Y116_A1;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X5Y116_A2;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X5Y116_A3;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X5Y116_A4;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X5Y116_A5;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X5Y116_A6;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X5Y116_AO5;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X5Y116_AO6;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X5Y116_A_CY;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X5Y116_A_XOR;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X5Y116_B;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X5Y116_B1;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X5Y116_B2;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X5Y116_B3;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X5Y116_B4;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X5Y116_B5;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X5Y116_B6;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X5Y116_BO5;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X5Y116_BO6;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X5Y116_B_CY;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X5Y116_B_XOR;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X5Y116_C;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X5Y116_C1;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X5Y116_C2;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X5Y116_C3;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X5Y116_C4;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X5Y116_C5;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X5Y116_C6;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X5Y116_CO5;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X5Y116_CO6;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X5Y116_C_CY;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X5Y116_C_XOR;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X5Y116_D;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X5Y116_D1;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X5Y116_D2;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X5Y116_D3;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X5Y116_D4;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X5Y116_D5;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X5Y116_D6;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X5Y116_DO5;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X5Y116_DO6;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X5Y116_D_CY;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X5Y116_D_XOR;
  wire [0:0] CLBLM_L_X10Y102_SLICE_X12Y102_A;
  wire [0:0] CLBLM_L_X10Y102_SLICE_X12Y102_A1;
  wire [0:0] CLBLM_L_X10Y102_SLICE_X12Y102_A2;
  wire [0:0] CLBLM_L_X10Y102_SLICE_X12Y102_A3;
  wire [0:0] CLBLM_L_X10Y102_SLICE_X12Y102_A4;
  wire [0:0] CLBLM_L_X10Y102_SLICE_X12Y102_A5;
  wire [0:0] CLBLM_L_X10Y102_SLICE_X12Y102_A6;
  wire [0:0] CLBLM_L_X10Y102_SLICE_X12Y102_AMUX;
  wire [0:0] CLBLM_L_X10Y102_SLICE_X12Y102_AO5;
  wire [0:0] CLBLM_L_X10Y102_SLICE_X12Y102_AO6;
  wire [0:0] CLBLM_L_X10Y102_SLICE_X12Y102_A_CY;
  wire [0:0] CLBLM_L_X10Y102_SLICE_X12Y102_A_XOR;
  wire [0:0] CLBLM_L_X10Y102_SLICE_X12Y102_B;
  wire [0:0] CLBLM_L_X10Y102_SLICE_X12Y102_B1;
  wire [0:0] CLBLM_L_X10Y102_SLICE_X12Y102_B2;
  wire [0:0] CLBLM_L_X10Y102_SLICE_X12Y102_B3;
  wire [0:0] CLBLM_L_X10Y102_SLICE_X12Y102_B4;
  wire [0:0] CLBLM_L_X10Y102_SLICE_X12Y102_B5;
  wire [0:0] CLBLM_L_X10Y102_SLICE_X12Y102_B6;
  wire [0:0] CLBLM_L_X10Y102_SLICE_X12Y102_BMUX;
  wire [0:0] CLBLM_L_X10Y102_SLICE_X12Y102_BO5;
  wire [0:0] CLBLM_L_X10Y102_SLICE_X12Y102_BO6;
  wire [0:0] CLBLM_L_X10Y102_SLICE_X12Y102_B_CY;
  wire [0:0] CLBLM_L_X10Y102_SLICE_X12Y102_B_XOR;
  wire [0:0] CLBLM_L_X10Y102_SLICE_X12Y102_C;
  wire [0:0] CLBLM_L_X10Y102_SLICE_X12Y102_C1;
  wire [0:0] CLBLM_L_X10Y102_SLICE_X12Y102_C2;
  wire [0:0] CLBLM_L_X10Y102_SLICE_X12Y102_C3;
  wire [0:0] CLBLM_L_X10Y102_SLICE_X12Y102_C4;
  wire [0:0] CLBLM_L_X10Y102_SLICE_X12Y102_C5;
  wire [0:0] CLBLM_L_X10Y102_SLICE_X12Y102_C6;
  wire [0:0] CLBLM_L_X10Y102_SLICE_X12Y102_CO5;
  wire [0:0] CLBLM_L_X10Y102_SLICE_X12Y102_CO6;
  wire [0:0] CLBLM_L_X10Y102_SLICE_X12Y102_C_CY;
  wire [0:0] CLBLM_L_X10Y102_SLICE_X12Y102_C_XOR;
  wire [0:0] CLBLM_L_X10Y102_SLICE_X12Y102_D;
  wire [0:0] CLBLM_L_X10Y102_SLICE_X12Y102_D1;
  wire [0:0] CLBLM_L_X10Y102_SLICE_X12Y102_D2;
  wire [0:0] CLBLM_L_X10Y102_SLICE_X12Y102_D3;
  wire [0:0] CLBLM_L_X10Y102_SLICE_X12Y102_D4;
  wire [0:0] CLBLM_L_X10Y102_SLICE_X12Y102_D5;
  wire [0:0] CLBLM_L_X10Y102_SLICE_X12Y102_D6;
  wire [0:0] CLBLM_L_X10Y102_SLICE_X12Y102_DO5;
  wire [0:0] CLBLM_L_X10Y102_SLICE_X12Y102_DO6;
  wire [0:0] CLBLM_L_X10Y102_SLICE_X12Y102_D_CY;
  wire [0:0] CLBLM_L_X10Y102_SLICE_X12Y102_D_XOR;
  wire [0:0] CLBLM_L_X10Y102_SLICE_X13Y102_A;
  wire [0:0] CLBLM_L_X10Y102_SLICE_X13Y102_A1;
  wire [0:0] CLBLM_L_X10Y102_SLICE_X13Y102_A2;
  wire [0:0] CLBLM_L_X10Y102_SLICE_X13Y102_A3;
  wire [0:0] CLBLM_L_X10Y102_SLICE_X13Y102_A4;
  wire [0:0] CLBLM_L_X10Y102_SLICE_X13Y102_A5;
  wire [0:0] CLBLM_L_X10Y102_SLICE_X13Y102_A6;
  wire [0:0] CLBLM_L_X10Y102_SLICE_X13Y102_AO5;
  wire [0:0] CLBLM_L_X10Y102_SLICE_X13Y102_AO6;
  wire [0:0] CLBLM_L_X10Y102_SLICE_X13Y102_A_CY;
  wire [0:0] CLBLM_L_X10Y102_SLICE_X13Y102_A_XOR;
  wire [0:0] CLBLM_L_X10Y102_SLICE_X13Y102_B;
  wire [0:0] CLBLM_L_X10Y102_SLICE_X13Y102_B1;
  wire [0:0] CLBLM_L_X10Y102_SLICE_X13Y102_B2;
  wire [0:0] CLBLM_L_X10Y102_SLICE_X13Y102_B3;
  wire [0:0] CLBLM_L_X10Y102_SLICE_X13Y102_B4;
  wire [0:0] CLBLM_L_X10Y102_SLICE_X13Y102_B5;
  wire [0:0] CLBLM_L_X10Y102_SLICE_X13Y102_B6;
  wire [0:0] CLBLM_L_X10Y102_SLICE_X13Y102_BO5;
  wire [0:0] CLBLM_L_X10Y102_SLICE_X13Y102_BO6;
  wire [0:0] CLBLM_L_X10Y102_SLICE_X13Y102_B_CY;
  wire [0:0] CLBLM_L_X10Y102_SLICE_X13Y102_B_XOR;
  wire [0:0] CLBLM_L_X10Y102_SLICE_X13Y102_C;
  wire [0:0] CLBLM_L_X10Y102_SLICE_X13Y102_C1;
  wire [0:0] CLBLM_L_X10Y102_SLICE_X13Y102_C2;
  wire [0:0] CLBLM_L_X10Y102_SLICE_X13Y102_C3;
  wire [0:0] CLBLM_L_X10Y102_SLICE_X13Y102_C4;
  wire [0:0] CLBLM_L_X10Y102_SLICE_X13Y102_C5;
  wire [0:0] CLBLM_L_X10Y102_SLICE_X13Y102_C6;
  wire [0:0] CLBLM_L_X10Y102_SLICE_X13Y102_CO5;
  wire [0:0] CLBLM_L_X10Y102_SLICE_X13Y102_CO6;
  wire [0:0] CLBLM_L_X10Y102_SLICE_X13Y102_C_CY;
  wire [0:0] CLBLM_L_X10Y102_SLICE_X13Y102_C_XOR;
  wire [0:0] CLBLM_L_X10Y102_SLICE_X13Y102_D;
  wire [0:0] CLBLM_L_X10Y102_SLICE_X13Y102_D1;
  wire [0:0] CLBLM_L_X10Y102_SLICE_X13Y102_D2;
  wire [0:0] CLBLM_L_X10Y102_SLICE_X13Y102_D3;
  wire [0:0] CLBLM_L_X10Y102_SLICE_X13Y102_D4;
  wire [0:0] CLBLM_L_X10Y102_SLICE_X13Y102_D5;
  wire [0:0] CLBLM_L_X10Y102_SLICE_X13Y102_D6;
  wire [0:0] CLBLM_L_X10Y102_SLICE_X13Y102_DO5;
  wire [0:0] CLBLM_L_X10Y102_SLICE_X13Y102_DO6;
  wire [0:0] CLBLM_L_X10Y102_SLICE_X13Y102_D_CY;
  wire [0:0] CLBLM_L_X10Y102_SLICE_X13Y102_D_XOR;
  wire [0:0] CLBLM_L_X10Y103_SLICE_X12Y103_A;
  wire [0:0] CLBLM_L_X10Y103_SLICE_X12Y103_A1;
  wire [0:0] CLBLM_L_X10Y103_SLICE_X12Y103_A2;
  wire [0:0] CLBLM_L_X10Y103_SLICE_X12Y103_A3;
  wire [0:0] CLBLM_L_X10Y103_SLICE_X12Y103_A4;
  wire [0:0] CLBLM_L_X10Y103_SLICE_X12Y103_A5;
  wire [0:0] CLBLM_L_X10Y103_SLICE_X12Y103_A6;
  wire [0:0] CLBLM_L_X10Y103_SLICE_X12Y103_AMUX;
  wire [0:0] CLBLM_L_X10Y103_SLICE_X12Y103_AO5;
  wire [0:0] CLBLM_L_X10Y103_SLICE_X12Y103_AO6;
  wire [0:0] CLBLM_L_X10Y103_SLICE_X12Y103_A_CY;
  wire [0:0] CLBLM_L_X10Y103_SLICE_X12Y103_A_XOR;
  wire [0:0] CLBLM_L_X10Y103_SLICE_X12Y103_B;
  wire [0:0] CLBLM_L_X10Y103_SLICE_X12Y103_B1;
  wire [0:0] CLBLM_L_X10Y103_SLICE_X12Y103_B2;
  wire [0:0] CLBLM_L_X10Y103_SLICE_X12Y103_B3;
  wire [0:0] CLBLM_L_X10Y103_SLICE_X12Y103_B4;
  wire [0:0] CLBLM_L_X10Y103_SLICE_X12Y103_B5;
  wire [0:0] CLBLM_L_X10Y103_SLICE_X12Y103_B6;
  wire [0:0] CLBLM_L_X10Y103_SLICE_X12Y103_BO5;
  wire [0:0] CLBLM_L_X10Y103_SLICE_X12Y103_BO6;
  wire [0:0] CLBLM_L_X10Y103_SLICE_X12Y103_B_CY;
  wire [0:0] CLBLM_L_X10Y103_SLICE_X12Y103_B_XOR;
  wire [0:0] CLBLM_L_X10Y103_SLICE_X12Y103_C;
  wire [0:0] CLBLM_L_X10Y103_SLICE_X12Y103_C1;
  wire [0:0] CLBLM_L_X10Y103_SLICE_X12Y103_C2;
  wire [0:0] CLBLM_L_X10Y103_SLICE_X12Y103_C3;
  wire [0:0] CLBLM_L_X10Y103_SLICE_X12Y103_C4;
  wire [0:0] CLBLM_L_X10Y103_SLICE_X12Y103_C5;
  wire [0:0] CLBLM_L_X10Y103_SLICE_X12Y103_C6;
  wire [0:0] CLBLM_L_X10Y103_SLICE_X12Y103_CO5;
  wire [0:0] CLBLM_L_X10Y103_SLICE_X12Y103_CO6;
  wire [0:0] CLBLM_L_X10Y103_SLICE_X12Y103_C_CY;
  wire [0:0] CLBLM_L_X10Y103_SLICE_X12Y103_C_XOR;
  wire [0:0] CLBLM_L_X10Y103_SLICE_X12Y103_D;
  wire [0:0] CLBLM_L_X10Y103_SLICE_X12Y103_D1;
  wire [0:0] CLBLM_L_X10Y103_SLICE_X12Y103_D2;
  wire [0:0] CLBLM_L_X10Y103_SLICE_X12Y103_D3;
  wire [0:0] CLBLM_L_X10Y103_SLICE_X12Y103_D4;
  wire [0:0] CLBLM_L_X10Y103_SLICE_X12Y103_D5;
  wire [0:0] CLBLM_L_X10Y103_SLICE_X12Y103_D6;
  wire [0:0] CLBLM_L_X10Y103_SLICE_X12Y103_DO5;
  wire [0:0] CLBLM_L_X10Y103_SLICE_X12Y103_DO6;
  wire [0:0] CLBLM_L_X10Y103_SLICE_X12Y103_D_CY;
  wire [0:0] CLBLM_L_X10Y103_SLICE_X12Y103_D_XOR;
  wire [0:0] CLBLM_L_X10Y103_SLICE_X13Y103_A;
  wire [0:0] CLBLM_L_X10Y103_SLICE_X13Y103_A1;
  wire [0:0] CLBLM_L_X10Y103_SLICE_X13Y103_A2;
  wire [0:0] CLBLM_L_X10Y103_SLICE_X13Y103_A3;
  wire [0:0] CLBLM_L_X10Y103_SLICE_X13Y103_A4;
  wire [0:0] CLBLM_L_X10Y103_SLICE_X13Y103_A5;
  wire [0:0] CLBLM_L_X10Y103_SLICE_X13Y103_A6;
  wire [0:0] CLBLM_L_X10Y103_SLICE_X13Y103_AO5;
  wire [0:0] CLBLM_L_X10Y103_SLICE_X13Y103_AO6;
  wire [0:0] CLBLM_L_X10Y103_SLICE_X13Y103_A_CY;
  wire [0:0] CLBLM_L_X10Y103_SLICE_X13Y103_A_XOR;
  wire [0:0] CLBLM_L_X10Y103_SLICE_X13Y103_B;
  wire [0:0] CLBLM_L_X10Y103_SLICE_X13Y103_B1;
  wire [0:0] CLBLM_L_X10Y103_SLICE_X13Y103_B2;
  wire [0:0] CLBLM_L_X10Y103_SLICE_X13Y103_B3;
  wire [0:0] CLBLM_L_X10Y103_SLICE_X13Y103_B4;
  wire [0:0] CLBLM_L_X10Y103_SLICE_X13Y103_B5;
  wire [0:0] CLBLM_L_X10Y103_SLICE_X13Y103_B6;
  wire [0:0] CLBLM_L_X10Y103_SLICE_X13Y103_BO5;
  wire [0:0] CLBLM_L_X10Y103_SLICE_X13Y103_BO6;
  wire [0:0] CLBLM_L_X10Y103_SLICE_X13Y103_B_CY;
  wire [0:0] CLBLM_L_X10Y103_SLICE_X13Y103_B_XOR;
  wire [0:0] CLBLM_L_X10Y103_SLICE_X13Y103_C;
  wire [0:0] CLBLM_L_X10Y103_SLICE_X13Y103_C1;
  wire [0:0] CLBLM_L_X10Y103_SLICE_X13Y103_C2;
  wire [0:0] CLBLM_L_X10Y103_SLICE_X13Y103_C3;
  wire [0:0] CLBLM_L_X10Y103_SLICE_X13Y103_C4;
  wire [0:0] CLBLM_L_X10Y103_SLICE_X13Y103_C5;
  wire [0:0] CLBLM_L_X10Y103_SLICE_X13Y103_C6;
  wire [0:0] CLBLM_L_X10Y103_SLICE_X13Y103_CO5;
  wire [0:0] CLBLM_L_X10Y103_SLICE_X13Y103_CO6;
  wire [0:0] CLBLM_L_X10Y103_SLICE_X13Y103_C_CY;
  wire [0:0] CLBLM_L_X10Y103_SLICE_X13Y103_C_XOR;
  wire [0:0] CLBLM_L_X10Y103_SLICE_X13Y103_D;
  wire [0:0] CLBLM_L_X10Y103_SLICE_X13Y103_D1;
  wire [0:0] CLBLM_L_X10Y103_SLICE_X13Y103_D2;
  wire [0:0] CLBLM_L_X10Y103_SLICE_X13Y103_D3;
  wire [0:0] CLBLM_L_X10Y103_SLICE_X13Y103_D4;
  wire [0:0] CLBLM_L_X10Y103_SLICE_X13Y103_D5;
  wire [0:0] CLBLM_L_X10Y103_SLICE_X13Y103_D6;
  wire [0:0] CLBLM_L_X10Y103_SLICE_X13Y103_DO5;
  wire [0:0] CLBLM_L_X10Y103_SLICE_X13Y103_DO6;
  wire [0:0] CLBLM_L_X10Y103_SLICE_X13Y103_D_CY;
  wire [0:0] CLBLM_L_X10Y103_SLICE_X13Y103_D_XOR;
  wire [0:0] CLBLM_L_X10Y104_SLICE_X12Y104_A;
  wire [0:0] CLBLM_L_X10Y104_SLICE_X12Y104_A1;
  wire [0:0] CLBLM_L_X10Y104_SLICE_X12Y104_A2;
  wire [0:0] CLBLM_L_X10Y104_SLICE_X12Y104_A3;
  wire [0:0] CLBLM_L_X10Y104_SLICE_X12Y104_A4;
  wire [0:0] CLBLM_L_X10Y104_SLICE_X12Y104_A5;
  wire [0:0] CLBLM_L_X10Y104_SLICE_X12Y104_A6;
  wire [0:0] CLBLM_L_X10Y104_SLICE_X12Y104_AO5;
  wire [0:0] CLBLM_L_X10Y104_SLICE_X12Y104_AO6;
  wire [0:0] CLBLM_L_X10Y104_SLICE_X12Y104_A_CY;
  wire [0:0] CLBLM_L_X10Y104_SLICE_X12Y104_A_XOR;
  wire [0:0] CLBLM_L_X10Y104_SLICE_X12Y104_B;
  wire [0:0] CLBLM_L_X10Y104_SLICE_X12Y104_B1;
  wire [0:0] CLBLM_L_X10Y104_SLICE_X12Y104_B2;
  wire [0:0] CLBLM_L_X10Y104_SLICE_X12Y104_B3;
  wire [0:0] CLBLM_L_X10Y104_SLICE_X12Y104_B4;
  wire [0:0] CLBLM_L_X10Y104_SLICE_X12Y104_B5;
  wire [0:0] CLBLM_L_X10Y104_SLICE_X12Y104_B6;
  wire [0:0] CLBLM_L_X10Y104_SLICE_X12Y104_BMUX;
  wire [0:0] CLBLM_L_X10Y104_SLICE_X12Y104_BO5;
  wire [0:0] CLBLM_L_X10Y104_SLICE_X12Y104_BO6;
  wire [0:0] CLBLM_L_X10Y104_SLICE_X12Y104_B_CY;
  wire [0:0] CLBLM_L_X10Y104_SLICE_X12Y104_B_XOR;
  wire [0:0] CLBLM_L_X10Y104_SLICE_X12Y104_C;
  wire [0:0] CLBLM_L_X10Y104_SLICE_X12Y104_C1;
  wire [0:0] CLBLM_L_X10Y104_SLICE_X12Y104_C2;
  wire [0:0] CLBLM_L_X10Y104_SLICE_X12Y104_C3;
  wire [0:0] CLBLM_L_X10Y104_SLICE_X12Y104_C4;
  wire [0:0] CLBLM_L_X10Y104_SLICE_X12Y104_C5;
  wire [0:0] CLBLM_L_X10Y104_SLICE_X12Y104_C6;
  wire [0:0] CLBLM_L_X10Y104_SLICE_X12Y104_CO5;
  wire [0:0] CLBLM_L_X10Y104_SLICE_X12Y104_CO6;
  wire [0:0] CLBLM_L_X10Y104_SLICE_X12Y104_C_CY;
  wire [0:0] CLBLM_L_X10Y104_SLICE_X12Y104_C_XOR;
  wire [0:0] CLBLM_L_X10Y104_SLICE_X12Y104_D;
  wire [0:0] CLBLM_L_X10Y104_SLICE_X12Y104_D1;
  wire [0:0] CLBLM_L_X10Y104_SLICE_X12Y104_D2;
  wire [0:0] CLBLM_L_X10Y104_SLICE_X12Y104_D3;
  wire [0:0] CLBLM_L_X10Y104_SLICE_X12Y104_D4;
  wire [0:0] CLBLM_L_X10Y104_SLICE_X12Y104_D5;
  wire [0:0] CLBLM_L_X10Y104_SLICE_X12Y104_D6;
  wire [0:0] CLBLM_L_X10Y104_SLICE_X12Y104_DO5;
  wire [0:0] CLBLM_L_X10Y104_SLICE_X12Y104_DO6;
  wire [0:0] CLBLM_L_X10Y104_SLICE_X12Y104_D_CY;
  wire [0:0] CLBLM_L_X10Y104_SLICE_X12Y104_D_XOR;
  wire [0:0] CLBLM_L_X10Y104_SLICE_X13Y104_A;
  wire [0:0] CLBLM_L_X10Y104_SLICE_X13Y104_A1;
  wire [0:0] CLBLM_L_X10Y104_SLICE_X13Y104_A2;
  wire [0:0] CLBLM_L_X10Y104_SLICE_X13Y104_A3;
  wire [0:0] CLBLM_L_X10Y104_SLICE_X13Y104_A4;
  wire [0:0] CLBLM_L_X10Y104_SLICE_X13Y104_A5;
  wire [0:0] CLBLM_L_X10Y104_SLICE_X13Y104_A6;
  wire [0:0] CLBLM_L_X10Y104_SLICE_X13Y104_AMUX;
  wire [0:0] CLBLM_L_X10Y104_SLICE_X13Y104_AO5;
  wire [0:0] CLBLM_L_X10Y104_SLICE_X13Y104_AO6;
  wire [0:0] CLBLM_L_X10Y104_SLICE_X13Y104_A_CY;
  wire [0:0] CLBLM_L_X10Y104_SLICE_X13Y104_A_XOR;
  wire [0:0] CLBLM_L_X10Y104_SLICE_X13Y104_B;
  wire [0:0] CLBLM_L_X10Y104_SLICE_X13Y104_B1;
  wire [0:0] CLBLM_L_X10Y104_SLICE_X13Y104_B2;
  wire [0:0] CLBLM_L_X10Y104_SLICE_X13Y104_B3;
  wire [0:0] CLBLM_L_X10Y104_SLICE_X13Y104_B4;
  wire [0:0] CLBLM_L_X10Y104_SLICE_X13Y104_B5;
  wire [0:0] CLBLM_L_X10Y104_SLICE_X13Y104_B6;
  wire [0:0] CLBLM_L_X10Y104_SLICE_X13Y104_BO5;
  wire [0:0] CLBLM_L_X10Y104_SLICE_X13Y104_BO6;
  wire [0:0] CLBLM_L_X10Y104_SLICE_X13Y104_B_CY;
  wire [0:0] CLBLM_L_X10Y104_SLICE_X13Y104_B_XOR;
  wire [0:0] CLBLM_L_X10Y104_SLICE_X13Y104_C;
  wire [0:0] CLBLM_L_X10Y104_SLICE_X13Y104_C1;
  wire [0:0] CLBLM_L_X10Y104_SLICE_X13Y104_C2;
  wire [0:0] CLBLM_L_X10Y104_SLICE_X13Y104_C3;
  wire [0:0] CLBLM_L_X10Y104_SLICE_X13Y104_C4;
  wire [0:0] CLBLM_L_X10Y104_SLICE_X13Y104_C5;
  wire [0:0] CLBLM_L_X10Y104_SLICE_X13Y104_C6;
  wire [0:0] CLBLM_L_X10Y104_SLICE_X13Y104_CO5;
  wire [0:0] CLBLM_L_X10Y104_SLICE_X13Y104_CO6;
  wire [0:0] CLBLM_L_X10Y104_SLICE_X13Y104_C_CY;
  wire [0:0] CLBLM_L_X10Y104_SLICE_X13Y104_C_XOR;
  wire [0:0] CLBLM_L_X10Y104_SLICE_X13Y104_D;
  wire [0:0] CLBLM_L_X10Y104_SLICE_X13Y104_D1;
  wire [0:0] CLBLM_L_X10Y104_SLICE_X13Y104_D2;
  wire [0:0] CLBLM_L_X10Y104_SLICE_X13Y104_D3;
  wire [0:0] CLBLM_L_X10Y104_SLICE_X13Y104_D4;
  wire [0:0] CLBLM_L_X10Y104_SLICE_X13Y104_D5;
  wire [0:0] CLBLM_L_X10Y104_SLICE_X13Y104_D6;
  wire [0:0] CLBLM_L_X10Y104_SLICE_X13Y104_DO5;
  wire [0:0] CLBLM_L_X10Y104_SLICE_X13Y104_DO6;
  wire [0:0] CLBLM_L_X10Y104_SLICE_X13Y104_D_CY;
  wire [0:0] CLBLM_L_X10Y104_SLICE_X13Y104_D_XOR;
  wire [0:0] CLBLM_L_X10Y105_SLICE_X12Y105_A;
  wire [0:0] CLBLM_L_X10Y105_SLICE_X12Y105_A1;
  wire [0:0] CLBLM_L_X10Y105_SLICE_X12Y105_A2;
  wire [0:0] CLBLM_L_X10Y105_SLICE_X12Y105_A3;
  wire [0:0] CLBLM_L_X10Y105_SLICE_X12Y105_A4;
  wire [0:0] CLBLM_L_X10Y105_SLICE_X12Y105_A5;
  wire [0:0] CLBLM_L_X10Y105_SLICE_X12Y105_A6;
  wire [0:0] CLBLM_L_X10Y105_SLICE_X12Y105_AMUX;
  wire [0:0] CLBLM_L_X10Y105_SLICE_X12Y105_AO5;
  wire [0:0] CLBLM_L_X10Y105_SLICE_X12Y105_AO6;
  wire [0:0] CLBLM_L_X10Y105_SLICE_X12Y105_A_CY;
  wire [0:0] CLBLM_L_X10Y105_SLICE_X12Y105_A_XOR;
  wire [0:0] CLBLM_L_X10Y105_SLICE_X12Y105_B;
  wire [0:0] CLBLM_L_X10Y105_SLICE_X12Y105_B1;
  wire [0:0] CLBLM_L_X10Y105_SLICE_X12Y105_B2;
  wire [0:0] CLBLM_L_X10Y105_SLICE_X12Y105_B3;
  wire [0:0] CLBLM_L_X10Y105_SLICE_X12Y105_B4;
  wire [0:0] CLBLM_L_X10Y105_SLICE_X12Y105_B5;
  wire [0:0] CLBLM_L_X10Y105_SLICE_X12Y105_B6;
  wire [0:0] CLBLM_L_X10Y105_SLICE_X12Y105_BO5;
  wire [0:0] CLBLM_L_X10Y105_SLICE_X12Y105_BO6;
  wire [0:0] CLBLM_L_X10Y105_SLICE_X12Y105_B_CY;
  wire [0:0] CLBLM_L_X10Y105_SLICE_X12Y105_B_XOR;
  wire [0:0] CLBLM_L_X10Y105_SLICE_X12Y105_C;
  wire [0:0] CLBLM_L_X10Y105_SLICE_X12Y105_C1;
  wire [0:0] CLBLM_L_X10Y105_SLICE_X12Y105_C2;
  wire [0:0] CLBLM_L_X10Y105_SLICE_X12Y105_C3;
  wire [0:0] CLBLM_L_X10Y105_SLICE_X12Y105_C4;
  wire [0:0] CLBLM_L_X10Y105_SLICE_X12Y105_C5;
  wire [0:0] CLBLM_L_X10Y105_SLICE_X12Y105_C6;
  wire [0:0] CLBLM_L_X10Y105_SLICE_X12Y105_CO5;
  wire [0:0] CLBLM_L_X10Y105_SLICE_X12Y105_CO6;
  wire [0:0] CLBLM_L_X10Y105_SLICE_X12Y105_C_CY;
  wire [0:0] CLBLM_L_X10Y105_SLICE_X12Y105_C_XOR;
  wire [0:0] CLBLM_L_X10Y105_SLICE_X12Y105_D;
  wire [0:0] CLBLM_L_X10Y105_SLICE_X12Y105_D1;
  wire [0:0] CLBLM_L_X10Y105_SLICE_X12Y105_D2;
  wire [0:0] CLBLM_L_X10Y105_SLICE_X12Y105_D3;
  wire [0:0] CLBLM_L_X10Y105_SLICE_X12Y105_D4;
  wire [0:0] CLBLM_L_X10Y105_SLICE_X12Y105_D5;
  wire [0:0] CLBLM_L_X10Y105_SLICE_X12Y105_D6;
  wire [0:0] CLBLM_L_X10Y105_SLICE_X12Y105_DO5;
  wire [0:0] CLBLM_L_X10Y105_SLICE_X12Y105_DO6;
  wire [0:0] CLBLM_L_X10Y105_SLICE_X12Y105_D_CY;
  wire [0:0] CLBLM_L_X10Y105_SLICE_X12Y105_D_XOR;
  wire [0:0] CLBLM_L_X10Y105_SLICE_X13Y105_A;
  wire [0:0] CLBLM_L_X10Y105_SLICE_X13Y105_A1;
  wire [0:0] CLBLM_L_X10Y105_SLICE_X13Y105_A2;
  wire [0:0] CLBLM_L_X10Y105_SLICE_X13Y105_A3;
  wire [0:0] CLBLM_L_X10Y105_SLICE_X13Y105_A4;
  wire [0:0] CLBLM_L_X10Y105_SLICE_X13Y105_A5;
  wire [0:0] CLBLM_L_X10Y105_SLICE_X13Y105_A6;
  wire [0:0] CLBLM_L_X10Y105_SLICE_X13Y105_AMUX;
  wire [0:0] CLBLM_L_X10Y105_SLICE_X13Y105_AO5;
  wire [0:0] CLBLM_L_X10Y105_SLICE_X13Y105_AO6;
  wire [0:0] CLBLM_L_X10Y105_SLICE_X13Y105_A_CY;
  wire [0:0] CLBLM_L_X10Y105_SLICE_X13Y105_A_XOR;
  wire [0:0] CLBLM_L_X10Y105_SLICE_X13Y105_B;
  wire [0:0] CLBLM_L_X10Y105_SLICE_X13Y105_B1;
  wire [0:0] CLBLM_L_X10Y105_SLICE_X13Y105_B2;
  wire [0:0] CLBLM_L_X10Y105_SLICE_X13Y105_B3;
  wire [0:0] CLBLM_L_X10Y105_SLICE_X13Y105_B4;
  wire [0:0] CLBLM_L_X10Y105_SLICE_X13Y105_B5;
  wire [0:0] CLBLM_L_X10Y105_SLICE_X13Y105_B6;
  wire [0:0] CLBLM_L_X10Y105_SLICE_X13Y105_BO5;
  wire [0:0] CLBLM_L_X10Y105_SLICE_X13Y105_BO6;
  wire [0:0] CLBLM_L_X10Y105_SLICE_X13Y105_B_CY;
  wire [0:0] CLBLM_L_X10Y105_SLICE_X13Y105_B_XOR;
  wire [0:0] CLBLM_L_X10Y105_SLICE_X13Y105_C;
  wire [0:0] CLBLM_L_X10Y105_SLICE_X13Y105_C1;
  wire [0:0] CLBLM_L_X10Y105_SLICE_X13Y105_C2;
  wire [0:0] CLBLM_L_X10Y105_SLICE_X13Y105_C3;
  wire [0:0] CLBLM_L_X10Y105_SLICE_X13Y105_C4;
  wire [0:0] CLBLM_L_X10Y105_SLICE_X13Y105_C5;
  wire [0:0] CLBLM_L_X10Y105_SLICE_X13Y105_C6;
  wire [0:0] CLBLM_L_X10Y105_SLICE_X13Y105_CO5;
  wire [0:0] CLBLM_L_X10Y105_SLICE_X13Y105_CO6;
  wire [0:0] CLBLM_L_X10Y105_SLICE_X13Y105_C_CY;
  wire [0:0] CLBLM_L_X10Y105_SLICE_X13Y105_C_XOR;
  wire [0:0] CLBLM_L_X10Y105_SLICE_X13Y105_D;
  wire [0:0] CLBLM_L_X10Y105_SLICE_X13Y105_D1;
  wire [0:0] CLBLM_L_X10Y105_SLICE_X13Y105_D2;
  wire [0:0] CLBLM_L_X10Y105_SLICE_X13Y105_D3;
  wire [0:0] CLBLM_L_X10Y105_SLICE_X13Y105_D4;
  wire [0:0] CLBLM_L_X10Y105_SLICE_X13Y105_D5;
  wire [0:0] CLBLM_L_X10Y105_SLICE_X13Y105_D6;
  wire [0:0] CLBLM_L_X10Y105_SLICE_X13Y105_DO5;
  wire [0:0] CLBLM_L_X10Y105_SLICE_X13Y105_DO6;
  wire [0:0] CLBLM_L_X10Y105_SLICE_X13Y105_D_CY;
  wire [0:0] CLBLM_L_X10Y105_SLICE_X13Y105_D_XOR;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X12Y106_A;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X12Y106_A1;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X12Y106_A2;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X12Y106_A3;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X12Y106_A4;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X12Y106_A5;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X12Y106_A6;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X12Y106_AO5;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X12Y106_AO6;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X12Y106_A_CY;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X12Y106_A_XOR;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X12Y106_B;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X12Y106_B1;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X12Y106_B2;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X12Y106_B3;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X12Y106_B4;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X12Y106_B5;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X12Y106_B6;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X12Y106_BO5;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X12Y106_BO6;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X12Y106_B_CY;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X12Y106_B_XOR;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X12Y106_C;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X12Y106_C1;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X12Y106_C2;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X12Y106_C3;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X12Y106_C4;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X12Y106_C5;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X12Y106_C6;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X12Y106_CO5;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X12Y106_CO6;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X12Y106_C_CY;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X12Y106_C_XOR;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X12Y106_D;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X12Y106_D1;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X12Y106_D2;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X12Y106_D3;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X12Y106_D4;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X12Y106_D5;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X12Y106_D6;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X12Y106_DO5;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X12Y106_DO6;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X12Y106_D_CY;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X12Y106_D_XOR;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X13Y106_A;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X13Y106_A1;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X13Y106_A2;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X13Y106_A3;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X13Y106_A4;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X13Y106_A5;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X13Y106_A6;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X13Y106_AO5;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X13Y106_AO6;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X13Y106_A_CY;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X13Y106_A_XOR;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X13Y106_B;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X13Y106_B1;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X13Y106_B2;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X13Y106_B3;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X13Y106_B4;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X13Y106_B5;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X13Y106_B6;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X13Y106_BO5;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X13Y106_BO6;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X13Y106_B_CY;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X13Y106_B_XOR;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X13Y106_C;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X13Y106_C1;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X13Y106_C2;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X13Y106_C3;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X13Y106_C4;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X13Y106_C5;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X13Y106_C6;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X13Y106_CO5;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X13Y106_CO6;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X13Y106_C_CY;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X13Y106_C_XOR;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X13Y106_D;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X13Y106_D1;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X13Y106_D2;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X13Y106_D3;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X13Y106_D4;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X13Y106_D5;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X13Y106_D6;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X13Y106_DO5;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X13Y106_DO6;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X13Y106_D_CY;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X13Y106_D_XOR;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X12Y107_A;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X12Y107_A1;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X12Y107_A2;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X12Y107_A3;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X12Y107_A4;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X12Y107_A5;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X12Y107_A6;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X12Y107_AO5;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X12Y107_AO6;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X12Y107_A_CY;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X12Y107_A_XOR;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X12Y107_B;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X12Y107_B1;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X12Y107_B2;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X12Y107_B3;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X12Y107_B4;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X12Y107_B5;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X12Y107_B6;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X12Y107_BO5;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X12Y107_BO6;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X12Y107_B_CY;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X12Y107_B_XOR;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X12Y107_C;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X12Y107_C1;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X12Y107_C2;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X12Y107_C3;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X12Y107_C4;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X12Y107_C5;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X12Y107_C6;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X12Y107_CO5;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X12Y107_CO6;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X12Y107_C_CY;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X12Y107_C_XOR;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X12Y107_D;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X12Y107_D1;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X12Y107_D2;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X12Y107_D3;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X12Y107_D4;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X12Y107_D5;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X12Y107_D6;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X12Y107_DO5;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X12Y107_DO6;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X12Y107_D_CY;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X12Y107_D_XOR;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X13Y107_A;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X13Y107_A1;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X13Y107_A2;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X13Y107_A3;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X13Y107_A4;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X13Y107_A5;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X13Y107_A6;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X13Y107_AMUX;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X13Y107_AO5;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X13Y107_AO6;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X13Y107_A_CY;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X13Y107_A_XOR;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X13Y107_B;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X13Y107_B1;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X13Y107_B2;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X13Y107_B3;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X13Y107_B4;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X13Y107_B5;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X13Y107_B6;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X13Y107_BO5;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X13Y107_BO6;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X13Y107_B_CY;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X13Y107_B_XOR;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X13Y107_C;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X13Y107_C1;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X13Y107_C2;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X13Y107_C3;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X13Y107_C4;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X13Y107_C5;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X13Y107_C6;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X13Y107_CO5;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X13Y107_CO6;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X13Y107_C_CY;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X13Y107_C_XOR;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X13Y107_D;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X13Y107_D1;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X13Y107_D2;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X13Y107_D3;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X13Y107_D4;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X13Y107_D5;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X13Y107_D6;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X13Y107_DO5;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X13Y107_DO6;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X13Y107_D_CY;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X13Y107_D_XOR;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X12Y108_A;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X12Y108_A1;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X12Y108_A2;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X12Y108_A3;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X12Y108_A4;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X12Y108_A5;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X12Y108_A6;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X12Y108_AO5;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X12Y108_AO6;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X12Y108_A_CY;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X12Y108_A_XOR;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X12Y108_B;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X12Y108_B1;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X12Y108_B2;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X12Y108_B3;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X12Y108_B4;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X12Y108_B5;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X12Y108_B6;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X12Y108_BO5;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X12Y108_BO6;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X12Y108_B_CY;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X12Y108_B_XOR;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X12Y108_C;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X12Y108_C1;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X12Y108_C2;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X12Y108_C3;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X12Y108_C4;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X12Y108_C5;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X12Y108_C6;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X12Y108_CO5;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X12Y108_CO6;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X12Y108_C_CY;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X12Y108_C_XOR;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X12Y108_D;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X12Y108_D1;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X12Y108_D2;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X12Y108_D3;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X12Y108_D4;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X12Y108_D5;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X12Y108_D6;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X12Y108_DO5;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X12Y108_DO6;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X12Y108_D_CY;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X12Y108_D_XOR;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X13Y108_A;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X13Y108_A1;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X13Y108_A2;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X13Y108_A3;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X13Y108_A4;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X13Y108_A5;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X13Y108_A6;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X13Y108_AMUX;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X13Y108_AO5;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X13Y108_AO6;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X13Y108_A_CY;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X13Y108_A_XOR;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X13Y108_B;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X13Y108_B1;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X13Y108_B2;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X13Y108_B3;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X13Y108_B4;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X13Y108_B5;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X13Y108_B6;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X13Y108_BMUX;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X13Y108_BO5;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X13Y108_BO6;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X13Y108_B_CY;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X13Y108_B_XOR;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X13Y108_C;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X13Y108_C1;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X13Y108_C2;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X13Y108_C3;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X13Y108_C4;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X13Y108_C5;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X13Y108_C6;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X13Y108_CMUX;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X13Y108_CO5;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X13Y108_CO6;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X13Y108_C_CY;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X13Y108_C_XOR;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X13Y108_D;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X13Y108_D1;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X13Y108_D2;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X13Y108_D3;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X13Y108_D4;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X13Y108_D5;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X13Y108_D6;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X13Y108_DO5;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X13Y108_DO6;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X13Y108_D_CY;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X13Y108_D_XOR;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X12Y109_A;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X12Y109_A1;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X12Y109_A2;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X12Y109_A3;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X12Y109_A4;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X12Y109_A5;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X12Y109_A6;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X12Y109_AMUX;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X12Y109_AO5;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X12Y109_AO6;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X12Y109_A_CY;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X12Y109_A_XOR;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X12Y109_B;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X12Y109_B1;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X12Y109_B2;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X12Y109_B3;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X12Y109_B4;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X12Y109_B5;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X12Y109_B6;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X12Y109_BO5;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X12Y109_BO6;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X12Y109_B_CY;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X12Y109_B_XOR;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X12Y109_C;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X12Y109_C1;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X12Y109_C2;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X12Y109_C3;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X12Y109_C4;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X12Y109_C5;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X12Y109_C6;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X12Y109_CO5;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X12Y109_CO6;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X12Y109_C_CY;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X12Y109_C_XOR;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X12Y109_D;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X12Y109_D1;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X12Y109_D2;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X12Y109_D3;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X12Y109_D4;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X12Y109_D5;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X12Y109_D6;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X12Y109_DO5;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X12Y109_DO6;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X12Y109_D_CY;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X12Y109_D_XOR;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X13Y109_A;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X13Y109_A1;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X13Y109_A2;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X13Y109_A3;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X13Y109_A4;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X13Y109_A5;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X13Y109_A6;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X13Y109_AMUX;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X13Y109_AO5;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X13Y109_AO6;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X13Y109_A_CY;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X13Y109_A_XOR;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X13Y109_B;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X13Y109_B1;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X13Y109_B2;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X13Y109_B3;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X13Y109_B4;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X13Y109_B5;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X13Y109_B6;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X13Y109_BO5;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X13Y109_BO6;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X13Y109_B_CY;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X13Y109_B_XOR;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X13Y109_C;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X13Y109_C1;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X13Y109_C2;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X13Y109_C3;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X13Y109_C4;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X13Y109_C5;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X13Y109_C6;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X13Y109_CO5;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X13Y109_CO6;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X13Y109_C_CY;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X13Y109_C_XOR;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X13Y109_D;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X13Y109_D1;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X13Y109_D2;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X13Y109_D3;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X13Y109_D4;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X13Y109_D5;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X13Y109_D6;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X13Y109_DO5;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X13Y109_DO6;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X13Y109_D_CY;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X13Y109_D_XOR;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X12Y110_A;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X12Y110_A1;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X12Y110_A2;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X12Y110_A3;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X12Y110_A4;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X12Y110_A5;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X12Y110_A6;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X12Y110_AO5;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X12Y110_AO6;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X12Y110_A_CY;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X12Y110_A_XOR;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X12Y110_B;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X12Y110_B1;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X12Y110_B2;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X12Y110_B3;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X12Y110_B4;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X12Y110_B5;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X12Y110_B6;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X12Y110_BO5;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X12Y110_BO6;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X12Y110_B_CY;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X12Y110_B_XOR;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X12Y110_C;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X12Y110_C1;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X12Y110_C2;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X12Y110_C3;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X12Y110_C4;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X12Y110_C5;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X12Y110_C6;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X12Y110_CO5;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X12Y110_CO6;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X12Y110_C_CY;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X12Y110_C_XOR;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X12Y110_D;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X12Y110_D1;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X12Y110_D2;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X12Y110_D3;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X12Y110_D4;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X12Y110_D5;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X12Y110_D6;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X12Y110_DO5;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X12Y110_DO6;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X12Y110_D_CY;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X12Y110_D_XOR;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X13Y110_A;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X13Y110_A1;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X13Y110_A2;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X13Y110_A3;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X13Y110_A4;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X13Y110_A5;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X13Y110_A6;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X13Y110_AMUX;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X13Y110_AO5;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X13Y110_AO6;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X13Y110_A_CY;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X13Y110_A_XOR;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X13Y110_B;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X13Y110_B1;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X13Y110_B2;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X13Y110_B3;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X13Y110_B4;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X13Y110_B5;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X13Y110_B6;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X13Y110_BO5;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X13Y110_BO6;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X13Y110_B_CY;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X13Y110_B_XOR;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X13Y110_C;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X13Y110_C1;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X13Y110_C2;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X13Y110_C3;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X13Y110_C4;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X13Y110_C5;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X13Y110_C6;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X13Y110_CO5;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X13Y110_CO6;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X13Y110_C_CY;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X13Y110_C_XOR;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X13Y110_D;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X13Y110_D1;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X13Y110_D2;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X13Y110_D3;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X13Y110_D4;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X13Y110_D5;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X13Y110_D6;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X13Y110_DO5;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X13Y110_DO6;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X13Y110_D_CY;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X13Y110_D_XOR;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X12Y111_A;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X12Y111_A1;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X12Y111_A2;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X12Y111_A3;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X12Y111_A4;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X12Y111_A5;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X12Y111_A6;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X12Y111_AO5;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X12Y111_AO6;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X12Y111_A_CY;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X12Y111_A_XOR;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X12Y111_B;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X12Y111_B1;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X12Y111_B2;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X12Y111_B3;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X12Y111_B4;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X12Y111_B5;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X12Y111_B6;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X12Y111_BO5;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X12Y111_BO6;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X12Y111_B_CY;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X12Y111_B_XOR;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X12Y111_C;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X12Y111_C1;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X12Y111_C2;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X12Y111_C3;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X12Y111_C4;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X12Y111_C5;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X12Y111_C6;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X12Y111_CO5;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X12Y111_CO6;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X12Y111_C_CY;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X12Y111_C_XOR;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X12Y111_D;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X12Y111_D1;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X12Y111_D2;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X12Y111_D3;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X12Y111_D4;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X12Y111_D5;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X12Y111_D6;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X12Y111_DO5;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X12Y111_DO6;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X12Y111_D_CY;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X12Y111_D_XOR;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X13Y111_A;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X13Y111_A1;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X13Y111_A2;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X13Y111_A3;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X13Y111_A4;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X13Y111_A5;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X13Y111_A6;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X13Y111_AMUX;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X13Y111_AO5;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X13Y111_AO6;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X13Y111_A_CY;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X13Y111_A_XOR;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X13Y111_B;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X13Y111_B1;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X13Y111_B2;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X13Y111_B3;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X13Y111_B4;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X13Y111_B5;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X13Y111_B6;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X13Y111_BMUX;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X13Y111_BO5;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X13Y111_BO6;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X13Y111_B_CY;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X13Y111_B_XOR;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X13Y111_C;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X13Y111_C1;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X13Y111_C2;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X13Y111_C3;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X13Y111_C4;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X13Y111_C5;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X13Y111_C6;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X13Y111_CO5;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X13Y111_CO6;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X13Y111_C_CY;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X13Y111_C_XOR;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X13Y111_D;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X13Y111_D1;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X13Y111_D2;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X13Y111_D3;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X13Y111_D4;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X13Y111_D5;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X13Y111_D6;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X13Y111_DO5;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X13Y111_DO6;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X13Y111_D_CY;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X13Y111_D_XOR;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X12Y112_A;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X12Y112_A1;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X12Y112_A2;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X12Y112_A3;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X12Y112_A4;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X12Y112_A5;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X12Y112_A6;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X12Y112_AO5;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X12Y112_AO6;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X12Y112_A_CY;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X12Y112_A_XOR;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X12Y112_B;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X12Y112_B1;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X12Y112_B2;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X12Y112_B3;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X12Y112_B4;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X12Y112_B5;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X12Y112_B6;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X12Y112_BO5;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X12Y112_BO6;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X12Y112_B_CY;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X12Y112_B_XOR;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X12Y112_C;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X12Y112_C1;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X12Y112_C2;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X12Y112_C3;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X12Y112_C4;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X12Y112_C5;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X12Y112_C6;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X12Y112_CO5;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X12Y112_CO6;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X12Y112_C_CY;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X12Y112_C_XOR;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X12Y112_D;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X12Y112_D1;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X12Y112_D2;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X12Y112_D3;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X12Y112_D4;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X12Y112_D5;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X12Y112_D6;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X12Y112_DO5;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X12Y112_DO6;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X12Y112_D_CY;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X12Y112_D_XOR;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X13Y112_A;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X13Y112_A1;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X13Y112_A2;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X13Y112_A3;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X13Y112_A4;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X13Y112_A5;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X13Y112_A6;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X13Y112_AMUX;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X13Y112_AO5;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X13Y112_AO6;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X13Y112_A_CY;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X13Y112_A_XOR;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X13Y112_B;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X13Y112_B1;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X13Y112_B2;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X13Y112_B3;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X13Y112_B4;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X13Y112_B5;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X13Y112_B6;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X13Y112_BO5;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X13Y112_BO6;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X13Y112_B_CY;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X13Y112_B_XOR;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X13Y112_C;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X13Y112_C1;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X13Y112_C2;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X13Y112_C3;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X13Y112_C4;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X13Y112_C5;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X13Y112_C6;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X13Y112_CO5;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X13Y112_CO6;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X13Y112_C_CY;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X13Y112_C_XOR;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X13Y112_D;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X13Y112_D1;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X13Y112_D2;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X13Y112_D3;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X13Y112_D4;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X13Y112_D5;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X13Y112_D6;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X13Y112_DO5;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X13Y112_DO6;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X13Y112_D_CY;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X13Y112_D_XOR;
  wire [0:0] CLBLM_L_X12Y104_SLICE_X16Y104_A;
  wire [0:0] CLBLM_L_X12Y104_SLICE_X16Y104_A1;
  wire [0:0] CLBLM_L_X12Y104_SLICE_X16Y104_A2;
  wire [0:0] CLBLM_L_X12Y104_SLICE_X16Y104_A3;
  wire [0:0] CLBLM_L_X12Y104_SLICE_X16Y104_A4;
  wire [0:0] CLBLM_L_X12Y104_SLICE_X16Y104_A5;
  wire [0:0] CLBLM_L_X12Y104_SLICE_X16Y104_A6;
  wire [0:0] CLBLM_L_X12Y104_SLICE_X16Y104_AMUX;
  wire [0:0] CLBLM_L_X12Y104_SLICE_X16Y104_AO5;
  wire [0:0] CLBLM_L_X12Y104_SLICE_X16Y104_AO6;
  wire [0:0] CLBLM_L_X12Y104_SLICE_X16Y104_A_CY;
  wire [0:0] CLBLM_L_X12Y104_SLICE_X16Y104_A_XOR;
  wire [0:0] CLBLM_L_X12Y104_SLICE_X16Y104_B;
  wire [0:0] CLBLM_L_X12Y104_SLICE_X16Y104_B1;
  wire [0:0] CLBLM_L_X12Y104_SLICE_X16Y104_B2;
  wire [0:0] CLBLM_L_X12Y104_SLICE_X16Y104_B3;
  wire [0:0] CLBLM_L_X12Y104_SLICE_X16Y104_B4;
  wire [0:0] CLBLM_L_X12Y104_SLICE_X16Y104_B5;
  wire [0:0] CLBLM_L_X12Y104_SLICE_X16Y104_B6;
  wire [0:0] CLBLM_L_X12Y104_SLICE_X16Y104_BO5;
  wire [0:0] CLBLM_L_X12Y104_SLICE_X16Y104_BO6;
  wire [0:0] CLBLM_L_X12Y104_SLICE_X16Y104_B_CY;
  wire [0:0] CLBLM_L_X12Y104_SLICE_X16Y104_B_XOR;
  wire [0:0] CLBLM_L_X12Y104_SLICE_X16Y104_C;
  wire [0:0] CLBLM_L_X12Y104_SLICE_X16Y104_C1;
  wire [0:0] CLBLM_L_X12Y104_SLICE_X16Y104_C2;
  wire [0:0] CLBLM_L_X12Y104_SLICE_X16Y104_C3;
  wire [0:0] CLBLM_L_X12Y104_SLICE_X16Y104_C4;
  wire [0:0] CLBLM_L_X12Y104_SLICE_X16Y104_C5;
  wire [0:0] CLBLM_L_X12Y104_SLICE_X16Y104_C6;
  wire [0:0] CLBLM_L_X12Y104_SLICE_X16Y104_CO5;
  wire [0:0] CLBLM_L_X12Y104_SLICE_X16Y104_CO6;
  wire [0:0] CLBLM_L_X12Y104_SLICE_X16Y104_C_CY;
  wire [0:0] CLBLM_L_X12Y104_SLICE_X16Y104_C_XOR;
  wire [0:0] CLBLM_L_X12Y104_SLICE_X16Y104_D;
  wire [0:0] CLBLM_L_X12Y104_SLICE_X16Y104_D1;
  wire [0:0] CLBLM_L_X12Y104_SLICE_X16Y104_D2;
  wire [0:0] CLBLM_L_X12Y104_SLICE_X16Y104_D3;
  wire [0:0] CLBLM_L_X12Y104_SLICE_X16Y104_D4;
  wire [0:0] CLBLM_L_X12Y104_SLICE_X16Y104_D5;
  wire [0:0] CLBLM_L_X12Y104_SLICE_X16Y104_D6;
  wire [0:0] CLBLM_L_X12Y104_SLICE_X16Y104_DO5;
  wire [0:0] CLBLM_L_X12Y104_SLICE_X16Y104_DO6;
  wire [0:0] CLBLM_L_X12Y104_SLICE_X16Y104_D_CY;
  wire [0:0] CLBLM_L_X12Y104_SLICE_X16Y104_D_XOR;
  wire [0:0] CLBLM_L_X12Y104_SLICE_X17Y104_A;
  wire [0:0] CLBLM_L_X12Y104_SLICE_X17Y104_A1;
  wire [0:0] CLBLM_L_X12Y104_SLICE_X17Y104_A2;
  wire [0:0] CLBLM_L_X12Y104_SLICE_X17Y104_A3;
  wire [0:0] CLBLM_L_X12Y104_SLICE_X17Y104_A4;
  wire [0:0] CLBLM_L_X12Y104_SLICE_X17Y104_A5;
  wire [0:0] CLBLM_L_X12Y104_SLICE_X17Y104_A6;
  wire [0:0] CLBLM_L_X12Y104_SLICE_X17Y104_AO5;
  wire [0:0] CLBLM_L_X12Y104_SLICE_X17Y104_AO6;
  wire [0:0] CLBLM_L_X12Y104_SLICE_X17Y104_A_CY;
  wire [0:0] CLBLM_L_X12Y104_SLICE_X17Y104_A_XOR;
  wire [0:0] CLBLM_L_X12Y104_SLICE_X17Y104_B;
  wire [0:0] CLBLM_L_X12Y104_SLICE_X17Y104_B1;
  wire [0:0] CLBLM_L_X12Y104_SLICE_X17Y104_B2;
  wire [0:0] CLBLM_L_X12Y104_SLICE_X17Y104_B3;
  wire [0:0] CLBLM_L_X12Y104_SLICE_X17Y104_B4;
  wire [0:0] CLBLM_L_X12Y104_SLICE_X17Y104_B5;
  wire [0:0] CLBLM_L_X12Y104_SLICE_X17Y104_B6;
  wire [0:0] CLBLM_L_X12Y104_SLICE_X17Y104_BO5;
  wire [0:0] CLBLM_L_X12Y104_SLICE_X17Y104_BO6;
  wire [0:0] CLBLM_L_X12Y104_SLICE_X17Y104_B_CY;
  wire [0:0] CLBLM_L_X12Y104_SLICE_X17Y104_B_XOR;
  wire [0:0] CLBLM_L_X12Y104_SLICE_X17Y104_C;
  wire [0:0] CLBLM_L_X12Y104_SLICE_X17Y104_C1;
  wire [0:0] CLBLM_L_X12Y104_SLICE_X17Y104_C2;
  wire [0:0] CLBLM_L_X12Y104_SLICE_X17Y104_C3;
  wire [0:0] CLBLM_L_X12Y104_SLICE_X17Y104_C4;
  wire [0:0] CLBLM_L_X12Y104_SLICE_X17Y104_C5;
  wire [0:0] CLBLM_L_X12Y104_SLICE_X17Y104_C6;
  wire [0:0] CLBLM_L_X12Y104_SLICE_X17Y104_CO5;
  wire [0:0] CLBLM_L_X12Y104_SLICE_X17Y104_CO6;
  wire [0:0] CLBLM_L_X12Y104_SLICE_X17Y104_C_CY;
  wire [0:0] CLBLM_L_X12Y104_SLICE_X17Y104_C_XOR;
  wire [0:0] CLBLM_L_X12Y104_SLICE_X17Y104_D;
  wire [0:0] CLBLM_L_X12Y104_SLICE_X17Y104_D1;
  wire [0:0] CLBLM_L_X12Y104_SLICE_X17Y104_D2;
  wire [0:0] CLBLM_L_X12Y104_SLICE_X17Y104_D3;
  wire [0:0] CLBLM_L_X12Y104_SLICE_X17Y104_D4;
  wire [0:0] CLBLM_L_X12Y104_SLICE_X17Y104_D5;
  wire [0:0] CLBLM_L_X12Y104_SLICE_X17Y104_D6;
  wire [0:0] CLBLM_L_X12Y104_SLICE_X17Y104_DO5;
  wire [0:0] CLBLM_L_X12Y104_SLICE_X17Y104_DO6;
  wire [0:0] CLBLM_L_X12Y104_SLICE_X17Y104_D_CY;
  wire [0:0] CLBLM_L_X12Y104_SLICE_X17Y104_D_XOR;
  wire [0:0] CLBLM_L_X12Y105_SLICE_X16Y105_A;
  wire [0:0] CLBLM_L_X12Y105_SLICE_X16Y105_A1;
  wire [0:0] CLBLM_L_X12Y105_SLICE_X16Y105_A2;
  wire [0:0] CLBLM_L_X12Y105_SLICE_X16Y105_A3;
  wire [0:0] CLBLM_L_X12Y105_SLICE_X16Y105_A4;
  wire [0:0] CLBLM_L_X12Y105_SLICE_X16Y105_A5;
  wire [0:0] CLBLM_L_X12Y105_SLICE_X16Y105_A6;
  wire [0:0] CLBLM_L_X12Y105_SLICE_X16Y105_AMUX;
  wire [0:0] CLBLM_L_X12Y105_SLICE_X16Y105_AO5;
  wire [0:0] CLBLM_L_X12Y105_SLICE_X16Y105_AO6;
  wire [0:0] CLBLM_L_X12Y105_SLICE_X16Y105_A_CY;
  wire [0:0] CLBLM_L_X12Y105_SLICE_X16Y105_A_XOR;
  wire [0:0] CLBLM_L_X12Y105_SLICE_X16Y105_B;
  wire [0:0] CLBLM_L_X12Y105_SLICE_X16Y105_B1;
  wire [0:0] CLBLM_L_X12Y105_SLICE_X16Y105_B2;
  wire [0:0] CLBLM_L_X12Y105_SLICE_X16Y105_B3;
  wire [0:0] CLBLM_L_X12Y105_SLICE_X16Y105_B4;
  wire [0:0] CLBLM_L_X12Y105_SLICE_X16Y105_B5;
  wire [0:0] CLBLM_L_X12Y105_SLICE_X16Y105_B6;
  wire [0:0] CLBLM_L_X12Y105_SLICE_X16Y105_BO5;
  wire [0:0] CLBLM_L_X12Y105_SLICE_X16Y105_BO6;
  wire [0:0] CLBLM_L_X12Y105_SLICE_X16Y105_B_CY;
  wire [0:0] CLBLM_L_X12Y105_SLICE_X16Y105_B_XOR;
  wire [0:0] CLBLM_L_X12Y105_SLICE_X16Y105_C;
  wire [0:0] CLBLM_L_X12Y105_SLICE_X16Y105_C1;
  wire [0:0] CLBLM_L_X12Y105_SLICE_X16Y105_C2;
  wire [0:0] CLBLM_L_X12Y105_SLICE_X16Y105_C3;
  wire [0:0] CLBLM_L_X12Y105_SLICE_X16Y105_C4;
  wire [0:0] CLBLM_L_X12Y105_SLICE_X16Y105_C5;
  wire [0:0] CLBLM_L_X12Y105_SLICE_X16Y105_C6;
  wire [0:0] CLBLM_L_X12Y105_SLICE_X16Y105_CO5;
  wire [0:0] CLBLM_L_X12Y105_SLICE_X16Y105_CO6;
  wire [0:0] CLBLM_L_X12Y105_SLICE_X16Y105_C_CY;
  wire [0:0] CLBLM_L_X12Y105_SLICE_X16Y105_C_XOR;
  wire [0:0] CLBLM_L_X12Y105_SLICE_X16Y105_D;
  wire [0:0] CLBLM_L_X12Y105_SLICE_X16Y105_D1;
  wire [0:0] CLBLM_L_X12Y105_SLICE_X16Y105_D2;
  wire [0:0] CLBLM_L_X12Y105_SLICE_X16Y105_D3;
  wire [0:0] CLBLM_L_X12Y105_SLICE_X16Y105_D4;
  wire [0:0] CLBLM_L_X12Y105_SLICE_X16Y105_D5;
  wire [0:0] CLBLM_L_X12Y105_SLICE_X16Y105_D6;
  wire [0:0] CLBLM_L_X12Y105_SLICE_X16Y105_DO5;
  wire [0:0] CLBLM_L_X12Y105_SLICE_X16Y105_DO6;
  wire [0:0] CLBLM_L_X12Y105_SLICE_X16Y105_D_CY;
  wire [0:0] CLBLM_L_X12Y105_SLICE_X16Y105_D_XOR;
  wire [0:0] CLBLM_L_X12Y105_SLICE_X17Y105_A;
  wire [0:0] CLBLM_L_X12Y105_SLICE_X17Y105_A1;
  wire [0:0] CLBLM_L_X12Y105_SLICE_X17Y105_A2;
  wire [0:0] CLBLM_L_X12Y105_SLICE_X17Y105_A3;
  wire [0:0] CLBLM_L_X12Y105_SLICE_X17Y105_A4;
  wire [0:0] CLBLM_L_X12Y105_SLICE_X17Y105_A5;
  wire [0:0] CLBLM_L_X12Y105_SLICE_X17Y105_A6;
  wire [0:0] CLBLM_L_X12Y105_SLICE_X17Y105_AO5;
  wire [0:0] CLBLM_L_X12Y105_SLICE_X17Y105_AO6;
  wire [0:0] CLBLM_L_X12Y105_SLICE_X17Y105_A_CY;
  wire [0:0] CLBLM_L_X12Y105_SLICE_X17Y105_A_XOR;
  wire [0:0] CLBLM_L_X12Y105_SLICE_X17Y105_B;
  wire [0:0] CLBLM_L_X12Y105_SLICE_X17Y105_B1;
  wire [0:0] CLBLM_L_X12Y105_SLICE_X17Y105_B2;
  wire [0:0] CLBLM_L_X12Y105_SLICE_X17Y105_B3;
  wire [0:0] CLBLM_L_X12Y105_SLICE_X17Y105_B4;
  wire [0:0] CLBLM_L_X12Y105_SLICE_X17Y105_B5;
  wire [0:0] CLBLM_L_X12Y105_SLICE_X17Y105_B6;
  wire [0:0] CLBLM_L_X12Y105_SLICE_X17Y105_BO5;
  wire [0:0] CLBLM_L_X12Y105_SLICE_X17Y105_BO6;
  wire [0:0] CLBLM_L_X12Y105_SLICE_X17Y105_B_CY;
  wire [0:0] CLBLM_L_X12Y105_SLICE_X17Y105_B_XOR;
  wire [0:0] CLBLM_L_X12Y105_SLICE_X17Y105_C;
  wire [0:0] CLBLM_L_X12Y105_SLICE_X17Y105_C1;
  wire [0:0] CLBLM_L_X12Y105_SLICE_X17Y105_C2;
  wire [0:0] CLBLM_L_X12Y105_SLICE_X17Y105_C3;
  wire [0:0] CLBLM_L_X12Y105_SLICE_X17Y105_C4;
  wire [0:0] CLBLM_L_X12Y105_SLICE_X17Y105_C5;
  wire [0:0] CLBLM_L_X12Y105_SLICE_X17Y105_C6;
  wire [0:0] CLBLM_L_X12Y105_SLICE_X17Y105_CO5;
  wire [0:0] CLBLM_L_X12Y105_SLICE_X17Y105_CO6;
  wire [0:0] CLBLM_L_X12Y105_SLICE_X17Y105_C_CY;
  wire [0:0] CLBLM_L_X12Y105_SLICE_X17Y105_C_XOR;
  wire [0:0] CLBLM_L_X12Y105_SLICE_X17Y105_D;
  wire [0:0] CLBLM_L_X12Y105_SLICE_X17Y105_D1;
  wire [0:0] CLBLM_L_X12Y105_SLICE_X17Y105_D2;
  wire [0:0] CLBLM_L_X12Y105_SLICE_X17Y105_D3;
  wire [0:0] CLBLM_L_X12Y105_SLICE_X17Y105_D4;
  wire [0:0] CLBLM_L_X12Y105_SLICE_X17Y105_D5;
  wire [0:0] CLBLM_L_X12Y105_SLICE_X17Y105_D6;
  wire [0:0] CLBLM_L_X12Y105_SLICE_X17Y105_DO5;
  wire [0:0] CLBLM_L_X12Y105_SLICE_X17Y105_DO6;
  wire [0:0] CLBLM_L_X12Y105_SLICE_X17Y105_D_CY;
  wire [0:0] CLBLM_L_X12Y105_SLICE_X17Y105_D_XOR;
  wire [0:0] CLBLM_L_X12Y106_SLICE_X16Y106_A;
  wire [0:0] CLBLM_L_X12Y106_SLICE_X16Y106_A1;
  wire [0:0] CLBLM_L_X12Y106_SLICE_X16Y106_A2;
  wire [0:0] CLBLM_L_X12Y106_SLICE_X16Y106_A3;
  wire [0:0] CLBLM_L_X12Y106_SLICE_X16Y106_A4;
  wire [0:0] CLBLM_L_X12Y106_SLICE_X16Y106_A5;
  wire [0:0] CLBLM_L_X12Y106_SLICE_X16Y106_A6;
  wire [0:0] CLBLM_L_X12Y106_SLICE_X16Y106_AMUX;
  wire [0:0] CLBLM_L_X12Y106_SLICE_X16Y106_AO5;
  wire [0:0] CLBLM_L_X12Y106_SLICE_X16Y106_AO6;
  wire [0:0] CLBLM_L_X12Y106_SLICE_X16Y106_A_CY;
  wire [0:0] CLBLM_L_X12Y106_SLICE_X16Y106_A_XOR;
  wire [0:0] CLBLM_L_X12Y106_SLICE_X16Y106_B;
  wire [0:0] CLBLM_L_X12Y106_SLICE_X16Y106_B1;
  wire [0:0] CLBLM_L_X12Y106_SLICE_X16Y106_B2;
  wire [0:0] CLBLM_L_X12Y106_SLICE_X16Y106_B3;
  wire [0:0] CLBLM_L_X12Y106_SLICE_X16Y106_B4;
  wire [0:0] CLBLM_L_X12Y106_SLICE_X16Y106_B5;
  wire [0:0] CLBLM_L_X12Y106_SLICE_X16Y106_B6;
  wire [0:0] CLBLM_L_X12Y106_SLICE_X16Y106_BMUX;
  wire [0:0] CLBLM_L_X12Y106_SLICE_X16Y106_BO5;
  wire [0:0] CLBLM_L_X12Y106_SLICE_X16Y106_BO6;
  wire [0:0] CLBLM_L_X12Y106_SLICE_X16Y106_B_CY;
  wire [0:0] CLBLM_L_X12Y106_SLICE_X16Y106_B_XOR;
  wire [0:0] CLBLM_L_X12Y106_SLICE_X16Y106_C;
  wire [0:0] CLBLM_L_X12Y106_SLICE_X16Y106_C1;
  wire [0:0] CLBLM_L_X12Y106_SLICE_X16Y106_C2;
  wire [0:0] CLBLM_L_X12Y106_SLICE_X16Y106_C3;
  wire [0:0] CLBLM_L_X12Y106_SLICE_X16Y106_C4;
  wire [0:0] CLBLM_L_X12Y106_SLICE_X16Y106_C5;
  wire [0:0] CLBLM_L_X12Y106_SLICE_X16Y106_C6;
  wire [0:0] CLBLM_L_X12Y106_SLICE_X16Y106_CO5;
  wire [0:0] CLBLM_L_X12Y106_SLICE_X16Y106_CO6;
  wire [0:0] CLBLM_L_X12Y106_SLICE_X16Y106_C_CY;
  wire [0:0] CLBLM_L_X12Y106_SLICE_X16Y106_C_XOR;
  wire [0:0] CLBLM_L_X12Y106_SLICE_X16Y106_D;
  wire [0:0] CLBLM_L_X12Y106_SLICE_X16Y106_D1;
  wire [0:0] CLBLM_L_X12Y106_SLICE_X16Y106_D2;
  wire [0:0] CLBLM_L_X12Y106_SLICE_X16Y106_D3;
  wire [0:0] CLBLM_L_X12Y106_SLICE_X16Y106_D4;
  wire [0:0] CLBLM_L_X12Y106_SLICE_X16Y106_D5;
  wire [0:0] CLBLM_L_X12Y106_SLICE_X16Y106_D6;
  wire [0:0] CLBLM_L_X12Y106_SLICE_X16Y106_DO5;
  wire [0:0] CLBLM_L_X12Y106_SLICE_X16Y106_DO6;
  wire [0:0] CLBLM_L_X12Y106_SLICE_X16Y106_D_CY;
  wire [0:0] CLBLM_L_X12Y106_SLICE_X16Y106_D_XOR;
  wire [0:0] CLBLM_L_X12Y106_SLICE_X17Y106_A;
  wire [0:0] CLBLM_L_X12Y106_SLICE_X17Y106_A1;
  wire [0:0] CLBLM_L_X12Y106_SLICE_X17Y106_A2;
  wire [0:0] CLBLM_L_X12Y106_SLICE_X17Y106_A3;
  wire [0:0] CLBLM_L_X12Y106_SLICE_X17Y106_A4;
  wire [0:0] CLBLM_L_X12Y106_SLICE_X17Y106_A5;
  wire [0:0] CLBLM_L_X12Y106_SLICE_X17Y106_A6;
  wire [0:0] CLBLM_L_X12Y106_SLICE_X17Y106_AMUX;
  wire [0:0] CLBLM_L_X12Y106_SLICE_X17Y106_AO5;
  wire [0:0] CLBLM_L_X12Y106_SLICE_X17Y106_AO6;
  wire [0:0] CLBLM_L_X12Y106_SLICE_X17Y106_A_CY;
  wire [0:0] CLBLM_L_X12Y106_SLICE_X17Y106_A_XOR;
  wire [0:0] CLBLM_L_X12Y106_SLICE_X17Y106_B;
  wire [0:0] CLBLM_L_X12Y106_SLICE_X17Y106_B1;
  wire [0:0] CLBLM_L_X12Y106_SLICE_X17Y106_B2;
  wire [0:0] CLBLM_L_X12Y106_SLICE_X17Y106_B3;
  wire [0:0] CLBLM_L_X12Y106_SLICE_X17Y106_B4;
  wire [0:0] CLBLM_L_X12Y106_SLICE_X17Y106_B5;
  wire [0:0] CLBLM_L_X12Y106_SLICE_X17Y106_B6;
  wire [0:0] CLBLM_L_X12Y106_SLICE_X17Y106_BO5;
  wire [0:0] CLBLM_L_X12Y106_SLICE_X17Y106_BO6;
  wire [0:0] CLBLM_L_X12Y106_SLICE_X17Y106_B_CY;
  wire [0:0] CLBLM_L_X12Y106_SLICE_X17Y106_B_XOR;
  wire [0:0] CLBLM_L_X12Y106_SLICE_X17Y106_C;
  wire [0:0] CLBLM_L_X12Y106_SLICE_X17Y106_C1;
  wire [0:0] CLBLM_L_X12Y106_SLICE_X17Y106_C2;
  wire [0:0] CLBLM_L_X12Y106_SLICE_X17Y106_C3;
  wire [0:0] CLBLM_L_X12Y106_SLICE_X17Y106_C4;
  wire [0:0] CLBLM_L_X12Y106_SLICE_X17Y106_C5;
  wire [0:0] CLBLM_L_X12Y106_SLICE_X17Y106_C6;
  wire [0:0] CLBLM_L_X12Y106_SLICE_X17Y106_CO5;
  wire [0:0] CLBLM_L_X12Y106_SLICE_X17Y106_CO6;
  wire [0:0] CLBLM_L_X12Y106_SLICE_X17Y106_C_CY;
  wire [0:0] CLBLM_L_X12Y106_SLICE_X17Y106_C_XOR;
  wire [0:0] CLBLM_L_X12Y106_SLICE_X17Y106_D;
  wire [0:0] CLBLM_L_X12Y106_SLICE_X17Y106_D1;
  wire [0:0] CLBLM_L_X12Y106_SLICE_X17Y106_D2;
  wire [0:0] CLBLM_L_X12Y106_SLICE_X17Y106_D3;
  wire [0:0] CLBLM_L_X12Y106_SLICE_X17Y106_D4;
  wire [0:0] CLBLM_L_X12Y106_SLICE_X17Y106_D5;
  wire [0:0] CLBLM_L_X12Y106_SLICE_X17Y106_D6;
  wire [0:0] CLBLM_L_X12Y106_SLICE_X17Y106_DO5;
  wire [0:0] CLBLM_L_X12Y106_SLICE_X17Y106_DO6;
  wire [0:0] CLBLM_L_X12Y106_SLICE_X17Y106_D_CY;
  wire [0:0] CLBLM_L_X12Y106_SLICE_X17Y106_D_XOR;
  wire [0:0] CLBLM_L_X12Y107_SLICE_X16Y107_A;
  wire [0:0] CLBLM_L_X12Y107_SLICE_X16Y107_A1;
  wire [0:0] CLBLM_L_X12Y107_SLICE_X16Y107_A2;
  wire [0:0] CLBLM_L_X12Y107_SLICE_X16Y107_A3;
  wire [0:0] CLBLM_L_X12Y107_SLICE_X16Y107_A4;
  wire [0:0] CLBLM_L_X12Y107_SLICE_X16Y107_A5;
  wire [0:0] CLBLM_L_X12Y107_SLICE_X16Y107_A6;
  wire [0:0] CLBLM_L_X12Y107_SLICE_X16Y107_AO5;
  wire [0:0] CLBLM_L_X12Y107_SLICE_X16Y107_AO6;
  wire [0:0] CLBLM_L_X12Y107_SLICE_X16Y107_A_CY;
  wire [0:0] CLBLM_L_X12Y107_SLICE_X16Y107_A_XOR;
  wire [0:0] CLBLM_L_X12Y107_SLICE_X16Y107_B;
  wire [0:0] CLBLM_L_X12Y107_SLICE_X16Y107_B1;
  wire [0:0] CLBLM_L_X12Y107_SLICE_X16Y107_B2;
  wire [0:0] CLBLM_L_X12Y107_SLICE_X16Y107_B3;
  wire [0:0] CLBLM_L_X12Y107_SLICE_X16Y107_B4;
  wire [0:0] CLBLM_L_X12Y107_SLICE_X16Y107_B5;
  wire [0:0] CLBLM_L_X12Y107_SLICE_X16Y107_B6;
  wire [0:0] CLBLM_L_X12Y107_SLICE_X16Y107_BO5;
  wire [0:0] CLBLM_L_X12Y107_SLICE_X16Y107_BO6;
  wire [0:0] CLBLM_L_X12Y107_SLICE_X16Y107_B_CY;
  wire [0:0] CLBLM_L_X12Y107_SLICE_X16Y107_B_XOR;
  wire [0:0] CLBLM_L_X12Y107_SLICE_X16Y107_C;
  wire [0:0] CLBLM_L_X12Y107_SLICE_X16Y107_C1;
  wire [0:0] CLBLM_L_X12Y107_SLICE_X16Y107_C2;
  wire [0:0] CLBLM_L_X12Y107_SLICE_X16Y107_C3;
  wire [0:0] CLBLM_L_X12Y107_SLICE_X16Y107_C4;
  wire [0:0] CLBLM_L_X12Y107_SLICE_X16Y107_C5;
  wire [0:0] CLBLM_L_X12Y107_SLICE_X16Y107_C6;
  wire [0:0] CLBLM_L_X12Y107_SLICE_X16Y107_CO5;
  wire [0:0] CLBLM_L_X12Y107_SLICE_X16Y107_CO6;
  wire [0:0] CLBLM_L_X12Y107_SLICE_X16Y107_C_CY;
  wire [0:0] CLBLM_L_X12Y107_SLICE_X16Y107_C_XOR;
  wire [0:0] CLBLM_L_X12Y107_SLICE_X16Y107_D;
  wire [0:0] CLBLM_L_X12Y107_SLICE_X16Y107_D1;
  wire [0:0] CLBLM_L_X12Y107_SLICE_X16Y107_D2;
  wire [0:0] CLBLM_L_X12Y107_SLICE_X16Y107_D3;
  wire [0:0] CLBLM_L_X12Y107_SLICE_X16Y107_D4;
  wire [0:0] CLBLM_L_X12Y107_SLICE_X16Y107_D5;
  wire [0:0] CLBLM_L_X12Y107_SLICE_X16Y107_D6;
  wire [0:0] CLBLM_L_X12Y107_SLICE_X16Y107_DO5;
  wire [0:0] CLBLM_L_X12Y107_SLICE_X16Y107_DO6;
  wire [0:0] CLBLM_L_X12Y107_SLICE_X16Y107_D_CY;
  wire [0:0] CLBLM_L_X12Y107_SLICE_X16Y107_D_XOR;
  wire [0:0] CLBLM_L_X12Y107_SLICE_X17Y107_A;
  wire [0:0] CLBLM_L_X12Y107_SLICE_X17Y107_A1;
  wire [0:0] CLBLM_L_X12Y107_SLICE_X17Y107_A2;
  wire [0:0] CLBLM_L_X12Y107_SLICE_X17Y107_A3;
  wire [0:0] CLBLM_L_X12Y107_SLICE_X17Y107_A4;
  wire [0:0] CLBLM_L_X12Y107_SLICE_X17Y107_A5;
  wire [0:0] CLBLM_L_X12Y107_SLICE_X17Y107_A6;
  wire [0:0] CLBLM_L_X12Y107_SLICE_X17Y107_AMUX;
  wire [0:0] CLBLM_L_X12Y107_SLICE_X17Y107_AO5;
  wire [0:0] CLBLM_L_X12Y107_SLICE_X17Y107_AO6;
  wire [0:0] CLBLM_L_X12Y107_SLICE_X17Y107_A_CY;
  wire [0:0] CLBLM_L_X12Y107_SLICE_X17Y107_A_XOR;
  wire [0:0] CLBLM_L_X12Y107_SLICE_X17Y107_B;
  wire [0:0] CLBLM_L_X12Y107_SLICE_X17Y107_B1;
  wire [0:0] CLBLM_L_X12Y107_SLICE_X17Y107_B2;
  wire [0:0] CLBLM_L_X12Y107_SLICE_X17Y107_B3;
  wire [0:0] CLBLM_L_X12Y107_SLICE_X17Y107_B4;
  wire [0:0] CLBLM_L_X12Y107_SLICE_X17Y107_B5;
  wire [0:0] CLBLM_L_X12Y107_SLICE_X17Y107_B6;
  wire [0:0] CLBLM_L_X12Y107_SLICE_X17Y107_BO5;
  wire [0:0] CLBLM_L_X12Y107_SLICE_X17Y107_BO6;
  wire [0:0] CLBLM_L_X12Y107_SLICE_X17Y107_B_CY;
  wire [0:0] CLBLM_L_X12Y107_SLICE_X17Y107_B_XOR;
  wire [0:0] CLBLM_L_X12Y107_SLICE_X17Y107_C;
  wire [0:0] CLBLM_L_X12Y107_SLICE_X17Y107_C1;
  wire [0:0] CLBLM_L_X12Y107_SLICE_X17Y107_C2;
  wire [0:0] CLBLM_L_X12Y107_SLICE_X17Y107_C3;
  wire [0:0] CLBLM_L_X12Y107_SLICE_X17Y107_C4;
  wire [0:0] CLBLM_L_X12Y107_SLICE_X17Y107_C5;
  wire [0:0] CLBLM_L_X12Y107_SLICE_X17Y107_C6;
  wire [0:0] CLBLM_L_X12Y107_SLICE_X17Y107_CO5;
  wire [0:0] CLBLM_L_X12Y107_SLICE_X17Y107_CO6;
  wire [0:0] CLBLM_L_X12Y107_SLICE_X17Y107_C_CY;
  wire [0:0] CLBLM_L_X12Y107_SLICE_X17Y107_C_XOR;
  wire [0:0] CLBLM_L_X12Y107_SLICE_X17Y107_D;
  wire [0:0] CLBLM_L_X12Y107_SLICE_X17Y107_D1;
  wire [0:0] CLBLM_L_X12Y107_SLICE_X17Y107_D2;
  wire [0:0] CLBLM_L_X12Y107_SLICE_X17Y107_D3;
  wire [0:0] CLBLM_L_X12Y107_SLICE_X17Y107_D4;
  wire [0:0] CLBLM_L_X12Y107_SLICE_X17Y107_D5;
  wire [0:0] CLBLM_L_X12Y107_SLICE_X17Y107_D6;
  wire [0:0] CLBLM_L_X12Y107_SLICE_X17Y107_DO5;
  wire [0:0] CLBLM_L_X12Y107_SLICE_X17Y107_DO6;
  wire [0:0] CLBLM_L_X12Y107_SLICE_X17Y107_D_CY;
  wire [0:0] CLBLM_L_X12Y107_SLICE_X17Y107_D_XOR;
  wire [0:0] CLBLM_L_X12Y108_SLICE_X16Y108_A;
  wire [0:0] CLBLM_L_X12Y108_SLICE_X16Y108_A1;
  wire [0:0] CLBLM_L_X12Y108_SLICE_X16Y108_A2;
  wire [0:0] CLBLM_L_X12Y108_SLICE_X16Y108_A3;
  wire [0:0] CLBLM_L_X12Y108_SLICE_X16Y108_A4;
  wire [0:0] CLBLM_L_X12Y108_SLICE_X16Y108_A5;
  wire [0:0] CLBLM_L_X12Y108_SLICE_X16Y108_A6;
  wire [0:0] CLBLM_L_X12Y108_SLICE_X16Y108_AMUX;
  wire [0:0] CLBLM_L_X12Y108_SLICE_X16Y108_AO5;
  wire [0:0] CLBLM_L_X12Y108_SLICE_X16Y108_AO6;
  wire [0:0] CLBLM_L_X12Y108_SLICE_X16Y108_A_CY;
  wire [0:0] CLBLM_L_X12Y108_SLICE_X16Y108_A_XOR;
  wire [0:0] CLBLM_L_X12Y108_SLICE_X16Y108_B;
  wire [0:0] CLBLM_L_X12Y108_SLICE_X16Y108_B1;
  wire [0:0] CLBLM_L_X12Y108_SLICE_X16Y108_B2;
  wire [0:0] CLBLM_L_X12Y108_SLICE_X16Y108_B3;
  wire [0:0] CLBLM_L_X12Y108_SLICE_X16Y108_B4;
  wire [0:0] CLBLM_L_X12Y108_SLICE_X16Y108_B5;
  wire [0:0] CLBLM_L_X12Y108_SLICE_X16Y108_B6;
  wire [0:0] CLBLM_L_X12Y108_SLICE_X16Y108_BO5;
  wire [0:0] CLBLM_L_X12Y108_SLICE_X16Y108_BO6;
  wire [0:0] CLBLM_L_X12Y108_SLICE_X16Y108_B_CY;
  wire [0:0] CLBLM_L_X12Y108_SLICE_X16Y108_B_XOR;
  wire [0:0] CLBLM_L_X12Y108_SLICE_X16Y108_C;
  wire [0:0] CLBLM_L_X12Y108_SLICE_X16Y108_C1;
  wire [0:0] CLBLM_L_X12Y108_SLICE_X16Y108_C2;
  wire [0:0] CLBLM_L_X12Y108_SLICE_X16Y108_C3;
  wire [0:0] CLBLM_L_X12Y108_SLICE_X16Y108_C4;
  wire [0:0] CLBLM_L_X12Y108_SLICE_X16Y108_C5;
  wire [0:0] CLBLM_L_X12Y108_SLICE_X16Y108_C6;
  wire [0:0] CLBLM_L_X12Y108_SLICE_X16Y108_CO5;
  wire [0:0] CLBLM_L_X12Y108_SLICE_X16Y108_CO6;
  wire [0:0] CLBLM_L_X12Y108_SLICE_X16Y108_C_CY;
  wire [0:0] CLBLM_L_X12Y108_SLICE_X16Y108_C_XOR;
  wire [0:0] CLBLM_L_X12Y108_SLICE_X16Y108_D;
  wire [0:0] CLBLM_L_X12Y108_SLICE_X16Y108_D1;
  wire [0:0] CLBLM_L_X12Y108_SLICE_X16Y108_D2;
  wire [0:0] CLBLM_L_X12Y108_SLICE_X16Y108_D3;
  wire [0:0] CLBLM_L_X12Y108_SLICE_X16Y108_D4;
  wire [0:0] CLBLM_L_X12Y108_SLICE_X16Y108_D5;
  wire [0:0] CLBLM_L_X12Y108_SLICE_X16Y108_D6;
  wire [0:0] CLBLM_L_X12Y108_SLICE_X16Y108_DO5;
  wire [0:0] CLBLM_L_X12Y108_SLICE_X16Y108_DO6;
  wire [0:0] CLBLM_L_X12Y108_SLICE_X16Y108_D_CY;
  wire [0:0] CLBLM_L_X12Y108_SLICE_X16Y108_D_XOR;
  wire [0:0] CLBLM_L_X12Y108_SLICE_X17Y108_A;
  wire [0:0] CLBLM_L_X12Y108_SLICE_X17Y108_A1;
  wire [0:0] CLBLM_L_X12Y108_SLICE_X17Y108_A2;
  wire [0:0] CLBLM_L_X12Y108_SLICE_X17Y108_A3;
  wire [0:0] CLBLM_L_X12Y108_SLICE_X17Y108_A4;
  wire [0:0] CLBLM_L_X12Y108_SLICE_X17Y108_A5;
  wire [0:0] CLBLM_L_X12Y108_SLICE_X17Y108_A6;
  wire [0:0] CLBLM_L_X12Y108_SLICE_X17Y108_AO5;
  wire [0:0] CLBLM_L_X12Y108_SLICE_X17Y108_AO6;
  wire [0:0] CLBLM_L_X12Y108_SLICE_X17Y108_A_CY;
  wire [0:0] CLBLM_L_X12Y108_SLICE_X17Y108_A_XOR;
  wire [0:0] CLBLM_L_X12Y108_SLICE_X17Y108_B;
  wire [0:0] CLBLM_L_X12Y108_SLICE_X17Y108_B1;
  wire [0:0] CLBLM_L_X12Y108_SLICE_X17Y108_B2;
  wire [0:0] CLBLM_L_X12Y108_SLICE_X17Y108_B3;
  wire [0:0] CLBLM_L_X12Y108_SLICE_X17Y108_B4;
  wire [0:0] CLBLM_L_X12Y108_SLICE_X17Y108_B5;
  wire [0:0] CLBLM_L_X12Y108_SLICE_X17Y108_B6;
  wire [0:0] CLBLM_L_X12Y108_SLICE_X17Y108_BO5;
  wire [0:0] CLBLM_L_X12Y108_SLICE_X17Y108_BO6;
  wire [0:0] CLBLM_L_X12Y108_SLICE_X17Y108_B_CY;
  wire [0:0] CLBLM_L_X12Y108_SLICE_X17Y108_B_XOR;
  wire [0:0] CLBLM_L_X12Y108_SLICE_X17Y108_C;
  wire [0:0] CLBLM_L_X12Y108_SLICE_X17Y108_C1;
  wire [0:0] CLBLM_L_X12Y108_SLICE_X17Y108_C2;
  wire [0:0] CLBLM_L_X12Y108_SLICE_X17Y108_C3;
  wire [0:0] CLBLM_L_X12Y108_SLICE_X17Y108_C4;
  wire [0:0] CLBLM_L_X12Y108_SLICE_X17Y108_C5;
  wire [0:0] CLBLM_L_X12Y108_SLICE_X17Y108_C6;
  wire [0:0] CLBLM_L_X12Y108_SLICE_X17Y108_CO5;
  wire [0:0] CLBLM_L_X12Y108_SLICE_X17Y108_CO6;
  wire [0:0] CLBLM_L_X12Y108_SLICE_X17Y108_C_CY;
  wire [0:0] CLBLM_L_X12Y108_SLICE_X17Y108_C_XOR;
  wire [0:0] CLBLM_L_X12Y108_SLICE_X17Y108_D;
  wire [0:0] CLBLM_L_X12Y108_SLICE_X17Y108_D1;
  wire [0:0] CLBLM_L_X12Y108_SLICE_X17Y108_D2;
  wire [0:0] CLBLM_L_X12Y108_SLICE_X17Y108_D3;
  wire [0:0] CLBLM_L_X12Y108_SLICE_X17Y108_D4;
  wire [0:0] CLBLM_L_X12Y108_SLICE_X17Y108_D5;
  wire [0:0] CLBLM_L_X12Y108_SLICE_X17Y108_D6;
  wire [0:0] CLBLM_L_X12Y108_SLICE_X17Y108_DO5;
  wire [0:0] CLBLM_L_X12Y108_SLICE_X17Y108_DO6;
  wire [0:0] CLBLM_L_X12Y108_SLICE_X17Y108_D_CY;
  wire [0:0] CLBLM_L_X12Y108_SLICE_X17Y108_D_XOR;
  wire [0:0] CLBLM_L_X12Y109_SLICE_X16Y109_A;
  wire [0:0] CLBLM_L_X12Y109_SLICE_X16Y109_A1;
  wire [0:0] CLBLM_L_X12Y109_SLICE_X16Y109_A2;
  wire [0:0] CLBLM_L_X12Y109_SLICE_X16Y109_A3;
  wire [0:0] CLBLM_L_X12Y109_SLICE_X16Y109_A4;
  wire [0:0] CLBLM_L_X12Y109_SLICE_X16Y109_A5;
  wire [0:0] CLBLM_L_X12Y109_SLICE_X16Y109_A6;
  wire [0:0] CLBLM_L_X12Y109_SLICE_X16Y109_AMUX;
  wire [0:0] CLBLM_L_X12Y109_SLICE_X16Y109_AO5;
  wire [0:0] CLBLM_L_X12Y109_SLICE_X16Y109_AO6;
  wire [0:0] CLBLM_L_X12Y109_SLICE_X16Y109_A_CY;
  wire [0:0] CLBLM_L_X12Y109_SLICE_X16Y109_A_XOR;
  wire [0:0] CLBLM_L_X12Y109_SLICE_X16Y109_B;
  wire [0:0] CLBLM_L_X12Y109_SLICE_X16Y109_B1;
  wire [0:0] CLBLM_L_X12Y109_SLICE_X16Y109_B2;
  wire [0:0] CLBLM_L_X12Y109_SLICE_X16Y109_B3;
  wire [0:0] CLBLM_L_X12Y109_SLICE_X16Y109_B4;
  wire [0:0] CLBLM_L_X12Y109_SLICE_X16Y109_B5;
  wire [0:0] CLBLM_L_X12Y109_SLICE_X16Y109_B6;
  wire [0:0] CLBLM_L_X12Y109_SLICE_X16Y109_BO5;
  wire [0:0] CLBLM_L_X12Y109_SLICE_X16Y109_BO6;
  wire [0:0] CLBLM_L_X12Y109_SLICE_X16Y109_B_CY;
  wire [0:0] CLBLM_L_X12Y109_SLICE_X16Y109_B_XOR;
  wire [0:0] CLBLM_L_X12Y109_SLICE_X16Y109_C;
  wire [0:0] CLBLM_L_X12Y109_SLICE_X16Y109_C1;
  wire [0:0] CLBLM_L_X12Y109_SLICE_X16Y109_C2;
  wire [0:0] CLBLM_L_X12Y109_SLICE_X16Y109_C3;
  wire [0:0] CLBLM_L_X12Y109_SLICE_X16Y109_C4;
  wire [0:0] CLBLM_L_X12Y109_SLICE_X16Y109_C5;
  wire [0:0] CLBLM_L_X12Y109_SLICE_X16Y109_C6;
  wire [0:0] CLBLM_L_X12Y109_SLICE_X16Y109_CO5;
  wire [0:0] CLBLM_L_X12Y109_SLICE_X16Y109_CO6;
  wire [0:0] CLBLM_L_X12Y109_SLICE_X16Y109_C_CY;
  wire [0:0] CLBLM_L_X12Y109_SLICE_X16Y109_C_XOR;
  wire [0:0] CLBLM_L_X12Y109_SLICE_X16Y109_D;
  wire [0:0] CLBLM_L_X12Y109_SLICE_X16Y109_D1;
  wire [0:0] CLBLM_L_X12Y109_SLICE_X16Y109_D2;
  wire [0:0] CLBLM_L_X12Y109_SLICE_X16Y109_D3;
  wire [0:0] CLBLM_L_X12Y109_SLICE_X16Y109_D4;
  wire [0:0] CLBLM_L_X12Y109_SLICE_X16Y109_D5;
  wire [0:0] CLBLM_L_X12Y109_SLICE_X16Y109_D6;
  wire [0:0] CLBLM_L_X12Y109_SLICE_X16Y109_DO5;
  wire [0:0] CLBLM_L_X12Y109_SLICE_X16Y109_DO6;
  wire [0:0] CLBLM_L_X12Y109_SLICE_X16Y109_D_CY;
  wire [0:0] CLBLM_L_X12Y109_SLICE_X16Y109_D_XOR;
  wire [0:0] CLBLM_L_X12Y109_SLICE_X17Y109_A;
  wire [0:0] CLBLM_L_X12Y109_SLICE_X17Y109_A1;
  wire [0:0] CLBLM_L_X12Y109_SLICE_X17Y109_A2;
  wire [0:0] CLBLM_L_X12Y109_SLICE_X17Y109_A3;
  wire [0:0] CLBLM_L_X12Y109_SLICE_X17Y109_A4;
  wire [0:0] CLBLM_L_X12Y109_SLICE_X17Y109_A5;
  wire [0:0] CLBLM_L_X12Y109_SLICE_X17Y109_A6;
  wire [0:0] CLBLM_L_X12Y109_SLICE_X17Y109_AO5;
  wire [0:0] CLBLM_L_X12Y109_SLICE_X17Y109_AO6;
  wire [0:0] CLBLM_L_X12Y109_SLICE_X17Y109_A_CY;
  wire [0:0] CLBLM_L_X12Y109_SLICE_X17Y109_A_XOR;
  wire [0:0] CLBLM_L_X12Y109_SLICE_X17Y109_B;
  wire [0:0] CLBLM_L_X12Y109_SLICE_X17Y109_B1;
  wire [0:0] CLBLM_L_X12Y109_SLICE_X17Y109_B2;
  wire [0:0] CLBLM_L_X12Y109_SLICE_X17Y109_B3;
  wire [0:0] CLBLM_L_X12Y109_SLICE_X17Y109_B4;
  wire [0:0] CLBLM_L_X12Y109_SLICE_X17Y109_B5;
  wire [0:0] CLBLM_L_X12Y109_SLICE_X17Y109_B6;
  wire [0:0] CLBLM_L_X12Y109_SLICE_X17Y109_BMUX;
  wire [0:0] CLBLM_L_X12Y109_SLICE_X17Y109_BO5;
  wire [0:0] CLBLM_L_X12Y109_SLICE_X17Y109_BO6;
  wire [0:0] CLBLM_L_X12Y109_SLICE_X17Y109_B_CY;
  wire [0:0] CLBLM_L_X12Y109_SLICE_X17Y109_B_XOR;
  wire [0:0] CLBLM_L_X12Y109_SLICE_X17Y109_C;
  wire [0:0] CLBLM_L_X12Y109_SLICE_X17Y109_C1;
  wire [0:0] CLBLM_L_X12Y109_SLICE_X17Y109_C2;
  wire [0:0] CLBLM_L_X12Y109_SLICE_X17Y109_C3;
  wire [0:0] CLBLM_L_X12Y109_SLICE_X17Y109_C4;
  wire [0:0] CLBLM_L_X12Y109_SLICE_X17Y109_C5;
  wire [0:0] CLBLM_L_X12Y109_SLICE_X17Y109_C6;
  wire [0:0] CLBLM_L_X12Y109_SLICE_X17Y109_CO5;
  wire [0:0] CLBLM_L_X12Y109_SLICE_X17Y109_CO6;
  wire [0:0] CLBLM_L_X12Y109_SLICE_X17Y109_C_CY;
  wire [0:0] CLBLM_L_X12Y109_SLICE_X17Y109_C_XOR;
  wire [0:0] CLBLM_L_X12Y109_SLICE_X17Y109_D;
  wire [0:0] CLBLM_L_X12Y109_SLICE_X17Y109_D1;
  wire [0:0] CLBLM_L_X12Y109_SLICE_X17Y109_D2;
  wire [0:0] CLBLM_L_X12Y109_SLICE_X17Y109_D3;
  wire [0:0] CLBLM_L_X12Y109_SLICE_X17Y109_D4;
  wire [0:0] CLBLM_L_X12Y109_SLICE_X17Y109_D5;
  wire [0:0] CLBLM_L_X12Y109_SLICE_X17Y109_D6;
  wire [0:0] CLBLM_L_X12Y109_SLICE_X17Y109_DO5;
  wire [0:0] CLBLM_L_X12Y109_SLICE_X17Y109_DO6;
  wire [0:0] CLBLM_L_X12Y109_SLICE_X17Y109_D_CY;
  wire [0:0] CLBLM_L_X12Y109_SLICE_X17Y109_D_XOR;
  wire [0:0] CLBLM_L_X12Y110_SLICE_X16Y110_A;
  wire [0:0] CLBLM_L_X12Y110_SLICE_X16Y110_A1;
  wire [0:0] CLBLM_L_X12Y110_SLICE_X16Y110_A2;
  wire [0:0] CLBLM_L_X12Y110_SLICE_X16Y110_A3;
  wire [0:0] CLBLM_L_X12Y110_SLICE_X16Y110_A4;
  wire [0:0] CLBLM_L_X12Y110_SLICE_X16Y110_A5;
  wire [0:0] CLBLM_L_X12Y110_SLICE_X16Y110_A6;
  wire [0:0] CLBLM_L_X12Y110_SLICE_X16Y110_AMUX;
  wire [0:0] CLBLM_L_X12Y110_SLICE_X16Y110_AO5;
  wire [0:0] CLBLM_L_X12Y110_SLICE_X16Y110_AO6;
  wire [0:0] CLBLM_L_X12Y110_SLICE_X16Y110_A_CY;
  wire [0:0] CLBLM_L_X12Y110_SLICE_X16Y110_A_XOR;
  wire [0:0] CLBLM_L_X12Y110_SLICE_X16Y110_B;
  wire [0:0] CLBLM_L_X12Y110_SLICE_X16Y110_B1;
  wire [0:0] CLBLM_L_X12Y110_SLICE_X16Y110_B2;
  wire [0:0] CLBLM_L_X12Y110_SLICE_X16Y110_B3;
  wire [0:0] CLBLM_L_X12Y110_SLICE_X16Y110_B4;
  wire [0:0] CLBLM_L_X12Y110_SLICE_X16Y110_B5;
  wire [0:0] CLBLM_L_X12Y110_SLICE_X16Y110_B6;
  wire [0:0] CLBLM_L_X12Y110_SLICE_X16Y110_BO5;
  wire [0:0] CLBLM_L_X12Y110_SLICE_X16Y110_BO6;
  wire [0:0] CLBLM_L_X12Y110_SLICE_X16Y110_B_CY;
  wire [0:0] CLBLM_L_X12Y110_SLICE_X16Y110_B_XOR;
  wire [0:0] CLBLM_L_X12Y110_SLICE_X16Y110_C;
  wire [0:0] CLBLM_L_X12Y110_SLICE_X16Y110_C1;
  wire [0:0] CLBLM_L_X12Y110_SLICE_X16Y110_C2;
  wire [0:0] CLBLM_L_X12Y110_SLICE_X16Y110_C3;
  wire [0:0] CLBLM_L_X12Y110_SLICE_X16Y110_C4;
  wire [0:0] CLBLM_L_X12Y110_SLICE_X16Y110_C5;
  wire [0:0] CLBLM_L_X12Y110_SLICE_X16Y110_C6;
  wire [0:0] CLBLM_L_X12Y110_SLICE_X16Y110_CO5;
  wire [0:0] CLBLM_L_X12Y110_SLICE_X16Y110_CO6;
  wire [0:0] CLBLM_L_X12Y110_SLICE_X16Y110_C_CY;
  wire [0:0] CLBLM_L_X12Y110_SLICE_X16Y110_C_XOR;
  wire [0:0] CLBLM_L_X12Y110_SLICE_X16Y110_D;
  wire [0:0] CLBLM_L_X12Y110_SLICE_X16Y110_D1;
  wire [0:0] CLBLM_L_X12Y110_SLICE_X16Y110_D2;
  wire [0:0] CLBLM_L_X12Y110_SLICE_X16Y110_D3;
  wire [0:0] CLBLM_L_X12Y110_SLICE_X16Y110_D4;
  wire [0:0] CLBLM_L_X12Y110_SLICE_X16Y110_D5;
  wire [0:0] CLBLM_L_X12Y110_SLICE_X16Y110_D6;
  wire [0:0] CLBLM_L_X12Y110_SLICE_X16Y110_DO5;
  wire [0:0] CLBLM_L_X12Y110_SLICE_X16Y110_DO6;
  wire [0:0] CLBLM_L_X12Y110_SLICE_X16Y110_D_CY;
  wire [0:0] CLBLM_L_X12Y110_SLICE_X16Y110_D_XOR;
  wire [0:0] CLBLM_L_X12Y110_SLICE_X17Y110_A;
  wire [0:0] CLBLM_L_X12Y110_SLICE_X17Y110_A1;
  wire [0:0] CLBLM_L_X12Y110_SLICE_X17Y110_A2;
  wire [0:0] CLBLM_L_X12Y110_SLICE_X17Y110_A3;
  wire [0:0] CLBLM_L_X12Y110_SLICE_X17Y110_A4;
  wire [0:0] CLBLM_L_X12Y110_SLICE_X17Y110_A5;
  wire [0:0] CLBLM_L_X12Y110_SLICE_X17Y110_A6;
  wire [0:0] CLBLM_L_X12Y110_SLICE_X17Y110_AO5;
  wire [0:0] CLBLM_L_X12Y110_SLICE_X17Y110_AO6;
  wire [0:0] CLBLM_L_X12Y110_SLICE_X17Y110_A_CY;
  wire [0:0] CLBLM_L_X12Y110_SLICE_X17Y110_A_XOR;
  wire [0:0] CLBLM_L_X12Y110_SLICE_X17Y110_B;
  wire [0:0] CLBLM_L_X12Y110_SLICE_X17Y110_B1;
  wire [0:0] CLBLM_L_X12Y110_SLICE_X17Y110_B2;
  wire [0:0] CLBLM_L_X12Y110_SLICE_X17Y110_B3;
  wire [0:0] CLBLM_L_X12Y110_SLICE_X17Y110_B4;
  wire [0:0] CLBLM_L_X12Y110_SLICE_X17Y110_B5;
  wire [0:0] CLBLM_L_X12Y110_SLICE_X17Y110_B6;
  wire [0:0] CLBLM_L_X12Y110_SLICE_X17Y110_BO5;
  wire [0:0] CLBLM_L_X12Y110_SLICE_X17Y110_BO6;
  wire [0:0] CLBLM_L_X12Y110_SLICE_X17Y110_B_CY;
  wire [0:0] CLBLM_L_X12Y110_SLICE_X17Y110_B_XOR;
  wire [0:0] CLBLM_L_X12Y110_SLICE_X17Y110_C;
  wire [0:0] CLBLM_L_X12Y110_SLICE_X17Y110_C1;
  wire [0:0] CLBLM_L_X12Y110_SLICE_X17Y110_C2;
  wire [0:0] CLBLM_L_X12Y110_SLICE_X17Y110_C3;
  wire [0:0] CLBLM_L_X12Y110_SLICE_X17Y110_C4;
  wire [0:0] CLBLM_L_X12Y110_SLICE_X17Y110_C5;
  wire [0:0] CLBLM_L_X12Y110_SLICE_X17Y110_C6;
  wire [0:0] CLBLM_L_X12Y110_SLICE_X17Y110_CO5;
  wire [0:0] CLBLM_L_X12Y110_SLICE_X17Y110_CO6;
  wire [0:0] CLBLM_L_X12Y110_SLICE_X17Y110_C_CY;
  wire [0:0] CLBLM_L_X12Y110_SLICE_X17Y110_C_XOR;
  wire [0:0] CLBLM_L_X12Y110_SLICE_X17Y110_D;
  wire [0:0] CLBLM_L_X12Y110_SLICE_X17Y110_D1;
  wire [0:0] CLBLM_L_X12Y110_SLICE_X17Y110_D2;
  wire [0:0] CLBLM_L_X12Y110_SLICE_X17Y110_D3;
  wire [0:0] CLBLM_L_X12Y110_SLICE_X17Y110_D4;
  wire [0:0] CLBLM_L_X12Y110_SLICE_X17Y110_D5;
  wire [0:0] CLBLM_L_X12Y110_SLICE_X17Y110_D6;
  wire [0:0] CLBLM_L_X12Y110_SLICE_X17Y110_DO5;
  wire [0:0] CLBLM_L_X12Y110_SLICE_X17Y110_DO6;
  wire [0:0] CLBLM_L_X12Y110_SLICE_X17Y110_D_CY;
  wire [0:0] CLBLM_L_X12Y110_SLICE_X17Y110_D_XOR;
  wire [0:0] CLBLM_L_X8Y103_SLICE_X10Y103_A;
  wire [0:0] CLBLM_L_X8Y103_SLICE_X10Y103_A1;
  wire [0:0] CLBLM_L_X8Y103_SLICE_X10Y103_A2;
  wire [0:0] CLBLM_L_X8Y103_SLICE_X10Y103_A3;
  wire [0:0] CLBLM_L_X8Y103_SLICE_X10Y103_A4;
  wire [0:0] CLBLM_L_X8Y103_SLICE_X10Y103_A5;
  wire [0:0] CLBLM_L_X8Y103_SLICE_X10Y103_A6;
  wire [0:0] CLBLM_L_X8Y103_SLICE_X10Y103_AMUX;
  wire [0:0] CLBLM_L_X8Y103_SLICE_X10Y103_AO5;
  wire [0:0] CLBLM_L_X8Y103_SLICE_X10Y103_AO6;
  wire [0:0] CLBLM_L_X8Y103_SLICE_X10Y103_A_CY;
  wire [0:0] CLBLM_L_X8Y103_SLICE_X10Y103_A_XOR;
  wire [0:0] CLBLM_L_X8Y103_SLICE_X10Y103_B;
  wire [0:0] CLBLM_L_X8Y103_SLICE_X10Y103_B1;
  wire [0:0] CLBLM_L_X8Y103_SLICE_X10Y103_B2;
  wire [0:0] CLBLM_L_X8Y103_SLICE_X10Y103_B3;
  wire [0:0] CLBLM_L_X8Y103_SLICE_X10Y103_B4;
  wire [0:0] CLBLM_L_X8Y103_SLICE_X10Y103_B5;
  wire [0:0] CLBLM_L_X8Y103_SLICE_X10Y103_B6;
  wire [0:0] CLBLM_L_X8Y103_SLICE_X10Y103_BO5;
  wire [0:0] CLBLM_L_X8Y103_SLICE_X10Y103_BO6;
  wire [0:0] CLBLM_L_X8Y103_SLICE_X10Y103_B_CY;
  wire [0:0] CLBLM_L_X8Y103_SLICE_X10Y103_B_XOR;
  wire [0:0] CLBLM_L_X8Y103_SLICE_X10Y103_C;
  wire [0:0] CLBLM_L_X8Y103_SLICE_X10Y103_C1;
  wire [0:0] CLBLM_L_X8Y103_SLICE_X10Y103_C2;
  wire [0:0] CLBLM_L_X8Y103_SLICE_X10Y103_C3;
  wire [0:0] CLBLM_L_X8Y103_SLICE_X10Y103_C4;
  wire [0:0] CLBLM_L_X8Y103_SLICE_X10Y103_C5;
  wire [0:0] CLBLM_L_X8Y103_SLICE_X10Y103_C6;
  wire [0:0] CLBLM_L_X8Y103_SLICE_X10Y103_CO5;
  wire [0:0] CLBLM_L_X8Y103_SLICE_X10Y103_CO6;
  wire [0:0] CLBLM_L_X8Y103_SLICE_X10Y103_C_CY;
  wire [0:0] CLBLM_L_X8Y103_SLICE_X10Y103_C_XOR;
  wire [0:0] CLBLM_L_X8Y103_SLICE_X10Y103_D;
  wire [0:0] CLBLM_L_X8Y103_SLICE_X10Y103_D1;
  wire [0:0] CLBLM_L_X8Y103_SLICE_X10Y103_D2;
  wire [0:0] CLBLM_L_X8Y103_SLICE_X10Y103_D3;
  wire [0:0] CLBLM_L_X8Y103_SLICE_X10Y103_D4;
  wire [0:0] CLBLM_L_X8Y103_SLICE_X10Y103_D5;
  wire [0:0] CLBLM_L_X8Y103_SLICE_X10Y103_D6;
  wire [0:0] CLBLM_L_X8Y103_SLICE_X10Y103_DO5;
  wire [0:0] CLBLM_L_X8Y103_SLICE_X10Y103_DO6;
  wire [0:0] CLBLM_L_X8Y103_SLICE_X10Y103_D_CY;
  wire [0:0] CLBLM_L_X8Y103_SLICE_X10Y103_D_XOR;
  wire [0:0] CLBLM_L_X8Y103_SLICE_X11Y103_A;
  wire [0:0] CLBLM_L_X8Y103_SLICE_X11Y103_A1;
  wire [0:0] CLBLM_L_X8Y103_SLICE_X11Y103_A2;
  wire [0:0] CLBLM_L_X8Y103_SLICE_X11Y103_A3;
  wire [0:0] CLBLM_L_X8Y103_SLICE_X11Y103_A4;
  wire [0:0] CLBLM_L_X8Y103_SLICE_X11Y103_A5;
  wire [0:0] CLBLM_L_X8Y103_SLICE_X11Y103_A6;
  wire [0:0] CLBLM_L_X8Y103_SLICE_X11Y103_AMUX;
  wire [0:0] CLBLM_L_X8Y103_SLICE_X11Y103_AO5;
  wire [0:0] CLBLM_L_X8Y103_SLICE_X11Y103_AO6;
  wire [0:0] CLBLM_L_X8Y103_SLICE_X11Y103_A_CY;
  wire [0:0] CLBLM_L_X8Y103_SLICE_X11Y103_A_XOR;
  wire [0:0] CLBLM_L_X8Y103_SLICE_X11Y103_B;
  wire [0:0] CLBLM_L_X8Y103_SLICE_X11Y103_B1;
  wire [0:0] CLBLM_L_X8Y103_SLICE_X11Y103_B2;
  wire [0:0] CLBLM_L_X8Y103_SLICE_X11Y103_B3;
  wire [0:0] CLBLM_L_X8Y103_SLICE_X11Y103_B4;
  wire [0:0] CLBLM_L_X8Y103_SLICE_X11Y103_B5;
  wire [0:0] CLBLM_L_X8Y103_SLICE_X11Y103_B6;
  wire [0:0] CLBLM_L_X8Y103_SLICE_X11Y103_BO5;
  wire [0:0] CLBLM_L_X8Y103_SLICE_X11Y103_BO6;
  wire [0:0] CLBLM_L_X8Y103_SLICE_X11Y103_B_CY;
  wire [0:0] CLBLM_L_X8Y103_SLICE_X11Y103_B_XOR;
  wire [0:0] CLBLM_L_X8Y103_SLICE_X11Y103_C;
  wire [0:0] CLBLM_L_X8Y103_SLICE_X11Y103_C1;
  wire [0:0] CLBLM_L_X8Y103_SLICE_X11Y103_C2;
  wire [0:0] CLBLM_L_X8Y103_SLICE_X11Y103_C3;
  wire [0:0] CLBLM_L_X8Y103_SLICE_X11Y103_C4;
  wire [0:0] CLBLM_L_X8Y103_SLICE_X11Y103_C5;
  wire [0:0] CLBLM_L_X8Y103_SLICE_X11Y103_C6;
  wire [0:0] CLBLM_L_X8Y103_SLICE_X11Y103_CO5;
  wire [0:0] CLBLM_L_X8Y103_SLICE_X11Y103_CO6;
  wire [0:0] CLBLM_L_X8Y103_SLICE_X11Y103_C_CY;
  wire [0:0] CLBLM_L_X8Y103_SLICE_X11Y103_C_XOR;
  wire [0:0] CLBLM_L_X8Y103_SLICE_X11Y103_D;
  wire [0:0] CLBLM_L_X8Y103_SLICE_X11Y103_D1;
  wire [0:0] CLBLM_L_X8Y103_SLICE_X11Y103_D2;
  wire [0:0] CLBLM_L_X8Y103_SLICE_X11Y103_D3;
  wire [0:0] CLBLM_L_X8Y103_SLICE_X11Y103_D4;
  wire [0:0] CLBLM_L_X8Y103_SLICE_X11Y103_D5;
  wire [0:0] CLBLM_L_X8Y103_SLICE_X11Y103_D6;
  wire [0:0] CLBLM_L_X8Y103_SLICE_X11Y103_DO5;
  wire [0:0] CLBLM_L_X8Y103_SLICE_X11Y103_DO6;
  wire [0:0] CLBLM_L_X8Y103_SLICE_X11Y103_D_CY;
  wire [0:0] CLBLM_L_X8Y103_SLICE_X11Y103_D_XOR;
  wire [0:0] CLBLM_L_X8Y104_SLICE_X10Y104_A;
  wire [0:0] CLBLM_L_X8Y104_SLICE_X10Y104_A1;
  wire [0:0] CLBLM_L_X8Y104_SLICE_X10Y104_A2;
  wire [0:0] CLBLM_L_X8Y104_SLICE_X10Y104_A3;
  wire [0:0] CLBLM_L_X8Y104_SLICE_X10Y104_A4;
  wire [0:0] CLBLM_L_X8Y104_SLICE_X10Y104_A5;
  wire [0:0] CLBLM_L_X8Y104_SLICE_X10Y104_A6;
  wire [0:0] CLBLM_L_X8Y104_SLICE_X10Y104_AMUX;
  wire [0:0] CLBLM_L_X8Y104_SLICE_X10Y104_AO5;
  wire [0:0] CLBLM_L_X8Y104_SLICE_X10Y104_AO6;
  wire [0:0] CLBLM_L_X8Y104_SLICE_X10Y104_A_CY;
  wire [0:0] CLBLM_L_X8Y104_SLICE_X10Y104_A_XOR;
  wire [0:0] CLBLM_L_X8Y104_SLICE_X10Y104_B;
  wire [0:0] CLBLM_L_X8Y104_SLICE_X10Y104_B1;
  wire [0:0] CLBLM_L_X8Y104_SLICE_X10Y104_B2;
  wire [0:0] CLBLM_L_X8Y104_SLICE_X10Y104_B3;
  wire [0:0] CLBLM_L_X8Y104_SLICE_X10Y104_B4;
  wire [0:0] CLBLM_L_X8Y104_SLICE_X10Y104_B5;
  wire [0:0] CLBLM_L_X8Y104_SLICE_X10Y104_B6;
  wire [0:0] CLBLM_L_X8Y104_SLICE_X10Y104_BO5;
  wire [0:0] CLBLM_L_X8Y104_SLICE_X10Y104_BO6;
  wire [0:0] CLBLM_L_X8Y104_SLICE_X10Y104_B_CY;
  wire [0:0] CLBLM_L_X8Y104_SLICE_X10Y104_B_XOR;
  wire [0:0] CLBLM_L_X8Y104_SLICE_X10Y104_C;
  wire [0:0] CLBLM_L_X8Y104_SLICE_X10Y104_C1;
  wire [0:0] CLBLM_L_X8Y104_SLICE_X10Y104_C2;
  wire [0:0] CLBLM_L_X8Y104_SLICE_X10Y104_C3;
  wire [0:0] CLBLM_L_X8Y104_SLICE_X10Y104_C4;
  wire [0:0] CLBLM_L_X8Y104_SLICE_X10Y104_C5;
  wire [0:0] CLBLM_L_X8Y104_SLICE_X10Y104_C6;
  wire [0:0] CLBLM_L_X8Y104_SLICE_X10Y104_CMUX;
  wire [0:0] CLBLM_L_X8Y104_SLICE_X10Y104_CO5;
  wire [0:0] CLBLM_L_X8Y104_SLICE_X10Y104_CO6;
  wire [0:0] CLBLM_L_X8Y104_SLICE_X10Y104_C_CY;
  wire [0:0] CLBLM_L_X8Y104_SLICE_X10Y104_C_XOR;
  wire [0:0] CLBLM_L_X8Y104_SLICE_X10Y104_D;
  wire [0:0] CLBLM_L_X8Y104_SLICE_X10Y104_D1;
  wire [0:0] CLBLM_L_X8Y104_SLICE_X10Y104_D2;
  wire [0:0] CLBLM_L_X8Y104_SLICE_X10Y104_D3;
  wire [0:0] CLBLM_L_X8Y104_SLICE_X10Y104_D4;
  wire [0:0] CLBLM_L_X8Y104_SLICE_X10Y104_D5;
  wire [0:0] CLBLM_L_X8Y104_SLICE_X10Y104_D6;
  wire [0:0] CLBLM_L_X8Y104_SLICE_X10Y104_DO5;
  wire [0:0] CLBLM_L_X8Y104_SLICE_X10Y104_DO6;
  wire [0:0] CLBLM_L_X8Y104_SLICE_X10Y104_D_CY;
  wire [0:0] CLBLM_L_X8Y104_SLICE_X10Y104_D_XOR;
  wire [0:0] CLBLM_L_X8Y104_SLICE_X11Y104_A;
  wire [0:0] CLBLM_L_X8Y104_SLICE_X11Y104_A1;
  wire [0:0] CLBLM_L_X8Y104_SLICE_X11Y104_A2;
  wire [0:0] CLBLM_L_X8Y104_SLICE_X11Y104_A3;
  wire [0:0] CLBLM_L_X8Y104_SLICE_X11Y104_A4;
  wire [0:0] CLBLM_L_X8Y104_SLICE_X11Y104_A5;
  wire [0:0] CLBLM_L_X8Y104_SLICE_X11Y104_A6;
  wire [0:0] CLBLM_L_X8Y104_SLICE_X11Y104_AO5;
  wire [0:0] CLBLM_L_X8Y104_SLICE_X11Y104_AO6;
  wire [0:0] CLBLM_L_X8Y104_SLICE_X11Y104_A_CY;
  wire [0:0] CLBLM_L_X8Y104_SLICE_X11Y104_A_XOR;
  wire [0:0] CLBLM_L_X8Y104_SLICE_X11Y104_B;
  wire [0:0] CLBLM_L_X8Y104_SLICE_X11Y104_B1;
  wire [0:0] CLBLM_L_X8Y104_SLICE_X11Y104_B2;
  wire [0:0] CLBLM_L_X8Y104_SLICE_X11Y104_B3;
  wire [0:0] CLBLM_L_X8Y104_SLICE_X11Y104_B4;
  wire [0:0] CLBLM_L_X8Y104_SLICE_X11Y104_B5;
  wire [0:0] CLBLM_L_X8Y104_SLICE_X11Y104_B6;
  wire [0:0] CLBLM_L_X8Y104_SLICE_X11Y104_BO5;
  wire [0:0] CLBLM_L_X8Y104_SLICE_X11Y104_BO6;
  wire [0:0] CLBLM_L_X8Y104_SLICE_X11Y104_B_CY;
  wire [0:0] CLBLM_L_X8Y104_SLICE_X11Y104_B_XOR;
  wire [0:0] CLBLM_L_X8Y104_SLICE_X11Y104_C;
  wire [0:0] CLBLM_L_X8Y104_SLICE_X11Y104_C1;
  wire [0:0] CLBLM_L_X8Y104_SLICE_X11Y104_C2;
  wire [0:0] CLBLM_L_X8Y104_SLICE_X11Y104_C3;
  wire [0:0] CLBLM_L_X8Y104_SLICE_X11Y104_C4;
  wire [0:0] CLBLM_L_X8Y104_SLICE_X11Y104_C5;
  wire [0:0] CLBLM_L_X8Y104_SLICE_X11Y104_C6;
  wire [0:0] CLBLM_L_X8Y104_SLICE_X11Y104_CO5;
  wire [0:0] CLBLM_L_X8Y104_SLICE_X11Y104_CO6;
  wire [0:0] CLBLM_L_X8Y104_SLICE_X11Y104_C_CY;
  wire [0:0] CLBLM_L_X8Y104_SLICE_X11Y104_C_XOR;
  wire [0:0] CLBLM_L_X8Y104_SLICE_X11Y104_D;
  wire [0:0] CLBLM_L_X8Y104_SLICE_X11Y104_D1;
  wire [0:0] CLBLM_L_X8Y104_SLICE_X11Y104_D2;
  wire [0:0] CLBLM_L_X8Y104_SLICE_X11Y104_D3;
  wire [0:0] CLBLM_L_X8Y104_SLICE_X11Y104_D4;
  wire [0:0] CLBLM_L_X8Y104_SLICE_X11Y104_D5;
  wire [0:0] CLBLM_L_X8Y104_SLICE_X11Y104_D6;
  wire [0:0] CLBLM_L_X8Y104_SLICE_X11Y104_DO5;
  wire [0:0] CLBLM_L_X8Y104_SLICE_X11Y104_DO6;
  wire [0:0] CLBLM_L_X8Y104_SLICE_X11Y104_D_CY;
  wire [0:0] CLBLM_L_X8Y104_SLICE_X11Y104_D_XOR;
  wire [0:0] CLBLM_L_X8Y105_SLICE_X10Y105_A;
  wire [0:0] CLBLM_L_X8Y105_SLICE_X10Y105_A1;
  wire [0:0] CLBLM_L_X8Y105_SLICE_X10Y105_A2;
  wire [0:0] CLBLM_L_X8Y105_SLICE_X10Y105_A3;
  wire [0:0] CLBLM_L_X8Y105_SLICE_X10Y105_A4;
  wire [0:0] CLBLM_L_X8Y105_SLICE_X10Y105_A5;
  wire [0:0] CLBLM_L_X8Y105_SLICE_X10Y105_A6;
  wire [0:0] CLBLM_L_X8Y105_SLICE_X10Y105_AMUX;
  wire [0:0] CLBLM_L_X8Y105_SLICE_X10Y105_AO5;
  wire [0:0] CLBLM_L_X8Y105_SLICE_X10Y105_AO6;
  wire [0:0] CLBLM_L_X8Y105_SLICE_X10Y105_A_CY;
  wire [0:0] CLBLM_L_X8Y105_SLICE_X10Y105_A_XOR;
  wire [0:0] CLBLM_L_X8Y105_SLICE_X10Y105_B;
  wire [0:0] CLBLM_L_X8Y105_SLICE_X10Y105_B1;
  wire [0:0] CLBLM_L_X8Y105_SLICE_X10Y105_B2;
  wire [0:0] CLBLM_L_X8Y105_SLICE_X10Y105_B3;
  wire [0:0] CLBLM_L_X8Y105_SLICE_X10Y105_B4;
  wire [0:0] CLBLM_L_X8Y105_SLICE_X10Y105_B5;
  wire [0:0] CLBLM_L_X8Y105_SLICE_X10Y105_B6;
  wire [0:0] CLBLM_L_X8Y105_SLICE_X10Y105_BO5;
  wire [0:0] CLBLM_L_X8Y105_SLICE_X10Y105_BO6;
  wire [0:0] CLBLM_L_X8Y105_SLICE_X10Y105_B_CY;
  wire [0:0] CLBLM_L_X8Y105_SLICE_X10Y105_B_XOR;
  wire [0:0] CLBLM_L_X8Y105_SLICE_X10Y105_C;
  wire [0:0] CLBLM_L_X8Y105_SLICE_X10Y105_C1;
  wire [0:0] CLBLM_L_X8Y105_SLICE_X10Y105_C2;
  wire [0:0] CLBLM_L_X8Y105_SLICE_X10Y105_C3;
  wire [0:0] CLBLM_L_X8Y105_SLICE_X10Y105_C4;
  wire [0:0] CLBLM_L_X8Y105_SLICE_X10Y105_C5;
  wire [0:0] CLBLM_L_X8Y105_SLICE_X10Y105_C6;
  wire [0:0] CLBLM_L_X8Y105_SLICE_X10Y105_CO5;
  wire [0:0] CLBLM_L_X8Y105_SLICE_X10Y105_CO6;
  wire [0:0] CLBLM_L_X8Y105_SLICE_X10Y105_C_CY;
  wire [0:0] CLBLM_L_X8Y105_SLICE_X10Y105_C_XOR;
  wire [0:0] CLBLM_L_X8Y105_SLICE_X10Y105_D;
  wire [0:0] CLBLM_L_X8Y105_SLICE_X10Y105_D1;
  wire [0:0] CLBLM_L_X8Y105_SLICE_X10Y105_D2;
  wire [0:0] CLBLM_L_X8Y105_SLICE_X10Y105_D3;
  wire [0:0] CLBLM_L_X8Y105_SLICE_X10Y105_D4;
  wire [0:0] CLBLM_L_X8Y105_SLICE_X10Y105_D5;
  wire [0:0] CLBLM_L_X8Y105_SLICE_X10Y105_D6;
  wire [0:0] CLBLM_L_X8Y105_SLICE_X10Y105_DO5;
  wire [0:0] CLBLM_L_X8Y105_SLICE_X10Y105_DO6;
  wire [0:0] CLBLM_L_X8Y105_SLICE_X10Y105_D_CY;
  wire [0:0] CLBLM_L_X8Y105_SLICE_X10Y105_D_XOR;
  wire [0:0] CLBLM_L_X8Y105_SLICE_X11Y105_A;
  wire [0:0] CLBLM_L_X8Y105_SLICE_X11Y105_A1;
  wire [0:0] CLBLM_L_X8Y105_SLICE_X11Y105_A2;
  wire [0:0] CLBLM_L_X8Y105_SLICE_X11Y105_A3;
  wire [0:0] CLBLM_L_X8Y105_SLICE_X11Y105_A4;
  wire [0:0] CLBLM_L_X8Y105_SLICE_X11Y105_A5;
  wire [0:0] CLBLM_L_X8Y105_SLICE_X11Y105_A6;
  wire [0:0] CLBLM_L_X8Y105_SLICE_X11Y105_AMUX;
  wire [0:0] CLBLM_L_X8Y105_SLICE_X11Y105_AO5;
  wire [0:0] CLBLM_L_X8Y105_SLICE_X11Y105_AO6;
  wire [0:0] CLBLM_L_X8Y105_SLICE_X11Y105_A_CY;
  wire [0:0] CLBLM_L_X8Y105_SLICE_X11Y105_A_XOR;
  wire [0:0] CLBLM_L_X8Y105_SLICE_X11Y105_B;
  wire [0:0] CLBLM_L_X8Y105_SLICE_X11Y105_B1;
  wire [0:0] CLBLM_L_X8Y105_SLICE_X11Y105_B2;
  wire [0:0] CLBLM_L_X8Y105_SLICE_X11Y105_B3;
  wire [0:0] CLBLM_L_X8Y105_SLICE_X11Y105_B4;
  wire [0:0] CLBLM_L_X8Y105_SLICE_X11Y105_B5;
  wire [0:0] CLBLM_L_X8Y105_SLICE_X11Y105_B6;
  wire [0:0] CLBLM_L_X8Y105_SLICE_X11Y105_BMUX;
  wire [0:0] CLBLM_L_X8Y105_SLICE_X11Y105_BO5;
  wire [0:0] CLBLM_L_X8Y105_SLICE_X11Y105_BO6;
  wire [0:0] CLBLM_L_X8Y105_SLICE_X11Y105_B_CY;
  wire [0:0] CLBLM_L_X8Y105_SLICE_X11Y105_B_XOR;
  wire [0:0] CLBLM_L_X8Y105_SLICE_X11Y105_C;
  wire [0:0] CLBLM_L_X8Y105_SLICE_X11Y105_C1;
  wire [0:0] CLBLM_L_X8Y105_SLICE_X11Y105_C2;
  wire [0:0] CLBLM_L_X8Y105_SLICE_X11Y105_C3;
  wire [0:0] CLBLM_L_X8Y105_SLICE_X11Y105_C4;
  wire [0:0] CLBLM_L_X8Y105_SLICE_X11Y105_C5;
  wire [0:0] CLBLM_L_X8Y105_SLICE_X11Y105_C6;
  wire [0:0] CLBLM_L_X8Y105_SLICE_X11Y105_CO5;
  wire [0:0] CLBLM_L_X8Y105_SLICE_X11Y105_CO6;
  wire [0:0] CLBLM_L_X8Y105_SLICE_X11Y105_C_CY;
  wire [0:0] CLBLM_L_X8Y105_SLICE_X11Y105_C_XOR;
  wire [0:0] CLBLM_L_X8Y105_SLICE_X11Y105_D;
  wire [0:0] CLBLM_L_X8Y105_SLICE_X11Y105_D1;
  wire [0:0] CLBLM_L_X8Y105_SLICE_X11Y105_D2;
  wire [0:0] CLBLM_L_X8Y105_SLICE_X11Y105_D3;
  wire [0:0] CLBLM_L_X8Y105_SLICE_X11Y105_D4;
  wire [0:0] CLBLM_L_X8Y105_SLICE_X11Y105_D5;
  wire [0:0] CLBLM_L_X8Y105_SLICE_X11Y105_D6;
  wire [0:0] CLBLM_L_X8Y105_SLICE_X11Y105_DO5;
  wire [0:0] CLBLM_L_X8Y105_SLICE_X11Y105_DO6;
  wire [0:0] CLBLM_L_X8Y105_SLICE_X11Y105_D_CY;
  wire [0:0] CLBLM_L_X8Y105_SLICE_X11Y105_D_XOR;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X10Y106_A;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X10Y106_A1;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X10Y106_A2;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X10Y106_A3;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X10Y106_A4;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X10Y106_A5;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X10Y106_A6;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X10Y106_AMUX;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X10Y106_AO5;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X10Y106_AO6;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X10Y106_A_CY;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X10Y106_A_XOR;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X10Y106_B;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X10Y106_B1;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X10Y106_B2;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X10Y106_B3;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X10Y106_B4;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X10Y106_B5;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X10Y106_B6;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X10Y106_BMUX;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X10Y106_BO5;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X10Y106_BO6;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X10Y106_B_CY;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X10Y106_B_XOR;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X10Y106_C;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X10Y106_C1;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X10Y106_C2;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X10Y106_C3;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X10Y106_C4;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X10Y106_C5;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X10Y106_C6;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X10Y106_CO5;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X10Y106_CO6;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X10Y106_C_CY;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X10Y106_C_XOR;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X10Y106_D;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X10Y106_D1;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X10Y106_D2;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X10Y106_D3;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X10Y106_D4;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X10Y106_D5;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X10Y106_D6;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X10Y106_DO5;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X10Y106_DO6;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X10Y106_D_CY;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X10Y106_D_XOR;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X11Y106_A;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X11Y106_A1;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X11Y106_A2;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X11Y106_A3;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X11Y106_A4;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X11Y106_A5;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X11Y106_A6;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X11Y106_AO5;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X11Y106_AO6;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X11Y106_A_CY;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X11Y106_A_XOR;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X11Y106_B;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X11Y106_B1;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X11Y106_B2;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X11Y106_B3;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X11Y106_B4;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X11Y106_B5;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X11Y106_B6;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X11Y106_BO5;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X11Y106_BO6;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X11Y106_B_CY;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X11Y106_B_XOR;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X11Y106_C;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X11Y106_C1;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X11Y106_C2;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X11Y106_C3;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X11Y106_C4;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X11Y106_C5;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X11Y106_C6;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X11Y106_CO5;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X11Y106_CO6;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X11Y106_C_CY;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X11Y106_C_XOR;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X11Y106_D;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X11Y106_D1;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X11Y106_D2;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X11Y106_D3;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X11Y106_D4;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X11Y106_D5;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X11Y106_D6;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X11Y106_DO5;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X11Y106_DO6;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X11Y106_D_CY;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X11Y106_D_XOR;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X10Y107_A;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X10Y107_A1;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X10Y107_A2;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X10Y107_A3;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X10Y107_A4;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X10Y107_A5;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X10Y107_A6;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X10Y107_AO5;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X10Y107_AO6;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X10Y107_A_CY;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X10Y107_A_XOR;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X10Y107_B;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X10Y107_B1;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X10Y107_B2;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X10Y107_B3;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X10Y107_B4;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X10Y107_B5;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X10Y107_B6;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X10Y107_BO5;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X10Y107_BO6;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X10Y107_B_CY;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X10Y107_B_XOR;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X10Y107_C;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X10Y107_C1;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X10Y107_C2;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X10Y107_C3;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X10Y107_C4;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X10Y107_C5;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X10Y107_C6;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X10Y107_CO5;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X10Y107_CO6;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X10Y107_C_CY;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X10Y107_C_XOR;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X10Y107_D;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X10Y107_D1;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X10Y107_D2;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X10Y107_D3;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X10Y107_D4;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X10Y107_D5;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X10Y107_D6;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X10Y107_DO5;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X10Y107_DO6;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X10Y107_D_CY;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X10Y107_D_XOR;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X11Y107_A;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X11Y107_A1;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X11Y107_A2;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X11Y107_A3;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X11Y107_A4;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X11Y107_A5;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X11Y107_A6;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X11Y107_AMUX;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X11Y107_AO5;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X11Y107_AO6;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X11Y107_A_CY;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X11Y107_A_XOR;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X11Y107_B;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X11Y107_B1;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X11Y107_B2;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X11Y107_B3;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X11Y107_B4;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X11Y107_B5;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X11Y107_B6;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X11Y107_BMUX;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X11Y107_BO5;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X11Y107_BO6;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X11Y107_B_CY;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X11Y107_B_XOR;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X11Y107_C;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X11Y107_C1;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X11Y107_C2;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X11Y107_C3;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X11Y107_C4;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X11Y107_C5;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X11Y107_C6;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X11Y107_CMUX;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X11Y107_CO5;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X11Y107_CO6;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X11Y107_C_CY;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X11Y107_C_XOR;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X11Y107_D;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X11Y107_D1;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X11Y107_D2;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X11Y107_D3;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X11Y107_D4;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X11Y107_D5;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X11Y107_D6;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X11Y107_DO5;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X11Y107_DO6;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X11Y107_D_CY;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X11Y107_D_XOR;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X10Y108_A;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X10Y108_A1;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X10Y108_A2;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X10Y108_A3;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X10Y108_A4;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X10Y108_A5;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X10Y108_A6;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X10Y108_AMUX;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X10Y108_AO5;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X10Y108_AO6;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X10Y108_A_CY;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X10Y108_A_XOR;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X10Y108_B;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X10Y108_B1;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X10Y108_B2;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X10Y108_B3;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X10Y108_B4;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X10Y108_B5;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X10Y108_B6;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X10Y108_BO5;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X10Y108_BO6;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X10Y108_B_CY;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X10Y108_B_XOR;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X10Y108_C;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X10Y108_C1;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X10Y108_C2;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X10Y108_C3;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X10Y108_C4;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X10Y108_C5;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X10Y108_C6;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X10Y108_CO5;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X10Y108_CO6;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X10Y108_C_CY;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X10Y108_C_XOR;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X10Y108_D;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X10Y108_D1;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X10Y108_D2;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X10Y108_D3;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X10Y108_D4;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X10Y108_D5;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X10Y108_D6;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X10Y108_DO5;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X10Y108_DO6;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X10Y108_D_CY;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X10Y108_D_XOR;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X11Y108_A;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X11Y108_A1;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X11Y108_A2;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X11Y108_A3;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X11Y108_A4;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X11Y108_A5;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X11Y108_A6;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X11Y108_AO5;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X11Y108_AO6;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X11Y108_A_CY;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X11Y108_A_XOR;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X11Y108_B;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X11Y108_B1;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X11Y108_B2;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X11Y108_B3;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X11Y108_B4;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X11Y108_B5;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X11Y108_B6;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X11Y108_BO5;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X11Y108_BO6;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X11Y108_B_CY;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X11Y108_B_XOR;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X11Y108_C;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X11Y108_C1;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X11Y108_C2;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X11Y108_C3;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X11Y108_C4;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X11Y108_C5;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X11Y108_C6;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X11Y108_CO5;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X11Y108_CO6;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X11Y108_C_CY;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X11Y108_C_XOR;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X11Y108_D;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X11Y108_D1;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X11Y108_D2;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X11Y108_D3;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X11Y108_D4;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X11Y108_D5;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X11Y108_D6;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X11Y108_DO5;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X11Y108_DO6;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X11Y108_D_CY;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X11Y108_D_XOR;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X10Y109_A;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X10Y109_A1;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X10Y109_A2;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X10Y109_A3;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X10Y109_A4;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X10Y109_A5;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X10Y109_A6;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X10Y109_AO5;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X10Y109_AO6;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X10Y109_A_CY;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X10Y109_A_XOR;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X10Y109_B;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X10Y109_B1;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X10Y109_B2;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X10Y109_B3;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X10Y109_B4;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X10Y109_B5;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X10Y109_B6;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X10Y109_BO5;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X10Y109_BO6;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X10Y109_B_CY;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X10Y109_B_XOR;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X10Y109_C;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X10Y109_C1;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X10Y109_C2;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X10Y109_C3;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X10Y109_C4;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X10Y109_C5;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X10Y109_C6;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X10Y109_CO5;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X10Y109_CO6;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X10Y109_C_CY;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X10Y109_C_XOR;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X10Y109_D;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X10Y109_D1;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X10Y109_D2;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X10Y109_D3;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X10Y109_D4;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X10Y109_D5;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X10Y109_D6;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X10Y109_DO5;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X10Y109_DO6;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X10Y109_D_CY;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X10Y109_D_XOR;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X11Y109_A;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X11Y109_A1;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X11Y109_A2;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X11Y109_A3;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X11Y109_A4;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X11Y109_A5;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X11Y109_A6;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X11Y109_AO5;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X11Y109_AO6;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X11Y109_A_CY;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X11Y109_A_XOR;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X11Y109_B;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X11Y109_B1;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X11Y109_B2;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X11Y109_B3;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X11Y109_B4;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X11Y109_B5;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X11Y109_B6;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X11Y109_BO5;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X11Y109_BO6;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X11Y109_B_CY;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X11Y109_B_XOR;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X11Y109_C;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X11Y109_C1;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X11Y109_C2;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X11Y109_C3;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X11Y109_C4;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X11Y109_C5;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X11Y109_C6;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X11Y109_CO5;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X11Y109_CO6;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X11Y109_C_CY;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X11Y109_C_XOR;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X11Y109_D;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X11Y109_D1;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X11Y109_D2;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X11Y109_D3;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X11Y109_D4;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X11Y109_D5;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X11Y109_D6;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X11Y109_DO5;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X11Y109_DO6;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X11Y109_D_CY;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X11Y109_D_XOR;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X10Y110_A;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X10Y110_A1;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X10Y110_A2;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X10Y110_A3;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X10Y110_A4;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X10Y110_A5;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X10Y110_A6;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X10Y110_AO5;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X10Y110_AO6;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X10Y110_A_CY;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X10Y110_A_XOR;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X10Y110_B;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X10Y110_B1;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X10Y110_B2;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X10Y110_B3;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X10Y110_B4;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X10Y110_B5;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X10Y110_B6;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X10Y110_BO5;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X10Y110_BO6;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X10Y110_B_CY;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X10Y110_B_XOR;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X10Y110_C;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X10Y110_C1;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X10Y110_C2;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X10Y110_C3;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X10Y110_C4;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X10Y110_C5;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X10Y110_C6;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X10Y110_CMUX;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X10Y110_CO5;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X10Y110_CO6;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X10Y110_C_CY;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X10Y110_C_XOR;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X10Y110_D;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X10Y110_D1;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X10Y110_D2;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X10Y110_D3;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X10Y110_D4;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X10Y110_D5;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X10Y110_D6;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X10Y110_DO5;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X10Y110_DO6;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X10Y110_D_CY;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X10Y110_D_XOR;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X11Y110_A;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X11Y110_A1;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X11Y110_A2;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X11Y110_A3;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X11Y110_A4;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X11Y110_A5;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X11Y110_A6;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X11Y110_AMUX;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X11Y110_AO5;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X11Y110_AO6;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X11Y110_A_CY;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X11Y110_A_XOR;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X11Y110_B;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X11Y110_B1;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X11Y110_B2;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X11Y110_B3;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X11Y110_B4;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X11Y110_B5;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X11Y110_B6;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X11Y110_BMUX;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X11Y110_BO5;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X11Y110_BO6;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X11Y110_B_CY;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X11Y110_B_XOR;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X11Y110_C;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X11Y110_C1;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X11Y110_C2;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X11Y110_C3;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X11Y110_C4;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X11Y110_C5;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X11Y110_C6;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X11Y110_CO5;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X11Y110_CO6;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X11Y110_C_CY;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X11Y110_C_XOR;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X11Y110_D;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X11Y110_D1;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X11Y110_D2;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X11Y110_D3;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X11Y110_D4;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X11Y110_D5;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X11Y110_D6;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X11Y110_DO5;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X11Y110_DO6;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X11Y110_D_CY;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X11Y110_D_XOR;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X10Y111_A;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X10Y111_A1;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X10Y111_A2;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X10Y111_A3;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X10Y111_A4;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X10Y111_A5;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X10Y111_A6;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X10Y111_AMUX;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X10Y111_AO5;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X10Y111_AO6;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X10Y111_A_CY;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X10Y111_A_XOR;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X10Y111_B;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X10Y111_B1;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X10Y111_B2;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X10Y111_B3;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X10Y111_B4;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X10Y111_B5;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X10Y111_B6;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X10Y111_BO5;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X10Y111_BO6;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X10Y111_B_CY;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X10Y111_B_XOR;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X10Y111_C;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X10Y111_C1;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X10Y111_C2;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X10Y111_C3;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X10Y111_C4;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X10Y111_C5;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X10Y111_C6;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X10Y111_CO5;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X10Y111_CO6;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X10Y111_C_CY;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X10Y111_C_XOR;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X10Y111_D;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X10Y111_D1;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X10Y111_D2;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X10Y111_D3;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X10Y111_D4;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X10Y111_D5;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X10Y111_D6;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X10Y111_DO5;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X10Y111_DO6;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X10Y111_D_CY;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X10Y111_D_XOR;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X11Y111_A;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X11Y111_A1;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X11Y111_A2;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X11Y111_A3;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X11Y111_A4;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X11Y111_A5;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X11Y111_A6;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X11Y111_AMUX;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X11Y111_AO5;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X11Y111_AO6;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X11Y111_A_CY;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X11Y111_A_XOR;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X11Y111_B;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X11Y111_B1;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X11Y111_B2;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X11Y111_B3;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X11Y111_B4;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X11Y111_B5;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X11Y111_B6;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X11Y111_BO5;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X11Y111_BO6;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X11Y111_B_CY;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X11Y111_B_XOR;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X11Y111_C;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X11Y111_C1;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X11Y111_C2;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X11Y111_C3;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X11Y111_C4;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X11Y111_C5;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X11Y111_C6;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X11Y111_CO5;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X11Y111_CO6;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X11Y111_C_CY;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X11Y111_C_XOR;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X11Y111_D;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X11Y111_D1;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X11Y111_D2;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X11Y111_D3;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X11Y111_D4;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X11Y111_D5;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X11Y111_D6;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X11Y111_DO5;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X11Y111_DO6;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X11Y111_D_CY;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X11Y111_D_XOR;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X10Y112_A;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X10Y112_A1;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X10Y112_A2;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X10Y112_A3;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X10Y112_A4;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X10Y112_A5;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X10Y112_A6;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X10Y112_AMUX;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X10Y112_AO5;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X10Y112_AO6;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X10Y112_A_CY;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X10Y112_A_XOR;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X10Y112_B;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X10Y112_B1;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X10Y112_B2;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X10Y112_B3;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X10Y112_B4;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X10Y112_B5;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X10Y112_B6;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X10Y112_BO5;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X10Y112_BO6;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X10Y112_B_CY;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X10Y112_B_XOR;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X10Y112_C;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X10Y112_C1;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X10Y112_C2;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X10Y112_C3;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X10Y112_C4;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X10Y112_C5;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X10Y112_C6;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X10Y112_CO5;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X10Y112_CO6;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X10Y112_C_CY;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X10Y112_C_XOR;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X10Y112_D;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X10Y112_D1;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X10Y112_D2;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X10Y112_D3;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X10Y112_D4;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X10Y112_D5;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X10Y112_D6;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X10Y112_DO5;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X10Y112_DO6;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X10Y112_D_CY;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X10Y112_D_XOR;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X11Y112_A;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X11Y112_A1;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X11Y112_A2;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X11Y112_A3;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X11Y112_A4;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X11Y112_A5;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X11Y112_A6;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X11Y112_AO5;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X11Y112_AO6;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X11Y112_A_CY;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X11Y112_A_XOR;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X11Y112_B;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X11Y112_B1;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X11Y112_B2;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X11Y112_B3;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X11Y112_B4;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X11Y112_B5;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X11Y112_B6;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X11Y112_BO5;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X11Y112_BO6;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X11Y112_B_CY;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X11Y112_B_XOR;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X11Y112_C;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X11Y112_C1;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X11Y112_C2;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X11Y112_C3;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X11Y112_C4;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X11Y112_C5;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X11Y112_C6;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X11Y112_CO5;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X11Y112_CO6;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X11Y112_C_CY;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X11Y112_C_XOR;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X11Y112_D;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X11Y112_D1;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X11Y112_D2;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X11Y112_D3;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X11Y112_D4;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X11Y112_D5;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X11Y112_D6;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X11Y112_DO5;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X11Y112_DO6;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X11Y112_D_CY;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X11Y112_D_XOR;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X10Y113_A;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X10Y113_A1;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X10Y113_A2;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X10Y113_A3;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X10Y113_A4;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X10Y113_A5;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X10Y113_A6;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X10Y113_AMUX;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X10Y113_AO5;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X10Y113_AO6;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X10Y113_A_CY;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X10Y113_A_XOR;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X10Y113_B;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X10Y113_B1;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X10Y113_B2;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X10Y113_B3;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X10Y113_B4;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X10Y113_B5;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X10Y113_B6;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X10Y113_BO5;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X10Y113_BO6;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X10Y113_B_CY;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X10Y113_B_XOR;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X10Y113_C;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X10Y113_C1;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X10Y113_C2;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X10Y113_C3;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X10Y113_C4;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X10Y113_C5;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X10Y113_C6;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X10Y113_CO5;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X10Y113_CO6;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X10Y113_C_CY;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X10Y113_C_XOR;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X10Y113_D;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X10Y113_D1;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X10Y113_D2;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X10Y113_D3;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X10Y113_D4;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X10Y113_D5;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X10Y113_D6;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X10Y113_DO5;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X10Y113_DO6;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X10Y113_D_CY;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X10Y113_D_XOR;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X11Y113_A;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X11Y113_A1;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X11Y113_A2;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X11Y113_A3;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X11Y113_A4;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X11Y113_A5;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X11Y113_A6;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X11Y113_AO5;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X11Y113_AO6;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X11Y113_A_CY;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X11Y113_A_XOR;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X11Y113_B;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X11Y113_B1;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X11Y113_B2;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X11Y113_B3;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X11Y113_B4;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X11Y113_B5;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X11Y113_B6;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X11Y113_BO5;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X11Y113_BO6;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X11Y113_B_CY;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X11Y113_B_XOR;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X11Y113_C;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X11Y113_C1;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X11Y113_C2;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X11Y113_C3;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X11Y113_C4;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X11Y113_C5;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X11Y113_C6;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X11Y113_CO5;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X11Y113_CO6;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X11Y113_C_CY;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X11Y113_C_XOR;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X11Y113_D;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X11Y113_D1;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X11Y113_D2;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X11Y113_D3;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X11Y113_D4;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X11Y113_D5;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X11Y113_D6;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X11Y113_DO5;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X11Y113_DO6;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X11Y113_D_CY;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X11Y113_D_XOR;
  wire [0:0] CLBLM_R_X11Y104_SLICE_X14Y104_A;
  wire [0:0] CLBLM_R_X11Y104_SLICE_X14Y104_A1;
  wire [0:0] CLBLM_R_X11Y104_SLICE_X14Y104_A2;
  wire [0:0] CLBLM_R_X11Y104_SLICE_X14Y104_A3;
  wire [0:0] CLBLM_R_X11Y104_SLICE_X14Y104_A4;
  wire [0:0] CLBLM_R_X11Y104_SLICE_X14Y104_A5;
  wire [0:0] CLBLM_R_X11Y104_SLICE_X14Y104_A6;
  wire [0:0] CLBLM_R_X11Y104_SLICE_X14Y104_AMUX;
  wire [0:0] CLBLM_R_X11Y104_SLICE_X14Y104_AO5;
  wire [0:0] CLBLM_R_X11Y104_SLICE_X14Y104_AO6;
  wire [0:0] CLBLM_R_X11Y104_SLICE_X14Y104_A_CY;
  wire [0:0] CLBLM_R_X11Y104_SLICE_X14Y104_A_XOR;
  wire [0:0] CLBLM_R_X11Y104_SLICE_X14Y104_B;
  wire [0:0] CLBLM_R_X11Y104_SLICE_X14Y104_B1;
  wire [0:0] CLBLM_R_X11Y104_SLICE_X14Y104_B2;
  wire [0:0] CLBLM_R_X11Y104_SLICE_X14Y104_B3;
  wire [0:0] CLBLM_R_X11Y104_SLICE_X14Y104_B4;
  wire [0:0] CLBLM_R_X11Y104_SLICE_X14Y104_B5;
  wire [0:0] CLBLM_R_X11Y104_SLICE_X14Y104_B6;
  wire [0:0] CLBLM_R_X11Y104_SLICE_X14Y104_BO5;
  wire [0:0] CLBLM_R_X11Y104_SLICE_X14Y104_BO6;
  wire [0:0] CLBLM_R_X11Y104_SLICE_X14Y104_B_CY;
  wire [0:0] CLBLM_R_X11Y104_SLICE_X14Y104_B_XOR;
  wire [0:0] CLBLM_R_X11Y104_SLICE_X14Y104_C;
  wire [0:0] CLBLM_R_X11Y104_SLICE_X14Y104_C1;
  wire [0:0] CLBLM_R_X11Y104_SLICE_X14Y104_C2;
  wire [0:0] CLBLM_R_X11Y104_SLICE_X14Y104_C3;
  wire [0:0] CLBLM_R_X11Y104_SLICE_X14Y104_C4;
  wire [0:0] CLBLM_R_X11Y104_SLICE_X14Y104_C5;
  wire [0:0] CLBLM_R_X11Y104_SLICE_X14Y104_C6;
  wire [0:0] CLBLM_R_X11Y104_SLICE_X14Y104_CO5;
  wire [0:0] CLBLM_R_X11Y104_SLICE_X14Y104_CO6;
  wire [0:0] CLBLM_R_X11Y104_SLICE_X14Y104_C_CY;
  wire [0:0] CLBLM_R_X11Y104_SLICE_X14Y104_C_XOR;
  wire [0:0] CLBLM_R_X11Y104_SLICE_X14Y104_D;
  wire [0:0] CLBLM_R_X11Y104_SLICE_X14Y104_D1;
  wire [0:0] CLBLM_R_X11Y104_SLICE_X14Y104_D2;
  wire [0:0] CLBLM_R_X11Y104_SLICE_X14Y104_D3;
  wire [0:0] CLBLM_R_X11Y104_SLICE_X14Y104_D4;
  wire [0:0] CLBLM_R_X11Y104_SLICE_X14Y104_D5;
  wire [0:0] CLBLM_R_X11Y104_SLICE_X14Y104_D6;
  wire [0:0] CLBLM_R_X11Y104_SLICE_X14Y104_DO5;
  wire [0:0] CLBLM_R_X11Y104_SLICE_X14Y104_DO6;
  wire [0:0] CLBLM_R_X11Y104_SLICE_X14Y104_D_CY;
  wire [0:0] CLBLM_R_X11Y104_SLICE_X14Y104_D_XOR;
  wire [0:0] CLBLM_R_X11Y104_SLICE_X15Y104_A;
  wire [0:0] CLBLM_R_X11Y104_SLICE_X15Y104_A1;
  wire [0:0] CLBLM_R_X11Y104_SLICE_X15Y104_A2;
  wire [0:0] CLBLM_R_X11Y104_SLICE_X15Y104_A3;
  wire [0:0] CLBLM_R_X11Y104_SLICE_X15Y104_A4;
  wire [0:0] CLBLM_R_X11Y104_SLICE_X15Y104_A5;
  wire [0:0] CLBLM_R_X11Y104_SLICE_X15Y104_A6;
  wire [0:0] CLBLM_R_X11Y104_SLICE_X15Y104_AMUX;
  wire [0:0] CLBLM_R_X11Y104_SLICE_X15Y104_AO5;
  wire [0:0] CLBLM_R_X11Y104_SLICE_X15Y104_AO6;
  wire [0:0] CLBLM_R_X11Y104_SLICE_X15Y104_A_CY;
  wire [0:0] CLBLM_R_X11Y104_SLICE_X15Y104_A_XOR;
  wire [0:0] CLBLM_R_X11Y104_SLICE_X15Y104_B;
  wire [0:0] CLBLM_R_X11Y104_SLICE_X15Y104_B1;
  wire [0:0] CLBLM_R_X11Y104_SLICE_X15Y104_B2;
  wire [0:0] CLBLM_R_X11Y104_SLICE_X15Y104_B3;
  wire [0:0] CLBLM_R_X11Y104_SLICE_X15Y104_B4;
  wire [0:0] CLBLM_R_X11Y104_SLICE_X15Y104_B5;
  wire [0:0] CLBLM_R_X11Y104_SLICE_X15Y104_B6;
  wire [0:0] CLBLM_R_X11Y104_SLICE_X15Y104_BMUX;
  wire [0:0] CLBLM_R_X11Y104_SLICE_X15Y104_BO5;
  wire [0:0] CLBLM_R_X11Y104_SLICE_X15Y104_BO6;
  wire [0:0] CLBLM_R_X11Y104_SLICE_X15Y104_B_CY;
  wire [0:0] CLBLM_R_X11Y104_SLICE_X15Y104_B_XOR;
  wire [0:0] CLBLM_R_X11Y104_SLICE_X15Y104_C;
  wire [0:0] CLBLM_R_X11Y104_SLICE_X15Y104_C1;
  wire [0:0] CLBLM_R_X11Y104_SLICE_X15Y104_C2;
  wire [0:0] CLBLM_R_X11Y104_SLICE_X15Y104_C3;
  wire [0:0] CLBLM_R_X11Y104_SLICE_X15Y104_C4;
  wire [0:0] CLBLM_R_X11Y104_SLICE_X15Y104_C5;
  wire [0:0] CLBLM_R_X11Y104_SLICE_X15Y104_C6;
  wire [0:0] CLBLM_R_X11Y104_SLICE_X15Y104_CO5;
  wire [0:0] CLBLM_R_X11Y104_SLICE_X15Y104_CO6;
  wire [0:0] CLBLM_R_X11Y104_SLICE_X15Y104_C_CY;
  wire [0:0] CLBLM_R_X11Y104_SLICE_X15Y104_C_XOR;
  wire [0:0] CLBLM_R_X11Y104_SLICE_X15Y104_D;
  wire [0:0] CLBLM_R_X11Y104_SLICE_X15Y104_D1;
  wire [0:0] CLBLM_R_X11Y104_SLICE_X15Y104_D2;
  wire [0:0] CLBLM_R_X11Y104_SLICE_X15Y104_D3;
  wire [0:0] CLBLM_R_X11Y104_SLICE_X15Y104_D4;
  wire [0:0] CLBLM_R_X11Y104_SLICE_X15Y104_D5;
  wire [0:0] CLBLM_R_X11Y104_SLICE_X15Y104_D6;
  wire [0:0] CLBLM_R_X11Y104_SLICE_X15Y104_DO5;
  wire [0:0] CLBLM_R_X11Y104_SLICE_X15Y104_DO6;
  wire [0:0] CLBLM_R_X11Y104_SLICE_X15Y104_D_CY;
  wire [0:0] CLBLM_R_X11Y104_SLICE_X15Y104_D_XOR;
  wire [0:0] CLBLM_R_X11Y105_SLICE_X14Y105_A;
  wire [0:0] CLBLM_R_X11Y105_SLICE_X14Y105_A1;
  wire [0:0] CLBLM_R_X11Y105_SLICE_X14Y105_A2;
  wire [0:0] CLBLM_R_X11Y105_SLICE_X14Y105_A3;
  wire [0:0] CLBLM_R_X11Y105_SLICE_X14Y105_A4;
  wire [0:0] CLBLM_R_X11Y105_SLICE_X14Y105_A5;
  wire [0:0] CLBLM_R_X11Y105_SLICE_X14Y105_A6;
  wire [0:0] CLBLM_R_X11Y105_SLICE_X14Y105_AMUX;
  wire [0:0] CLBLM_R_X11Y105_SLICE_X14Y105_AO5;
  wire [0:0] CLBLM_R_X11Y105_SLICE_X14Y105_AO6;
  wire [0:0] CLBLM_R_X11Y105_SLICE_X14Y105_A_CY;
  wire [0:0] CLBLM_R_X11Y105_SLICE_X14Y105_A_XOR;
  wire [0:0] CLBLM_R_X11Y105_SLICE_X14Y105_B;
  wire [0:0] CLBLM_R_X11Y105_SLICE_X14Y105_B1;
  wire [0:0] CLBLM_R_X11Y105_SLICE_X14Y105_B2;
  wire [0:0] CLBLM_R_X11Y105_SLICE_X14Y105_B3;
  wire [0:0] CLBLM_R_X11Y105_SLICE_X14Y105_B4;
  wire [0:0] CLBLM_R_X11Y105_SLICE_X14Y105_B5;
  wire [0:0] CLBLM_R_X11Y105_SLICE_X14Y105_B6;
  wire [0:0] CLBLM_R_X11Y105_SLICE_X14Y105_BO5;
  wire [0:0] CLBLM_R_X11Y105_SLICE_X14Y105_BO6;
  wire [0:0] CLBLM_R_X11Y105_SLICE_X14Y105_B_CY;
  wire [0:0] CLBLM_R_X11Y105_SLICE_X14Y105_B_XOR;
  wire [0:0] CLBLM_R_X11Y105_SLICE_X14Y105_C;
  wire [0:0] CLBLM_R_X11Y105_SLICE_X14Y105_C1;
  wire [0:0] CLBLM_R_X11Y105_SLICE_X14Y105_C2;
  wire [0:0] CLBLM_R_X11Y105_SLICE_X14Y105_C3;
  wire [0:0] CLBLM_R_X11Y105_SLICE_X14Y105_C4;
  wire [0:0] CLBLM_R_X11Y105_SLICE_X14Y105_C5;
  wire [0:0] CLBLM_R_X11Y105_SLICE_X14Y105_C6;
  wire [0:0] CLBLM_R_X11Y105_SLICE_X14Y105_CO5;
  wire [0:0] CLBLM_R_X11Y105_SLICE_X14Y105_CO6;
  wire [0:0] CLBLM_R_X11Y105_SLICE_X14Y105_C_CY;
  wire [0:0] CLBLM_R_X11Y105_SLICE_X14Y105_C_XOR;
  wire [0:0] CLBLM_R_X11Y105_SLICE_X14Y105_D;
  wire [0:0] CLBLM_R_X11Y105_SLICE_X14Y105_D1;
  wire [0:0] CLBLM_R_X11Y105_SLICE_X14Y105_D2;
  wire [0:0] CLBLM_R_X11Y105_SLICE_X14Y105_D3;
  wire [0:0] CLBLM_R_X11Y105_SLICE_X14Y105_D4;
  wire [0:0] CLBLM_R_X11Y105_SLICE_X14Y105_D5;
  wire [0:0] CLBLM_R_X11Y105_SLICE_X14Y105_D6;
  wire [0:0] CLBLM_R_X11Y105_SLICE_X14Y105_DO5;
  wire [0:0] CLBLM_R_X11Y105_SLICE_X14Y105_DO6;
  wire [0:0] CLBLM_R_X11Y105_SLICE_X14Y105_D_CY;
  wire [0:0] CLBLM_R_X11Y105_SLICE_X14Y105_D_XOR;
  wire [0:0] CLBLM_R_X11Y105_SLICE_X15Y105_A;
  wire [0:0] CLBLM_R_X11Y105_SLICE_X15Y105_A1;
  wire [0:0] CLBLM_R_X11Y105_SLICE_X15Y105_A2;
  wire [0:0] CLBLM_R_X11Y105_SLICE_X15Y105_A3;
  wire [0:0] CLBLM_R_X11Y105_SLICE_X15Y105_A4;
  wire [0:0] CLBLM_R_X11Y105_SLICE_X15Y105_A5;
  wire [0:0] CLBLM_R_X11Y105_SLICE_X15Y105_A6;
  wire [0:0] CLBLM_R_X11Y105_SLICE_X15Y105_AMUX;
  wire [0:0] CLBLM_R_X11Y105_SLICE_X15Y105_AO5;
  wire [0:0] CLBLM_R_X11Y105_SLICE_X15Y105_AO6;
  wire [0:0] CLBLM_R_X11Y105_SLICE_X15Y105_A_CY;
  wire [0:0] CLBLM_R_X11Y105_SLICE_X15Y105_A_XOR;
  wire [0:0] CLBLM_R_X11Y105_SLICE_X15Y105_B;
  wire [0:0] CLBLM_R_X11Y105_SLICE_X15Y105_B1;
  wire [0:0] CLBLM_R_X11Y105_SLICE_X15Y105_B2;
  wire [0:0] CLBLM_R_X11Y105_SLICE_X15Y105_B3;
  wire [0:0] CLBLM_R_X11Y105_SLICE_X15Y105_B4;
  wire [0:0] CLBLM_R_X11Y105_SLICE_X15Y105_B5;
  wire [0:0] CLBLM_R_X11Y105_SLICE_X15Y105_B6;
  wire [0:0] CLBLM_R_X11Y105_SLICE_X15Y105_BO5;
  wire [0:0] CLBLM_R_X11Y105_SLICE_X15Y105_BO6;
  wire [0:0] CLBLM_R_X11Y105_SLICE_X15Y105_B_CY;
  wire [0:0] CLBLM_R_X11Y105_SLICE_X15Y105_B_XOR;
  wire [0:0] CLBLM_R_X11Y105_SLICE_X15Y105_C;
  wire [0:0] CLBLM_R_X11Y105_SLICE_X15Y105_C1;
  wire [0:0] CLBLM_R_X11Y105_SLICE_X15Y105_C2;
  wire [0:0] CLBLM_R_X11Y105_SLICE_X15Y105_C3;
  wire [0:0] CLBLM_R_X11Y105_SLICE_X15Y105_C4;
  wire [0:0] CLBLM_R_X11Y105_SLICE_X15Y105_C5;
  wire [0:0] CLBLM_R_X11Y105_SLICE_X15Y105_C6;
  wire [0:0] CLBLM_R_X11Y105_SLICE_X15Y105_CO5;
  wire [0:0] CLBLM_R_X11Y105_SLICE_X15Y105_CO6;
  wire [0:0] CLBLM_R_X11Y105_SLICE_X15Y105_C_CY;
  wire [0:0] CLBLM_R_X11Y105_SLICE_X15Y105_C_XOR;
  wire [0:0] CLBLM_R_X11Y105_SLICE_X15Y105_D;
  wire [0:0] CLBLM_R_X11Y105_SLICE_X15Y105_D1;
  wire [0:0] CLBLM_R_X11Y105_SLICE_X15Y105_D2;
  wire [0:0] CLBLM_R_X11Y105_SLICE_X15Y105_D3;
  wire [0:0] CLBLM_R_X11Y105_SLICE_X15Y105_D4;
  wire [0:0] CLBLM_R_X11Y105_SLICE_X15Y105_D5;
  wire [0:0] CLBLM_R_X11Y105_SLICE_X15Y105_D6;
  wire [0:0] CLBLM_R_X11Y105_SLICE_X15Y105_DO5;
  wire [0:0] CLBLM_R_X11Y105_SLICE_X15Y105_DO6;
  wire [0:0] CLBLM_R_X11Y105_SLICE_X15Y105_D_CY;
  wire [0:0] CLBLM_R_X11Y105_SLICE_X15Y105_D_XOR;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X14Y106_A;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X14Y106_A1;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X14Y106_A2;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X14Y106_A3;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X14Y106_A4;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X14Y106_A5;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X14Y106_A6;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X14Y106_AO5;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X14Y106_AO6;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X14Y106_A_CY;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X14Y106_A_XOR;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X14Y106_B;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X14Y106_B1;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X14Y106_B2;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X14Y106_B3;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X14Y106_B4;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X14Y106_B5;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X14Y106_B6;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X14Y106_BMUX;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X14Y106_BO5;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X14Y106_BO6;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X14Y106_B_CY;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X14Y106_B_XOR;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X14Y106_C;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X14Y106_C1;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X14Y106_C2;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X14Y106_C3;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X14Y106_C4;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X14Y106_C5;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X14Y106_C6;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X14Y106_CO5;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X14Y106_CO6;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X14Y106_C_CY;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X14Y106_C_XOR;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X14Y106_D;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X14Y106_D1;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X14Y106_D2;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X14Y106_D3;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X14Y106_D4;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X14Y106_D5;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X14Y106_D6;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X14Y106_DO5;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X14Y106_DO6;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X14Y106_D_CY;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X14Y106_D_XOR;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X15Y106_A;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X15Y106_A1;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X15Y106_A2;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X15Y106_A3;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X15Y106_A4;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X15Y106_A5;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X15Y106_A6;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X15Y106_AMUX;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X15Y106_AO5;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X15Y106_AO6;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X15Y106_A_CY;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X15Y106_A_XOR;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X15Y106_B;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X15Y106_B1;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X15Y106_B2;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X15Y106_B3;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X15Y106_B4;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X15Y106_B5;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X15Y106_B6;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X15Y106_BO5;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X15Y106_BO6;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X15Y106_B_CY;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X15Y106_B_XOR;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X15Y106_C;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X15Y106_C1;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X15Y106_C2;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X15Y106_C3;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X15Y106_C4;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X15Y106_C5;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X15Y106_C6;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X15Y106_CO5;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X15Y106_CO6;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X15Y106_C_CY;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X15Y106_C_XOR;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X15Y106_D;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X15Y106_D1;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X15Y106_D2;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X15Y106_D3;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X15Y106_D4;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X15Y106_D5;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X15Y106_D6;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X15Y106_DO5;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X15Y106_DO6;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X15Y106_D_CY;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X15Y106_D_XOR;
  wire [0:0] CLBLM_R_X11Y107_SLICE_X14Y107_A;
  wire [0:0] CLBLM_R_X11Y107_SLICE_X14Y107_A1;
  wire [0:0] CLBLM_R_X11Y107_SLICE_X14Y107_A2;
  wire [0:0] CLBLM_R_X11Y107_SLICE_X14Y107_A3;
  wire [0:0] CLBLM_R_X11Y107_SLICE_X14Y107_A4;
  wire [0:0] CLBLM_R_X11Y107_SLICE_X14Y107_A5;
  wire [0:0] CLBLM_R_X11Y107_SLICE_X14Y107_A6;
  wire [0:0] CLBLM_R_X11Y107_SLICE_X14Y107_AMUX;
  wire [0:0] CLBLM_R_X11Y107_SLICE_X14Y107_AO5;
  wire [0:0] CLBLM_R_X11Y107_SLICE_X14Y107_AO6;
  wire [0:0] CLBLM_R_X11Y107_SLICE_X14Y107_A_CY;
  wire [0:0] CLBLM_R_X11Y107_SLICE_X14Y107_A_XOR;
  wire [0:0] CLBLM_R_X11Y107_SLICE_X14Y107_B;
  wire [0:0] CLBLM_R_X11Y107_SLICE_X14Y107_B1;
  wire [0:0] CLBLM_R_X11Y107_SLICE_X14Y107_B2;
  wire [0:0] CLBLM_R_X11Y107_SLICE_X14Y107_B3;
  wire [0:0] CLBLM_R_X11Y107_SLICE_X14Y107_B4;
  wire [0:0] CLBLM_R_X11Y107_SLICE_X14Y107_B5;
  wire [0:0] CLBLM_R_X11Y107_SLICE_X14Y107_B6;
  wire [0:0] CLBLM_R_X11Y107_SLICE_X14Y107_BMUX;
  wire [0:0] CLBLM_R_X11Y107_SLICE_X14Y107_BO5;
  wire [0:0] CLBLM_R_X11Y107_SLICE_X14Y107_BO6;
  wire [0:0] CLBLM_R_X11Y107_SLICE_X14Y107_B_CY;
  wire [0:0] CLBLM_R_X11Y107_SLICE_X14Y107_B_XOR;
  wire [0:0] CLBLM_R_X11Y107_SLICE_X14Y107_C;
  wire [0:0] CLBLM_R_X11Y107_SLICE_X14Y107_C1;
  wire [0:0] CLBLM_R_X11Y107_SLICE_X14Y107_C2;
  wire [0:0] CLBLM_R_X11Y107_SLICE_X14Y107_C3;
  wire [0:0] CLBLM_R_X11Y107_SLICE_X14Y107_C4;
  wire [0:0] CLBLM_R_X11Y107_SLICE_X14Y107_C5;
  wire [0:0] CLBLM_R_X11Y107_SLICE_X14Y107_C6;
  wire [0:0] CLBLM_R_X11Y107_SLICE_X14Y107_CMUX;
  wire [0:0] CLBLM_R_X11Y107_SLICE_X14Y107_CO5;
  wire [0:0] CLBLM_R_X11Y107_SLICE_X14Y107_CO6;
  wire [0:0] CLBLM_R_X11Y107_SLICE_X14Y107_C_CY;
  wire [0:0] CLBLM_R_X11Y107_SLICE_X14Y107_C_XOR;
  wire [0:0] CLBLM_R_X11Y107_SLICE_X14Y107_D;
  wire [0:0] CLBLM_R_X11Y107_SLICE_X14Y107_D1;
  wire [0:0] CLBLM_R_X11Y107_SLICE_X14Y107_D2;
  wire [0:0] CLBLM_R_X11Y107_SLICE_X14Y107_D3;
  wire [0:0] CLBLM_R_X11Y107_SLICE_X14Y107_D4;
  wire [0:0] CLBLM_R_X11Y107_SLICE_X14Y107_D5;
  wire [0:0] CLBLM_R_X11Y107_SLICE_X14Y107_D6;
  wire [0:0] CLBLM_R_X11Y107_SLICE_X14Y107_DMUX;
  wire [0:0] CLBLM_R_X11Y107_SLICE_X14Y107_DO5;
  wire [0:0] CLBLM_R_X11Y107_SLICE_X14Y107_DO6;
  wire [0:0] CLBLM_R_X11Y107_SLICE_X14Y107_D_CY;
  wire [0:0] CLBLM_R_X11Y107_SLICE_X14Y107_D_XOR;
  wire [0:0] CLBLM_R_X11Y107_SLICE_X15Y107_A;
  wire [0:0] CLBLM_R_X11Y107_SLICE_X15Y107_A1;
  wire [0:0] CLBLM_R_X11Y107_SLICE_X15Y107_A2;
  wire [0:0] CLBLM_R_X11Y107_SLICE_X15Y107_A3;
  wire [0:0] CLBLM_R_X11Y107_SLICE_X15Y107_A4;
  wire [0:0] CLBLM_R_X11Y107_SLICE_X15Y107_A5;
  wire [0:0] CLBLM_R_X11Y107_SLICE_X15Y107_A6;
  wire [0:0] CLBLM_R_X11Y107_SLICE_X15Y107_AMUX;
  wire [0:0] CLBLM_R_X11Y107_SLICE_X15Y107_AO5;
  wire [0:0] CLBLM_R_X11Y107_SLICE_X15Y107_AO6;
  wire [0:0] CLBLM_R_X11Y107_SLICE_X15Y107_A_CY;
  wire [0:0] CLBLM_R_X11Y107_SLICE_X15Y107_A_XOR;
  wire [0:0] CLBLM_R_X11Y107_SLICE_X15Y107_B;
  wire [0:0] CLBLM_R_X11Y107_SLICE_X15Y107_B1;
  wire [0:0] CLBLM_R_X11Y107_SLICE_X15Y107_B2;
  wire [0:0] CLBLM_R_X11Y107_SLICE_X15Y107_B3;
  wire [0:0] CLBLM_R_X11Y107_SLICE_X15Y107_B4;
  wire [0:0] CLBLM_R_X11Y107_SLICE_X15Y107_B5;
  wire [0:0] CLBLM_R_X11Y107_SLICE_X15Y107_B6;
  wire [0:0] CLBLM_R_X11Y107_SLICE_X15Y107_BO5;
  wire [0:0] CLBLM_R_X11Y107_SLICE_X15Y107_BO6;
  wire [0:0] CLBLM_R_X11Y107_SLICE_X15Y107_B_CY;
  wire [0:0] CLBLM_R_X11Y107_SLICE_X15Y107_B_XOR;
  wire [0:0] CLBLM_R_X11Y107_SLICE_X15Y107_C;
  wire [0:0] CLBLM_R_X11Y107_SLICE_X15Y107_C1;
  wire [0:0] CLBLM_R_X11Y107_SLICE_X15Y107_C2;
  wire [0:0] CLBLM_R_X11Y107_SLICE_X15Y107_C3;
  wire [0:0] CLBLM_R_X11Y107_SLICE_X15Y107_C4;
  wire [0:0] CLBLM_R_X11Y107_SLICE_X15Y107_C5;
  wire [0:0] CLBLM_R_X11Y107_SLICE_X15Y107_C6;
  wire [0:0] CLBLM_R_X11Y107_SLICE_X15Y107_CO5;
  wire [0:0] CLBLM_R_X11Y107_SLICE_X15Y107_CO6;
  wire [0:0] CLBLM_R_X11Y107_SLICE_X15Y107_C_CY;
  wire [0:0] CLBLM_R_X11Y107_SLICE_X15Y107_C_XOR;
  wire [0:0] CLBLM_R_X11Y107_SLICE_X15Y107_D;
  wire [0:0] CLBLM_R_X11Y107_SLICE_X15Y107_D1;
  wire [0:0] CLBLM_R_X11Y107_SLICE_X15Y107_D2;
  wire [0:0] CLBLM_R_X11Y107_SLICE_X15Y107_D3;
  wire [0:0] CLBLM_R_X11Y107_SLICE_X15Y107_D4;
  wire [0:0] CLBLM_R_X11Y107_SLICE_X15Y107_D5;
  wire [0:0] CLBLM_R_X11Y107_SLICE_X15Y107_D6;
  wire [0:0] CLBLM_R_X11Y107_SLICE_X15Y107_DO5;
  wire [0:0] CLBLM_R_X11Y107_SLICE_X15Y107_DO6;
  wire [0:0] CLBLM_R_X11Y107_SLICE_X15Y107_D_CY;
  wire [0:0] CLBLM_R_X11Y107_SLICE_X15Y107_D_XOR;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X14Y108_A;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X14Y108_A1;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X14Y108_A2;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X14Y108_A3;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X14Y108_A4;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X14Y108_A5;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X14Y108_A6;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X14Y108_AO5;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X14Y108_AO6;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X14Y108_A_CY;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X14Y108_A_XOR;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X14Y108_B;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X14Y108_B1;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X14Y108_B2;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X14Y108_B3;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X14Y108_B4;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X14Y108_B5;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X14Y108_B6;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X14Y108_BO5;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X14Y108_BO6;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X14Y108_B_CY;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X14Y108_B_XOR;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X14Y108_C;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X14Y108_C1;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X14Y108_C2;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X14Y108_C3;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X14Y108_C4;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X14Y108_C5;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X14Y108_C6;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X14Y108_CO5;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X14Y108_CO6;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X14Y108_C_CY;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X14Y108_C_XOR;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X14Y108_D;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X14Y108_D1;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X14Y108_D2;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X14Y108_D3;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X14Y108_D4;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X14Y108_D5;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X14Y108_D6;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X14Y108_DO5;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X14Y108_DO6;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X14Y108_D_CY;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X14Y108_D_XOR;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X15Y108_A;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X15Y108_A1;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X15Y108_A2;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X15Y108_A3;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X15Y108_A4;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X15Y108_A5;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X15Y108_A6;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X15Y108_AO5;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X15Y108_AO6;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X15Y108_A_CY;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X15Y108_A_XOR;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X15Y108_B;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X15Y108_B1;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X15Y108_B2;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X15Y108_B3;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X15Y108_B4;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X15Y108_B5;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X15Y108_B6;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X15Y108_BO5;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X15Y108_BO6;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X15Y108_B_CY;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X15Y108_B_XOR;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X15Y108_C;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X15Y108_C1;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X15Y108_C2;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X15Y108_C3;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X15Y108_C4;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X15Y108_C5;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X15Y108_C6;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X15Y108_CMUX;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X15Y108_CO5;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X15Y108_CO6;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X15Y108_C_CY;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X15Y108_C_XOR;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X15Y108_D;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X15Y108_D1;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X15Y108_D2;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X15Y108_D3;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X15Y108_D4;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X15Y108_D5;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X15Y108_D6;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X15Y108_DO5;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X15Y108_DO6;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X15Y108_D_CY;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X15Y108_D_XOR;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X14Y109_A;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X14Y109_A1;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X14Y109_A2;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X14Y109_A3;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X14Y109_A4;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X14Y109_A5;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X14Y109_A6;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X14Y109_AMUX;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X14Y109_AO5;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X14Y109_AO6;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X14Y109_A_CY;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X14Y109_A_XOR;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X14Y109_B;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X14Y109_B1;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X14Y109_B2;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X14Y109_B3;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X14Y109_B4;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X14Y109_B5;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X14Y109_B6;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X14Y109_BO5;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X14Y109_BO6;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X14Y109_B_CY;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X14Y109_B_XOR;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X14Y109_C;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X14Y109_C1;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X14Y109_C2;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X14Y109_C3;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X14Y109_C4;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X14Y109_C5;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X14Y109_C6;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X14Y109_CO5;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X14Y109_CO6;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X14Y109_C_CY;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X14Y109_C_XOR;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X14Y109_D;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X14Y109_D1;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X14Y109_D2;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X14Y109_D3;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X14Y109_D4;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X14Y109_D5;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X14Y109_D6;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X14Y109_DO5;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X14Y109_DO6;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X14Y109_D_CY;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X14Y109_D_XOR;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X15Y109_A;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X15Y109_A1;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X15Y109_A2;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X15Y109_A3;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X15Y109_A4;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X15Y109_A5;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X15Y109_A6;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X15Y109_AO5;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X15Y109_AO6;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X15Y109_A_CY;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X15Y109_A_XOR;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X15Y109_B;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X15Y109_B1;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X15Y109_B2;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X15Y109_B3;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X15Y109_B4;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X15Y109_B5;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X15Y109_B6;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X15Y109_BMUX;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X15Y109_BO5;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X15Y109_BO6;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X15Y109_B_CY;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X15Y109_B_XOR;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X15Y109_C;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X15Y109_C1;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X15Y109_C2;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X15Y109_C3;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X15Y109_C4;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X15Y109_C5;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X15Y109_C6;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X15Y109_CO5;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X15Y109_CO6;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X15Y109_C_CY;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X15Y109_C_XOR;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X15Y109_D;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X15Y109_D1;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X15Y109_D2;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X15Y109_D3;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X15Y109_D4;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X15Y109_D5;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X15Y109_D6;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X15Y109_DO5;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X15Y109_DO6;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X15Y109_D_CY;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X15Y109_D_XOR;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X14Y110_A;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X14Y110_A1;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X14Y110_A2;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X14Y110_A3;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X14Y110_A4;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X14Y110_A5;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X14Y110_A6;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X14Y110_AMUX;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X14Y110_AO5;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X14Y110_AO6;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X14Y110_A_CY;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X14Y110_A_XOR;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X14Y110_B;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X14Y110_B1;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X14Y110_B2;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X14Y110_B3;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X14Y110_B4;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X14Y110_B5;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X14Y110_B6;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X14Y110_BO5;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X14Y110_BO6;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X14Y110_B_CY;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X14Y110_B_XOR;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X14Y110_C;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X14Y110_C1;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X14Y110_C2;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X14Y110_C3;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X14Y110_C4;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X14Y110_C5;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X14Y110_C6;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X14Y110_CO5;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X14Y110_CO6;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X14Y110_C_CY;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X14Y110_C_XOR;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X14Y110_D;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X14Y110_D1;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X14Y110_D2;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X14Y110_D3;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X14Y110_D4;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X14Y110_D5;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X14Y110_D6;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X14Y110_DO5;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X14Y110_DO6;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X14Y110_D_CY;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X14Y110_D_XOR;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X15Y110_A;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X15Y110_A1;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X15Y110_A2;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X15Y110_A3;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X15Y110_A4;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X15Y110_A5;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X15Y110_A6;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X15Y110_AMUX;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X15Y110_AO5;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X15Y110_AO6;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X15Y110_A_CY;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X15Y110_A_XOR;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X15Y110_B;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X15Y110_B1;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X15Y110_B2;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X15Y110_B3;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X15Y110_B4;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X15Y110_B5;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X15Y110_B6;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X15Y110_BMUX;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X15Y110_BO5;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X15Y110_BO6;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X15Y110_B_CY;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X15Y110_B_XOR;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X15Y110_C;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X15Y110_C1;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X15Y110_C2;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X15Y110_C3;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X15Y110_C4;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X15Y110_C5;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X15Y110_C6;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X15Y110_CO5;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X15Y110_CO6;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X15Y110_C_CY;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X15Y110_C_XOR;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X15Y110_D;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X15Y110_D1;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X15Y110_D2;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X15Y110_D3;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X15Y110_D4;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X15Y110_D5;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X15Y110_D6;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X15Y110_DO5;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X15Y110_DO6;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X15Y110_D_CY;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X15Y110_D_XOR;
  wire [0:0] CLBLM_R_X11Y111_SLICE_X14Y111_A;
  wire [0:0] CLBLM_R_X11Y111_SLICE_X14Y111_A1;
  wire [0:0] CLBLM_R_X11Y111_SLICE_X14Y111_A2;
  wire [0:0] CLBLM_R_X11Y111_SLICE_X14Y111_A3;
  wire [0:0] CLBLM_R_X11Y111_SLICE_X14Y111_A4;
  wire [0:0] CLBLM_R_X11Y111_SLICE_X14Y111_A5;
  wire [0:0] CLBLM_R_X11Y111_SLICE_X14Y111_A6;
  wire [0:0] CLBLM_R_X11Y111_SLICE_X14Y111_AMUX;
  wire [0:0] CLBLM_R_X11Y111_SLICE_X14Y111_AO5;
  wire [0:0] CLBLM_R_X11Y111_SLICE_X14Y111_AO6;
  wire [0:0] CLBLM_R_X11Y111_SLICE_X14Y111_A_CY;
  wire [0:0] CLBLM_R_X11Y111_SLICE_X14Y111_A_XOR;
  wire [0:0] CLBLM_R_X11Y111_SLICE_X14Y111_B;
  wire [0:0] CLBLM_R_X11Y111_SLICE_X14Y111_B1;
  wire [0:0] CLBLM_R_X11Y111_SLICE_X14Y111_B2;
  wire [0:0] CLBLM_R_X11Y111_SLICE_X14Y111_B3;
  wire [0:0] CLBLM_R_X11Y111_SLICE_X14Y111_B4;
  wire [0:0] CLBLM_R_X11Y111_SLICE_X14Y111_B5;
  wire [0:0] CLBLM_R_X11Y111_SLICE_X14Y111_B6;
  wire [0:0] CLBLM_R_X11Y111_SLICE_X14Y111_BMUX;
  wire [0:0] CLBLM_R_X11Y111_SLICE_X14Y111_BO5;
  wire [0:0] CLBLM_R_X11Y111_SLICE_X14Y111_BO6;
  wire [0:0] CLBLM_R_X11Y111_SLICE_X14Y111_B_CY;
  wire [0:0] CLBLM_R_X11Y111_SLICE_X14Y111_B_XOR;
  wire [0:0] CLBLM_R_X11Y111_SLICE_X14Y111_C;
  wire [0:0] CLBLM_R_X11Y111_SLICE_X14Y111_C1;
  wire [0:0] CLBLM_R_X11Y111_SLICE_X14Y111_C2;
  wire [0:0] CLBLM_R_X11Y111_SLICE_X14Y111_C3;
  wire [0:0] CLBLM_R_X11Y111_SLICE_X14Y111_C4;
  wire [0:0] CLBLM_R_X11Y111_SLICE_X14Y111_C5;
  wire [0:0] CLBLM_R_X11Y111_SLICE_X14Y111_C6;
  wire [0:0] CLBLM_R_X11Y111_SLICE_X14Y111_CO5;
  wire [0:0] CLBLM_R_X11Y111_SLICE_X14Y111_CO6;
  wire [0:0] CLBLM_R_X11Y111_SLICE_X14Y111_C_CY;
  wire [0:0] CLBLM_R_X11Y111_SLICE_X14Y111_C_XOR;
  wire [0:0] CLBLM_R_X11Y111_SLICE_X14Y111_D;
  wire [0:0] CLBLM_R_X11Y111_SLICE_X14Y111_D1;
  wire [0:0] CLBLM_R_X11Y111_SLICE_X14Y111_D2;
  wire [0:0] CLBLM_R_X11Y111_SLICE_X14Y111_D3;
  wire [0:0] CLBLM_R_X11Y111_SLICE_X14Y111_D4;
  wire [0:0] CLBLM_R_X11Y111_SLICE_X14Y111_D5;
  wire [0:0] CLBLM_R_X11Y111_SLICE_X14Y111_D6;
  wire [0:0] CLBLM_R_X11Y111_SLICE_X14Y111_DO5;
  wire [0:0] CLBLM_R_X11Y111_SLICE_X14Y111_DO6;
  wire [0:0] CLBLM_R_X11Y111_SLICE_X14Y111_D_CY;
  wire [0:0] CLBLM_R_X11Y111_SLICE_X14Y111_D_XOR;
  wire [0:0] CLBLM_R_X11Y111_SLICE_X15Y111_A;
  wire [0:0] CLBLM_R_X11Y111_SLICE_X15Y111_A1;
  wire [0:0] CLBLM_R_X11Y111_SLICE_X15Y111_A2;
  wire [0:0] CLBLM_R_X11Y111_SLICE_X15Y111_A3;
  wire [0:0] CLBLM_R_X11Y111_SLICE_X15Y111_A4;
  wire [0:0] CLBLM_R_X11Y111_SLICE_X15Y111_A5;
  wire [0:0] CLBLM_R_X11Y111_SLICE_X15Y111_A6;
  wire [0:0] CLBLM_R_X11Y111_SLICE_X15Y111_AMUX;
  wire [0:0] CLBLM_R_X11Y111_SLICE_X15Y111_AO5;
  wire [0:0] CLBLM_R_X11Y111_SLICE_X15Y111_AO6;
  wire [0:0] CLBLM_R_X11Y111_SLICE_X15Y111_A_CY;
  wire [0:0] CLBLM_R_X11Y111_SLICE_X15Y111_A_XOR;
  wire [0:0] CLBLM_R_X11Y111_SLICE_X15Y111_B;
  wire [0:0] CLBLM_R_X11Y111_SLICE_X15Y111_B1;
  wire [0:0] CLBLM_R_X11Y111_SLICE_X15Y111_B2;
  wire [0:0] CLBLM_R_X11Y111_SLICE_X15Y111_B3;
  wire [0:0] CLBLM_R_X11Y111_SLICE_X15Y111_B4;
  wire [0:0] CLBLM_R_X11Y111_SLICE_X15Y111_B5;
  wire [0:0] CLBLM_R_X11Y111_SLICE_X15Y111_B6;
  wire [0:0] CLBLM_R_X11Y111_SLICE_X15Y111_BMUX;
  wire [0:0] CLBLM_R_X11Y111_SLICE_X15Y111_BO5;
  wire [0:0] CLBLM_R_X11Y111_SLICE_X15Y111_BO6;
  wire [0:0] CLBLM_R_X11Y111_SLICE_X15Y111_B_CY;
  wire [0:0] CLBLM_R_X11Y111_SLICE_X15Y111_B_XOR;
  wire [0:0] CLBLM_R_X11Y111_SLICE_X15Y111_C;
  wire [0:0] CLBLM_R_X11Y111_SLICE_X15Y111_C1;
  wire [0:0] CLBLM_R_X11Y111_SLICE_X15Y111_C2;
  wire [0:0] CLBLM_R_X11Y111_SLICE_X15Y111_C3;
  wire [0:0] CLBLM_R_X11Y111_SLICE_X15Y111_C4;
  wire [0:0] CLBLM_R_X11Y111_SLICE_X15Y111_C5;
  wire [0:0] CLBLM_R_X11Y111_SLICE_X15Y111_C6;
  wire [0:0] CLBLM_R_X11Y111_SLICE_X15Y111_CO5;
  wire [0:0] CLBLM_R_X11Y111_SLICE_X15Y111_CO6;
  wire [0:0] CLBLM_R_X11Y111_SLICE_X15Y111_C_CY;
  wire [0:0] CLBLM_R_X11Y111_SLICE_X15Y111_C_XOR;
  wire [0:0] CLBLM_R_X11Y111_SLICE_X15Y111_D;
  wire [0:0] CLBLM_R_X11Y111_SLICE_X15Y111_D1;
  wire [0:0] CLBLM_R_X11Y111_SLICE_X15Y111_D2;
  wire [0:0] CLBLM_R_X11Y111_SLICE_X15Y111_D3;
  wire [0:0] CLBLM_R_X11Y111_SLICE_X15Y111_D4;
  wire [0:0] CLBLM_R_X11Y111_SLICE_X15Y111_D5;
  wire [0:0] CLBLM_R_X11Y111_SLICE_X15Y111_D6;
  wire [0:0] CLBLM_R_X11Y111_SLICE_X15Y111_DO5;
  wire [0:0] CLBLM_R_X11Y111_SLICE_X15Y111_DO6;
  wire [0:0] CLBLM_R_X11Y111_SLICE_X15Y111_D_CY;
  wire [0:0] CLBLM_R_X11Y111_SLICE_X15Y111_D_XOR;
  wire [0:0] CLBLM_R_X13Y105_SLICE_X18Y105_A;
  wire [0:0] CLBLM_R_X13Y105_SLICE_X18Y105_A1;
  wire [0:0] CLBLM_R_X13Y105_SLICE_X18Y105_A2;
  wire [0:0] CLBLM_R_X13Y105_SLICE_X18Y105_A3;
  wire [0:0] CLBLM_R_X13Y105_SLICE_X18Y105_A4;
  wire [0:0] CLBLM_R_X13Y105_SLICE_X18Y105_A5;
  wire [0:0] CLBLM_R_X13Y105_SLICE_X18Y105_A6;
  wire [0:0] CLBLM_R_X13Y105_SLICE_X18Y105_AO5;
  wire [0:0] CLBLM_R_X13Y105_SLICE_X18Y105_AO6;
  wire [0:0] CLBLM_R_X13Y105_SLICE_X18Y105_A_CY;
  wire [0:0] CLBLM_R_X13Y105_SLICE_X18Y105_A_XOR;
  wire [0:0] CLBLM_R_X13Y105_SLICE_X18Y105_B;
  wire [0:0] CLBLM_R_X13Y105_SLICE_X18Y105_B1;
  wire [0:0] CLBLM_R_X13Y105_SLICE_X18Y105_B2;
  wire [0:0] CLBLM_R_X13Y105_SLICE_X18Y105_B3;
  wire [0:0] CLBLM_R_X13Y105_SLICE_X18Y105_B4;
  wire [0:0] CLBLM_R_X13Y105_SLICE_X18Y105_B5;
  wire [0:0] CLBLM_R_X13Y105_SLICE_X18Y105_B6;
  wire [0:0] CLBLM_R_X13Y105_SLICE_X18Y105_BO5;
  wire [0:0] CLBLM_R_X13Y105_SLICE_X18Y105_BO6;
  wire [0:0] CLBLM_R_X13Y105_SLICE_X18Y105_B_CY;
  wire [0:0] CLBLM_R_X13Y105_SLICE_X18Y105_B_XOR;
  wire [0:0] CLBLM_R_X13Y105_SLICE_X18Y105_C;
  wire [0:0] CLBLM_R_X13Y105_SLICE_X18Y105_C1;
  wire [0:0] CLBLM_R_X13Y105_SLICE_X18Y105_C2;
  wire [0:0] CLBLM_R_X13Y105_SLICE_X18Y105_C3;
  wire [0:0] CLBLM_R_X13Y105_SLICE_X18Y105_C4;
  wire [0:0] CLBLM_R_X13Y105_SLICE_X18Y105_C5;
  wire [0:0] CLBLM_R_X13Y105_SLICE_X18Y105_C6;
  wire [0:0] CLBLM_R_X13Y105_SLICE_X18Y105_CO5;
  wire [0:0] CLBLM_R_X13Y105_SLICE_X18Y105_CO6;
  wire [0:0] CLBLM_R_X13Y105_SLICE_X18Y105_C_CY;
  wire [0:0] CLBLM_R_X13Y105_SLICE_X18Y105_C_XOR;
  wire [0:0] CLBLM_R_X13Y105_SLICE_X18Y105_D;
  wire [0:0] CLBLM_R_X13Y105_SLICE_X18Y105_D1;
  wire [0:0] CLBLM_R_X13Y105_SLICE_X18Y105_D2;
  wire [0:0] CLBLM_R_X13Y105_SLICE_X18Y105_D3;
  wire [0:0] CLBLM_R_X13Y105_SLICE_X18Y105_D4;
  wire [0:0] CLBLM_R_X13Y105_SLICE_X18Y105_D5;
  wire [0:0] CLBLM_R_X13Y105_SLICE_X18Y105_D6;
  wire [0:0] CLBLM_R_X13Y105_SLICE_X18Y105_DO5;
  wire [0:0] CLBLM_R_X13Y105_SLICE_X18Y105_DO6;
  wire [0:0] CLBLM_R_X13Y105_SLICE_X18Y105_D_CY;
  wire [0:0] CLBLM_R_X13Y105_SLICE_X18Y105_D_XOR;
  wire [0:0] CLBLM_R_X13Y105_SLICE_X19Y105_A;
  wire [0:0] CLBLM_R_X13Y105_SLICE_X19Y105_A1;
  wire [0:0] CLBLM_R_X13Y105_SLICE_X19Y105_A2;
  wire [0:0] CLBLM_R_X13Y105_SLICE_X19Y105_A3;
  wire [0:0] CLBLM_R_X13Y105_SLICE_X19Y105_A4;
  wire [0:0] CLBLM_R_X13Y105_SLICE_X19Y105_A5;
  wire [0:0] CLBLM_R_X13Y105_SLICE_X19Y105_A6;
  wire [0:0] CLBLM_R_X13Y105_SLICE_X19Y105_AO5;
  wire [0:0] CLBLM_R_X13Y105_SLICE_X19Y105_AO6;
  wire [0:0] CLBLM_R_X13Y105_SLICE_X19Y105_A_CY;
  wire [0:0] CLBLM_R_X13Y105_SLICE_X19Y105_A_XOR;
  wire [0:0] CLBLM_R_X13Y105_SLICE_X19Y105_B;
  wire [0:0] CLBLM_R_X13Y105_SLICE_X19Y105_B1;
  wire [0:0] CLBLM_R_X13Y105_SLICE_X19Y105_B2;
  wire [0:0] CLBLM_R_X13Y105_SLICE_X19Y105_B3;
  wire [0:0] CLBLM_R_X13Y105_SLICE_X19Y105_B4;
  wire [0:0] CLBLM_R_X13Y105_SLICE_X19Y105_B5;
  wire [0:0] CLBLM_R_X13Y105_SLICE_X19Y105_B6;
  wire [0:0] CLBLM_R_X13Y105_SLICE_X19Y105_BO5;
  wire [0:0] CLBLM_R_X13Y105_SLICE_X19Y105_BO6;
  wire [0:0] CLBLM_R_X13Y105_SLICE_X19Y105_B_CY;
  wire [0:0] CLBLM_R_X13Y105_SLICE_X19Y105_B_XOR;
  wire [0:0] CLBLM_R_X13Y105_SLICE_X19Y105_C;
  wire [0:0] CLBLM_R_X13Y105_SLICE_X19Y105_C1;
  wire [0:0] CLBLM_R_X13Y105_SLICE_X19Y105_C2;
  wire [0:0] CLBLM_R_X13Y105_SLICE_X19Y105_C3;
  wire [0:0] CLBLM_R_X13Y105_SLICE_X19Y105_C4;
  wire [0:0] CLBLM_R_X13Y105_SLICE_X19Y105_C5;
  wire [0:0] CLBLM_R_X13Y105_SLICE_X19Y105_C6;
  wire [0:0] CLBLM_R_X13Y105_SLICE_X19Y105_CO5;
  wire [0:0] CLBLM_R_X13Y105_SLICE_X19Y105_CO6;
  wire [0:0] CLBLM_R_X13Y105_SLICE_X19Y105_C_CY;
  wire [0:0] CLBLM_R_X13Y105_SLICE_X19Y105_C_XOR;
  wire [0:0] CLBLM_R_X13Y105_SLICE_X19Y105_D;
  wire [0:0] CLBLM_R_X13Y105_SLICE_X19Y105_D1;
  wire [0:0] CLBLM_R_X13Y105_SLICE_X19Y105_D2;
  wire [0:0] CLBLM_R_X13Y105_SLICE_X19Y105_D3;
  wire [0:0] CLBLM_R_X13Y105_SLICE_X19Y105_D4;
  wire [0:0] CLBLM_R_X13Y105_SLICE_X19Y105_D5;
  wire [0:0] CLBLM_R_X13Y105_SLICE_X19Y105_D6;
  wire [0:0] CLBLM_R_X13Y105_SLICE_X19Y105_DO5;
  wire [0:0] CLBLM_R_X13Y105_SLICE_X19Y105_DO6;
  wire [0:0] CLBLM_R_X13Y105_SLICE_X19Y105_D_CY;
  wire [0:0] CLBLM_R_X13Y105_SLICE_X19Y105_D_XOR;
  wire [0:0] CLBLM_R_X13Y106_SLICE_X18Y106_A;
  wire [0:0] CLBLM_R_X13Y106_SLICE_X18Y106_A1;
  wire [0:0] CLBLM_R_X13Y106_SLICE_X18Y106_A2;
  wire [0:0] CLBLM_R_X13Y106_SLICE_X18Y106_A3;
  wire [0:0] CLBLM_R_X13Y106_SLICE_X18Y106_A4;
  wire [0:0] CLBLM_R_X13Y106_SLICE_X18Y106_A5;
  wire [0:0] CLBLM_R_X13Y106_SLICE_X18Y106_A6;
  wire [0:0] CLBLM_R_X13Y106_SLICE_X18Y106_AMUX;
  wire [0:0] CLBLM_R_X13Y106_SLICE_X18Y106_AO5;
  wire [0:0] CLBLM_R_X13Y106_SLICE_X18Y106_AO6;
  wire [0:0] CLBLM_R_X13Y106_SLICE_X18Y106_A_CY;
  wire [0:0] CLBLM_R_X13Y106_SLICE_X18Y106_A_XOR;
  wire [0:0] CLBLM_R_X13Y106_SLICE_X18Y106_B;
  wire [0:0] CLBLM_R_X13Y106_SLICE_X18Y106_B1;
  wire [0:0] CLBLM_R_X13Y106_SLICE_X18Y106_B2;
  wire [0:0] CLBLM_R_X13Y106_SLICE_X18Y106_B3;
  wire [0:0] CLBLM_R_X13Y106_SLICE_X18Y106_B4;
  wire [0:0] CLBLM_R_X13Y106_SLICE_X18Y106_B5;
  wire [0:0] CLBLM_R_X13Y106_SLICE_X18Y106_B6;
  wire [0:0] CLBLM_R_X13Y106_SLICE_X18Y106_BO5;
  wire [0:0] CLBLM_R_X13Y106_SLICE_X18Y106_BO6;
  wire [0:0] CLBLM_R_X13Y106_SLICE_X18Y106_B_CY;
  wire [0:0] CLBLM_R_X13Y106_SLICE_X18Y106_B_XOR;
  wire [0:0] CLBLM_R_X13Y106_SLICE_X18Y106_C;
  wire [0:0] CLBLM_R_X13Y106_SLICE_X18Y106_C1;
  wire [0:0] CLBLM_R_X13Y106_SLICE_X18Y106_C2;
  wire [0:0] CLBLM_R_X13Y106_SLICE_X18Y106_C3;
  wire [0:0] CLBLM_R_X13Y106_SLICE_X18Y106_C4;
  wire [0:0] CLBLM_R_X13Y106_SLICE_X18Y106_C5;
  wire [0:0] CLBLM_R_X13Y106_SLICE_X18Y106_C6;
  wire [0:0] CLBLM_R_X13Y106_SLICE_X18Y106_CO5;
  wire [0:0] CLBLM_R_X13Y106_SLICE_X18Y106_CO6;
  wire [0:0] CLBLM_R_X13Y106_SLICE_X18Y106_C_CY;
  wire [0:0] CLBLM_R_X13Y106_SLICE_X18Y106_C_XOR;
  wire [0:0] CLBLM_R_X13Y106_SLICE_X18Y106_D;
  wire [0:0] CLBLM_R_X13Y106_SLICE_X18Y106_D1;
  wire [0:0] CLBLM_R_X13Y106_SLICE_X18Y106_D2;
  wire [0:0] CLBLM_R_X13Y106_SLICE_X18Y106_D3;
  wire [0:0] CLBLM_R_X13Y106_SLICE_X18Y106_D4;
  wire [0:0] CLBLM_R_X13Y106_SLICE_X18Y106_D5;
  wire [0:0] CLBLM_R_X13Y106_SLICE_X18Y106_D6;
  wire [0:0] CLBLM_R_X13Y106_SLICE_X18Y106_DO5;
  wire [0:0] CLBLM_R_X13Y106_SLICE_X18Y106_DO6;
  wire [0:0] CLBLM_R_X13Y106_SLICE_X18Y106_D_CY;
  wire [0:0] CLBLM_R_X13Y106_SLICE_X18Y106_D_XOR;
  wire [0:0] CLBLM_R_X13Y106_SLICE_X19Y106_A;
  wire [0:0] CLBLM_R_X13Y106_SLICE_X19Y106_A1;
  wire [0:0] CLBLM_R_X13Y106_SLICE_X19Y106_A2;
  wire [0:0] CLBLM_R_X13Y106_SLICE_X19Y106_A3;
  wire [0:0] CLBLM_R_X13Y106_SLICE_X19Y106_A4;
  wire [0:0] CLBLM_R_X13Y106_SLICE_X19Y106_A5;
  wire [0:0] CLBLM_R_X13Y106_SLICE_X19Y106_A6;
  wire [0:0] CLBLM_R_X13Y106_SLICE_X19Y106_AMUX;
  wire [0:0] CLBLM_R_X13Y106_SLICE_X19Y106_AO5;
  wire [0:0] CLBLM_R_X13Y106_SLICE_X19Y106_AO6;
  wire [0:0] CLBLM_R_X13Y106_SLICE_X19Y106_A_CY;
  wire [0:0] CLBLM_R_X13Y106_SLICE_X19Y106_A_XOR;
  wire [0:0] CLBLM_R_X13Y106_SLICE_X19Y106_B;
  wire [0:0] CLBLM_R_X13Y106_SLICE_X19Y106_B1;
  wire [0:0] CLBLM_R_X13Y106_SLICE_X19Y106_B2;
  wire [0:0] CLBLM_R_X13Y106_SLICE_X19Y106_B3;
  wire [0:0] CLBLM_R_X13Y106_SLICE_X19Y106_B4;
  wire [0:0] CLBLM_R_X13Y106_SLICE_X19Y106_B5;
  wire [0:0] CLBLM_R_X13Y106_SLICE_X19Y106_B6;
  wire [0:0] CLBLM_R_X13Y106_SLICE_X19Y106_BMUX;
  wire [0:0] CLBLM_R_X13Y106_SLICE_X19Y106_BO5;
  wire [0:0] CLBLM_R_X13Y106_SLICE_X19Y106_BO6;
  wire [0:0] CLBLM_R_X13Y106_SLICE_X19Y106_B_CY;
  wire [0:0] CLBLM_R_X13Y106_SLICE_X19Y106_B_XOR;
  wire [0:0] CLBLM_R_X13Y106_SLICE_X19Y106_C;
  wire [0:0] CLBLM_R_X13Y106_SLICE_X19Y106_C1;
  wire [0:0] CLBLM_R_X13Y106_SLICE_X19Y106_C2;
  wire [0:0] CLBLM_R_X13Y106_SLICE_X19Y106_C3;
  wire [0:0] CLBLM_R_X13Y106_SLICE_X19Y106_C4;
  wire [0:0] CLBLM_R_X13Y106_SLICE_X19Y106_C5;
  wire [0:0] CLBLM_R_X13Y106_SLICE_X19Y106_C6;
  wire [0:0] CLBLM_R_X13Y106_SLICE_X19Y106_CMUX;
  wire [0:0] CLBLM_R_X13Y106_SLICE_X19Y106_CO5;
  wire [0:0] CLBLM_R_X13Y106_SLICE_X19Y106_CO6;
  wire [0:0] CLBLM_R_X13Y106_SLICE_X19Y106_C_CY;
  wire [0:0] CLBLM_R_X13Y106_SLICE_X19Y106_C_XOR;
  wire [0:0] CLBLM_R_X13Y106_SLICE_X19Y106_D;
  wire [0:0] CLBLM_R_X13Y106_SLICE_X19Y106_D1;
  wire [0:0] CLBLM_R_X13Y106_SLICE_X19Y106_D2;
  wire [0:0] CLBLM_R_X13Y106_SLICE_X19Y106_D3;
  wire [0:0] CLBLM_R_X13Y106_SLICE_X19Y106_D4;
  wire [0:0] CLBLM_R_X13Y106_SLICE_X19Y106_D5;
  wire [0:0] CLBLM_R_X13Y106_SLICE_X19Y106_D6;
  wire [0:0] CLBLM_R_X13Y106_SLICE_X19Y106_DO5;
  wire [0:0] CLBLM_R_X13Y106_SLICE_X19Y106_DO6;
  wire [0:0] CLBLM_R_X13Y106_SLICE_X19Y106_D_CY;
  wire [0:0] CLBLM_R_X13Y106_SLICE_X19Y106_D_XOR;
  wire [0:0] CLBLM_R_X13Y107_SLICE_X18Y107_A;
  wire [0:0] CLBLM_R_X13Y107_SLICE_X18Y107_A1;
  wire [0:0] CLBLM_R_X13Y107_SLICE_X18Y107_A2;
  wire [0:0] CLBLM_R_X13Y107_SLICE_X18Y107_A3;
  wire [0:0] CLBLM_R_X13Y107_SLICE_X18Y107_A4;
  wire [0:0] CLBLM_R_X13Y107_SLICE_X18Y107_A5;
  wire [0:0] CLBLM_R_X13Y107_SLICE_X18Y107_A6;
  wire [0:0] CLBLM_R_X13Y107_SLICE_X18Y107_AO5;
  wire [0:0] CLBLM_R_X13Y107_SLICE_X18Y107_AO6;
  wire [0:0] CLBLM_R_X13Y107_SLICE_X18Y107_A_CY;
  wire [0:0] CLBLM_R_X13Y107_SLICE_X18Y107_A_XOR;
  wire [0:0] CLBLM_R_X13Y107_SLICE_X18Y107_B;
  wire [0:0] CLBLM_R_X13Y107_SLICE_X18Y107_B1;
  wire [0:0] CLBLM_R_X13Y107_SLICE_X18Y107_B2;
  wire [0:0] CLBLM_R_X13Y107_SLICE_X18Y107_B3;
  wire [0:0] CLBLM_R_X13Y107_SLICE_X18Y107_B4;
  wire [0:0] CLBLM_R_X13Y107_SLICE_X18Y107_B5;
  wire [0:0] CLBLM_R_X13Y107_SLICE_X18Y107_B6;
  wire [0:0] CLBLM_R_X13Y107_SLICE_X18Y107_BO5;
  wire [0:0] CLBLM_R_X13Y107_SLICE_X18Y107_BO6;
  wire [0:0] CLBLM_R_X13Y107_SLICE_X18Y107_B_CY;
  wire [0:0] CLBLM_R_X13Y107_SLICE_X18Y107_B_XOR;
  wire [0:0] CLBLM_R_X13Y107_SLICE_X18Y107_C;
  wire [0:0] CLBLM_R_X13Y107_SLICE_X18Y107_C1;
  wire [0:0] CLBLM_R_X13Y107_SLICE_X18Y107_C2;
  wire [0:0] CLBLM_R_X13Y107_SLICE_X18Y107_C3;
  wire [0:0] CLBLM_R_X13Y107_SLICE_X18Y107_C4;
  wire [0:0] CLBLM_R_X13Y107_SLICE_X18Y107_C5;
  wire [0:0] CLBLM_R_X13Y107_SLICE_X18Y107_C6;
  wire [0:0] CLBLM_R_X13Y107_SLICE_X18Y107_CO5;
  wire [0:0] CLBLM_R_X13Y107_SLICE_X18Y107_CO6;
  wire [0:0] CLBLM_R_X13Y107_SLICE_X18Y107_C_CY;
  wire [0:0] CLBLM_R_X13Y107_SLICE_X18Y107_C_XOR;
  wire [0:0] CLBLM_R_X13Y107_SLICE_X18Y107_D;
  wire [0:0] CLBLM_R_X13Y107_SLICE_X18Y107_D1;
  wire [0:0] CLBLM_R_X13Y107_SLICE_X18Y107_D2;
  wire [0:0] CLBLM_R_X13Y107_SLICE_X18Y107_D3;
  wire [0:0] CLBLM_R_X13Y107_SLICE_X18Y107_D4;
  wire [0:0] CLBLM_R_X13Y107_SLICE_X18Y107_D5;
  wire [0:0] CLBLM_R_X13Y107_SLICE_X18Y107_D6;
  wire [0:0] CLBLM_R_X13Y107_SLICE_X18Y107_DO5;
  wire [0:0] CLBLM_R_X13Y107_SLICE_X18Y107_DO6;
  wire [0:0] CLBLM_R_X13Y107_SLICE_X18Y107_D_CY;
  wire [0:0] CLBLM_R_X13Y107_SLICE_X18Y107_D_XOR;
  wire [0:0] CLBLM_R_X13Y107_SLICE_X19Y107_A;
  wire [0:0] CLBLM_R_X13Y107_SLICE_X19Y107_A1;
  wire [0:0] CLBLM_R_X13Y107_SLICE_X19Y107_A2;
  wire [0:0] CLBLM_R_X13Y107_SLICE_X19Y107_A3;
  wire [0:0] CLBLM_R_X13Y107_SLICE_X19Y107_A4;
  wire [0:0] CLBLM_R_X13Y107_SLICE_X19Y107_A5;
  wire [0:0] CLBLM_R_X13Y107_SLICE_X19Y107_A6;
  wire [0:0] CLBLM_R_X13Y107_SLICE_X19Y107_AO5;
  wire [0:0] CLBLM_R_X13Y107_SLICE_X19Y107_AO6;
  wire [0:0] CLBLM_R_X13Y107_SLICE_X19Y107_A_CY;
  wire [0:0] CLBLM_R_X13Y107_SLICE_X19Y107_A_XOR;
  wire [0:0] CLBLM_R_X13Y107_SLICE_X19Y107_B;
  wire [0:0] CLBLM_R_X13Y107_SLICE_X19Y107_B1;
  wire [0:0] CLBLM_R_X13Y107_SLICE_X19Y107_B2;
  wire [0:0] CLBLM_R_X13Y107_SLICE_X19Y107_B3;
  wire [0:0] CLBLM_R_X13Y107_SLICE_X19Y107_B4;
  wire [0:0] CLBLM_R_X13Y107_SLICE_X19Y107_B5;
  wire [0:0] CLBLM_R_X13Y107_SLICE_X19Y107_B6;
  wire [0:0] CLBLM_R_X13Y107_SLICE_X19Y107_BO5;
  wire [0:0] CLBLM_R_X13Y107_SLICE_X19Y107_BO6;
  wire [0:0] CLBLM_R_X13Y107_SLICE_X19Y107_B_CY;
  wire [0:0] CLBLM_R_X13Y107_SLICE_X19Y107_B_XOR;
  wire [0:0] CLBLM_R_X13Y107_SLICE_X19Y107_C;
  wire [0:0] CLBLM_R_X13Y107_SLICE_X19Y107_C1;
  wire [0:0] CLBLM_R_X13Y107_SLICE_X19Y107_C2;
  wire [0:0] CLBLM_R_X13Y107_SLICE_X19Y107_C3;
  wire [0:0] CLBLM_R_X13Y107_SLICE_X19Y107_C4;
  wire [0:0] CLBLM_R_X13Y107_SLICE_X19Y107_C5;
  wire [0:0] CLBLM_R_X13Y107_SLICE_X19Y107_C6;
  wire [0:0] CLBLM_R_X13Y107_SLICE_X19Y107_CO5;
  wire [0:0] CLBLM_R_X13Y107_SLICE_X19Y107_CO6;
  wire [0:0] CLBLM_R_X13Y107_SLICE_X19Y107_C_CY;
  wire [0:0] CLBLM_R_X13Y107_SLICE_X19Y107_C_XOR;
  wire [0:0] CLBLM_R_X13Y107_SLICE_X19Y107_D;
  wire [0:0] CLBLM_R_X13Y107_SLICE_X19Y107_D1;
  wire [0:0] CLBLM_R_X13Y107_SLICE_X19Y107_D2;
  wire [0:0] CLBLM_R_X13Y107_SLICE_X19Y107_D3;
  wire [0:0] CLBLM_R_X13Y107_SLICE_X19Y107_D4;
  wire [0:0] CLBLM_R_X13Y107_SLICE_X19Y107_D5;
  wire [0:0] CLBLM_R_X13Y107_SLICE_X19Y107_D6;
  wire [0:0] CLBLM_R_X13Y107_SLICE_X19Y107_DO5;
  wire [0:0] CLBLM_R_X13Y107_SLICE_X19Y107_DO6;
  wire [0:0] CLBLM_R_X13Y107_SLICE_X19Y107_D_CY;
  wire [0:0] CLBLM_R_X13Y107_SLICE_X19Y107_D_XOR;
  wire [0:0] CLBLM_R_X3Y103_SLICE_X2Y103_A;
  wire [0:0] CLBLM_R_X3Y103_SLICE_X2Y103_A1;
  wire [0:0] CLBLM_R_X3Y103_SLICE_X2Y103_A2;
  wire [0:0] CLBLM_R_X3Y103_SLICE_X2Y103_A3;
  wire [0:0] CLBLM_R_X3Y103_SLICE_X2Y103_A4;
  wire [0:0] CLBLM_R_X3Y103_SLICE_X2Y103_A5;
  wire [0:0] CLBLM_R_X3Y103_SLICE_X2Y103_A6;
  wire [0:0] CLBLM_R_X3Y103_SLICE_X2Y103_AO5;
  wire [0:0] CLBLM_R_X3Y103_SLICE_X2Y103_AO6;
  wire [0:0] CLBLM_R_X3Y103_SLICE_X2Y103_A_CY;
  wire [0:0] CLBLM_R_X3Y103_SLICE_X2Y103_A_XOR;
  wire [0:0] CLBLM_R_X3Y103_SLICE_X2Y103_B;
  wire [0:0] CLBLM_R_X3Y103_SLICE_X2Y103_B1;
  wire [0:0] CLBLM_R_X3Y103_SLICE_X2Y103_B2;
  wire [0:0] CLBLM_R_X3Y103_SLICE_X2Y103_B3;
  wire [0:0] CLBLM_R_X3Y103_SLICE_X2Y103_B4;
  wire [0:0] CLBLM_R_X3Y103_SLICE_X2Y103_B5;
  wire [0:0] CLBLM_R_X3Y103_SLICE_X2Y103_B6;
  wire [0:0] CLBLM_R_X3Y103_SLICE_X2Y103_BO5;
  wire [0:0] CLBLM_R_X3Y103_SLICE_X2Y103_BO6;
  wire [0:0] CLBLM_R_X3Y103_SLICE_X2Y103_B_CY;
  wire [0:0] CLBLM_R_X3Y103_SLICE_X2Y103_B_XOR;
  wire [0:0] CLBLM_R_X3Y103_SLICE_X2Y103_C;
  wire [0:0] CLBLM_R_X3Y103_SLICE_X2Y103_C1;
  wire [0:0] CLBLM_R_X3Y103_SLICE_X2Y103_C2;
  wire [0:0] CLBLM_R_X3Y103_SLICE_X2Y103_C3;
  wire [0:0] CLBLM_R_X3Y103_SLICE_X2Y103_C4;
  wire [0:0] CLBLM_R_X3Y103_SLICE_X2Y103_C5;
  wire [0:0] CLBLM_R_X3Y103_SLICE_X2Y103_C6;
  wire [0:0] CLBLM_R_X3Y103_SLICE_X2Y103_CO5;
  wire [0:0] CLBLM_R_X3Y103_SLICE_X2Y103_CO6;
  wire [0:0] CLBLM_R_X3Y103_SLICE_X2Y103_C_CY;
  wire [0:0] CLBLM_R_X3Y103_SLICE_X2Y103_C_XOR;
  wire [0:0] CLBLM_R_X3Y103_SLICE_X2Y103_D;
  wire [0:0] CLBLM_R_X3Y103_SLICE_X2Y103_D1;
  wire [0:0] CLBLM_R_X3Y103_SLICE_X2Y103_D2;
  wire [0:0] CLBLM_R_X3Y103_SLICE_X2Y103_D3;
  wire [0:0] CLBLM_R_X3Y103_SLICE_X2Y103_D4;
  wire [0:0] CLBLM_R_X3Y103_SLICE_X2Y103_D5;
  wire [0:0] CLBLM_R_X3Y103_SLICE_X2Y103_D6;
  wire [0:0] CLBLM_R_X3Y103_SLICE_X2Y103_DO5;
  wire [0:0] CLBLM_R_X3Y103_SLICE_X2Y103_DO6;
  wire [0:0] CLBLM_R_X3Y103_SLICE_X2Y103_D_CY;
  wire [0:0] CLBLM_R_X3Y103_SLICE_X2Y103_D_XOR;
  wire [0:0] CLBLM_R_X3Y103_SLICE_X3Y103_A;
  wire [0:0] CLBLM_R_X3Y103_SLICE_X3Y103_A1;
  wire [0:0] CLBLM_R_X3Y103_SLICE_X3Y103_A2;
  wire [0:0] CLBLM_R_X3Y103_SLICE_X3Y103_A3;
  wire [0:0] CLBLM_R_X3Y103_SLICE_X3Y103_A4;
  wire [0:0] CLBLM_R_X3Y103_SLICE_X3Y103_A5;
  wire [0:0] CLBLM_R_X3Y103_SLICE_X3Y103_A6;
  wire [0:0] CLBLM_R_X3Y103_SLICE_X3Y103_AMUX;
  wire [0:0] CLBLM_R_X3Y103_SLICE_X3Y103_AO5;
  wire [0:0] CLBLM_R_X3Y103_SLICE_X3Y103_AO6;
  wire [0:0] CLBLM_R_X3Y103_SLICE_X3Y103_A_CY;
  wire [0:0] CLBLM_R_X3Y103_SLICE_X3Y103_A_XOR;
  wire [0:0] CLBLM_R_X3Y103_SLICE_X3Y103_B;
  wire [0:0] CLBLM_R_X3Y103_SLICE_X3Y103_B1;
  wire [0:0] CLBLM_R_X3Y103_SLICE_X3Y103_B2;
  wire [0:0] CLBLM_R_X3Y103_SLICE_X3Y103_B3;
  wire [0:0] CLBLM_R_X3Y103_SLICE_X3Y103_B4;
  wire [0:0] CLBLM_R_X3Y103_SLICE_X3Y103_B5;
  wire [0:0] CLBLM_R_X3Y103_SLICE_X3Y103_B6;
  wire [0:0] CLBLM_R_X3Y103_SLICE_X3Y103_BO5;
  wire [0:0] CLBLM_R_X3Y103_SLICE_X3Y103_BO6;
  wire [0:0] CLBLM_R_X3Y103_SLICE_X3Y103_B_CY;
  wire [0:0] CLBLM_R_X3Y103_SLICE_X3Y103_B_XOR;
  wire [0:0] CLBLM_R_X3Y103_SLICE_X3Y103_C;
  wire [0:0] CLBLM_R_X3Y103_SLICE_X3Y103_C1;
  wire [0:0] CLBLM_R_X3Y103_SLICE_X3Y103_C2;
  wire [0:0] CLBLM_R_X3Y103_SLICE_X3Y103_C3;
  wire [0:0] CLBLM_R_X3Y103_SLICE_X3Y103_C4;
  wire [0:0] CLBLM_R_X3Y103_SLICE_X3Y103_C5;
  wire [0:0] CLBLM_R_X3Y103_SLICE_X3Y103_C6;
  wire [0:0] CLBLM_R_X3Y103_SLICE_X3Y103_CO5;
  wire [0:0] CLBLM_R_X3Y103_SLICE_X3Y103_CO6;
  wire [0:0] CLBLM_R_X3Y103_SLICE_X3Y103_C_CY;
  wire [0:0] CLBLM_R_X3Y103_SLICE_X3Y103_C_XOR;
  wire [0:0] CLBLM_R_X3Y103_SLICE_X3Y103_D;
  wire [0:0] CLBLM_R_X3Y103_SLICE_X3Y103_D1;
  wire [0:0] CLBLM_R_X3Y103_SLICE_X3Y103_D2;
  wire [0:0] CLBLM_R_X3Y103_SLICE_X3Y103_D3;
  wire [0:0] CLBLM_R_X3Y103_SLICE_X3Y103_D4;
  wire [0:0] CLBLM_R_X3Y103_SLICE_X3Y103_D5;
  wire [0:0] CLBLM_R_X3Y103_SLICE_X3Y103_D6;
  wire [0:0] CLBLM_R_X3Y103_SLICE_X3Y103_DO5;
  wire [0:0] CLBLM_R_X3Y103_SLICE_X3Y103_DO6;
  wire [0:0] CLBLM_R_X3Y103_SLICE_X3Y103_D_CY;
  wire [0:0] CLBLM_R_X3Y103_SLICE_X3Y103_D_XOR;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X2Y104_A;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X2Y104_A1;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X2Y104_A2;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X2Y104_A3;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X2Y104_A4;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X2Y104_A5;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X2Y104_A6;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X2Y104_AMUX;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X2Y104_AO5;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X2Y104_AO6;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X2Y104_A_CY;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X2Y104_A_XOR;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X2Y104_B;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X2Y104_B1;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X2Y104_B2;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X2Y104_B3;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X2Y104_B4;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X2Y104_B5;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X2Y104_B6;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X2Y104_BO5;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X2Y104_BO6;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X2Y104_B_CY;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X2Y104_B_XOR;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X2Y104_C;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X2Y104_C1;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X2Y104_C2;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X2Y104_C3;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X2Y104_C4;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X2Y104_C5;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X2Y104_C6;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X2Y104_CO5;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X2Y104_CO6;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X2Y104_C_CY;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X2Y104_C_XOR;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X2Y104_D;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X2Y104_D1;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X2Y104_D2;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X2Y104_D3;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X2Y104_D4;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X2Y104_D5;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X2Y104_D6;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X2Y104_DO5;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X2Y104_DO6;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X2Y104_D_CY;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X2Y104_D_XOR;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X3Y104_A;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X3Y104_A1;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X3Y104_A2;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X3Y104_A3;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X3Y104_A4;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X3Y104_A5;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X3Y104_A6;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X3Y104_AMUX;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X3Y104_AO5;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X3Y104_AO6;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X3Y104_A_CY;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X3Y104_A_XOR;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X3Y104_B;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X3Y104_B1;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X3Y104_B2;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X3Y104_B3;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X3Y104_B4;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X3Y104_B5;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X3Y104_B6;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X3Y104_BO5;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X3Y104_BO6;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X3Y104_B_CY;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X3Y104_B_XOR;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X3Y104_C;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X3Y104_C1;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X3Y104_C2;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X3Y104_C3;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X3Y104_C4;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X3Y104_C5;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X3Y104_C6;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X3Y104_CO5;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X3Y104_CO6;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X3Y104_C_CY;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X3Y104_C_XOR;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X3Y104_D;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X3Y104_D1;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X3Y104_D2;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X3Y104_D3;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X3Y104_D4;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X3Y104_D5;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X3Y104_D6;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X3Y104_DO5;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X3Y104_DO6;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X3Y104_D_CY;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X3Y104_D_XOR;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X2Y105_A;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X2Y105_A1;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X2Y105_A2;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X2Y105_A3;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X2Y105_A4;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X2Y105_A5;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X2Y105_A6;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X2Y105_AO5;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X2Y105_AO6;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X2Y105_A_CY;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X2Y105_A_XOR;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X2Y105_B;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X2Y105_B1;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X2Y105_B2;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X2Y105_B3;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X2Y105_B4;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X2Y105_B5;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X2Y105_B6;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X2Y105_BO5;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X2Y105_BO6;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X2Y105_B_CY;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X2Y105_B_XOR;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X2Y105_C;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X2Y105_C1;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X2Y105_C2;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X2Y105_C3;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X2Y105_C4;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X2Y105_C5;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X2Y105_C6;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X2Y105_CO5;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X2Y105_CO6;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X2Y105_C_CY;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X2Y105_C_XOR;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X2Y105_D;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X2Y105_D1;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X2Y105_D2;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X2Y105_D3;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X2Y105_D4;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X2Y105_D5;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X2Y105_D6;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X2Y105_DO5;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X2Y105_DO6;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X2Y105_D_CY;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X2Y105_D_XOR;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X3Y105_A;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X3Y105_A1;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X3Y105_A2;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X3Y105_A3;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X3Y105_A4;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X3Y105_A5;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X3Y105_A6;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X3Y105_AO5;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X3Y105_AO6;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X3Y105_A_CY;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X3Y105_A_XOR;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X3Y105_B;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X3Y105_B1;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X3Y105_B2;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X3Y105_B3;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X3Y105_B4;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X3Y105_B5;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X3Y105_B6;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X3Y105_BO5;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X3Y105_BO6;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X3Y105_B_CY;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X3Y105_B_XOR;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X3Y105_C;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X3Y105_C1;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X3Y105_C2;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X3Y105_C3;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X3Y105_C4;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X3Y105_C5;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X3Y105_C6;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X3Y105_CO5;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X3Y105_CO6;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X3Y105_C_CY;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X3Y105_C_XOR;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X3Y105_D;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X3Y105_D1;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X3Y105_D2;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X3Y105_D3;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X3Y105_D4;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X3Y105_D5;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X3Y105_D6;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X3Y105_DO5;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X3Y105_DO6;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X3Y105_D_CY;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X3Y105_D_XOR;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X2Y106_A;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X2Y106_A1;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X2Y106_A2;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X2Y106_A3;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X2Y106_A4;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X2Y106_A5;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X2Y106_A6;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X2Y106_AMUX;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X2Y106_AO5;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X2Y106_AO6;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X2Y106_A_CY;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X2Y106_A_XOR;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X2Y106_B;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X2Y106_B1;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X2Y106_B2;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X2Y106_B3;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X2Y106_B4;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X2Y106_B5;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X2Y106_B6;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X2Y106_BMUX;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X2Y106_BO5;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X2Y106_BO6;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X2Y106_B_CY;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X2Y106_B_XOR;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X2Y106_C;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X2Y106_C1;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X2Y106_C2;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X2Y106_C3;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X2Y106_C4;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X2Y106_C5;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X2Y106_C6;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X2Y106_CO5;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X2Y106_CO6;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X2Y106_C_CY;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X2Y106_C_XOR;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X2Y106_D;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X2Y106_D1;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X2Y106_D2;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X2Y106_D3;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X2Y106_D4;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X2Y106_D5;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X2Y106_D6;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X2Y106_DO5;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X2Y106_DO6;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X2Y106_D_CY;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X2Y106_D_XOR;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X3Y106_A;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X3Y106_A1;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X3Y106_A2;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X3Y106_A3;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X3Y106_A4;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X3Y106_A5;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X3Y106_A6;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X3Y106_AMUX;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X3Y106_AO5;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X3Y106_AO6;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X3Y106_A_CY;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X3Y106_A_XOR;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X3Y106_B;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X3Y106_B1;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X3Y106_B2;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X3Y106_B3;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X3Y106_B4;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X3Y106_B5;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X3Y106_B6;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X3Y106_BO5;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X3Y106_BO6;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X3Y106_B_CY;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X3Y106_B_XOR;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X3Y106_C;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X3Y106_C1;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X3Y106_C2;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X3Y106_C3;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X3Y106_C4;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X3Y106_C5;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X3Y106_C6;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X3Y106_CO5;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X3Y106_CO6;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X3Y106_C_CY;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X3Y106_C_XOR;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X3Y106_D;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X3Y106_D1;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X3Y106_D2;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X3Y106_D3;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X3Y106_D4;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X3Y106_D5;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X3Y106_D6;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X3Y106_DO5;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X3Y106_DO6;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X3Y106_D_CY;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X3Y106_D_XOR;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X2Y107_A;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X2Y107_A1;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X2Y107_A2;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X2Y107_A3;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X2Y107_A4;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X2Y107_A5;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X2Y107_A6;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X2Y107_AMUX;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X2Y107_AO5;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X2Y107_AO6;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X2Y107_A_CY;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X2Y107_A_XOR;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X2Y107_B;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X2Y107_B1;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X2Y107_B2;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X2Y107_B3;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X2Y107_B4;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X2Y107_B5;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X2Y107_B6;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X2Y107_BO5;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X2Y107_BO6;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X2Y107_B_CY;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X2Y107_B_XOR;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X2Y107_C;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X2Y107_C1;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X2Y107_C2;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X2Y107_C3;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X2Y107_C4;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X2Y107_C5;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X2Y107_C6;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X2Y107_CO5;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X2Y107_CO6;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X2Y107_C_CY;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X2Y107_C_XOR;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X2Y107_D;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X2Y107_D1;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X2Y107_D2;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X2Y107_D3;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X2Y107_D4;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X2Y107_D5;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X2Y107_D6;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X2Y107_DO5;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X2Y107_DO6;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X2Y107_D_CY;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X2Y107_D_XOR;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X3Y107_A;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X3Y107_A1;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X3Y107_A2;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X3Y107_A3;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X3Y107_A4;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X3Y107_A5;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X3Y107_A6;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X3Y107_AMUX;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X3Y107_AO5;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X3Y107_AO6;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X3Y107_A_CY;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X3Y107_A_XOR;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X3Y107_B;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X3Y107_B1;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X3Y107_B2;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X3Y107_B3;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X3Y107_B4;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X3Y107_B5;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X3Y107_B6;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X3Y107_BMUX;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X3Y107_BO5;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X3Y107_BO6;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X3Y107_B_CY;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X3Y107_B_XOR;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X3Y107_C;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X3Y107_C1;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X3Y107_C2;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X3Y107_C3;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X3Y107_C4;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X3Y107_C5;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X3Y107_C6;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X3Y107_CMUX;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X3Y107_CO5;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X3Y107_CO6;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X3Y107_C_CY;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X3Y107_C_XOR;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X3Y107_D;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X3Y107_D1;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X3Y107_D2;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X3Y107_D3;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X3Y107_D4;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X3Y107_D5;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X3Y107_D6;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X3Y107_DO5;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X3Y107_DO6;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X3Y107_D_CY;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X3Y107_D_XOR;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X2Y108_A;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X2Y108_A1;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X2Y108_A2;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X2Y108_A3;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X2Y108_A4;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X2Y108_A5;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X2Y108_A6;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X2Y108_AO5;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X2Y108_AO6;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X2Y108_A_CY;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X2Y108_A_XOR;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X2Y108_B;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X2Y108_B1;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X2Y108_B2;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X2Y108_B3;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X2Y108_B4;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X2Y108_B5;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X2Y108_B6;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X2Y108_BO5;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X2Y108_BO6;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X2Y108_B_CY;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X2Y108_B_XOR;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X2Y108_C;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X2Y108_C1;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X2Y108_C2;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X2Y108_C3;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X2Y108_C4;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X2Y108_C5;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X2Y108_C6;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X2Y108_CO5;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X2Y108_CO6;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X2Y108_C_CY;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X2Y108_C_XOR;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X2Y108_D;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X2Y108_D1;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X2Y108_D2;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X2Y108_D3;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X2Y108_D4;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X2Y108_D5;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X2Y108_D6;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X2Y108_DO5;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X2Y108_DO6;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X2Y108_D_CY;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X2Y108_D_XOR;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X3Y108_A;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X3Y108_A1;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X3Y108_A2;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X3Y108_A3;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X3Y108_A4;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X3Y108_A5;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X3Y108_A6;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X3Y108_AO5;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X3Y108_AO6;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X3Y108_A_CY;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X3Y108_A_XOR;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X3Y108_B;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X3Y108_B1;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X3Y108_B2;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X3Y108_B3;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X3Y108_B4;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X3Y108_B5;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X3Y108_B6;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X3Y108_BO5;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X3Y108_BO6;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X3Y108_B_CY;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X3Y108_B_XOR;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X3Y108_C;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X3Y108_C1;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X3Y108_C2;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X3Y108_C3;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X3Y108_C4;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X3Y108_C5;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X3Y108_C6;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X3Y108_CO5;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X3Y108_CO6;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X3Y108_C_CY;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X3Y108_C_XOR;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X3Y108_D;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X3Y108_D1;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X3Y108_D2;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X3Y108_D3;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X3Y108_D4;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X3Y108_D5;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X3Y108_D6;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X3Y108_DO5;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X3Y108_DO6;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X3Y108_D_CY;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X3Y108_D_XOR;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X2Y109_A;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X2Y109_A1;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X2Y109_A2;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X2Y109_A3;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X2Y109_A4;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X2Y109_A5;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X2Y109_A6;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X2Y109_AO5;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X2Y109_AO6;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X2Y109_A_CY;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X2Y109_A_XOR;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X2Y109_B;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X2Y109_B1;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X2Y109_B2;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X2Y109_B3;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X2Y109_B4;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X2Y109_B5;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X2Y109_B6;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X2Y109_BO5;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X2Y109_BO6;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X2Y109_B_CY;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X2Y109_B_XOR;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X2Y109_C;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X2Y109_C1;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X2Y109_C2;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X2Y109_C3;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X2Y109_C4;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X2Y109_C5;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X2Y109_C6;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X2Y109_CO5;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X2Y109_CO6;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X2Y109_C_CY;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X2Y109_C_XOR;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X2Y109_D;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X2Y109_D1;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X2Y109_D2;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X2Y109_D3;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X2Y109_D4;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X2Y109_D5;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X2Y109_D6;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X2Y109_DO5;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X2Y109_DO6;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X2Y109_D_CY;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X2Y109_D_XOR;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X3Y109_A;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X3Y109_A1;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X3Y109_A2;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X3Y109_A3;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X3Y109_A4;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X3Y109_A5;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X3Y109_A6;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X3Y109_AO5;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X3Y109_AO6;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X3Y109_A_CY;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X3Y109_A_XOR;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X3Y109_B;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X3Y109_B1;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X3Y109_B2;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X3Y109_B3;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X3Y109_B4;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X3Y109_B5;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X3Y109_B6;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X3Y109_BO5;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X3Y109_BO6;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X3Y109_B_CY;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X3Y109_B_XOR;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X3Y109_C;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X3Y109_C1;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X3Y109_C2;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X3Y109_C3;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X3Y109_C4;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X3Y109_C5;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X3Y109_C6;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X3Y109_CO5;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X3Y109_CO6;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X3Y109_C_CY;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X3Y109_C_XOR;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X3Y109_D;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X3Y109_D1;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X3Y109_D2;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X3Y109_D3;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X3Y109_D4;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X3Y109_D5;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X3Y109_D6;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X3Y109_DO5;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X3Y109_DO6;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X3Y109_D_CY;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X3Y109_D_XOR;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X2Y112_A;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X2Y112_A1;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X2Y112_A2;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X2Y112_A3;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X2Y112_A4;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X2Y112_A5;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X2Y112_A6;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X2Y112_AMUX;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X2Y112_AO5;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X2Y112_AO6;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X2Y112_A_CY;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X2Y112_A_XOR;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X2Y112_B;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X2Y112_B1;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X2Y112_B2;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X2Y112_B3;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X2Y112_B4;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X2Y112_B5;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X2Y112_B6;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X2Y112_BMUX;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X2Y112_BO5;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X2Y112_BO6;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X2Y112_B_CY;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X2Y112_B_XOR;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X2Y112_C;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X2Y112_C1;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X2Y112_C2;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X2Y112_C3;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X2Y112_C4;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X2Y112_C5;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X2Y112_C6;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X2Y112_CO5;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X2Y112_CO6;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X2Y112_C_CY;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X2Y112_C_XOR;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X2Y112_D;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X2Y112_D1;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X2Y112_D2;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X2Y112_D3;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X2Y112_D4;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X2Y112_D5;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X2Y112_D6;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X2Y112_DO5;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X2Y112_DO6;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X2Y112_D_CY;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X2Y112_D_XOR;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X3Y112_A;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X3Y112_A1;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X3Y112_A2;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X3Y112_A3;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X3Y112_A4;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X3Y112_A5;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X3Y112_A6;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X3Y112_AMUX;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X3Y112_AO5;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X3Y112_AO6;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X3Y112_A_CY;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X3Y112_A_XOR;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X3Y112_B;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X3Y112_B1;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X3Y112_B2;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X3Y112_B3;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X3Y112_B4;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X3Y112_B5;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X3Y112_B6;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X3Y112_BO5;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X3Y112_BO6;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X3Y112_B_CY;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X3Y112_B_XOR;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X3Y112_C;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X3Y112_C1;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X3Y112_C2;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X3Y112_C3;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X3Y112_C4;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X3Y112_C5;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X3Y112_C6;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X3Y112_CO5;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X3Y112_CO6;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X3Y112_C_CY;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X3Y112_C_XOR;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X3Y112_D;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X3Y112_D1;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X3Y112_D2;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X3Y112_D3;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X3Y112_D4;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X3Y112_D5;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X3Y112_D6;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X3Y112_DO5;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X3Y112_DO6;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X3Y112_D_CY;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X3Y112_D_XOR;
  wire [0:0] CLBLM_R_X5Y104_SLICE_X6Y104_A;
  wire [0:0] CLBLM_R_X5Y104_SLICE_X6Y104_A1;
  wire [0:0] CLBLM_R_X5Y104_SLICE_X6Y104_A2;
  wire [0:0] CLBLM_R_X5Y104_SLICE_X6Y104_A3;
  wire [0:0] CLBLM_R_X5Y104_SLICE_X6Y104_A4;
  wire [0:0] CLBLM_R_X5Y104_SLICE_X6Y104_A5;
  wire [0:0] CLBLM_R_X5Y104_SLICE_X6Y104_A6;
  wire [0:0] CLBLM_R_X5Y104_SLICE_X6Y104_AMUX;
  wire [0:0] CLBLM_R_X5Y104_SLICE_X6Y104_AO5;
  wire [0:0] CLBLM_R_X5Y104_SLICE_X6Y104_AO6;
  wire [0:0] CLBLM_R_X5Y104_SLICE_X6Y104_A_CY;
  wire [0:0] CLBLM_R_X5Y104_SLICE_X6Y104_A_XOR;
  wire [0:0] CLBLM_R_X5Y104_SLICE_X6Y104_B;
  wire [0:0] CLBLM_R_X5Y104_SLICE_X6Y104_B1;
  wire [0:0] CLBLM_R_X5Y104_SLICE_X6Y104_B2;
  wire [0:0] CLBLM_R_X5Y104_SLICE_X6Y104_B3;
  wire [0:0] CLBLM_R_X5Y104_SLICE_X6Y104_B4;
  wire [0:0] CLBLM_R_X5Y104_SLICE_X6Y104_B5;
  wire [0:0] CLBLM_R_X5Y104_SLICE_X6Y104_B6;
  wire [0:0] CLBLM_R_X5Y104_SLICE_X6Y104_BO5;
  wire [0:0] CLBLM_R_X5Y104_SLICE_X6Y104_BO6;
  wire [0:0] CLBLM_R_X5Y104_SLICE_X6Y104_B_CY;
  wire [0:0] CLBLM_R_X5Y104_SLICE_X6Y104_B_XOR;
  wire [0:0] CLBLM_R_X5Y104_SLICE_X6Y104_C;
  wire [0:0] CLBLM_R_X5Y104_SLICE_X6Y104_C1;
  wire [0:0] CLBLM_R_X5Y104_SLICE_X6Y104_C2;
  wire [0:0] CLBLM_R_X5Y104_SLICE_X6Y104_C3;
  wire [0:0] CLBLM_R_X5Y104_SLICE_X6Y104_C4;
  wire [0:0] CLBLM_R_X5Y104_SLICE_X6Y104_C5;
  wire [0:0] CLBLM_R_X5Y104_SLICE_X6Y104_C6;
  wire [0:0] CLBLM_R_X5Y104_SLICE_X6Y104_CO5;
  wire [0:0] CLBLM_R_X5Y104_SLICE_X6Y104_CO6;
  wire [0:0] CLBLM_R_X5Y104_SLICE_X6Y104_C_CY;
  wire [0:0] CLBLM_R_X5Y104_SLICE_X6Y104_C_XOR;
  wire [0:0] CLBLM_R_X5Y104_SLICE_X6Y104_D;
  wire [0:0] CLBLM_R_X5Y104_SLICE_X6Y104_D1;
  wire [0:0] CLBLM_R_X5Y104_SLICE_X6Y104_D2;
  wire [0:0] CLBLM_R_X5Y104_SLICE_X6Y104_D3;
  wire [0:0] CLBLM_R_X5Y104_SLICE_X6Y104_D4;
  wire [0:0] CLBLM_R_X5Y104_SLICE_X6Y104_D5;
  wire [0:0] CLBLM_R_X5Y104_SLICE_X6Y104_D6;
  wire [0:0] CLBLM_R_X5Y104_SLICE_X6Y104_DO5;
  wire [0:0] CLBLM_R_X5Y104_SLICE_X6Y104_DO6;
  wire [0:0] CLBLM_R_X5Y104_SLICE_X6Y104_D_CY;
  wire [0:0] CLBLM_R_X5Y104_SLICE_X6Y104_D_XOR;
  wire [0:0] CLBLM_R_X5Y104_SLICE_X7Y104_A;
  wire [0:0] CLBLM_R_X5Y104_SLICE_X7Y104_A1;
  wire [0:0] CLBLM_R_X5Y104_SLICE_X7Y104_A2;
  wire [0:0] CLBLM_R_X5Y104_SLICE_X7Y104_A3;
  wire [0:0] CLBLM_R_X5Y104_SLICE_X7Y104_A4;
  wire [0:0] CLBLM_R_X5Y104_SLICE_X7Y104_A5;
  wire [0:0] CLBLM_R_X5Y104_SLICE_X7Y104_A6;
  wire [0:0] CLBLM_R_X5Y104_SLICE_X7Y104_AO5;
  wire [0:0] CLBLM_R_X5Y104_SLICE_X7Y104_AO6;
  wire [0:0] CLBLM_R_X5Y104_SLICE_X7Y104_A_CY;
  wire [0:0] CLBLM_R_X5Y104_SLICE_X7Y104_A_XOR;
  wire [0:0] CLBLM_R_X5Y104_SLICE_X7Y104_B;
  wire [0:0] CLBLM_R_X5Y104_SLICE_X7Y104_B1;
  wire [0:0] CLBLM_R_X5Y104_SLICE_X7Y104_B2;
  wire [0:0] CLBLM_R_X5Y104_SLICE_X7Y104_B3;
  wire [0:0] CLBLM_R_X5Y104_SLICE_X7Y104_B4;
  wire [0:0] CLBLM_R_X5Y104_SLICE_X7Y104_B5;
  wire [0:0] CLBLM_R_X5Y104_SLICE_X7Y104_B6;
  wire [0:0] CLBLM_R_X5Y104_SLICE_X7Y104_BO5;
  wire [0:0] CLBLM_R_X5Y104_SLICE_X7Y104_BO6;
  wire [0:0] CLBLM_R_X5Y104_SLICE_X7Y104_B_CY;
  wire [0:0] CLBLM_R_X5Y104_SLICE_X7Y104_B_XOR;
  wire [0:0] CLBLM_R_X5Y104_SLICE_X7Y104_C;
  wire [0:0] CLBLM_R_X5Y104_SLICE_X7Y104_C1;
  wire [0:0] CLBLM_R_X5Y104_SLICE_X7Y104_C2;
  wire [0:0] CLBLM_R_X5Y104_SLICE_X7Y104_C3;
  wire [0:0] CLBLM_R_X5Y104_SLICE_X7Y104_C4;
  wire [0:0] CLBLM_R_X5Y104_SLICE_X7Y104_C5;
  wire [0:0] CLBLM_R_X5Y104_SLICE_X7Y104_C6;
  wire [0:0] CLBLM_R_X5Y104_SLICE_X7Y104_CO5;
  wire [0:0] CLBLM_R_X5Y104_SLICE_X7Y104_CO6;
  wire [0:0] CLBLM_R_X5Y104_SLICE_X7Y104_C_CY;
  wire [0:0] CLBLM_R_X5Y104_SLICE_X7Y104_C_XOR;
  wire [0:0] CLBLM_R_X5Y104_SLICE_X7Y104_D;
  wire [0:0] CLBLM_R_X5Y104_SLICE_X7Y104_D1;
  wire [0:0] CLBLM_R_X5Y104_SLICE_X7Y104_D2;
  wire [0:0] CLBLM_R_X5Y104_SLICE_X7Y104_D3;
  wire [0:0] CLBLM_R_X5Y104_SLICE_X7Y104_D4;
  wire [0:0] CLBLM_R_X5Y104_SLICE_X7Y104_D5;
  wire [0:0] CLBLM_R_X5Y104_SLICE_X7Y104_D6;
  wire [0:0] CLBLM_R_X5Y104_SLICE_X7Y104_DO5;
  wire [0:0] CLBLM_R_X5Y104_SLICE_X7Y104_DO6;
  wire [0:0] CLBLM_R_X5Y104_SLICE_X7Y104_D_CY;
  wire [0:0] CLBLM_R_X5Y104_SLICE_X7Y104_D_XOR;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X6Y105_A;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X6Y105_A1;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X6Y105_A2;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X6Y105_A3;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X6Y105_A4;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X6Y105_A5;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X6Y105_A6;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X6Y105_AO5;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X6Y105_AO6;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X6Y105_A_CY;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X6Y105_A_XOR;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X6Y105_B;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X6Y105_B1;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X6Y105_B2;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X6Y105_B3;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X6Y105_B4;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X6Y105_B5;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X6Y105_B6;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X6Y105_BO5;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X6Y105_BO6;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X6Y105_B_CY;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X6Y105_B_XOR;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X6Y105_C;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X6Y105_C1;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X6Y105_C2;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X6Y105_C3;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X6Y105_C4;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X6Y105_C5;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X6Y105_C6;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X6Y105_CO5;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X6Y105_CO6;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X6Y105_C_CY;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X6Y105_C_XOR;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X6Y105_D;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X6Y105_D1;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X6Y105_D2;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X6Y105_D3;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X6Y105_D4;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X6Y105_D5;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X6Y105_D6;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X6Y105_DO5;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X6Y105_DO6;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X6Y105_D_CY;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X6Y105_D_XOR;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X7Y105_A;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X7Y105_A1;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X7Y105_A2;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X7Y105_A3;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X7Y105_A4;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X7Y105_A5;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X7Y105_A6;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X7Y105_AMUX;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X7Y105_AO5;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X7Y105_AO6;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X7Y105_A_CY;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X7Y105_A_XOR;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X7Y105_B;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X7Y105_B1;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X7Y105_B2;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X7Y105_B3;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X7Y105_B4;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X7Y105_B5;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X7Y105_B6;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X7Y105_BO5;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X7Y105_BO6;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X7Y105_B_CY;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X7Y105_B_XOR;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X7Y105_C;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X7Y105_C1;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X7Y105_C2;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X7Y105_C3;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X7Y105_C4;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X7Y105_C5;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X7Y105_C6;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X7Y105_CO5;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X7Y105_CO6;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X7Y105_C_CY;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X7Y105_C_XOR;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X7Y105_D;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X7Y105_D1;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X7Y105_D2;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X7Y105_D3;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X7Y105_D4;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X7Y105_D5;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X7Y105_D6;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X7Y105_DO5;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X7Y105_DO6;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X7Y105_D_CY;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X7Y105_D_XOR;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X6Y106_A;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X6Y106_A1;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X6Y106_A2;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X6Y106_A3;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X6Y106_A4;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X6Y106_A5;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X6Y106_A6;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X6Y106_AMUX;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X6Y106_AO5;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X6Y106_AO6;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X6Y106_A_CY;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X6Y106_A_XOR;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X6Y106_B;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X6Y106_B1;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X6Y106_B2;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X6Y106_B3;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X6Y106_B4;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X6Y106_B5;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X6Y106_B6;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X6Y106_BO5;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X6Y106_BO6;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X6Y106_B_CY;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X6Y106_B_XOR;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X6Y106_C;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X6Y106_C1;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X6Y106_C2;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X6Y106_C3;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X6Y106_C4;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X6Y106_C5;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X6Y106_C6;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X6Y106_CO5;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X6Y106_CO6;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X6Y106_C_CY;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X6Y106_C_XOR;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X6Y106_D;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X6Y106_D1;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X6Y106_D2;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X6Y106_D3;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X6Y106_D4;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X6Y106_D5;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X6Y106_D6;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X6Y106_DO5;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X6Y106_DO6;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X6Y106_D_CY;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X6Y106_D_XOR;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X7Y106_A;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X7Y106_A1;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X7Y106_A2;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X7Y106_A3;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X7Y106_A4;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X7Y106_A5;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X7Y106_A6;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X7Y106_AMUX;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X7Y106_AO5;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X7Y106_AO6;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X7Y106_A_CY;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X7Y106_A_XOR;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X7Y106_B;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X7Y106_B1;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X7Y106_B2;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X7Y106_B3;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X7Y106_B4;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X7Y106_B5;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X7Y106_B6;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X7Y106_BMUX;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X7Y106_BO5;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X7Y106_BO6;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X7Y106_B_CY;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X7Y106_B_XOR;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X7Y106_C;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X7Y106_C1;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X7Y106_C2;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X7Y106_C3;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X7Y106_C4;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X7Y106_C5;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X7Y106_C6;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X7Y106_CO5;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X7Y106_CO6;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X7Y106_C_CY;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X7Y106_C_XOR;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X7Y106_D;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X7Y106_D1;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X7Y106_D2;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X7Y106_D3;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X7Y106_D4;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X7Y106_D5;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X7Y106_D6;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X7Y106_DO5;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X7Y106_DO6;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X7Y106_D_CY;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X7Y106_D_XOR;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X6Y107_A;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X6Y107_A1;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X6Y107_A2;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X6Y107_A3;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X6Y107_A4;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X6Y107_A5;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X6Y107_A6;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X6Y107_AO5;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X6Y107_AO6;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X6Y107_A_CY;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X6Y107_A_XOR;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X6Y107_B;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X6Y107_B1;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X6Y107_B2;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X6Y107_B3;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X6Y107_B4;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X6Y107_B5;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X6Y107_B6;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X6Y107_BO5;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X6Y107_BO6;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X6Y107_B_CY;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X6Y107_B_XOR;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X6Y107_C;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X6Y107_C1;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X6Y107_C2;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X6Y107_C3;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X6Y107_C4;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X6Y107_C5;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X6Y107_C6;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X6Y107_CO5;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X6Y107_CO6;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X6Y107_C_CY;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X6Y107_C_XOR;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X6Y107_D;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X6Y107_D1;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X6Y107_D2;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X6Y107_D3;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X6Y107_D4;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X6Y107_D5;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X6Y107_D6;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X6Y107_DO5;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X6Y107_DO6;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X6Y107_D_CY;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X6Y107_D_XOR;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X7Y107_A;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X7Y107_A1;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X7Y107_A2;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X7Y107_A3;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X7Y107_A4;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X7Y107_A5;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X7Y107_A6;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X7Y107_AMUX;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X7Y107_AO5;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X7Y107_AO6;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X7Y107_A_CY;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X7Y107_A_XOR;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X7Y107_B;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X7Y107_B1;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X7Y107_B2;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X7Y107_B3;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X7Y107_B4;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X7Y107_B5;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X7Y107_B6;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X7Y107_BO5;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X7Y107_BO6;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X7Y107_B_CY;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X7Y107_B_XOR;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X7Y107_C;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X7Y107_C1;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X7Y107_C2;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X7Y107_C3;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X7Y107_C4;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X7Y107_C5;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X7Y107_C6;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X7Y107_CO5;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X7Y107_CO6;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X7Y107_C_CY;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X7Y107_C_XOR;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X7Y107_D;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X7Y107_D1;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X7Y107_D2;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X7Y107_D3;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X7Y107_D4;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X7Y107_D5;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X7Y107_D6;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X7Y107_DO5;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X7Y107_DO6;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X7Y107_D_CY;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X7Y107_D_XOR;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X6Y108_A;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X6Y108_A1;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X6Y108_A2;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X6Y108_A3;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X6Y108_A4;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X6Y108_A5;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X6Y108_A6;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X6Y108_AO5;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X6Y108_AO6;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X6Y108_A_CY;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X6Y108_A_XOR;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X6Y108_B;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X6Y108_B1;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X6Y108_B2;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X6Y108_B3;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X6Y108_B4;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X6Y108_B5;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X6Y108_B6;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X6Y108_BMUX;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X6Y108_BO5;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X6Y108_BO6;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X6Y108_B_CY;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X6Y108_B_XOR;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X6Y108_C;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X6Y108_C1;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X6Y108_C2;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X6Y108_C3;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X6Y108_C4;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X6Y108_C5;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X6Y108_C6;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X6Y108_CO5;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X6Y108_CO6;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X6Y108_C_CY;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X6Y108_C_XOR;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X6Y108_D;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X6Y108_D1;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X6Y108_D2;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X6Y108_D3;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X6Y108_D4;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X6Y108_D5;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X6Y108_D6;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X6Y108_DO5;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X6Y108_DO6;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X6Y108_D_CY;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X6Y108_D_XOR;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X7Y108_A;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X7Y108_A1;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X7Y108_A2;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X7Y108_A3;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X7Y108_A4;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X7Y108_A5;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X7Y108_A6;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X7Y108_AMUX;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X7Y108_AO5;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X7Y108_AO6;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X7Y108_A_CY;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X7Y108_A_XOR;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X7Y108_B;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X7Y108_B1;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X7Y108_B2;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X7Y108_B3;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X7Y108_B4;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X7Y108_B5;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X7Y108_B6;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X7Y108_BO5;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X7Y108_BO6;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X7Y108_B_CY;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X7Y108_B_XOR;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X7Y108_C;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X7Y108_C1;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X7Y108_C2;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X7Y108_C3;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X7Y108_C4;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X7Y108_C5;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X7Y108_C6;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X7Y108_CO5;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X7Y108_CO6;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X7Y108_C_CY;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X7Y108_C_XOR;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X7Y108_D;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X7Y108_D1;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X7Y108_D2;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X7Y108_D3;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X7Y108_D4;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X7Y108_D5;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X7Y108_D6;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X7Y108_DO5;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X7Y108_DO6;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X7Y108_D_CY;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X7Y108_D_XOR;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X6Y109_A;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X6Y109_A1;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X6Y109_A2;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X6Y109_A3;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X6Y109_A4;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X6Y109_A5;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X6Y109_A6;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X6Y109_AO5;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X6Y109_AO6;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X6Y109_A_CY;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X6Y109_A_XOR;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X6Y109_B;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X6Y109_B1;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X6Y109_B2;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X6Y109_B3;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X6Y109_B4;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X6Y109_B5;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X6Y109_B6;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X6Y109_BO5;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X6Y109_BO6;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X6Y109_B_CY;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X6Y109_B_XOR;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X6Y109_C;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X6Y109_C1;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X6Y109_C2;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X6Y109_C3;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X6Y109_C4;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X6Y109_C5;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X6Y109_C6;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X6Y109_CO5;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X6Y109_CO6;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X6Y109_C_CY;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X6Y109_C_XOR;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X6Y109_D;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X6Y109_D1;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X6Y109_D2;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X6Y109_D3;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X6Y109_D4;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X6Y109_D5;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X6Y109_D6;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X6Y109_DO5;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X6Y109_DO6;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X6Y109_D_CY;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X6Y109_D_XOR;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X7Y109_A;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X7Y109_A1;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X7Y109_A2;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X7Y109_A3;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X7Y109_A4;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X7Y109_A5;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X7Y109_A6;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X7Y109_AO5;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X7Y109_AO6;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X7Y109_A_CY;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X7Y109_A_XOR;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X7Y109_B;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X7Y109_B1;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X7Y109_B2;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X7Y109_B3;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X7Y109_B4;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X7Y109_B5;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X7Y109_B6;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X7Y109_BO5;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X7Y109_BO6;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X7Y109_B_CY;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X7Y109_B_XOR;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X7Y109_C;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X7Y109_C1;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X7Y109_C2;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X7Y109_C3;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X7Y109_C4;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X7Y109_C5;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X7Y109_C6;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X7Y109_CO5;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X7Y109_CO6;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X7Y109_C_CY;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X7Y109_C_XOR;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X7Y109_D;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X7Y109_D1;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X7Y109_D2;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X7Y109_D3;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X7Y109_D4;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X7Y109_D5;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X7Y109_D6;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X7Y109_DO5;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X7Y109_DO6;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X7Y109_D_CY;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X7Y109_D_XOR;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X6Y110_A;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X6Y110_A1;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X6Y110_A2;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X6Y110_A3;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X6Y110_A4;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X6Y110_A5;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X6Y110_A6;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X6Y110_AMUX;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X6Y110_AO5;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X6Y110_AO6;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X6Y110_A_CY;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X6Y110_A_XOR;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X6Y110_B;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X6Y110_B1;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X6Y110_B2;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X6Y110_B3;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X6Y110_B4;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X6Y110_B5;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X6Y110_B6;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X6Y110_BMUX;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X6Y110_BO5;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X6Y110_BO6;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X6Y110_B_CY;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X6Y110_B_XOR;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X6Y110_C;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X6Y110_C1;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X6Y110_C2;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X6Y110_C3;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X6Y110_C4;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X6Y110_C5;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X6Y110_C6;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X6Y110_CO5;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X6Y110_CO6;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X6Y110_C_CY;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X6Y110_C_XOR;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X6Y110_D;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X6Y110_D1;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X6Y110_D2;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X6Y110_D3;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X6Y110_D4;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X6Y110_D5;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X6Y110_D6;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X6Y110_DO5;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X6Y110_DO6;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X6Y110_D_CY;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X6Y110_D_XOR;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X7Y110_A;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X7Y110_A1;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X7Y110_A2;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X7Y110_A3;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X7Y110_A4;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X7Y110_A5;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X7Y110_A6;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X7Y110_AMUX;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X7Y110_AO5;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X7Y110_AO6;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X7Y110_A_CY;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X7Y110_A_XOR;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X7Y110_B;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X7Y110_B1;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X7Y110_B2;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X7Y110_B3;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X7Y110_B4;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X7Y110_B5;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X7Y110_B6;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X7Y110_BMUX;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X7Y110_BO5;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X7Y110_BO6;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X7Y110_B_CY;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X7Y110_B_XOR;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X7Y110_C;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X7Y110_C1;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X7Y110_C2;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X7Y110_C3;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X7Y110_C4;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X7Y110_C5;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X7Y110_C6;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X7Y110_CMUX;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X7Y110_CO5;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X7Y110_CO6;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X7Y110_C_CY;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X7Y110_C_XOR;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X7Y110_D;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X7Y110_D1;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X7Y110_D2;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X7Y110_D3;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X7Y110_D4;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X7Y110_D5;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X7Y110_D6;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X7Y110_DO5;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X7Y110_DO6;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X7Y110_D_CY;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X7Y110_D_XOR;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X6Y111_A;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X6Y111_A1;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X6Y111_A2;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X6Y111_A3;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X6Y111_A4;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X6Y111_A5;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X6Y111_A6;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X6Y111_AO5;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X6Y111_AO6;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X6Y111_A_CY;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X6Y111_A_XOR;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X6Y111_B;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X6Y111_B1;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X6Y111_B2;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X6Y111_B3;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X6Y111_B4;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X6Y111_B5;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X6Y111_B6;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X6Y111_BO5;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X6Y111_BO6;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X6Y111_B_CY;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X6Y111_B_XOR;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X6Y111_C;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X6Y111_C1;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X6Y111_C2;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X6Y111_C3;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X6Y111_C4;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X6Y111_C5;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X6Y111_C6;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X6Y111_CO5;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X6Y111_CO6;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X6Y111_C_CY;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X6Y111_C_XOR;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X6Y111_D;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X6Y111_D1;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X6Y111_D2;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X6Y111_D3;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X6Y111_D4;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X6Y111_D5;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X6Y111_D6;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X6Y111_DO5;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X6Y111_DO6;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X6Y111_D_CY;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X6Y111_D_XOR;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X7Y111_A;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X7Y111_A1;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X7Y111_A2;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X7Y111_A3;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X7Y111_A4;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X7Y111_A5;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X7Y111_A6;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X7Y111_AO5;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X7Y111_AO6;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X7Y111_A_CY;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X7Y111_A_XOR;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X7Y111_B;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X7Y111_B1;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X7Y111_B2;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X7Y111_B3;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X7Y111_B4;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X7Y111_B5;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X7Y111_B6;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X7Y111_BO5;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X7Y111_BO6;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X7Y111_B_CY;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X7Y111_B_XOR;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X7Y111_C;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X7Y111_C1;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X7Y111_C2;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X7Y111_C3;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X7Y111_C4;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X7Y111_C5;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X7Y111_C6;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X7Y111_CO5;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X7Y111_CO6;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X7Y111_C_CY;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X7Y111_C_XOR;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X7Y111_D;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X7Y111_D1;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X7Y111_D2;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X7Y111_D3;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X7Y111_D4;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X7Y111_D5;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X7Y111_D6;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X7Y111_DO5;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X7Y111_DO6;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X7Y111_D_CY;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X7Y111_D_XOR;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X6Y112_A;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X6Y112_A1;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X6Y112_A2;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X6Y112_A3;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X6Y112_A4;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X6Y112_A5;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X6Y112_A6;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X6Y112_AMUX;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X6Y112_AO5;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X6Y112_AO6;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X6Y112_A_CY;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X6Y112_A_XOR;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X6Y112_B;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X6Y112_B1;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X6Y112_B2;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X6Y112_B3;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X6Y112_B4;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X6Y112_B5;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X6Y112_B6;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X6Y112_BO5;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X6Y112_BO6;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X6Y112_B_CY;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X6Y112_B_XOR;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X6Y112_C;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X6Y112_C1;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X6Y112_C2;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X6Y112_C3;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X6Y112_C4;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X6Y112_C5;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X6Y112_C6;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X6Y112_CMUX;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X6Y112_CO5;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X6Y112_CO6;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X6Y112_C_CY;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X6Y112_C_XOR;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X6Y112_D;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X6Y112_D1;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X6Y112_D2;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X6Y112_D3;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X6Y112_D4;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X6Y112_D5;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X6Y112_D6;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X6Y112_DO5;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X6Y112_DO6;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X6Y112_D_CY;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X6Y112_D_XOR;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X7Y112_A;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X7Y112_A1;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X7Y112_A2;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X7Y112_A3;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X7Y112_A4;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X7Y112_A5;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X7Y112_A6;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X7Y112_AMUX;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X7Y112_AO5;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X7Y112_AO6;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X7Y112_A_CY;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X7Y112_A_XOR;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X7Y112_B;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X7Y112_B1;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X7Y112_B2;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X7Y112_B3;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X7Y112_B4;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X7Y112_B5;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X7Y112_B6;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X7Y112_BO5;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X7Y112_BO6;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X7Y112_B_CY;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X7Y112_B_XOR;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X7Y112_C;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X7Y112_C1;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X7Y112_C2;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X7Y112_C3;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X7Y112_C4;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X7Y112_C5;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X7Y112_C6;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X7Y112_CO5;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X7Y112_CO6;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X7Y112_C_CY;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X7Y112_C_XOR;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X7Y112_D;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X7Y112_D1;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X7Y112_D2;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X7Y112_D3;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X7Y112_D4;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X7Y112_D5;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X7Y112_D6;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X7Y112_DO5;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X7Y112_DO6;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X7Y112_D_CY;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X7Y112_D_XOR;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X6Y113_A;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X6Y113_A1;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X6Y113_A2;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X6Y113_A3;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X6Y113_A4;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X6Y113_A5;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X6Y113_A6;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X6Y113_AO5;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X6Y113_AO6;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X6Y113_A_CY;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X6Y113_A_XOR;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X6Y113_B;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X6Y113_B1;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X6Y113_B2;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X6Y113_B3;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X6Y113_B4;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X6Y113_B5;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X6Y113_B6;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X6Y113_BO5;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X6Y113_BO6;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X6Y113_B_CY;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X6Y113_B_XOR;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X6Y113_C;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X6Y113_C1;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X6Y113_C2;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X6Y113_C3;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X6Y113_C4;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X6Y113_C5;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X6Y113_C6;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X6Y113_CO5;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X6Y113_CO6;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X6Y113_C_CY;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X6Y113_C_XOR;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X6Y113_D;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X6Y113_D1;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X6Y113_D2;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X6Y113_D3;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X6Y113_D4;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X6Y113_D5;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X6Y113_D6;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X6Y113_DO5;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X6Y113_DO6;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X6Y113_D_CY;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X6Y113_D_XOR;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X7Y113_A;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X7Y113_A1;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X7Y113_A2;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X7Y113_A3;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X7Y113_A4;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X7Y113_A5;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X7Y113_A6;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X7Y113_AMUX;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X7Y113_AO5;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X7Y113_AO6;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X7Y113_A_CY;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X7Y113_A_XOR;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X7Y113_B;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X7Y113_B1;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X7Y113_B2;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X7Y113_B3;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X7Y113_B4;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X7Y113_B5;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X7Y113_B6;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X7Y113_BO5;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X7Y113_BO6;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X7Y113_B_CY;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X7Y113_B_XOR;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X7Y113_C;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X7Y113_C1;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X7Y113_C2;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X7Y113_C3;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X7Y113_C4;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X7Y113_C5;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X7Y113_C6;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X7Y113_CO5;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X7Y113_CO6;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X7Y113_C_CY;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X7Y113_C_XOR;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X7Y113_D;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X7Y113_D1;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X7Y113_D2;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X7Y113_D3;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X7Y113_D4;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X7Y113_D5;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X7Y113_D6;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X7Y113_DO5;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X7Y113_DO6;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X7Y113_D_CY;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X7Y113_D_XOR;
  wire [0:0] CLBLM_R_X7Y103_SLICE_X8Y103_A;
  wire [0:0] CLBLM_R_X7Y103_SLICE_X8Y103_A1;
  wire [0:0] CLBLM_R_X7Y103_SLICE_X8Y103_A2;
  wire [0:0] CLBLM_R_X7Y103_SLICE_X8Y103_A3;
  wire [0:0] CLBLM_R_X7Y103_SLICE_X8Y103_A4;
  wire [0:0] CLBLM_R_X7Y103_SLICE_X8Y103_A5;
  wire [0:0] CLBLM_R_X7Y103_SLICE_X8Y103_A6;
  wire [0:0] CLBLM_R_X7Y103_SLICE_X8Y103_AO5;
  wire [0:0] CLBLM_R_X7Y103_SLICE_X8Y103_AO6;
  wire [0:0] CLBLM_R_X7Y103_SLICE_X8Y103_A_CY;
  wire [0:0] CLBLM_R_X7Y103_SLICE_X8Y103_A_XOR;
  wire [0:0] CLBLM_R_X7Y103_SLICE_X8Y103_B;
  wire [0:0] CLBLM_R_X7Y103_SLICE_X8Y103_B1;
  wire [0:0] CLBLM_R_X7Y103_SLICE_X8Y103_B2;
  wire [0:0] CLBLM_R_X7Y103_SLICE_X8Y103_B3;
  wire [0:0] CLBLM_R_X7Y103_SLICE_X8Y103_B4;
  wire [0:0] CLBLM_R_X7Y103_SLICE_X8Y103_B5;
  wire [0:0] CLBLM_R_X7Y103_SLICE_X8Y103_B6;
  wire [0:0] CLBLM_R_X7Y103_SLICE_X8Y103_BO5;
  wire [0:0] CLBLM_R_X7Y103_SLICE_X8Y103_BO6;
  wire [0:0] CLBLM_R_X7Y103_SLICE_X8Y103_B_CY;
  wire [0:0] CLBLM_R_X7Y103_SLICE_X8Y103_B_XOR;
  wire [0:0] CLBLM_R_X7Y103_SLICE_X8Y103_C;
  wire [0:0] CLBLM_R_X7Y103_SLICE_X8Y103_C1;
  wire [0:0] CLBLM_R_X7Y103_SLICE_X8Y103_C2;
  wire [0:0] CLBLM_R_X7Y103_SLICE_X8Y103_C3;
  wire [0:0] CLBLM_R_X7Y103_SLICE_X8Y103_C4;
  wire [0:0] CLBLM_R_X7Y103_SLICE_X8Y103_C5;
  wire [0:0] CLBLM_R_X7Y103_SLICE_X8Y103_C6;
  wire [0:0] CLBLM_R_X7Y103_SLICE_X8Y103_CO5;
  wire [0:0] CLBLM_R_X7Y103_SLICE_X8Y103_CO6;
  wire [0:0] CLBLM_R_X7Y103_SLICE_X8Y103_C_CY;
  wire [0:0] CLBLM_R_X7Y103_SLICE_X8Y103_C_XOR;
  wire [0:0] CLBLM_R_X7Y103_SLICE_X8Y103_D;
  wire [0:0] CLBLM_R_X7Y103_SLICE_X8Y103_D1;
  wire [0:0] CLBLM_R_X7Y103_SLICE_X8Y103_D2;
  wire [0:0] CLBLM_R_X7Y103_SLICE_X8Y103_D3;
  wire [0:0] CLBLM_R_X7Y103_SLICE_X8Y103_D4;
  wire [0:0] CLBLM_R_X7Y103_SLICE_X8Y103_D5;
  wire [0:0] CLBLM_R_X7Y103_SLICE_X8Y103_D6;
  wire [0:0] CLBLM_R_X7Y103_SLICE_X8Y103_DO5;
  wire [0:0] CLBLM_R_X7Y103_SLICE_X8Y103_DO6;
  wire [0:0] CLBLM_R_X7Y103_SLICE_X8Y103_D_CY;
  wire [0:0] CLBLM_R_X7Y103_SLICE_X8Y103_D_XOR;
  wire [0:0] CLBLM_R_X7Y103_SLICE_X9Y103_A;
  wire [0:0] CLBLM_R_X7Y103_SLICE_X9Y103_A1;
  wire [0:0] CLBLM_R_X7Y103_SLICE_X9Y103_A2;
  wire [0:0] CLBLM_R_X7Y103_SLICE_X9Y103_A3;
  wire [0:0] CLBLM_R_X7Y103_SLICE_X9Y103_A4;
  wire [0:0] CLBLM_R_X7Y103_SLICE_X9Y103_A5;
  wire [0:0] CLBLM_R_X7Y103_SLICE_X9Y103_A6;
  wire [0:0] CLBLM_R_X7Y103_SLICE_X9Y103_AO5;
  wire [0:0] CLBLM_R_X7Y103_SLICE_X9Y103_AO6;
  wire [0:0] CLBLM_R_X7Y103_SLICE_X9Y103_A_CY;
  wire [0:0] CLBLM_R_X7Y103_SLICE_X9Y103_A_XOR;
  wire [0:0] CLBLM_R_X7Y103_SLICE_X9Y103_B;
  wire [0:0] CLBLM_R_X7Y103_SLICE_X9Y103_B1;
  wire [0:0] CLBLM_R_X7Y103_SLICE_X9Y103_B2;
  wire [0:0] CLBLM_R_X7Y103_SLICE_X9Y103_B3;
  wire [0:0] CLBLM_R_X7Y103_SLICE_X9Y103_B4;
  wire [0:0] CLBLM_R_X7Y103_SLICE_X9Y103_B5;
  wire [0:0] CLBLM_R_X7Y103_SLICE_X9Y103_B6;
  wire [0:0] CLBLM_R_X7Y103_SLICE_X9Y103_BO5;
  wire [0:0] CLBLM_R_X7Y103_SLICE_X9Y103_BO6;
  wire [0:0] CLBLM_R_X7Y103_SLICE_X9Y103_B_CY;
  wire [0:0] CLBLM_R_X7Y103_SLICE_X9Y103_B_XOR;
  wire [0:0] CLBLM_R_X7Y103_SLICE_X9Y103_C;
  wire [0:0] CLBLM_R_X7Y103_SLICE_X9Y103_C1;
  wire [0:0] CLBLM_R_X7Y103_SLICE_X9Y103_C2;
  wire [0:0] CLBLM_R_X7Y103_SLICE_X9Y103_C3;
  wire [0:0] CLBLM_R_X7Y103_SLICE_X9Y103_C4;
  wire [0:0] CLBLM_R_X7Y103_SLICE_X9Y103_C5;
  wire [0:0] CLBLM_R_X7Y103_SLICE_X9Y103_C6;
  wire [0:0] CLBLM_R_X7Y103_SLICE_X9Y103_CO5;
  wire [0:0] CLBLM_R_X7Y103_SLICE_X9Y103_CO6;
  wire [0:0] CLBLM_R_X7Y103_SLICE_X9Y103_C_CY;
  wire [0:0] CLBLM_R_X7Y103_SLICE_X9Y103_C_XOR;
  wire [0:0] CLBLM_R_X7Y103_SLICE_X9Y103_D;
  wire [0:0] CLBLM_R_X7Y103_SLICE_X9Y103_D1;
  wire [0:0] CLBLM_R_X7Y103_SLICE_X9Y103_D2;
  wire [0:0] CLBLM_R_X7Y103_SLICE_X9Y103_D3;
  wire [0:0] CLBLM_R_X7Y103_SLICE_X9Y103_D4;
  wire [0:0] CLBLM_R_X7Y103_SLICE_X9Y103_D5;
  wire [0:0] CLBLM_R_X7Y103_SLICE_X9Y103_D6;
  wire [0:0] CLBLM_R_X7Y103_SLICE_X9Y103_DO5;
  wire [0:0] CLBLM_R_X7Y103_SLICE_X9Y103_DO6;
  wire [0:0] CLBLM_R_X7Y103_SLICE_X9Y103_D_CY;
  wire [0:0] CLBLM_R_X7Y103_SLICE_X9Y103_D_XOR;
  wire [0:0] CLBLM_R_X7Y104_SLICE_X8Y104_A;
  wire [0:0] CLBLM_R_X7Y104_SLICE_X8Y104_A1;
  wire [0:0] CLBLM_R_X7Y104_SLICE_X8Y104_A2;
  wire [0:0] CLBLM_R_X7Y104_SLICE_X8Y104_A3;
  wire [0:0] CLBLM_R_X7Y104_SLICE_X8Y104_A4;
  wire [0:0] CLBLM_R_X7Y104_SLICE_X8Y104_A5;
  wire [0:0] CLBLM_R_X7Y104_SLICE_X8Y104_A6;
  wire [0:0] CLBLM_R_X7Y104_SLICE_X8Y104_AMUX;
  wire [0:0] CLBLM_R_X7Y104_SLICE_X8Y104_AO5;
  wire [0:0] CLBLM_R_X7Y104_SLICE_X8Y104_AO6;
  wire [0:0] CLBLM_R_X7Y104_SLICE_X8Y104_A_CY;
  wire [0:0] CLBLM_R_X7Y104_SLICE_X8Y104_A_XOR;
  wire [0:0] CLBLM_R_X7Y104_SLICE_X8Y104_B;
  wire [0:0] CLBLM_R_X7Y104_SLICE_X8Y104_B1;
  wire [0:0] CLBLM_R_X7Y104_SLICE_X8Y104_B2;
  wire [0:0] CLBLM_R_X7Y104_SLICE_X8Y104_B3;
  wire [0:0] CLBLM_R_X7Y104_SLICE_X8Y104_B4;
  wire [0:0] CLBLM_R_X7Y104_SLICE_X8Y104_B5;
  wire [0:0] CLBLM_R_X7Y104_SLICE_X8Y104_B6;
  wire [0:0] CLBLM_R_X7Y104_SLICE_X8Y104_BMUX;
  wire [0:0] CLBLM_R_X7Y104_SLICE_X8Y104_BO5;
  wire [0:0] CLBLM_R_X7Y104_SLICE_X8Y104_BO6;
  wire [0:0] CLBLM_R_X7Y104_SLICE_X8Y104_B_CY;
  wire [0:0] CLBLM_R_X7Y104_SLICE_X8Y104_B_XOR;
  wire [0:0] CLBLM_R_X7Y104_SLICE_X8Y104_C;
  wire [0:0] CLBLM_R_X7Y104_SLICE_X8Y104_C1;
  wire [0:0] CLBLM_R_X7Y104_SLICE_X8Y104_C2;
  wire [0:0] CLBLM_R_X7Y104_SLICE_X8Y104_C3;
  wire [0:0] CLBLM_R_X7Y104_SLICE_X8Y104_C4;
  wire [0:0] CLBLM_R_X7Y104_SLICE_X8Y104_C5;
  wire [0:0] CLBLM_R_X7Y104_SLICE_X8Y104_C6;
  wire [0:0] CLBLM_R_X7Y104_SLICE_X8Y104_CO5;
  wire [0:0] CLBLM_R_X7Y104_SLICE_X8Y104_CO6;
  wire [0:0] CLBLM_R_X7Y104_SLICE_X8Y104_C_CY;
  wire [0:0] CLBLM_R_X7Y104_SLICE_X8Y104_C_XOR;
  wire [0:0] CLBLM_R_X7Y104_SLICE_X8Y104_D;
  wire [0:0] CLBLM_R_X7Y104_SLICE_X8Y104_D1;
  wire [0:0] CLBLM_R_X7Y104_SLICE_X8Y104_D2;
  wire [0:0] CLBLM_R_X7Y104_SLICE_X8Y104_D3;
  wire [0:0] CLBLM_R_X7Y104_SLICE_X8Y104_D4;
  wire [0:0] CLBLM_R_X7Y104_SLICE_X8Y104_D5;
  wire [0:0] CLBLM_R_X7Y104_SLICE_X8Y104_D6;
  wire [0:0] CLBLM_R_X7Y104_SLICE_X8Y104_DO5;
  wire [0:0] CLBLM_R_X7Y104_SLICE_X8Y104_DO6;
  wire [0:0] CLBLM_R_X7Y104_SLICE_X8Y104_D_CY;
  wire [0:0] CLBLM_R_X7Y104_SLICE_X8Y104_D_XOR;
  wire [0:0] CLBLM_R_X7Y104_SLICE_X9Y104_A;
  wire [0:0] CLBLM_R_X7Y104_SLICE_X9Y104_A1;
  wire [0:0] CLBLM_R_X7Y104_SLICE_X9Y104_A2;
  wire [0:0] CLBLM_R_X7Y104_SLICE_X9Y104_A3;
  wire [0:0] CLBLM_R_X7Y104_SLICE_X9Y104_A4;
  wire [0:0] CLBLM_R_X7Y104_SLICE_X9Y104_A5;
  wire [0:0] CLBLM_R_X7Y104_SLICE_X9Y104_A6;
  wire [0:0] CLBLM_R_X7Y104_SLICE_X9Y104_AMUX;
  wire [0:0] CLBLM_R_X7Y104_SLICE_X9Y104_AO5;
  wire [0:0] CLBLM_R_X7Y104_SLICE_X9Y104_AO6;
  wire [0:0] CLBLM_R_X7Y104_SLICE_X9Y104_A_CY;
  wire [0:0] CLBLM_R_X7Y104_SLICE_X9Y104_A_XOR;
  wire [0:0] CLBLM_R_X7Y104_SLICE_X9Y104_B;
  wire [0:0] CLBLM_R_X7Y104_SLICE_X9Y104_B1;
  wire [0:0] CLBLM_R_X7Y104_SLICE_X9Y104_B2;
  wire [0:0] CLBLM_R_X7Y104_SLICE_X9Y104_B3;
  wire [0:0] CLBLM_R_X7Y104_SLICE_X9Y104_B4;
  wire [0:0] CLBLM_R_X7Y104_SLICE_X9Y104_B5;
  wire [0:0] CLBLM_R_X7Y104_SLICE_X9Y104_B6;
  wire [0:0] CLBLM_R_X7Y104_SLICE_X9Y104_BO5;
  wire [0:0] CLBLM_R_X7Y104_SLICE_X9Y104_BO6;
  wire [0:0] CLBLM_R_X7Y104_SLICE_X9Y104_B_CY;
  wire [0:0] CLBLM_R_X7Y104_SLICE_X9Y104_B_XOR;
  wire [0:0] CLBLM_R_X7Y104_SLICE_X9Y104_C;
  wire [0:0] CLBLM_R_X7Y104_SLICE_X9Y104_C1;
  wire [0:0] CLBLM_R_X7Y104_SLICE_X9Y104_C2;
  wire [0:0] CLBLM_R_X7Y104_SLICE_X9Y104_C3;
  wire [0:0] CLBLM_R_X7Y104_SLICE_X9Y104_C4;
  wire [0:0] CLBLM_R_X7Y104_SLICE_X9Y104_C5;
  wire [0:0] CLBLM_R_X7Y104_SLICE_X9Y104_C6;
  wire [0:0] CLBLM_R_X7Y104_SLICE_X9Y104_CO5;
  wire [0:0] CLBLM_R_X7Y104_SLICE_X9Y104_CO6;
  wire [0:0] CLBLM_R_X7Y104_SLICE_X9Y104_C_CY;
  wire [0:0] CLBLM_R_X7Y104_SLICE_X9Y104_C_XOR;
  wire [0:0] CLBLM_R_X7Y104_SLICE_X9Y104_D;
  wire [0:0] CLBLM_R_X7Y104_SLICE_X9Y104_D1;
  wire [0:0] CLBLM_R_X7Y104_SLICE_X9Y104_D2;
  wire [0:0] CLBLM_R_X7Y104_SLICE_X9Y104_D3;
  wire [0:0] CLBLM_R_X7Y104_SLICE_X9Y104_D4;
  wire [0:0] CLBLM_R_X7Y104_SLICE_X9Y104_D5;
  wire [0:0] CLBLM_R_X7Y104_SLICE_X9Y104_D6;
  wire [0:0] CLBLM_R_X7Y104_SLICE_X9Y104_DO5;
  wire [0:0] CLBLM_R_X7Y104_SLICE_X9Y104_DO6;
  wire [0:0] CLBLM_R_X7Y104_SLICE_X9Y104_D_CY;
  wire [0:0] CLBLM_R_X7Y104_SLICE_X9Y104_D_XOR;
  wire [0:0] CLBLM_R_X7Y105_SLICE_X8Y105_A;
  wire [0:0] CLBLM_R_X7Y105_SLICE_X8Y105_A1;
  wire [0:0] CLBLM_R_X7Y105_SLICE_X8Y105_A2;
  wire [0:0] CLBLM_R_X7Y105_SLICE_X8Y105_A3;
  wire [0:0] CLBLM_R_X7Y105_SLICE_X8Y105_A4;
  wire [0:0] CLBLM_R_X7Y105_SLICE_X8Y105_A5;
  wire [0:0] CLBLM_R_X7Y105_SLICE_X8Y105_A6;
  wire [0:0] CLBLM_R_X7Y105_SLICE_X8Y105_AMUX;
  wire [0:0] CLBLM_R_X7Y105_SLICE_X8Y105_AO5;
  wire [0:0] CLBLM_R_X7Y105_SLICE_X8Y105_AO6;
  wire [0:0] CLBLM_R_X7Y105_SLICE_X8Y105_A_CY;
  wire [0:0] CLBLM_R_X7Y105_SLICE_X8Y105_A_XOR;
  wire [0:0] CLBLM_R_X7Y105_SLICE_X8Y105_B;
  wire [0:0] CLBLM_R_X7Y105_SLICE_X8Y105_B1;
  wire [0:0] CLBLM_R_X7Y105_SLICE_X8Y105_B2;
  wire [0:0] CLBLM_R_X7Y105_SLICE_X8Y105_B3;
  wire [0:0] CLBLM_R_X7Y105_SLICE_X8Y105_B4;
  wire [0:0] CLBLM_R_X7Y105_SLICE_X8Y105_B5;
  wire [0:0] CLBLM_R_X7Y105_SLICE_X8Y105_B6;
  wire [0:0] CLBLM_R_X7Y105_SLICE_X8Y105_BO5;
  wire [0:0] CLBLM_R_X7Y105_SLICE_X8Y105_BO6;
  wire [0:0] CLBLM_R_X7Y105_SLICE_X8Y105_B_CY;
  wire [0:0] CLBLM_R_X7Y105_SLICE_X8Y105_B_XOR;
  wire [0:0] CLBLM_R_X7Y105_SLICE_X8Y105_C;
  wire [0:0] CLBLM_R_X7Y105_SLICE_X8Y105_C1;
  wire [0:0] CLBLM_R_X7Y105_SLICE_X8Y105_C2;
  wire [0:0] CLBLM_R_X7Y105_SLICE_X8Y105_C3;
  wire [0:0] CLBLM_R_X7Y105_SLICE_X8Y105_C4;
  wire [0:0] CLBLM_R_X7Y105_SLICE_X8Y105_C5;
  wire [0:0] CLBLM_R_X7Y105_SLICE_X8Y105_C6;
  wire [0:0] CLBLM_R_X7Y105_SLICE_X8Y105_CO5;
  wire [0:0] CLBLM_R_X7Y105_SLICE_X8Y105_CO6;
  wire [0:0] CLBLM_R_X7Y105_SLICE_X8Y105_C_CY;
  wire [0:0] CLBLM_R_X7Y105_SLICE_X8Y105_C_XOR;
  wire [0:0] CLBLM_R_X7Y105_SLICE_X8Y105_D;
  wire [0:0] CLBLM_R_X7Y105_SLICE_X8Y105_D1;
  wire [0:0] CLBLM_R_X7Y105_SLICE_X8Y105_D2;
  wire [0:0] CLBLM_R_X7Y105_SLICE_X8Y105_D3;
  wire [0:0] CLBLM_R_X7Y105_SLICE_X8Y105_D4;
  wire [0:0] CLBLM_R_X7Y105_SLICE_X8Y105_D5;
  wire [0:0] CLBLM_R_X7Y105_SLICE_X8Y105_D6;
  wire [0:0] CLBLM_R_X7Y105_SLICE_X8Y105_DO5;
  wire [0:0] CLBLM_R_X7Y105_SLICE_X8Y105_DO6;
  wire [0:0] CLBLM_R_X7Y105_SLICE_X8Y105_D_CY;
  wire [0:0] CLBLM_R_X7Y105_SLICE_X8Y105_D_XOR;
  wire [0:0] CLBLM_R_X7Y105_SLICE_X9Y105_A;
  wire [0:0] CLBLM_R_X7Y105_SLICE_X9Y105_A1;
  wire [0:0] CLBLM_R_X7Y105_SLICE_X9Y105_A2;
  wire [0:0] CLBLM_R_X7Y105_SLICE_X9Y105_A3;
  wire [0:0] CLBLM_R_X7Y105_SLICE_X9Y105_A4;
  wire [0:0] CLBLM_R_X7Y105_SLICE_X9Y105_A5;
  wire [0:0] CLBLM_R_X7Y105_SLICE_X9Y105_A6;
  wire [0:0] CLBLM_R_X7Y105_SLICE_X9Y105_AO5;
  wire [0:0] CLBLM_R_X7Y105_SLICE_X9Y105_AO6;
  wire [0:0] CLBLM_R_X7Y105_SLICE_X9Y105_A_CY;
  wire [0:0] CLBLM_R_X7Y105_SLICE_X9Y105_A_XOR;
  wire [0:0] CLBLM_R_X7Y105_SLICE_X9Y105_B;
  wire [0:0] CLBLM_R_X7Y105_SLICE_X9Y105_B1;
  wire [0:0] CLBLM_R_X7Y105_SLICE_X9Y105_B2;
  wire [0:0] CLBLM_R_X7Y105_SLICE_X9Y105_B3;
  wire [0:0] CLBLM_R_X7Y105_SLICE_X9Y105_B4;
  wire [0:0] CLBLM_R_X7Y105_SLICE_X9Y105_B5;
  wire [0:0] CLBLM_R_X7Y105_SLICE_X9Y105_B6;
  wire [0:0] CLBLM_R_X7Y105_SLICE_X9Y105_BO5;
  wire [0:0] CLBLM_R_X7Y105_SLICE_X9Y105_BO6;
  wire [0:0] CLBLM_R_X7Y105_SLICE_X9Y105_B_CY;
  wire [0:0] CLBLM_R_X7Y105_SLICE_X9Y105_B_XOR;
  wire [0:0] CLBLM_R_X7Y105_SLICE_X9Y105_C;
  wire [0:0] CLBLM_R_X7Y105_SLICE_X9Y105_C1;
  wire [0:0] CLBLM_R_X7Y105_SLICE_X9Y105_C2;
  wire [0:0] CLBLM_R_X7Y105_SLICE_X9Y105_C3;
  wire [0:0] CLBLM_R_X7Y105_SLICE_X9Y105_C4;
  wire [0:0] CLBLM_R_X7Y105_SLICE_X9Y105_C5;
  wire [0:0] CLBLM_R_X7Y105_SLICE_X9Y105_C6;
  wire [0:0] CLBLM_R_X7Y105_SLICE_X9Y105_CO5;
  wire [0:0] CLBLM_R_X7Y105_SLICE_X9Y105_CO6;
  wire [0:0] CLBLM_R_X7Y105_SLICE_X9Y105_C_CY;
  wire [0:0] CLBLM_R_X7Y105_SLICE_X9Y105_C_XOR;
  wire [0:0] CLBLM_R_X7Y105_SLICE_X9Y105_D;
  wire [0:0] CLBLM_R_X7Y105_SLICE_X9Y105_D1;
  wire [0:0] CLBLM_R_X7Y105_SLICE_X9Y105_D2;
  wire [0:0] CLBLM_R_X7Y105_SLICE_X9Y105_D3;
  wire [0:0] CLBLM_R_X7Y105_SLICE_X9Y105_D4;
  wire [0:0] CLBLM_R_X7Y105_SLICE_X9Y105_D5;
  wire [0:0] CLBLM_R_X7Y105_SLICE_X9Y105_D6;
  wire [0:0] CLBLM_R_X7Y105_SLICE_X9Y105_DO5;
  wire [0:0] CLBLM_R_X7Y105_SLICE_X9Y105_DO6;
  wire [0:0] CLBLM_R_X7Y105_SLICE_X9Y105_D_CY;
  wire [0:0] CLBLM_R_X7Y105_SLICE_X9Y105_D_XOR;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X8Y106_A;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X8Y106_A1;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X8Y106_A2;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X8Y106_A3;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X8Y106_A4;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X8Y106_A5;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X8Y106_A6;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X8Y106_AMUX;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X8Y106_AO5;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X8Y106_AO6;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X8Y106_A_CY;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X8Y106_A_XOR;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X8Y106_B;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X8Y106_B1;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X8Y106_B2;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X8Y106_B3;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X8Y106_B4;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X8Y106_B5;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X8Y106_B6;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X8Y106_BO5;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X8Y106_BO6;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X8Y106_B_CY;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X8Y106_B_XOR;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X8Y106_C;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X8Y106_C1;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X8Y106_C2;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X8Y106_C3;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X8Y106_C4;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X8Y106_C5;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X8Y106_C6;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X8Y106_CMUX;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X8Y106_CO5;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X8Y106_CO6;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X8Y106_C_CY;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X8Y106_C_XOR;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X8Y106_D;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X8Y106_D1;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X8Y106_D2;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X8Y106_D3;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X8Y106_D4;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X8Y106_D5;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X8Y106_D6;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X8Y106_DO5;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X8Y106_DO6;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X8Y106_D_CY;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X8Y106_D_XOR;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X9Y106_A;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X9Y106_A1;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X9Y106_A2;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X9Y106_A3;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X9Y106_A4;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X9Y106_A5;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X9Y106_A6;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X9Y106_AO5;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X9Y106_AO6;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X9Y106_A_CY;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X9Y106_A_XOR;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X9Y106_B;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X9Y106_B1;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X9Y106_B2;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X9Y106_B3;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X9Y106_B4;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X9Y106_B5;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X9Y106_B6;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X9Y106_BO5;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X9Y106_BO6;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X9Y106_B_CY;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X9Y106_B_XOR;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X9Y106_C;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X9Y106_C1;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X9Y106_C2;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X9Y106_C3;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X9Y106_C4;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X9Y106_C5;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X9Y106_C6;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X9Y106_CO5;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X9Y106_CO6;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X9Y106_C_CY;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X9Y106_C_XOR;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X9Y106_D;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X9Y106_D1;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X9Y106_D2;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X9Y106_D3;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X9Y106_D4;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X9Y106_D5;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X9Y106_D6;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X9Y106_DO5;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X9Y106_DO6;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X9Y106_D_CY;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X9Y106_D_XOR;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X8Y107_A;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X8Y107_A1;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X8Y107_A2;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X8Y107_A3;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X8Y107_A4;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X8Y107_A5;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X8Y107_A6;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X8Y107_AMUX;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X8Y107_AO5;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X8Y107_AO6;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X8Y107_A_CY;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X8Y107_A_XOR;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X8Y107_B;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X8Y107_B1;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X8Y107_B2;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X8Y107_B3;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X8Y107_B4;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X8Y107_B5;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X8Y107_B6;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X8Y107_BO5;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X8Y107_BO6;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X8Y107_B_CY;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X8Y107_B_XOR;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X8Y107_C;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X8Y107_C1;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X8Y107_C2;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X8Y107_C3;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X8Y107_C4;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X8Y107_C5;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X8Y107_C6;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X8Y107_CO5;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X8Y107_CO6;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X8Y107_C_CY;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X8Y107_C_XOR;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X8Y107_D;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X8Y107_D1;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X8Y107_D2;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X8Y107_D3;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X8Y107_D4;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X8Y107_D5;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X8Y107_D6;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X8Y107_DO5;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X8Y107_DO6;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X8Y107_D_CY;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X8Y107_D_XOR;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X9Y107_A;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X9Y107_A1;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X9Y107_A2;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X9Y107_A3;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X9Y107_A4;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X9Y107_A5;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X9Y107_A6;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X9Y107_AO5;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X9Y107_AO6;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X9Y107_A_CY;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X9Y107_A_XOR;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X9Y107_B;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X9Y107_B1;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X9Y107_B2;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X9Y107_B3;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X9Y107_B4;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X9Y107_B5;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X9Y107_B6;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X9Y107_BMUX;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X9Y107_BO5;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X9Y107_BO6;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X9Y107_B_CY;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X9Y107_B_XOR;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X9Y107_C;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X9Y107_C1;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X9Y107_C2;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X9Y107_C3;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X9Y107_C4;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X9Y107_C5;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X9Y107_C6;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X9Y107_CMUX;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X9Y107_CO5;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X9Y107_CO6;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X9Y107_C_CY;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X9Y107_C_XOR;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X9Y107_D;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X9Y107_D1;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X9Y107_D2;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X9Y107_D3;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X9Y107_D4;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X9Y107_D5;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X9Y107_D6;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X9Y107_DO5;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X9Y107_DO6;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X9Y107_D_CY;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X9Y107_D_XOR;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X8Y108_A;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X8Y108_A1;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X8Y108_A2;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X8Y108_A3;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X8Y108_A4;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X8Y108_A5;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X8Y108_A6;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X8Y108_AMUX;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X8Y108_AO5;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X8Y108_AO6;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X8Y108_A_CY;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X8Y108_A_XOR;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X8Y108_B;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X8Y108_B1;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X8Y108_B2;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X8Y108_B3;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X8Y108_B4;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X8Y108_B5;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X8Y108_B6;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X8Y108_BO5;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X8Y108_BO6;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X8Y108_B_CY;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X8Y108_B_XOR;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X8Y108_C;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X8Y108_C1;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X8Y108_C2;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X8Y108_C3;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X8Y108_C4;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X8Y108_C5;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X8Y108_C6;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X8Y108_CO5;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X8Y108_CO6;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X8Y108_C_CY;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X8Y108_C_XOR;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X8Y108_D;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X8Y108_D1;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X8Y108_D2;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X8Y108_D3;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X8Y108_D4;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X8Y108_D5;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X8Y108_D6;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X8Y108_DO5;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X8Y108_DO6;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X8Y108_D_CY;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X8Y108_D_XOR;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X9Y108_A;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X9Y108_A1;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X9Y108_A2;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X9Y108_A3;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X9Y108_A4;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X9Y108_A5;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X9Y108_A6;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X9Y108_AO5;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X9Y108_AO6;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X9Y108_A_CY;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X9Y108_A_XOR;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X9Y108_B;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X9Y108_B1;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X9Y108_B2;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X9Y108_B3;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X9Y108_B4;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X9Y108_B5;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X9Y108_B6;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X9Y108_BMUX;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X9Y108_BO5;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X9Y108_BO6;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X9Y108_B_CY;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X9Y108_B_XOR;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X9Y108_C;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X9Y108_C1;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X9Y108_C2;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X9Y108_C3;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X9Y108_C4;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X9Y108_C5;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X9Y108_C6;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X9Y108_CO5;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X9Y108_CO6;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X9Y108_C_CY;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X9Y108_C_XOR;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X9Y108_D;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X9Y108_D1;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X9Y108_D2;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X9Y108_D3;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X9Y108_D4;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X9Y108_D5;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X9Y108_D6;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X9Y108_DO5;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X9Y108_DO6;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X9Y108_D_CY;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X9Y108_D_XOR;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X8Y109_A;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X8Y109_A1;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X8Y109_A2;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X8Y109_A3;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X8Y109_A4;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X8Y109_A5;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X8Y109_A6;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X8Y109_AMUX;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X8Y109_AO5;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X8Y109_AO6;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X8Y109_A_CY;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X8Y109_A_XOR;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X8Y109_B;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X8Y109_B1;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X8Y109_B2;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X8Y109_B3;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X8Y109_B4;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X8Y109_B5;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X8Y109_B6;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X8Y109_BO5;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X8Y109_BO6;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X8Y109_B_CY;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X8Y109_B_XOR;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X8Y109_C;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X8Y109_C1;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X8Y109_C2;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X8Y109_C3;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X8Y109_C4;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X8Y109_C5;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X8Y109_C6;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X8Y109_CO5;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X8Y109_CO6;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X8Y109_C_CY;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X8Y109_C_XOR;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X8Y109_D;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X8Y109_D1;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X8Y109_D2;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X8Y109_D3;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X8Y109_D4;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X8Y109_D5;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X8Y109_D6;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X8Y109_DO5;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X8Y109_DO6;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X8Y109_D_CY;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X8Y109_D_XOR;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X9Y109_A;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X9Y109_A1;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X9Y109_A2;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X9Y109_A3;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X9Y109_A4;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X9Y109_A5;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X9Y109_A6;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X9Y109_AMUX;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X9Y109_AO5;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X9Y109_AO6;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X9Y109_A_CY;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X9Y109_A_XOR;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X9Y109_B;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X9Y109_B1;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X9Y109_B2;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X9Y109_B3;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X9Y109_B4;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X9Y109_B5;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X9Y109_B6;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X9Y109_BO5;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X9Y109_BO6;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X9Y109_B_CY;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X9Y109_B_XOR;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X9Y109_C;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X9Y109_C1;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X9Y109_C2;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X9Y109_C3;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X9Y109_C4;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X9Y109_C5;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X9Y109_C6;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X9Y109_CO5;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X9Y109_CO6;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X9Y109_C_CY;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X9Y109_C_XOR;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X9Y109_D;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X9Y109_D1;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X9Y109_D2;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X9Y109_D3;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X9Y109_D4;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X9Y109_D5;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X9Y109_D6;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X9Y109_DO5;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X9Y109_DO6;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X9Y109_D_CY;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X9Y109_D_XOR;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X8Y110_A;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X8Y110_A1;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X8Y110_A2;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X8Y110_A3;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X8Y110_A4;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X8Y110_A5;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X8Y110_A6;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X8Y110_AO5;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X8Y110_AO6;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X8Y110_A_CY;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X8Y110_A_XOR;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X8Y110_B;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X8Y110_B1;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X8Y110_B2;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X8Y110_B3;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X8Y110_B4;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X8Y110_B5;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X8Y110_B6;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X8Y110_BMUX;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X8Y110_BO5;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X8Y110_BO6;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X8Y110_B_CY;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X8Y110_B_XOR;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X8Y110_C;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X8Y110_C1;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X8Y110_C2;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X8Y110_C3;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X8Y110_C4;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X8Y110_C5;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X8Y110_C6;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X8Y110_CO5;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X8Y110_CO6;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X8Y110_C_CY;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X8Y110_C_XOR;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X8Y110_D;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X8Y110_D1;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X8Y110_D2;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X8Y110_D3;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X8Y110_D4;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X8Y110_D5;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X8Y110_D6;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X8Y110_DO5;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X8Y110_DO6;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X8Y110_D_CY;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X8Y110_D_XOR;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X9Y110_A;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X9Y110_A1;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X9Y110_A2;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X9Y110_A3;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X9Y110_A4;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X9Y110_A5;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X9Y110_A6;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X9Y110_AMUX;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X9Y110_AO5;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X9Y110_AO6;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X9Y110_A_CY;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X9Y110_A_XOR;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X9Y110_B;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X9Y110_B1;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X9Y110_B2;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X9Y110_B3;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X9Y110_B4;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X9Y110_B5;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X9Y110_B6;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X9Y110_BMUX;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X9Y110_BO5;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X9Y110_BO6;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X9Y110_B_CY;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X9Y110_B_XOR;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X9Y110_C;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X9Y110_C1;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X9Y110_C2;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X9Y110_C3;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X9Y110_C4;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X9Y110_C5;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X9Y110_C6;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X9Y110_CMUX;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X9Y110_CO5;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X9Y110_CO6;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X9Y110_C_CY;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X9Y110_C_XOR;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X9Y110_D;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X9Y110_D1;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X9Y110_D2;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X9Y110_D3;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X9Y110_D4;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X9Y110_D5;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X9Y110_D6;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X9Y110_DO5;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X9Y110_DO6;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X9Y110_D_CY;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X9Y110_D_XOR;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X8Y111_A;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X8Y111_A1;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X8Y111_A2;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X8Y111_A3;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X8Y111_A4;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X8Y111_A5;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X8Y111_A6;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X8Y111_AMUX;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X8Y111_AO5;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X8Y111_AO6;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X8Y111_A_CY;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X8Y111_A_XOR;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X8Y111_B;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X8Y111_B1;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X8Y111_B2;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X8Y111_B3;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X8Y111_B4;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X8Y111_B5;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X8Y111_B6;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X8Y111_BO5;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X8Y111_BO6;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X8Y111_B_CY;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X8Y111_B_XOR;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X8Y111_C;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X8Y111_C1;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X8Y111_C2;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X8Y111_C3;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X8Y111_C4;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X8Y111_C5;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X8Y111_C6;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X8Y111_CO5;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X8Y111_CO6;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X8Y111_C_CY;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X8Y111_C_XOR;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X8Y111_D;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X8Y111_D1;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X8Y111_D2;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X8Y111_D3;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X8Y111_D4;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X8Y111_D5;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X8Y111_D6;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X8Y111_DO5;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X8Y111_DO6;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X8Y111_D_CY;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X8Y111_D_XOR;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X9Y111_A;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X9Y111_A1;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X9Y111_A2;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X9Y111_A3;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X9Y111_A4;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X9Y111_A5;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X9Y111_A6;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X9Y111_AMUX;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X9Y111_AO5;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X9Y111_AO6;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X9Y111_A_CY;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X9Y111_A_XOR;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X9Y111_B;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X9Y111_B1;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X9Y111_B2;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X9Y111_B3;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X9Y111_B4;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X9Y111_B5;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X9Y111_B6;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X9Y111_BO5;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X9Y111_BO6;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X9Y111_B_CY;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X9Y111_B_XOR;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X9Y111_C;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X9Y111_C1;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X9Y111_C2;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X9Y111_C3;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X9Y111_C4;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X9Y111_C5;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X9Y111_C6;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X9Y111_CO5;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X9Y111_CO6;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X9Y111_C_CY;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X9Y111_C_XOR;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X9Y111_D;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X9Y111_D1;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X9Y111_D2;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X9Y111_D3;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X9Y111_D4;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X9Y111_D5;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X9Y111_D6;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X9Y111_DO5;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X9Y111_DO6;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X9Y111_D_CY;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X9Y111_D_XOR;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X8Y112_A;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X8Y112_A1;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X8Y112_A2;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X8Y112_A3;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X8Y112_A4;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X8Y112_A5;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X8Y112_A6;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X8Y112_AMUX;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X8Y112_AO5;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X8Y112_AO6;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X8Y112_A_CY;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X8Y112_A_XOR;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X8Y112_B;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X8Y112_B1;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X8Y112_B2;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X8Y112_B3;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X8Y112_B4;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X8Y112_B5;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X8Y112_B6;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X8Y112_BO5;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X8Y112_BO6;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X8Y112_B_CY;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X8Y112_B_XOR;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X8Y112_C;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X8Y112_C1;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X8Y112_C2;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X8Y112_C3;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X8Y112_C4;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X8Y112_C5;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X8Y112_C6;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X8Y112_CO5;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X8Y112_CO6;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X8Y112_C_CY;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X8Y112_C_XOR;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X8Y112_D;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X8Y112_D1;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X8Y112_D2;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X8Y112_D3;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X8Y112_D4;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X8Y112_D5;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X8Y112_D6;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X8Y112_DO5;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X8Y112_DO6;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X8Y112_D_CY;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X8Y112_D_XOR;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X9Y112_A;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X9Y112_A1;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X9Y112_A2;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X9Y112_A3;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X9Y112_A4;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X9Y112_A5;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X9Y112_A6;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X9Y112_AO5;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X9Y112_AO6;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X9Y112_A_CY;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X9Y112_A_XOR;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X9Y112_B;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X9Y112_B1;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X9Y112_B2;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X9Y112_B3;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X9Y112_B4;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X9Y112_B5;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X9Y112_B6;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X9Y112_BO5;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X9Y112_BO6;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X9Y112_B_CY;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X9Y112_B_XOR;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X9Y112_C;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X9Y112_C1;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X9Y112_C2;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X9Y112_C3;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X9Y112_C4;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X9Y112_C5;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X9Y112_C6;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X9Y112_CO5;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X9Y112_CO6;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X9Y112_C_CY;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X9Y112_C_XOR;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X9Y112_D;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X9Y112_D1;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X9Y112_D2;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X9Y112_D3;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X9Y112_D4;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X9Y112_D5;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X9Y112_D6;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X9Y112_DO5;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X9Y112_DO6;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X9Y112_D_CY;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X9Y112_D_XOR;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X8Y113_A;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X8Y113_A1;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X8Y113_A2;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X8Y113_A3;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X8Y113_A4;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X8Y113_A5;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X8Y113_A6;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X8Y113_AMUX;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X8Y113_AO5;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X8Y113_AO6;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X8Y113_A_CY;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X8Y113_A_XOR;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X8Y113_B;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X8Y113_B1;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X8Y113_B2;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X8Y113_B3;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X8Y113_B4;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X8Y113_B5;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X8Y113_B6;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X8Y113_BMUX;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X8Y113_BO5;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X8Y113_BO6;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X8Y113_B_CY;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X8Y113_B_XOR;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X8Y113_C;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X8Y113_C1;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X8Y113_C2;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X8Y113_C3;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X8Y113_C4;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X8Y113_C5;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X8Y113_C6;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X8Y113_CO5;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X8Y113_CO6;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X8Y113_C_CY;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X8Y113_C_XOR;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X8Y113_D;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X8Y113_D1;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X8Y113_D2;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X8Y113_D3;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X8Y113_D4;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X8Y113_D5;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X8Y113_D6;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X8Y113_DO5;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X8Y113_DO6;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X8Y113_D_CY;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X8Y113_D_XOR;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X9Y113_A;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X9Y113_A1;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X9Y113_A2;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X9Y113_A3;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X9Y113_A4;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X9Y113_A5;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X9Y113_A6;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X9Y113_AO5;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X9Y113_AO6;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X9Y113_A_CY;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X9Y113_A_XOR;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X9Y113_B;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X9Y113_B1;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X9Y113_B2;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X9Y113_B3;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X9Y113_B4;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X9Y113_B5;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X9Y113_B6;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X9Y113_BO5;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X9Y113_BO6;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X9Y113_B_CY;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X9Y113_B_XOR;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X9Y113_C;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X9Y113_C1;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X9Y113_C2;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X9Y113_C3;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X9Y113_C4;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X9Y113_C5;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X9Y113_C6;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X9Y113_CO5;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X9Y113_CO6;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X9Y113_C_CY;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X9Y113_C_XOR;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X9Y113_D;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X9Y113_D1;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X9Y113_D2;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X9Y113_D3;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X9Y113_D4;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X9Y113_D5;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X9Y113_D6;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X9Y113_DO5;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X9Y113_DO6;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X9Y113_D_CY;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X9Y113_D_XOR;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X8Y114_A;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X8Y114_A1;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X8Y114_A2;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X8Y114_A3;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X8Y114_A4;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X8Y114_A5;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X8Y114_A6;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X8Y114_AMUX;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X8Y114_AO5;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X8Y114_AO6;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X8Y114_A_CY;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X8Y114_A_XOR;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X8Y114_B;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X8Y114_B1;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X8Y114_B2;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X8Y114_B3;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X8Y114_B4;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X8Y114_B5;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X8Y114_B6;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X8Y114_BO5;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X8Y114_BO6;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X8Y114_B_CY;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X8Y114_B_XOR;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X8Y114_C;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X8Y114_C1;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X8Y114_C2;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X8Y114_C3;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X8Y114_C4;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X8Y114_C5;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X8Y114_C6;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X8Y114_CO5;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X8Y114_CO6;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X8Y114_C_CY;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X8Y114_C_XOR;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X8Y114_D;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X8Y114_D1;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X8Y114_D2;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X8Y114_D3;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X8Y114_D4;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X8Y114_D5;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X8Y114_D6;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X8Y114_DO5;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X8Y114_DO6;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X8Y114_D_CY;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X8Y114_D_XOR;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X9Y114_A;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X9Y114_A1;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X9Y114_A2;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X9Y114_A3;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X9Y114_A4;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X9Y114_A5;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X9Y114_A6;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X9Y114_AO5;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X9Y114_AO6;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X9Y114_A_CY;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X9Y114_A_XOR;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X9Y114_B;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X9Y114_B1;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X9Y114_B2;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X9Y114_B3;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X9Y114_B4;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X9Y114_B5;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X9Y114_B6;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X9Y114_BO5;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X9Y114_BO6;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X9Y114_B_CY;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X9Y114_B_XOR;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X9Y114_C;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X9Y114_C1;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X9Y114_C2;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X9Y114_C3;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X9Y114_C4;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X9Y114_C5;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X9Y114_C6;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X9Y114_CO5;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X9Y114_CO6;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X9Y114_C_CY;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X9Y114_C_XOR;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X9Y114_D;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X9Y114_D1;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X9Y114_D2;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X9Y114_D3;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X9Y114_D4;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X9Y114_D5;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X9Y114_D6;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X9Y114_DO5;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X9Y114_DO6;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X9Y114_D_CY;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X9Y114_D_XOR;
  wire [0:0] LIOB33_SING_X0Y100_IOB_X0Y100_I;
  wire [0:0] LIOB33_SING_X0Y149_IOB_X0Y149_O;
  wire [0:0] LIOB33_X0Y101_IOB_X0Y101_I;
  wire [0:0] LIOB33_X0Y101_IOB_X0Y102_I;
  wire [0:0] LIOB33_X0Y103_IOB_X0Y103_I;
  wire [0:0] LIOB33_X0Y103_IOB_X0Y104_I;
  wire [0:0] LIOB33_X0Y105_IOB_X0Y105_I;
  wire [0:0] LIOB33_X0Y105_IOB_X0Y106_I;
  wire [0:0] LIOB33_X0Y107_IOB_X0Y107_I;
  wire [0:0] LIOB33_X0Y107_IOB_X0Y108_I;
  wire [0:0] LIOB33_X0Y109_IOB_X0Y109_I;
  wire [0:0] LIOB33_X0Y109_IOB_X0Y110_I;
  wire [0:0] LIOB33_X0Y111_IOB_X0Y111_I;
  wire [0:0] LIOB33_X0Y111_IOB_X0Y112_I;
  wire [0:0] LIOB33_X0Y113_IOB_X0Y113_I;
  wire [0:0] LIOB33_X0Y113_IOB_X0Y114_I;
  wire [0:0] LIOB33_X0Y115_IOB_X0Y115_I;
  wire [0:0] LIOB33_X0Y115_IOB_X0Y116_I;
  wire [0:0] LIOB33_X0Y117_IOB_X0Y117_I;
  wire [0:0] LIOB33_X0Y117_IOB_X0Y118_O;
  wire [0:0] LIOB33_X0Y119_IOB_X0Y119_O;
  wire [0:0] LIOB33_X0Y119_IOB_X0Y120_O;
  wire [0:0] LIOB33_X0Y121_IOB_X0Y121_O;
  wire [0:0] LIOB33_X0Y121_IOB_X0Y122_O;
  wire [0:0] LIOB33_X0Y123_IOB_X0Y123_O;
  wire [0:0] LIOB33_X0Y123_IOB_X0Y124_O;
  wire [0:0] LIOB33_X0Y125_IOB_X0Y125_O;
  wire [0:0] LIOB33_X0Y125_IOB_X0Y126_O;
  wire [0:0] LIOB33_X0Y127_IOB_X0Y127_O;
  wire [0:0] LIOB33_X0Y127_IOB_X0Y128_O;
  wire [0:0] LIOB33_X0Y129_IOB_X0Y129_O;
  wire [0:0] LIOB33_X0Y129_IOB_X0Y130_O;
  wire [0:0] LIOB33_X0Y131_IOB_X0Y131_O;
  wire [0:0] LIOB33_X0Y131_IOB_X0Y132_O;
  wire [0:0] LIOB33_X0Y133_IOB_X0Y133_O;
  wire [0:0] LIOB33_X0Y133_IOB_X0Y134_O;
  wire [0:0] LIOB33_X0Y135_IOB_X0Y135_O;
  wire [0:0] LIOB33_X0Y135_IOB_X0Y136_O;
  wire [0:0] LIOB33_X0Y137_IOB_X0Y137_O;
  wire [0:0] LIOB33_X0Y137_IOB_X0Y138_O;
  wire [0:0] LIOB33_X0Y139_IOB_X0Y139_O;
  wire [0:0] LIOB33_X0Y139_IOB_X0Y140_O;
  wire [0:0] LIOB33_X0Y141_IOB_X0Y141_O;
  wire [0:0] LIOB33_X0Y141_IOB_X0Y142_O;
  wire [0:0] LIOB33_X0Y143_IOB_X0Y143_O;
  wire [0:0] LIOB33_X0Y145_IOB_X0Y145_O;
  wire [0:0] LIOB33_X0Y145_IOB_X0Y146_O;
  wire [0:0] LIOB33_X0Y147_IOB_X0Y147_O;
  wire [0:0] LIOB33_X0Y147_IOB_X0Y148_O;
  wire [0:0] LIOI3_SING_X0Y100_ILOGIC_X0Y100_D;
  wire [0:0] LIOI3_SING_X0Y100_ILOGIC_X0Y100_O;
  wire [0:0] LIOI3_SING_X0Y149_OLOGIC_X0Y149_D1;
  wire [0:0] LIOI3_SING_X0Y149_OLOGIC_X0Y149_OQ;
  wire [0:0] LIOI3_SING_X0Y149_OLOGIC_X0Y149_T1;
  wire [0:0] LIOI3_SING_X0Y149_OLOGIC_X0Y149_TQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y107_ILOGIC_X0Y107_D;
  wire [0:0] LIOI3_TBYTESRC_X0Y107_ILOGIC_X0Y107_O;
  wire [0:0] LIOI3_TBYTESRC_X0Y107_ILOGIC_X0Y108_D;
  wire [0:0] LIOI3_TBYTESRC_X0Y107_ILOGIC_X0Y108_O;
  wire [0:0] LIOI3_TBYTESRC_X0Y119_OLOGIC_X0Y119_D1;
  wire [0:0] LIOI3_TBYTESRC_X0Y119_OLOGIC_X0Y119_OQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y119_OLOGIC_X0Y119_T1;
  wire [0:0] LIOI3_TBYTESRC_X0Y119_OLOGIC_X0Y119_TQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y119_OLOGIC_X0Y120_D1;
  wire [0:0] LIOI3_TBYTESRC_X0Y119_OLOGIC_X0Y120_OQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y119_OLOGIC_X0Y120_T1;
  wire [0:0] LIOI3_TBYTESRC_X0Y119_OLOGIC_X0Y120_TQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y131_OLOGIC_X0Y131_D1;
  wire [0:0] LIOI3_TBYTESRC_X0Y131_OLOGIC_X0Y131_OQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y131_OLOGIC_X0Y131_T1;
  wire [0:0] LIOI3_TBYTESRC_X0Y131_OLOGIC_X0Y131_TQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y131_OLOGIC_X0Y132_D1;
  wire [0:0] LIOI3_TBYTESRC_X0Y131_OLOGIC_X0Y132_OQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y131_OLOGIC_X0Y132_T1;
  wire [0:0] LIOI3_TBYTESRC_X0Y131_OLOGIC_X0Y132_TQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y143_OLOGIC_X0Y143_D1;
  wire [0:0] LIOI3_TBYTESRC_X0Y143_OLOGIC_X0Y143_OQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y143_OLOGIC_X0Y143_T1;
  wire [0:0] LIOI3_TBYTESRC_X0Y143_OLOGIC_X0Y143_TQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y143_OLOGIC_X0Y144_D1;
  wire [0:0] LIOI3_TBYTESRC_X0Y143_OLOGIC_X0Y144_OQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y143_OLOGIC_X0Y144_T1;
  wire [0:0] LIOI3_TBYTESRC_X0Y143_OLOGIC_X0Y144_TQ;
  wire [0:0] LIOI3_TBYTETERM_X0Y113_ILOGIC_X0Y113_D;
  wire [0:0] LIOI3_TBYTETERM_X0Y113_ILOGIC_X0Y113_O;
  wire [0:0] LIOI3_TBYTETERM_X0Y113_ILOGIC_X0Y114_D;
  wire [0:0] LIOI3_TBYTETERM_X0Y113_ILOGIC_X0Y114_O;
  wire [0:0] LIOI3_TBYTETERM_X0Y137_OLOGIC_X0Y137_D1;
  wire [0:0] LIOI3_TBYTETERM_X0Y137_OLOGIC_X0Y137_OQ;
  wire [0:0] LIOI3_TBYTETERM_X0Y137_OLOGIC_X0Y137_T1;
  wire [0:0] LIOI3_TBYTETERM_X0Y137_OLOGIC_X0Y137_TQ;
  wire [0:0] LIOI3_TBYTETERM_X0Y137_OLOGIC_X0Y138_D1;
  wire [0:0] LIOI3_TBYTETERM_X0Y137_OLOGIC_X0Y138_OQ;
  wire [0:0] LIOI3_TBYTETERM_X0Y137_OLOGIC_X0Y138_T1;
  wire [0:0] LIOI3_TBYTETERM_X0Y137_OLOGIC_X0Y138_TQ;
  wire [0:0] LIOI3_X0Y101_ILOGIC_X0Y101_D;
  wire [0:0] LIOI3_X0Y101_ILOGIC_X0Y101_O;
  wire [0:0] LIOI3_X0Y101_ILOGIC_X0Y102_D;
  wire [0:0] LIOI3_X0Y101_ILOGIC_X0Y102_O;
  wire [0:0] LIOI3_X0Y103_ILOGIC_X0Y103_D;
  wire [0:0] LIOI3_X0Y103_ILOGIC_X0Y103_O;
  wire [0:0] LIOI3_X0Y103_ILOGIC_X0Y104_D;
  wire [0:0] LIOI3_X0Y103_ILOGIC_X0Y104_O;
  wire [0:0] LIOI3_X0Y105_ILOGIC_X0Y105_D;
  wire [0:0] LIOI3_X0Y105_ILOGIC_X0Y105_O;
  wire [0:0] LIOI3_X0Y105_ILOGIC_X0Y106_D;
  wire [0:0] LIOI3_X0Y105_ILOGIC_X0Y106_O;
  wire [0:0] LIOI3_X0Y109_ILOGIC_X0Y109_D;
  wire [0:0] LIOI3_X0Y109_ILOGIC_X0Y109_O;
  wire [0:0] LIOI3_X0Y109_ILOGIC_X0Y110_D;
  wire [0:0] LIOI3_X0Y109_ILOGIC_X0Y110_O;
  wire [0:0] LIOI3_X0Y111_ILOGIC_X0Y111_D;
  wire [0:0] LIOI3_X0Y111_ILOGIC_X0Y111_O;
  wire [0:0] LIOI3_X0Y111_ILOGIC_X0Y112_D;
  wire [0:0] LIOI3_X0Y111_ILOGIC_X0Y112_O;
  wire [0:0] LIOI3_X0Y115_ILOGIC_X0Y115_D;
  wire [0:0] LIOI3_X0Y115_ILOGIC_X0Y115_O;
  wire [0:0] LIOI3_X0Y115_ILOGIC_X0Y116_D;
  wire [0:0] LIOI3_X0Y115_ILOGIC_X0Y116_O;
  wire [0:0] LIOI3_X0Y117_ILOGIC_X0Y117_D;
  wire [0:0] LIOI3_X0Y117_ILOGIC_X0Y117_O;
  wire [0:0] LIOI3_X0Y117_OLOGIC_X0Y118_D1;
  wire [0:0] LIOI3_X0Y117_OLOGIC_X0Y118_OQ;
  wire [0:0] LIOI3_X0Y117_OLOGIC_X0Y118_T1;
  wire [0:0] LIOI3_X0Y117_OLOGIC_X0Y118_TQ;
  wire [0:0] LIOI3_X0Y121_OLOGIC_X0Y121_D1;
  wire [0:0] LIOI3_X0Y121_OLOGIC_X0Y121_OQ;
  wire [0:0] LIOI3_X0Y121_OLOGIC_X0Y121_T1;
  wire [0:0] LIOI3_X0Y121_OLOGIC_X0Y121_TQ;
  wire [0:0] LIOI3_X0Y121_OLOGIC_X0Y122_D1;
  wire [0:0] LIOI3_X0Y121_OLOGIC_X0Y122_OQ;
  wire [0:0] LIOI3_X0Y121_OLOGIC_X0Y122_T1;
  wire [0:0] LIOI3_X0Y121_OLOGIC_X0Y122_TQ;
  wire [0:0] LIOI3_X0Y123_OLOGIC_X0Y123_D1;
  wire [0:0] LIOI3_X0Y123_OLOGIC_X0Y123_OQ;
  wire [0:0] LIOI3_X0Y123_OLOGIC_X0Y123_T1;
  wire [0:0] LIOI3_X0Y123_OLOGIC_X0Y123_TQ;
  wire [0:0] LIOI3_X0Y123_OLOGIC_X0Y124_D1;
  wire [0:0] LIOI3_X0Y123_OLOGIC_X0Y124_OQ;
  wire [0:0] LIOI3_X0Y123_OLOGIC_X0Y124_T1;
  wire [0:0] LIOI3_X0Y123_OLOGIC_X0Y124_TQ;
  wire [0:0] LIOI3_X0Y125_OLOGIC_X0Y125_D1;
  wire [0:0] LIOI3_X0Y125_OLOGIC_X0Y125_OQ;
  wire [0:0] LIOI3_X0Y125_OLOGIC_X0Y125_T1;
  wire [0:0] LIOI3_X0Y125_OLOGIC_X0Y125_TQ;
  wire [0:0] LIOI3_X0Y125_OLOGIC_X0Y126_D1;
  wire [0:0] LIOI3_X0Y125_OLOGIC_X0Y126_OQ;
  wire [0:0] LIOI3_X0Y125_OLOGIC_X0Y126_T1;
  wire [0:0] LIOI3_X0Y125_OLOGIC_X0Y126_TQ;
  wire [0:0] LIOI3_X0Y127_OLOGIC_X0Y127_D1;
  wire [0:0] LIOI3_X0Y127_OLOGIC_X0Y127_OQ;
  wire [0:0] LIOI3_X0Y127_OLOGIC_X0Y127_T1;
  wire [0:0] LIOI3_X0Y127_OLOGIC_X0Y127_TQ;
  wire [0:0] LIOI3_X0Y127_OLOGIC_X0Y128_D1;
  wire [0:0] LIOI3_X0Y127_OLOGIC_X0Y128_OQ;
  wire [0:0] LIOI3_X0Y127_OLOGIC_X0Y128_T1;
  wire [0:0] LIOI3_X0Y127_OLOGIC_X0Y128_TQ;
  wire [0:0] LIOI3_X0Y129_OLOGIC_X0Y129_D1;
  wire [0:0] LIOI3_X0Y129_OLOGIC_X0Y129_OQ;
  wire [0:0] LIOI3_X0Y129_OLOGIC_X0Y129_T1;
  wire [0:0] LIOI3_X0Y129_OLOGIC_X0Y129_TQ;
  wire [0:0] LIOI3_X0Y129_OLOGIC_X0Y130_D1;
  wire [0:0] LIOI3_X0Y129_OLOGIC_X0Y130_OQ;
  wire [0:0] LIOI3_X0Y129_OLOGIC_X0Y130_T1;
  wire [0:0] LIOI3_X0Y129_OLOGIC_X0Y130_TQ;
  wire [0:0] LIOI3_X0Y133_OLOGIC_X0Y133_D1;
  wire [0:0] LIOI3_X0Y133_OLOGIC_X0Y133_OQ;
  wire [0:0] LIOI3_X0Y133_OLOGIC_X0Y133_T1;
  wire [0:0] LIOI3_X0Y133_OLOGIC_X0Y133_TQ;
  wire [0:0] LIOI3_X0Y133_OLOGIC_X0Y134_D1;
  wire [0:0] LIOI3_X0Y133_OLOGIC_X0Y134_OQ;
  wire [0:0] LIOI3_X0Y133_OLOGIC_X0Y134_T1;
  wire [0:0] LIOI3_X0Y133_OLOGIC_X0Y134_TQ;
  wire [0:0] LIOI3_X0Y135_OLOGIC_X0Y135_D1;
  wire [0:0] LIOI3_X0Y135_OLOGIC_X0Y135_OQ;
  wire [0:0] LIOI3_X0Y135_OLOGIC_X0Y135_T1;
  wire [0:0] LIOI3_X0Y135_OLOGIC_X0Y135_TQ;
  wire [0:0] LIOI3_X0Y135_OLOGIC_X0Y136_D1;
  wire [0:0] LIOI3_X0Y135_OLOGIC_X0Y136_OQ;
  wire [0:0] LIOI3_X0Y135_OLOGIC_X0Y136_T1;
  wire [0:0] LIOI3_X0Y135_OLOGIC_X0Y136_TQ;
  wire [0:0] LIOI3_X0Y139_OLOGIC_X0Y139_D1;
  wire [0:0] LIOI3_X0Y139_OLOGIC_X0Y139_OQ;
  wire [0:0] LIOI3_X0Y139_OLOGIC_X0Y139_T1;
  wire [0:0] LIOI3_X0Y139_OLOGIC_X0Y139_TQ;
  wire [0:0] LIOI3_X0Y139_OLOGIC_X0Y140_D1;
  wire [0:0] LIOI3_X0Y139_OLOGIC_X0Y140_OQ;
  wire [0:0] LIOI3_X0Y139_OLOGIC_X0Y140_T1;
  wire [0:0] LIOI3_X0Y139_OLOGIC_X0Y140_TQ;
  wire [0:0] LIOI3_X0Y141_OLOGIC_X0Y141_D1;
  wire [0:0] LIOI3_X0Y141_OLOGIC_X0Y141_OQ;
  wire [0:0] LIOI3_X0Y141_OLOGIC_X0Y141_T1;
  wire [0:0] LIOI3_X0Y141_OLOGIC_X0Y141_TQ;
  wire [0:0] LIOI3_X0Y141_OLOGIC_X0Y142_D1;
  wire [0:0] LIOI3_X0Y141_OLOGIC_X0Y142_OQ;
  wire [0:0] LIOI3_X0Y141_OLOGIC_X0Y142_T1;
  wire [0:0] LIOI3_X0Y141_OLOGIC_X0Y142_TQ;
  wire [0:0] LIOI3_X0Y145_OLOGIC_X0Y145_D1;
  wire [0:0] LIOI3_X0Y145_OLOGIC_X0Y145_OQ;
  wire [0:0] LIOI3_X0Y145_OLOGIC_X0Y145_T1;
  wire [0:0] LIOI3_X0Y145_OLOGIC_X0Y145_TQ;
  wire [0:0] LIOI3_X0Y145_OLOGIC_X0Y146_D1;
  wire [0:0] LIOI3_X0Y145_OLOGIC_X0Y146_OQ;
  wire [0:0] LIOI3_X0Y145_OLOGIC_X0Y146_T1;
  wire [0:0] LIOI3_X0Y145_OLOGIC_X0Y146_TQ;
  wire [0:0] LIOI3_X0Y147_OLOGIC_X0Y147_D1;
  wire [0:0] LIOI3_X0Y147_OLOGIC_X0Y147_OQ;
  wire [0:0] LIOI3_X0Y147_OLOGIC_X0Y147_T1;
  wire [0:0] LIOI3_X0Y147_OLOGIC_X0Y147_TQ;
  wire [0:0] LIOI3_X0Y147_OLOGIC_X0Y148_D1;
  wire [0:0] LIOI3_X0Y147_OLOGIC_X0Y148_OQ;
  wire [0:0] LIOI3_X0Y147_OLOGIC_X0Y148_T1;
  wire [0:0] LIOI3_X0Y147_OLOGIC_X0Y148_TQ;
  wire [0:0] RIOB33_SING_X105Y100_IOB_X1Y100_I;
  wire [0:0] RIOB33_X105Y101_IOB_X1Y101_I;
  wire [0:0] RIOB33_X105Y101_IOB_X1Y102_I;
  wire [0:0] RIOB33_X105Y103_IOB_X1Y103_I;
  wire [0:0] RIOB33_X105Y103_IOB_X1Y104_I;
  wire [0:0] RIOB33_X105Y105_IOB_X1Y105_I;
  wire [0:0] RIOB33_X105Y105_IOB_X1Y106_I;
  wire [0:0] RIOB33_X105Y107_IOB_X1Y107_I;
  wire [0:0] RIOB33_X105Y107_IOB_X1Y108_I;
  wire [0:0] RIOB33_X105Y109_IOB_X1Y109_I;
  wire [0:0] RIOB33_X105Y109_IOB_X1Y110_I;
  wire [0:0] RIOB33_X105Y111_IOB_X1Y111_I;
  wire [0:0] RIOB33_X105Y111_IOB_X1Y112_I;
  wire [0:0] RIOB33_X105Y113_IOB_X1Y113_I;
  wire [0:0] RIOI3_SING_X105Y100_ILOGIC_X1Y100_D;
  wire [0:0] RIOI3_SING_X105Y100_ILOGIC_X1Y100_O;
  wire [0:0] RIOI3_TBYTESRC_X105Y107_ILOGIC_X1Y107_D;
  wire [0:0] RIOI3_TBYTESRC_X105Y107_ILOGIC_X1Y107_O;
  wire [0:0] RIOI3_TBYTESRC_X105Y107_ILOGIC_X1Y108_D;
  wire [0:0] RIOI3_TBYTESRC_X105Y107_ILOGIC_X1Y108_O;
  wire [0:0] RIOI3_TBYTETERM_X105Y113_ILOGIC_X1Y113_D;
  wire [0:0] RIOI3_TBYTETERM_X105Y113_ILOGIC_X1Y113_O;
  wire [0:0] RIOI3_X105Y101_ILOGIC_X1Y101_D;
  wire [0:0] RIOI3_X105Y101_ILOGIC_X1Y101_O;
  wire [0:0] RIOI3_X105Y101_ILOGIC_X1Y102_D;
  wire [0:0] RIOI3_X105Y101_ILOGIC_X1Y102_O;
  wire [0:0] RIOI3_X105Y103_ILOGIC_X1Y103_D;
  wire [0:0] RIOI3_X105Y103_ILOGIC_X1Y103_O;
  wire [0:0] RIOI3_X105Y103_ILOGIC_X1Y104_D;
  wire [0:0] RIOI3_X105Y103_ILOGIC_X1Y104_O;
  wire [0:0] RIOI3_X105Y105_ILOGIC_X1Y105_D;
  wire [0:0] RIOI3_X105Y105_ILOGIC_X1Y105_O;
  wire [0:0] RIOI3_X105Y105_ILOGIC_X1Y106_D;
  wire [0:0] RIOI3_X105Y105_ILOGIC_X1Y106_O;
  wire [0:0] RIOI3_X105Y109_ILOGIC_X1Y109_D;
  wire [0:0] RIOI3_X105Y109_ILOGIC_X1Y109_O;
  wire [0:0] RIOI3_X105Y109_ILOGIC_X1Y110_D;
  wire [0:0] RIOI3_X105Y109_ILOGIC_X1Y110_O;
  wire [0:0] RIOI3_X105Y111_ILOGIC_X1Y111_D;
  wire [0:0] RIOI3_X105Y111_ILOGIC_X1Y111_O;
  wire [0:0] RIOI3_X105Y111_ILOGIC_X1Y112_D;
  wire [0:0] RIOI3_X105Y111_ILOGIC_X1Y112_O;


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y104_SLICE_X0Y104_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y104_SLICE_X0Y104_DO5),
.O6(CLBLL_L_X2Y104_SLICE_X0Y104_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h13b1220000aa2200)
  ) CLBLL_L_X2Y104_SLICE_X0Y104_CLUT (
.I0(LIOB33_X0Y103_IOB_X0Y103_I),
.I1(RIOB33_X105Y105_IOB_X1Y106_I),
.I2(RIOB33_X105Y111_IOB_X1Y112_I),
.I3(LIOB33_SING_X0Y100_IOB_X0Y100_I),
.I4(RIOB33_X105Y113_IOB_X1Y113_I),
.I5(LIOB33_X0Y113_IOB_X0Y114_I),
.O5(CLBLL_L_X2Y104_SLICE_X0Y104_CO5),
.O6(CLBLL_L_X2Y104_SLICE_X0Y104_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h13a03c3043f0ccc0)
  ) CLBLL_L_X2Y104_SLICE_X0Y104_BLUT (
.I0(RIOB33_X105Y111_IOB_X1Y112_I),
.I1(RIOB33_X105Y105_IOB_X1Y106_I),
.I2(RIOB33_X105Y113_IOB_X1Y113_I),
.I3(LIOB33_SING_X0Y100_IOB_X0Y100_I),
.I4(LIOB33_X0Y103_IOB_X0Y103_I),
.I5(LIOB33_X0Y113_IOB_X0Y114_I),
.O5(CLBLL_L_X2Y104_SLICE_X0Y104_BO5),
.O6(CLBLL_L_X2Y104_SLICE_X0Y104_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h939393930f0fffff)
  ) CLBLL_L_X2Y104_SLICE_X0Y104_ALUT (
.I0(RIOB33_SING_X105Y100_IOB_X1Y100_I),
.I1(CLBLL_L_X2Y104_SLICE_X1Y104_BO6),
.I2(LIOB33_X0Y103_IOB_X0Y104_I),
.I3(1'b1),
.I4(LIOB33_X0Y103_IOB_X0Y103_I),
.I5(1'b1),
.O5(CLBLL_L_X2Y104_SLICE_X0Y104_AO5),
.O6(CLBLL_L_X2Y104_SLICE_X0Y104_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hc3699999693ccccc)
  ) CLBLL_L_X2Y104_SLICE_X1Y104_DLUT (
.I0(CLBLL_L_X2Y104_SLICE_X1Y104_AO6),
.I1(CLBLM_R_X3Y104_SLICE_X2Y104_BO6),
.I2(LIOB33_X0Y103_IOB_X0Y103_I),
.I3(RIOB33_X105Y105_IOB_X1Y106_I),
.I4(LIOB33_X0Y101_IOB_X0Y102_I),
.I5(CLBLM_R_X3Y104_SLICE_X2Y104_AO6),
.O5(CLBLL_L_X2Y104_SLICE_X1Y104_DO5),
.O6(CLBLL_L_X2Y104_SLICE_X1Y104_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h67cd983265cf9a30)
  ) CLBLL_L_X2Y104_SLICE_X1Y104_CLUT (
.I0(LIOB33_X0Y101_IOB_X0Y101_I),
.I1(CLBLL_L_X2Y104_SLICE_X0Y104_CO6),
.I2(CLBLL_L_X2Y104_SLICE_X0Y104_BO6),
.I3(LIOB33_X0Y103_IOB_X0Y103_I),
.I4(CLBLM_R_X3Y105_SLICE_X2Y105_AO6),
.I5(RIOB33_X105Y105_IOB_X1Y106_I),
.O5(CLBLL_L_X2Y104_SLICE_X1Y104_CO5),
.O6(CLBLL_L_X2Y104_SLICE_X1Y104_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hc93969996c9c3ccc)
  ) CLBLL_L_X2Y104_SLICE_X1Y104_BLUT (
.I0(CLBLL_L_X2Y106_SLICE_X1Y106_AO5),
.I1(CLBLL_L_X2Y104_SLICE_X1Y104_CO6),
.I2(LIOB33_X0Y101_IOB_X0Y102_I),
.I3(RIOB33_X105Y105_IOB_X1Y106_I),
.I4(RIOB33_SING_X105Y100_IOB_X1Y100_I),
.I5(CLBLL_L_X2Y104_SLICE_X1Y104_AO5),
.O5(CLBLL_L_X2Y104_SLICE_X1Y104_BO5),
.O6(CLBLL_L_X2Y104_SLICE_X1Y104_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hf1f1f3f399993333)
  ) CLBLL_L_X2Y104_SLICE_X1Y104_ALUT (
.I0(RIOB33_X105Y105_IOB_X1Y106_I),
.I1(CLBLL_L_X2Y104_SLICE_X0Y104_BO6),
.I2(CLBLL_L_X2Y104_SLICE_X0Y104_CO6),
.I3(1'b1),
.I4(LIOB33_X0Y101_IOB_X0Y101_I),
.I5(1'b1),
.O5(CLBLL_L_X2Y104_SLICE_X1Y104_AO5),
.O6(CLBLL_L_X2Y104_SLICE_X1Y104_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y106_SLICE_X0Y106_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y106_SLICE_X0Y106_DO5),
.O6(CLBLL_L_X2Y106_SLICE_X0Y106_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y106_SLICE_X0Y106_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y106_SLICE_X0Y106_CO5),
.O6(CLBLL_L_X2Y106_SLICE_X0Y106_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h4d8eddeecf0cffcc)
  ) CLBLL_L_X2Y106_SLICE_X0Y106_BLUT (
.I0(RIOB33_X105Y105_IOB_X1Y106_I),
.I1(CLBLL_L_X2Y106_SLICE_X1Y106_DO6),
.I2(LIOB33_X0Y103_IOB_X0Y104_I),
.I3(CLBLL_L_X2Y104_SLICE_X1Y104_CO6),
.I4(RIOB33_SING_X105Y100_IOB_X1Y100_I),
.I5(LIOB33_X0Y101_IOB_X0Y102_I),
.O5(CLBLL_L_X2Y106_SLICE_X0Y106_BO5),
.O6(CLBLL_L_X2Y106_SLICE_X0Y106_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h33ff33ffc30fc30f)
  ) CLBLL_L_X2Y106_SLICE_X0Y106_ALUT (
.I0(1'b1),
.I1(RIOB33_SING_X105Y100_IOB_X1Y100_I),
.I2(CLBLL_L_X2Y106_SLICE_X1Y106_CO6),
.I3(LIOB33_X0Y101_IOB_X0Y102_I),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y106_SLICE_X0Y106_AO5),
.O6(CLBLL_L_X2Y106_SLICE_X0Y106_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hfcf3c030fefbc832)
  ) CLBLL_L_X2Y106_SLICE_X1Y106_DLUT (
.I0(CLBLL_L_X2Y106_SLICE_X1Y106_AO6),
.I1(CLBLM_R_X13Y106_SLICE_X18Y106_AO5),
.I2(CLBLM_R_X3Y106_SLICE_X2Y106_CO6),
.I3(CLBLL_L_X2Y104_SLICE_X0Y104_BO6),
.I4(CLBLL_L_X2Y106_SLICE_X0Y106_AO6),
.I5(CLBLL_L_X2Y106_SLICE_X1Y106_BO6),
.O5(CLBLL_L_X2Y106_SLICE_X1Y106_DO5),
.O6(CLBLL_L_X2Y106_SLICE_X1Y106_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h6c6c93937d5f82a0)
  ) CLBLL_L_X2Y106_SLICE_X1Y106_CLUT (
.I0(LIOB33_X0Y101_IOB_X0Y101_I),
.I1(CLBLM_R_X3Y106_SLICE_X2Y106_CO6),
.I2(RIOB33_X105Y105_IOB_X1Y106_I),
.I3(RIOB33_SING_X105Y100_IOB_X1Y100_I),
.I4(CLBLL_L_X2Y104_SLICE_X0Y104_BO6),
.I5(CLBLL_L_X2Y106_SLICE_X1Y106_BO6),
.O5(CLBLL_L_X2Y106_SLICE_X1Y106_CO5),
.O6(CLBLL_L_X2Y106_SLICE_X1Y106_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h087f50507d0aa0a0)
  ) CLBLL_L_X2Y106_SLICE_X1Y106_BLUT (
.I0(RIOB33_X105Y105_IOB_X1Y106_I),
.I1(RIOB33_X105Y111_IOB_X1Y112_I),
.I2(LIOB33_SING_X0Y100_IOB_X0Y100_I),
.I3(LIOB33_X0Y103_IOB_X0Y103_I),
.I4(RIOB33_X105Y113_IOB_X1Y113_I),
.I5(RIOB33_SING_X105Y100_IOB_X1Y100_I),
.O5(CLBLL_L_X2Y106_SLICE_X1Y106_BO5),
.O6(CLBLL_L_X2Y106_SLICE_X1Y106_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h5f5f5f5fccdfccdf)
  ) CLBLL_L_X2Y106_SLICE_X1Y106_ALUT (
.I0(RIOB33_SING_X105Y100_IOB_X1Y100_I),
.I1(CLBLM_R_X3Y106_SLICE_X2Y106_CO6),
.I2(LIOB33_X0Y101_IOB_X0Y101_I),
.I3(CLBLL_L_X2Y106_SLICE_X1Y106_BO6),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y106_SLICE_X1Y106_AO5),
.O6(CLBLL_L_X2Y106_SLICE_X1Y106_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y107_SLICE_X0Y107_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y107_SLICE_X0Y107_DO5),
.O6(CLBLL_L_X2Y107_SLICE_X0Y107_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y107_SLICE_X0Y107_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y107_SLICE_X0Y107_CO5),
.O6(CLBLL_L_X2Y107_SLICE_X0Y107_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h2abfbf2abf2abf2a)
  ) CLBLL_L_X2Y107_SLICE_X0Y107_BLUT (
.I0(CLBLL_L_X2Y106_SLICE_X0Y106_BO6),
.I1(RIOB33_SING_X105Y100_IOB_X1Y100_I),
.I2(LIOB33_X0Y105_IOB_X0Y105_I),
.I3(CLBLL_L_X2Y104_SLICE_X1Y104_DO6),
.I4(LIOB33_X0Y103_IOB_X0Y104_I),
.I5(RIOB33_X105Y105_IOB_X1Y106_I),
.O5(CLBLL_L_X2Y107_SLICE_X0Y107_BO5),
.O6(CLBLL_L_X2Y107_SLICE_X0Y107_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h6c939393936c6c6c)
  ) CLBLL_L_X2Y107_SLICE_X0Y107_ALUT (
.I0(RIOB33_X105Y105_IOB_X1Y106_I),
.I1(CLBLL_L_X2Y106_SLICE_X0Y106_BO6),
.I2(LIOB33_X0Y103_IOB_X0Y104_I),
.I3(RIOB33_SING_X105Y100_IOB_X1Y100_I),
.I4(LIOB33_X0Y105_IOB_X0Y105_I),
.I5(CLBLL_L_X2Y104_SLICE_X1Y104_DO6),
.O5(CLBLL_L_X2Y107_SLICE_X0Y107_AO5),
.O6(CLBLL_L_X2Y107_SLICE_X0Y107_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y107_SLICE_X1Y107_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y107_SLICE_X1Y107_DO5),
.O6(CLBLL_L_X2Y107_SLICE_X1Y107_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y107_SLICE_X1Y107_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y107_SLICE_X1Y107_CO5),
.O6(CLBLL_L_X2Y107_SLICE_X1Y107_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y107_SLICE_X1Y107_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y107_SLICE_X1Y107_BO5),
.O6(CLBLL_L_X2Y107_SLICE_X1Y107_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y107_SLICE_X1Y107_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y107_SLICE_X1Y107_AO5),
.O6(CLBLL_L_X2Y107_SLICE_X1Y107_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y109_SLICE_X0Y109_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y109_SLICE_X0Y109_DO5),
.O6(CLBLL_L_X2Y109_SLICE_X0Y109_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y109_SLICE_X0Y109_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y109_SLICE_X0Y109_CO5),
.O6(CLBLL_L_X2Y109_SLICE_X0Y109_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y109_SLICE_X0Y109_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y109_SLICE_X0Y109_BO5),
.O6(CLBLL_L_X2Y109_SLICE_X0Y109_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'ha2775d7755ff55ff)
  ) CLBLL_L_X2Y109_SLICE_X0Y109_ALUT (
.I0(RIOB33_X105Y113_IOB_X1Y113_I),
.I1(RIOB33_X105Y105_IOB_X1Y106_I),
.I2(RIOB33_X105Y111_IOB_X1Y112_I),
.I3(RIOB33_SING_X105Y100_IOB_X1Y100_I),
.I4(LIOB33_SING_X0Y100_IOB_X0Y100_I),
.I5(1'b1),
.O5(CLBLL_L_X2Y109_SLICE_X0Y109_AO5),
.O6(CLBLL_L_X2Y109_SLICE_X0Y109_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y109_SLICE_X1Y109_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y109_SLICE_X1Y109_DO5),
.O6(CLBLL_L_X2Y109_SLICE_X1Y109_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y109_SLICE_X1Y109_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y109_SLICE_X1Y109_CO5),
.O6(CLBLL_L_X2Y109_SLICE_X1Y109_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y109_SLICE_X1Y109_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y109_SLICE_X1Y109_BO5),
.O6(CLBLL_L_X2Y109_SLICE_X1Y109_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y109_SLICE_X1Y109_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y109_SLICE_X1Y109_AO5),
.O6(CLBLL_L_X2Y109_SLICE_X1Y109_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y110_SLICE_X0Y110_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y110_SLICE_X0Y110_DO5),
.O6(CLBLL_L_X2Y110_SLICE_X0Y110_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y110_SLICE_X0Y110_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y110_SLICE_X0Y110_CO5),
.O6(CLBLL_L_X2Y110_SLICE_X0Y110_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y110_SLICE_X0Y110_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y110_SLICE_X0Y110_BO5),
.O6(CLBLL_L_X2Y110_SLICE_X0Y110_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hcccc0000f00f00ff)
  ) CLBLL_L_X2Y110_SLICE_X0Y110_ALUT (
.I0(1'b1),
.I1(RIOB33_X105Y111_IOB_X1Y112_I),
.I2(LIOB33_X0Y113_IOB_X0Y113_I),
.I3(CLBLL_L_X4Y108_SLICE_X4Y108_CO6),
.I4(RIOB33_SING_X105Y100_IOB_X1Y100_I),
.I5(1'b1),
.O5(CLBLL_L_X2Y110_SLICE_X0Y110_AO5),
.O6(CLBLL_L_X2Y110_SLICE_X0Y110_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y110_SLICE_X1Y110_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y110_SLICE_X1Y110_DO5),
.O6(CLBLL_L_X2Y110_SLICE_X1Y110_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y110_SLICE_X1Y110_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y110_SLICE_X1Y110_CO5),
.O6(CLBLL_L_X2Y110_SLICE_X1Y110_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y110_SLICE_X1Y110_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y110_SLICE_X1Y110_BO5),
.O6(CLBLL_L_X2Y110_SLICE_X1Y110_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y110_SLICE_X1Y110_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y110_SLICE_X1Y110_AO5),
.O6(CLBLL_L_X2Y110_SLICE_X1Y110_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'he88ec00cfccfe88e)
  ) CLBLL_L_X4Y103_SLICE_X4Y103_DLUT (
.I0(CLBLM_R_X3Y103_SLICE_X3Y103_BO6),
.I1(CLBLL_L_X4Y103_SLICE_X5Y103_AO5),
.I2(CLBLL_L_X4Y104_SLICE_X5Y104_BO6),
.I3(CLBLL_L_X4Y103_SLICE_X4Y103_AO5),
.I4(CLBLM_R_X3Y106_SLICE_X2Y106_BO5),
.I5(CLBLM_R_X3Y103_SLICE_X2Y103_BO6),
.O5(CLBLL_L_X4Y103_SLICE_X4Y103_DO5),
.O6(CLBLL_L_X4Y103_SLICE_X4Y103_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h6996c33c3cc36996)
  ) CLBLL_L_X4Y103_SLICE_X4Y103_CLUT (
.I0(CLBLM_R_X3Y103_SLICE_X3Y103_BO6),
.I1(CLBLL_L_X4Y103_SLICE_X5Y103_AO5),
.I2(CLBLL_L_X4Y104_SLICE_X5Y104_BO6),
.I3(CLBLL_L_X4Y103_SLICE_X4Y103_AO5),
.I4(CLBLM_R_X3Y106_SLICE_X2Y106_BO5),
.I5(CLBLM_R_X3Y103_SLICE_X2Y103_BO6),
.O5(CLBLL_L_X4Y103_SLICE_X4Y103_CO5),
.O6(CLBLL_L_X4Y103_SLICE_X4Y103_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hc96c696663c6c3cc)
  ) CLBLL_L_X4Y103_SLICE_X4Y103_BLUT (
.I0(LIOB33_X0Y101_IOB_X0Y101_I),
.I1(CLBLL_L_X4Y104_SLICE_X5Y104_BO6),
.I2(CLBLM_R_X3Y103_SLICE_X3Y103_BO6),
.I3(CLBLM_R_X3Y103_SLICE_X2Y103_BO6),
.I4(LIOB33_X0Y113_IOB_X0Y114_I),
.I5(LIOB33_X0Y115_IOB_X0Y116_I),
.O5(CLBLL_L_X4Y103_SLICE_X4Y103_BO5),
.O6(CLBLL_L_X4Y103_SLICE_X4Y103_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h5555ffff55ff55ff)
  ) CLBLL_L_X4Y103_SLICE_X4Y103_ALUT (
.I0(LIOB33_X0Y101_IOB_X0Y101_I),
.I1(1'b1),
.I2(1'b1),
.I3(LIOB33_X0Y115_IOB_X0Y116_I),
.I4(LIOB33_X0Y103_IOB_X0Y103_I),
.I5(1'b1),
.O5(CLBLL_L_X4Y103_SLICE_X4Y103_AO5),
.O6(CLBLL_L_X4Y103_SLICE_X4Y103_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X4Y103_SLICE_X5Y103_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y103_SLICE_X5Y103_DO5),
.O6(CLBLL_L_X4Y103_SLICE_X5Y103_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'he8fa8eafe8e88e8e)
  ) CLBLL_L_X4Y103_SLICE_X5Y103_CLUT (
.I0(CLBLL_L_X4Y103_SLICE_X5Y103_AO6),
.I1(CLBLM_R_X5Y104_SLICE_X6Y104_BO6),
.I2(CLBLM_R_X7Y104_SLICE_X8Y104_AO6),
.I3(CLBLL_L_X4Y104_SLICE_X5Y104_BO6),
.I4(CLBLM_R_X7Y103_SLICE_X8Y103_AO6),
.I5(CLBLL_L_X4Y103_SLICE_X4Y103_AO5),
.O5(CLBLL_L_X4Y103_SLICE_X5Y103_CO5),
.O6(CLBLL_L_X4Y103_SLICE_X5Y103_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h6699996666699996)
  ) CLBLL_L_X4Y103_SLICE_X5Y103_BLUT (
.I0(CLBLM_R_X7Y103_SLICE_X8Y103_AO6),
.I1(CLBLM_R_X7Y104_SLICE_X8Y104_AO6),
.I2(CLBLL_L_X4Y103_SLICE_X4Y103_AO5),
.I3(CLBLM_R_X5Y104_SLICE_X6Y104_BO6),
.I4(CLBLL_L_X4Y103_SLICE_X5Y103_AO6),
.I5(CLBLL_L_X4Y104_SLICE_X5Y104_BO6),
.O5(CLBLL_L_X4Y103_SLICE_X5Y103_BO5),
.O6(CLBLL_L_X4Y103_SLICE_X5Y103_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h3f3f3f3f5f5f5f5f)
  ) CLBLL_L_X4Y103_SLICE_X5Y103_ALUT (
.I0(LIOB33_X0Y113_IOB_X0Y114_I),
.I1(LIOB33_X0Y115_IOB_X0Y116_I),
.I2(LIOB33_X0Y101_IOB_X0Y102_I),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y103_SLICE_X5Y103_AO5),
.O6(CLBLL_L_X4Y103_SLICE_X5Y103_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h9666cccc99963c3c)
  ) CLBLL_L_X4Y104_SLICE_X4Y104_DLUT (
.I0(LIOB33_X0Y115_IOB_X0Y116_I),
.I1(CLBLL_L_X4Y104_SLICE_X5Y104_CO6),
.I2(CLBLL_L_X4Y104_SLICE_X5Y104_AO6),
.I3(LIOB33_X0Y113_IOB_X0Y114_I),
.I4(LIOB33_X0Y101_IOB_X0Y102_I),
.I5(CLBLM_R_X3Y103_SLICE_X3Y103_AO5),
.O5(CLBLL_L_X4Y104_SLICE_X4Y104_DO5),
.O6(CLBLL_L_X4Y104_SLICE_X4Y104_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h78ffffff00787878)
  ) CLBLL_L_X4Y104_SLICE_X4Y104_CLUT (
.I0(LIOB33_X0Y101_IOB_X0Y102_I),
.I1(LIOB33_X0Y113_IOB_X0Y114_I),
.I2(CLBLL_L_X4Y103_SLICE_X4Y103_BO6),
.I3(LIOB33_X0Y103_IOB_X0Y104_I),
.I4(LIOB33_X0Y103_IOB_X0Y103_I),
.I5(CLBLM_R_X3Y104_SLICE_X3Y104_DO6),
.O5(CLBLL_L_X4Y104_SLICE_X4Y104_CO5),
.O6(CLBLL_L_X4Y104_SLICE_X4Y104_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h6a959595956a6a6a)
  ) CLBLL_L_X4Y104_SLICE_X4Y104_BLUT (
.I0(CLBLL_L_X4Y103_SLICE_X4Y103_BO6),
.I1(LIOB33_X0Y103_IOB_X0Y103_I),
.I2(LIOB33_X0Y103_IOB_X0Y104_I),
.I3(LIOB33_X0Y113_IOB_X0Y114_I),
.I4(LIOB33_X0Y101_IOB_X0Y102_I),
.I5(CLBLM_R_X3Y104_SLICE_X3Y104_DO6),
.O5(CLBLL_L_X4Y104_SLICE_X4Y104_BO5),
.O6(CLBLL_L_X4Y104_SLICE_X4Y104_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h639c9c63c63939c6)
  ) CLBLL_L_X4Y104_SLICE_X4Y104_ALUT (
.I0(CLBLL_L_X2Y104_SLICE_X0Y104_AO5),
.I1(CLBLM_R_X5Y104_SLICE_X6Y104_AO6),
.I2(CLBLL_L_X4Y103_SLICE_X4Y103_CO6),
.I3(CLBLL_L_X4Y103_SLICE_X4Y103_DO6),
.I4(CLBLL_L_X4Y103_SLICE_X5Y103_BO6),
.I5(CLBLM_R_X3Y104_SLICE_X3Y104_DO6),
.O5(CLBLL_L_X4Y104_SLICE_X4Y104_AO5),
.O6(CLBLL_L_X4Y104_SLICE_X4Y104_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h718e8e718e71718e)
  ) CLBLL_L_X4Y104_SLICE_X5Y104_DLUT (
.I0(CLBLM_R_X5Y104_SLICE_X6Y104_AO6),
.I1(CLBLL_L_X4Y103_SLICE_X4Y103_DO6),
.I2(CLBLL_L_X4Y103_SLICE_X5Y103_BO6),
.I3(CLBLL_L_X4Y103_SLICE_X5Y103_CO6),
.I4(CLBLM_R_X5Y104_SLICE_X6Y104_AO5),
.I5(CLBLM_R_X7Y104_SLICE_X8Y104_CO6),
.O5(CLBLL_L_X4Y104_SLICE_X5Y104_DO5),
.O6(CLBLL_L_X4Y104_SLICE_X5Y104_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h699969996c9c3ccc)
  ) CLBLL_L_X4Y104_SLICE_X5Y104_CLUT (
.I0(CLBLM_R_X5Y104_SLICE_X6Y104_BO6),
.I1(CLBLM_R_X7Y103_SLICE_X8Y103_AO6),
.I2(LIOB33_X0Y101_IOB_X0Y101_I),
.I3(LIOB33_X0Y117_IOB_X0Y117_I),
.I4(LIOB33_X0Y115_IOB_X0Y116_I),
.I5(CLBLL_L_X4Y104_SLICE_X5Y104_BO6),
.O5(CLBLL_L_X4Y104_SLICE_X5Y104_CO5),
.O6(CLBLL_L_X4Y104_SLICE_X5Y104_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h08507da07f500aa0)
  ) CLBLL_L_X4Y104_SLICE_X5Y104_BLUT (
.I0(LIOB33_X0Y117_IOB_X0Y117_I),
.I1(RIOB33_X105Y111_IOB_X1Y112_I),
.I2(LIOB33_SING_X0Y100_IOB_X0Y100_I),
.I3(RIOB33_X105Y113_IOB_X1Y113_I),
.I4(LIOB33_X0Y115_IOB_X0Y116_I),
.I5(RIOB33_X105Y101_IOB_X1Y101_I),
.O5(CLBLL_L_X4Y104_SLICE_X5Y104_BO5),
.O6(CLBLL_L_X4Y104_SLICE_X5Y104_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hc03fc03fffff003f)
  ) CLBLL_L_X4Y104_SLICE_X5Y104_ALUT (
.I0(1'b1),
.I1(LIOB33_X0Y101_IOB_X0Y101_I),
.I2(LIOB33_X0Y115_IOB_X0Y116_I),
.I3(CLBLL_L_X4Y104_SLICE_X5Y104_BO6),
.I4(CLBLM_R_X5Y104_SLICE_X6Y104_BO6),
.I5(1'b1),
.O5(CLBLL_L_X4Y104_SLICE_X5Y104_AO5),
.O6(CLBLL_L_X4Y104_SLICE_X5Y104_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X4Y105_SLICE_X4Y105_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y105_SLICE_X4Y105_DO5),
.O6(CLBLL_L_X4Y105_SLICE_X4Y105_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X4Y105_SLICE_X4Y105_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y105_SLICE_X4Y105_CO5),
.O6(CLBLL_L_X4Y105_SLICE_X4Y105_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h69a5c30f965a3cf0)
  ) CLBLL_L_X4Y105_SLICE_X4Y105_BLUT (
.I0(LIOB33_X0Y101_IOB_X0Y102_I),
.I1(LIOB33_X0Y103_IOB_X0Y104_I),
.I2(CLBLL_L_X4Y103_SLICE_X4Y103_DO6),
.I3(LIOB33_X0Y113_IOB_X0Y114_I),
.I4(LIOB33_X0Y115_IOB_X0Y116_I),
.I5(CLBLL_L_X4Y104_SLICE_X5Y104_CO6),
.O5(CLBLL_L_X4Y105_SLICE_X4Y105_BO5),
.O6(CLBLL_L_X4Y105_SLICE_X4Y105_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h9a6a6a6a959a956a)
  ) CLBLL_L_X4Y105_SLICE_X4Y105_ALUT (
.I0(CLBLL_L_X4Y104_SLICE_X5Y104_DO6),
.I1(LIOB33_X0Y113_IOB_X0Y114_I),
.I2(LIOB33_X0Y105_IOB_X0Y105_I),
.I3(CLBLL_L_X4Y105_SLICE_X4Y105_BO6),
.I4(LIOB33_X0Y103_IOB_X0Y103_I),
.I5(CLBLL_L_X4Y104_SLICE_X4Y104_CO6),
.O5(CLBLL_L_X4Y105_SLICE_X4Y105_AO5),
.O6(CLBLL_L_X4Y105_SLICE_X4Y105_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X4Y105_SLICE_X5Y105_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y105_SLICE_X5Y105_DO5),
.O6(CLBLL_L_X4Y105_SLICE_X5Y105_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X4Y105_SLICE_X5Y105_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y105_SLICE_X5Y105_CO5),
.O6(CLBLL_L_X4Y105_SLICE_X5Y105_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfbbaf775a2205110)
  ) CLBLL_L_X4Y105_SLICE_X5Y105_BLUT (
.I0(CLBLL_L_X4Y104_SLICE_X5Y104_DO6),
.I1(CLBLL_L_X4Y105_SLICE_X4Y105_BO6),
.I2(CLBLM_R_X3Y106_SLICE_X3Y106_AO6),
.I3(CLBLL_L_X4Y104_SLICE_X4Y104_CO6),
.I4(CLBLM_R_X5Y106_SLICE_X7Y106_AO5),
.I5(CLBLM_R_X5Y105_SLICE_X7Y105_AO5),
.O5(CLBLL_L_X4Y105_SLICE_X5Y105_BO5),
.O6(CLBLL_L_X4Y105_SLICE_X5Y105_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h7fff135fb3ff20a0)
  ) CLBLL_L_X4Y105_SLICE_X5Y105_ALUT (
.I0(LIOB33_X0Y101_IOB_X0Y102_I),
.I1(LIOB33_X0Y103_IOB_X0Y104_I),
.I2(LIOB33_X0Y115_IOB_X0Y116_I),
.I3(LIOB33_X0Y113_IOB_X0Y114_I),
.I4(CLBLL_L_X4Y103_SLICE_X4Y103_DO6),
.I5(CLBLL_L_X4Y104_SLICE_X5Y104_CO6),
.O5(CLBLL_L_X4Y105_SLICE_X5Y105_AO5),
.O6(CLBLL_L_X4Y105_SLICE_X5Y105_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h7f07f770f770f770)
  ) CLBLL_L_X4Y106_SLICE_X4Y106_DLUT (
.I0(LIOB33_X0Y105_IOB_X0Y105_I),
.I1(LIOB33_X0Y103_IOB_X0Y103_I),
.I2(CLBLL_L_X4Y104_SLICE_X4Y104_DO6),
.I3(CLBLL_L_X4Y104_SLICE_X4Y104_CO6),
.I4(LIOB33_X0Y103_IOB_X0Y104_I),
.I5(LIOB33_X0Y113_IOB_X0Y114_I),
.O5(CLBLL_L_X4Y106_SLICE_X4Y106_DO5),
.O6(CLBLL_L_X4Y106_SLICE_X4Y106_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h6fcfffff060c66cc)
  ) CLBLL_L_X4Y106_SLICE_X4Y106_CLUT (
.I0(LIOB33_X0Y103_IOB_X0Y103_I),
.I1(CLBLL_L_X4Y105_SLICE_X4Y105_AO6),
.I2(RIOB33_X105Y105_IOB_X1Y106_I),
.I3(LIOB33_X0Y105_IOB_X0Y106_I),
.I4(LIOB33_X0Y107_IOB_X0Y107_I),
.I5(CLBLM_R_X3Y106_SLICE_X3Y106_DO6),
.O5(CLBLL_L_X4Y106_SLICE_X4Y106_CO5),
.O6(CLBLL_L_X4Y106_SLICE_X4Y106_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hdb4b24b42bbbd444)
  ) CLBLL_L_X4Y106_SLICE_X4Y106_BLUT (
.I0(CLBLL_L_X4Y106_SLICE_X4Y106_DO6),
.I1(CLBLM_R_X5Y105_SLICE_X6Y105_BO6),
.I2(LIOB33_X0Y105_IOB_X0Y106_I),
.I3(LIOB33_X0Y103_IOB_X0Y103_I),
.I4(CLBLM_R_X5Y105_SLICE_X6Y105_AO6),
.I5(LIOB33_X0Y113_IOB_X0Y114_I),
.O5(CLBLL_L_X4Y106_SLICE_X4Y106_BO5),
.O6(CLBLL_L_X4Y106_SLICE_X4Y106_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h69a59955965a66aa)
  ) CLBLL_L_X4Y106_SLICE_X4Y106_ALUT (
.I0(CLBLL_L_X4Y104_SLICE_X4Y104_DO6),
.I1(LIOB33_X0Y103_IOB_X0Y104_I),
.I2(LIOB33_X0Y105_IOB_X0Y105_I),
.I3(LIOB33_X0Y113_IOB_X0Y114_I),
.I4(LIOB33_X0Y103_IOB_X0Y103_I),
.I5(CLBLL_L_X4Y104_SLICE_X4Y104_CO6),
.O5(CLBLL_L_X4Y106_SLICE_X4Y106_AO5),
.O6(CLBLL_L_X4Y106_SLICE_X4Y106_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h6cffffff006c6c6c)
  ) CLBLL_L_X4Y106_SLICE_X5Y106_DLUT (
.I0(LIOB33_X0Y113_IOB_X0Y114_I),
.I1(CLBLM_R_X5Y105_SLICE_X6Y105_CO6),
.I2(LIOB33_X0Y107_IOB_X0Y107_I),
.I3(LIOB33_X0Y107_IOB_X0Y108_I),
.I4(LIOB33_X0Y103_IOB_X0Y103_I),
.I5(CLBLL_L_X4Y106_SLICE_X5Y106_BO6),
.O5(CLBLL_L_X4Y106_SLICE_X5Y106_DO5),
.O6(CLBLL_L_X4Y106_SLICE_X5Y106_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h6c939393936c6c6c)
  ) CLBLL_L_X4Y106_SLICE_X5Y106_CLUT (
.I0(LIOB33_X0Y107_IOB_X0Y107_I),
.I1(CLBLM_R_X5Y105_SLICE_X6Y105_CO6),
.I2(LIOB33_X0Y113_IOB_X0Y114_I),
.I3(LIOB33_X0Y107_IOB_X0Y108_I),
.I4(LIOB33_X0Y103_IOB_X0Y103_I),
.I5(CLBLL_L_X4Y106_SLICE_X5Y106_BO6),
.O5(CLBLL_L_X4Y106_SLICE_X5Y106_CO5),
.O6(CLBLL_L_X4Y106_SLICE_X5Y106_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h48c0defcdefcdefc)
  ) CLBLL_L_X4Y106_SLICE_X5Y106_BLUT (
.I0(LIOB33_X0Y105_IOB_X0Y106_I),
.I1(CLBLL_L_X4Y105_SLICE_X5Y105_BO6),
.I2(CLBLM_R_X5Y105_SLICE_X6Y105_AO6),
.I3(LIOB33_X0Y113_IOB_X0Y114_I),
.I4(LIOB33_X0Y107_IOB_X0Y107_I),
.I5(LIOB33_X0Y103_IOB_X0Y103_I),
.O5(CLBLL_L_X4Y106_SLICE_X5Y106_BO5),
.O6(CLBLL_L_X4Y106_SLICE_X5Y106_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h7887877887788778)
  ) CLBLL_L_X4Y106_SLICE_X5Y106_ALUT (
.I0(LIOB33_X0Y105_IOB_X0Y106_I),
.I1(LIOB33_X0Y113_IOB_X0Y114_I),
.I2(CLBLM_R_X5Y105_SLICE_X6Y105_AO6),
.I3(CLBLL_L_X4Y105_SLICE_X5Y105_BO6),
.I4(LIOB33_X0Y107_IOB_X0Y107_I),
.I5(LIOB33_X0Y103_IOB_X0Y103_I),
.O5(CLBLL_L_X4Y106_SLICE_X5Y106_AO5),
.O6(CLBLL_L_X4Y106_SLICE_X5Y106_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X4Y107_SLICE_X4Y107_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y107_SLICE_X4Y107_DO5),
.O6(CLBLL_L_X4Y107_SLICE_X4Y107_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h4dddcfff8eee0ccc)
  ) CLBLL_L_X4Y107_SLICE_X4Y107_CLUT (
.I0(LIOB33_X0Y107_IOB_X0Y107_I),
.I1(CLBLL_L_X4Y106_SLICE_X4Y106_CO6),
.I2(RIOB33_X105Y105_IOB_X1Y106_I),
.I3(LIOB33_X0Y107_IOB_X0Y108_I),
.I4(LIOB33_X0Y103_IOB_X0Y103_I),
.I5(CLBLL_L_X4Y106_SLICE_X4Y106_BO6),
.O5(CLBLL_L_X4Y107_SLICE_X4Y107_CO5),
.O6(CLBLL_L_X4Y107_SLICE_X4Y107_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h454d5d5f4fcfdfff)
  ) CLBLL_L_X4Y107_SLICE_X4Y107_BLUT (
.I0(RIOB33_SING_X105Y100_IOB_X1Y100_I),
.I1(CLBLM_R_X3Y107_SLICE_X3Y107_CO6),
.I2(CLBLL_L_X4Y107_SLICE_X5Y107_CO6),
.I3(LIOB33_X0Y109_IOB_X0Y109_I),
.I4(CLBLL_L_X4Y107_SLICE_X4Y107_AO6),
.I5(LIOB33_X0Y109_IOB_X0Y110_I),
.O5(CLBLL_L_X4Y107_SLICE_X4Y107_BO5),
.O6(CLBLL_L_X4Y107_SLICE_X4Y107_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h6c93936c93936c6c)
  ) CLBLL_L_X4Y107_SLICE_X4Y107_ALUT (
.I0(LIOB33_X0Y103_IOB_X0Y103_I),
.I1(CLBLL_L_X4Y106_SLICE_X4Y106_CO6),
.I2(LIOB33_X0Y107_IOB_X0Y107_I),
.I3(RIOB33_X105Y105_IOB_X1Y106_I),
.I4(CLBLL_L_X4Y106_SLICE_X4Y106_BO6),
.I5(LIOB33_X0Y107_IOB_X0Y108_I),
.O5(CLBLL_L_X4Y107_SLICE_X4Y107_AO5),
.O6(CLBLL_L_X4Y107_SLICE_X4Y107_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hf990f9f99090f990)
  ) CLBLL_L_X4Y107_SLICE_X5Y107_DLUT (
.I0(CLBLL_L_X4Y107_SLICE_X5Y107_AO6),
.I1(CLBLM_R_X5Y106_SLICE_X7Y106_CO6),
.I2(CLBLM_R_X3Y107_SLICE_X3Y107_AO5),
.I3(CLBLL_L_X4Y107_SLICE_X5Y107_AO5),
.I4(CLBLL_L_X4Y106_SLICE_X5Y106_AO6),
.I5(CLBLL_L_X4Y106_SLICE_X4Y106_CO6),
.O5(CLBLL_L_X4Y107_SLICE_X5Y107_DO5),
.O6(CLBLL_L_X4Y107_SLICE_X5Y107_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h6996696996966996)
  ) CLBLL_L_X4Y107_SLICE_X5Y107_CLUT (
.I0(CLBLL_L_X4Y107_SLICE_X5Y107_AO6),
.I1(CLBLM_R_X5Y106_SLICE_X7Y106_CO6),
.I2(CLBLM_R_X3Y107_SLICE_X3Y107_AO5),
.I3(CLBLL_L_X4Y107_SLICE_X5Y107_AO5),
.I4(CLBLL_L_X4Y106_SLICE_X5Y106_AO6),
.I5(CLBLL_L_X4Y106_SLICE_X4Y106_CO6),
.O5(CLBLL_L_X4Y107_SLICE_X5Y107_CO5),
.O6(CLBLL_L_X4Y107_SLICE_X5Y107_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h9c936c9c6c936c6c)
  ) CLBLL_L_X4Y107_SLICE_X5Y107_BLUT (
.I0(LIOB33_X0Y103_IOB_X0Y103_I),
.I1(CLBLM_R_X5Y106_SLICE_X7Y106_CO6),
.I2(LIOB33_X0Y107_IOB_X0Y108_I),
.I3(CLBLL_L_X4Y106_SLICE_X4Y106_CO6),
.I4(CLBLL_L_X4Y106_SLICE_X5Y106_AO6),
.I5(RIOB33_X105Y105_IOB_X1Y106_I),
.O5(CLBLL_L_X4Y107_SLICE_X5Y107_BO5),
.O6(CLBLL_L_X4Y107_SLICE_X5Y107_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h55ff55ff33ff33ff)
  ) CLBLL_L_X4Y107_SLICE_X5Y107_ALUT (
.I0(LIOB33_X0Y103_IOB_X0Y103_I),
.I1(RIOB33_X105Y105_IOB_X1Y106_I),
.I2(1'b1),
.I3(LIOB33_X0Y107_IOB_X0Y108_I),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y107_SLICE_X5Y107_AO5),
.O6(CLBLL_L_X4Y107_SLICE_X5Y107_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h4dd4cffcd44dfccf)
  ) CLBLL_L_X4Y108_SLICE_X4Y108_DLUT (
.I0(RIOB33_SING_X105Y100_IOB_X1Y100_I),
.I1(CLBLM_R_X5Y108_SLICE_X6Y108_CO6),
.I2(CLBLM_R_X7Y107_SLICE_X8Y107_AO6),
.I3(CLBLL_L_X4Y108_SLICE_X4Y108_AO5),
.I4(LIOB33_X0Y113_IOB_X0Y113_I),
.I5(CLBLM_R_X5Y108_SLICE_X6Y108_BO6),
.O5(CLBLL_L_X4Y108_SLICE_X4Y108_DO5),
.O6(CLBLL_L_X4Y108_SLICE_X4Y108_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h69965aa5a55a6996)
  ) CLBLL_L_X4Y108_SLICE_X4Y108_CLUT (
.I0(CLBLM_R_X5Y108_SLICE_X6Y108_BO6),
.I1(CLBLM_R_X5Y110_SLICE_X7Y110_AO6),
.I2(CLBLM_R_X7Y107_SLICE_X8Y107_AO6),
.I3(CLBLL_L_X4Y108_SLICE_X4Y108_AO5),
.I4(CLBLM_R_X5Y108_SLICE_X6Y108_AO6),
.I5(CLBLL_L_X4Y108_SLICE_X4Y108_BO6),
.O5(CLBLL_L_X4Y108_SLICE_X4Y108_CO5),
.O6(CLBLL_L_X4Y108_SLICE_X4Y108_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h7f15d540ff3fffc0)
  ) CLBLL_L_X4Y108_SLICE_X4Y108_BLUT (
.I0(LIOB33_X0Y111_IOB_X0Y111_I),
.I1(LIOB33_X0Y109_IOB_X0Y110_I),
.I2(RIOB33_X105Y105_IOB_X1Y106_I),
.I3(CLBLL_L_X4Y107_SLICE_X4Y107_BO6),
.I4(CLBLM_R_X5Y107_SLICE_X6Y107_AO6),
.I5(RIOB33_SING_X105Y100_IOB_X1Y100_I),
.O5(CLBLL_L_X4Y108_SLICE_X4Y108_BO5),
.O6(CLBLL_L_X4Y108_SLICE_X4Y108_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h5aa5aa553f3f3f3f)
  ) CLBLL_L_X4Y108_SLICE_X4Y108_ALUT (
.I0(CLBLM_R_X5Y108_SLICE_X6Y108_AO6),
.I1(RIOB33_X105Y105_IOB_X1Y106_I),
.I2(LIOB33_X0Y111_IOB_X0Y112_I),
.I3(CLBLL_L_X4Y108_SLICE_X4Y108_BO6),
.I4(RIOB33_SING_X105Y100_IOB_X1Y100_I),
.I5(1'b1),
.O5(CLBLL_L_X4Y108_SLICE_X4Y108_AO5),
.O6(CLBLL_L_X4Y108_SLICE_X4Y108_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hac536c936f905fa0)
  ) CLBLL_L_X4Y108_SLICE_X5Y108_DLUT (
.I0(LIOB33_X0Y113_IOB_X0Y114_I),
.I1(CLBLM_R_X7Y107_SLICE_X8Y107_CO6),
.I2(LIOB33_X0Y111_IOB_X0Y112_I),
.I3(CLBLM_R_X7Y108_SLICE_X8Y108_CO6),
.I4(LIOB33_X0Y103_IOB_X0Y103_I),
.I5(CLBLM_R_X5Y108_SLICE_X7Y108_CO6),
.O5(CLBLL_L_X4Y108_SLICE_X5Y108_DO5),
.O6(CLBLL_L_X4Y108_SLICE_X5Y108_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h054ddddd4d5fffff)
  ) CLBLL_L_X4Y108_SLICE_X5Y108_CLUT (
.I0(CLBLM_R_X7Y108_SLICE_X8Y108_BO6),
.I1(CLBLM_R_X7Y107_SLICE_X8Y107_CO6),
.I2(LIOB33_X0Y113_IOB_X0Y113_I),
.I3(LIOB33_X0Y111_IOB_X0Y112_I),
.I4(LIOB33_X0Y103_IOB_X0Y103_I),
.I5(CLBLM_R_X5Y108_SLICE_X7Y108_CO6),
.O5(CLBLL_L_X4Y108_SLICE_X5Y108_CO5),
.O6(CLBLL_L_X4Y108_SLICE_X5Y108_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hac6f53906c5f93a0)
  ) CLBLL_L_X4Y108_SLICE_X5Y108_BLUT (
.I0(LIOB33_X0Y113_IOB_X0Y113_I),
.I1(CLBLM_R_X7Y107_SLICE_X8Y107_CO6),
.I2(LIOB33_X0Y103_IOB_X0Y103_I),
.I3(CLBLM_R_X5Y108_SLICE_X7Y108_CO6),
.I4(CLBLM_R_X7Y108_SLICE_X8Y108_BO6),
.I5(LIOB33_X0Y111_IOB_X0Y112_I),
.O5(CLBLL_L_X4Y108_SLICE_X5Y108_BO5),
.O6(CLBLL_L_X4Y108_SLICE_X5Y108_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hb7483fc0d12e956a)
  ) CLBLL_L_X4Y108_SLICE_X5Y108_ALUT (
.I0(CLBLM_R_X7Y107_SLICE_X8Y107_AO6),
.I1(LIOB33_X0Y111_IOB_X0Y112_I),
.I2(LIOB33_X0Y103_IOB_X0Y103_I),
.I3(CLBLM_R_X7Y107_SLICE_X8Y107_BO6),
.I4(RIOB33_X105Y105_IOB_X1Y106_I),
.I5(CLBLM_R_X5Y108_SLICE_X6Y108_BO6),
.O5(CLBLL_L_X4Y108_SLICE_X5Y108_AO5),
.O6(CLBLL_L_X4Y108_SLICE_X5Y108_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'he41b6c937d825fa0)
  ) CLBLL_L_X4Y109_SLICE_X4Y109_DLUT (
.I0(RIOB33_X105Y105_IOB_X1Y106_I),
.I1(CLBLM_R_X5Y108_SLICE_X6Y108_BO6),
.I2(LIOB33_X0Y113_IOB_X0Y113_I),
.I3(CLBLM_R_X7Y107_SLICE_X8Y107_DO6),
.I4(LIOB33_X0Y111_IOB_X0Y112_I),
.I5(CLBLM_R_X7Y107_SLICE_X8Y107_AO6),
.O5(CLBLL_L_X4Y109_SLICE_X4Y109_DO5),
.O6(CLBLL_L_X4Y109_SLICE_X4Y109_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h445f4cdf5ddf5fff)
  ) CLBLL_L_X4Y109_SLICE_X4Y109_CLUT (
.I0(RIOB33_X105Y105_IOB_X1Y106_I),
.I1(CLBLM_R_X5Y108_SLICE_X6Y108_BO6),
.I2(LIOB33_X0Y113_IOB_X0Y113_I),
.I3(CLBLM_R_X7Y107_SLICE_X8Y107_DO6),
.I4(LIOB33_X0Y111_IOB_X0Y112_I),
.I5(CLBLM_R_X7Y107_SLICE_X8Y107_AO6),
.O5(CLBLL_L_X4Y109_SLICE_X4Y109_CO5),
.O6(CLBLL_L_X4Y109_SLICE_X4Y109_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hc369693c3c9696c3)
  ) CLBLL_L_X4Y109_SLICE_X4Y109_BLUT (
.I0(CLBLL_L_X4Y109_SLICE_X4Y109_DO6),
.I1(CLBLL_L_X4Y109_SLICE_X4Y109_AO5),
.I2(CLBLL_L_X4Y108_SLICE_X5Y108_BO6),
.I3(CLBLL_L_X4Y108_SLICE_X4Y108_DO6),
.I4(CLBLL_L_X4Y109_SLICE_X4Y109_AO6),
.I5(CLBLL_L_X4Y109_SLICE_X4Y109_CO6),
.O5(CLBLL_L_X4Y109_SLICE_X4Y109_BO5),
.O6(CLBLL_L_X4Y109_SLICE_X4Y109_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h33ff33ff3f3f3f3f)
  ) CLBLL_L_X4Y109_SLICE_X4Y109_ALUT (
.I0(1'b1),
.I1(LIOB33_X0Y115_IOB_X0Y115_I),
.I2(RIOB33_X105Y105_IOB_X1Y106_I),
.I3(RIOB33_SING_X105Y100_IOB_X1Y100_I),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y109_SLICE_X4Y109_AO5),
.O6(CLBLL_L_X4Y109_SLICE_X4Y109_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h4dddcfffd444fccc)
  ) CLBLL_L_X4Y109_SLICE_X5Y109_DLUT (
.I0(LIOB33_X0Y115_IOB_X0Y115_I),
.I1(CLBLL_L_X4Y108_SLICE_X5Y108_CO6),
.I2(LIOB33_X0Y113_IOB_X0Y113_I),
.I3(LIOB33_X0Y113_IOB_X0Y114_I),
.I4(LIOB33_X0Y103_IOB_X0Y103_I),
.I5(CLBLM_R_X5Y109_SLICE_X7Y109_AO6),
.O5(CLBLL_L_X4Y109_SLICE_X5Y109_DO5),
.O6(CLBLL_L_X4Y109_SLICE_X5Y109_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h4dcfd4fcddff44cc)
  ) CLBLL_L_X4Y109_SLICE_X5Y109_CLUT (
.I0(LIOB33_X0Y115_IOB_X0Y115_I),
.I1(CLBLL_L_X4Y109_SLICE_X4Y109_CO6),
.I2(LIOB33_X0Y113_IOB_X0Y113_I),
.I3(RIOB33_X105Y105_IOB_X1Y106_I),
.I4(CLBLL_L_X4Y108_SLICE_X5Y108_DO6),
.I5(LIOB33_X0Y103_IOB_X0Y103_I),
.O5(CLBLL_L_X4Y109_SLICE_X5Y109_CO5),
.O6(CLBLL_L_X4Y109_SLICE_X5Y109_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h6c939393936c6c6c)
  ) CLBLL_L_X4Y109_SLICE_X5Y109_BLUT (
.I0(LIOB33_X0Y113_IOB_X0Y113_I),
.I1(CLBLM_R_X5Y109_SLICE_X7Y109_AO6),
.I2(LIOB33_X0Y113_IOB_X0Y114_I),
.I3(LIOB33_X0Y103_IOB_X0Y103_I),
.I4(LIOB33_X0Y115_IOB_X0Y115_I),
.I5(CLBLL_L_X4Y108_SLICE_X5Y108_CO6),
.O5(CLBLL_L_X4Y109_SLICE_X5Y109_BO5),
.O6(CLBLL_L_X4Y109_SLICE_X5Y109_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h93939393aa5500ff)
  ) CLBLL_L_X4Y109_SLICE_X5Y109_ALUT (
.I0(LIOB33_X0Y113_IOB_X0Y113_I),
.I1(CLBLM_R_X5Y109_SLICE_X7Y109_AO6),
.I2(LIOB33_X0Y113_IOB_X0Y114_I),
.I3(CLBLM_R_X5Y110_SLICE_X7Y110_CO6),
.I4(RIOB33_X105Y101_IOB_X1Y102_I),
.I5(1'b1),
.O5(CLBLL_L_X4Y109_SLICE_X5Y109_AO5),
.O6(CLBLL_L_X4Y109_SLICE_X5Y109_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X4Y110_SLICE_X4Y110_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y110_SLICE_X4Y110_DO5),
.O6(CLBLL_L_X4Y110_SLICE_X4Y110_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X4Y110_SLICE_X4Y110_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y110_SLICE_X4Y110_CO5),
.O6(CLBLL_L_X4Y110_SLICE_X4Y110_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h70f780f8f7f7f8f8)
  ) CLBLL_L_X4Y110_SLICE_X4Y110_BLUT (
.I0(LIOB33_X0Y113_IOB_X0Y113_I),
.I1(LIOB33_X0Y115_IOB_X0Y116_I),
.I2(CLBLM_R_X5Y109_SLICE_X7Y109_BO6),
.I3(LIOB33_X0Y113_IOB_X0Y114_I),
.I4(CLBLM_R_X7Y110_SLICE_X8Y110_AO6),
.I5(LIOB33_X0Y115_IOB_X0Y115_I),
.O5(CLBLL_L_X4Y110_SLICE_X4Y110_BO5),
.O6(CLBLL_L_X4Y110_SLICE_X4Y110_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h6996c33c96963c3c)
  ) CLBLL_L_X4Y110_SLICE_X4Y110_ALUT (
.I0(LIOB33_X0Y113_IOB_X0Y113_I),
.I1(CLBLM_R_X7Y110_SLICE_X8Y110_AO6),
.I2(CLBLM_R_X5Y109_SLICE_X7Y109_BO6),
.I3(LIOB33_X0Y113_IOB_X0Y114_I),
.I4(LIOB33_X0Y115_IOB_X0Y116_I),
.I5(LIOB33_X0Y115_IOB_X0Y115_I),
.O5(CLBLL_L_X4Y110_SLICE_X4Y110_AO5),
.O6(CLBLL_L_X4Y110_SLICE_X4Y110_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffdf0dffff4f04)
  ) CLBLL_L_X4Y110_SLICE_X5Y110_DLUT (
.I0(CLBLL_L_X4Y109_SLICE_X5Y109_CO6),
.I1(CLBLL_L_X4Y109_SLICE_X5Y109_BO6),
.I2(CLBLL_L_X4Y109_SLICE_X5Y109_DO6),
.I3(CLBLL_L_X4Y110_SLICE_X4Y110_AO6),
.I4(CLBLL_L_X4Y112_SLICE_X4Y112_DO6),
.I5(CLBLL_L_X4Y109_SLICE_X4Y109_BO6),
.O5(CLBLL_L_X4Y110_SLICE_X5Y110_DO5),
.O6(CLBLL_L_X4Y110_SLICE_X5Y110_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h4d04ffdf0400df4d)
  ) CLBLL_L_X4Y110_SLICE_X5Y110_CLUT (
.I0(CLBLL_L_X4Y109_SLICE_X5Y109_AO6),
.I1(CLBLL_L_X4Y108_SLICE_X5Y108_CO6),
.I2(CLBLL_L_X4Y109_SLICE_X4Y109_BO6),
.I3(CLBLL_L_X4Y109_SLICE_X5Y109_CO6),
.I4(CLBLL_L_X4Y110_SLICE_X4Y110_AO6),
.I5(CLBLL_L_X4Y110_SLICE_X5Y110_BO6),
.O5(CLBLL_L_X4Y110_SLICE_X5Y110_CO5),
.O6(CLBLL_L_X4Y110_SLICE_X5Y110_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h5555ffff77777777)
  ) CLBLL_L_X4Y110_SLICE_X5Y110_BLUT (
.I0(LIOB33_X0Y115_IOB_X0Y115_I),
.I1(LIOB33_X0Y113_IOB_X0Y114_I),
.I2(1'b1),
.I3(1'b1),
.I4(LIOB33_X0Y103_IOB_X0Y103_I),
.I5(1'b1),
.O5(CLBLL_L_X4Y110_SLICE_X5Y110_BO5),
.O6(CLBLL_L_X4Y110_SLICE_X5Y110_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h3cc33cc36a5695a9)
  ) CLBLL_L_X4Y110_SLICE_X5Y110_ALUT (
.I0(CLBLL_L_X4Y109_SLICE_X5Y109_DO6),
.I1(CLBLL_L_X4Y109_SLICE_X4Y109_BO6),
.I2(CLBLL_L_X4Y109_SLICE_X5Y109_BO6),
.I3(CLBLL_L_X4Y109_SLICE_X5Y109_CO6),
.I4(CLBLL_L_X4Y110_SLICE_X4Y110_AO6),
.I5(1'b1),
.O5(CLBLL_L_X4Y110_SLICE_X5Y110_AO5),
.O6(CLBLL_L_X4Y110_SLICE_X5Y110_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hd4404000fffdfdd4)
  ) CLBLL_L_X4Y111_SLICE_X4Y111_DLUT (
.I0(CLBLM_L_X8Y112_SLICE_X10Y112_DO6),
.I1(CLBLL_L_X4Y110_SLICE_X5Y110_CO6),
.I2(CLBLM_R_X7Y112_SLICE_X9Y112_BO6),
.I3(CLBLL_L_X4Y114_SLICE_X4Y114_AO6),
.I4(CLBLL_L_X4Y110_SLICE_X4Y110_BO6),
.I5(CLBLL_L_X4Y112_SLICE_X4Y112_BO6),
.O5(CLBLL_L_X4Y111_SLICE_X4Y111_DO5),
.O6(CLBLL_L_X4Y111_SLICE_X4Y111_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h7ddd1444ffff3ccc)
  ) CLBLL_L_X4Y111_SLICE_X4Y111_CLUT (
.I0(LIOB33_X0Y115_IOB_X0Y115_I),
.I1(CLBLM_R_X7Y112_SLICE_X9Y112_AO6),
.I2(LIOB33_X0Y117_IOB_X0Y117_I),
.I3(LIOB33_X0Y113_IOB_X0Y113_I),
.I4(CLBLM_R_X7Y112_SLICE_X9Y112_BO6),
.I5(LIOB33_X0Y115_IOB_X0Y116_I),
.O5(CLBLL_L_X4Y111_SLICE_X4Y111_CO5),
.O6(CLBLL_L_X4Y111_SLICE_X4Y111_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h69969966a55a55aa)
  ) CLBLL_L_X4Y111_SLICE_X4Y111_BLUT (
.I0(CLBLM_R_X7Y112_SLICE_X9Y112_BO6),
.I1(LIOB33_X0Y117_IOB_X0Y117_I),
.I2(LIOB33_X0Y115_IOB_X0Y116_I),
.I3(CLBLM_R_X7Y112_SLICE_X9Y112_AO6),
.I4(LIOB33_X0Y115_IOB_X0Y115_I),
.I5(LIOB33_X0Y113_IOB_X0Y113_I),
.O5(CLBLL_L_X4Y111_SLICE_X4Y111_BO5),
.O6(CLBLL_L_X4Y111_SLICE_X4Y111_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h96969696d42b2bd4)
  ) CLBLL_L_X4Y111_SLICE_X4Y111_ALUT (
.I0(CLBLL_L_X4Y111_SLICE_X4Y111_BO6),
.I1(CLBLL_L_X4Y110_SLICE_X4Y110_BO6),
.I2(CLBLL_L_X4Y110_SLICE_X5Y110_CO6),
.I3(CLBLL_L_X4Y112_SLICE_X4Y112_BO6),
.I4(CLBLL_L_X4Y111_SLICE_X4Y111_CO6),
.I5(1'b1),
.O5(CLBLL_L_X4Y111_SLICE_X4Y111_AO5),
.O6(CLBLL_L_X4Y111_SLICE_X4Y111_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hd450d4d4f5d4f5f5)
  ) CLBLL_L_X4Y111_SLICE_X5Y111_DLUT (
.I0(CLBLM_R_X5Y111_SLICE_X6Y111_AO6),
.I1(CLBLL_L_X4Y111_SLICE_X4Y111_CO6),
.I2(CLBLL_L_X4Y112_SLICE_X4Y112_CO6),
.I3(CLBLL_L_X4Y111_SLICE_X5Y111_CO6),
.I4(CLBLL_L_X4Y110_SLICE_X5Y110_DO6),
.I5(CLBLL_L_X4Y112_SLICE_X4Y112_BO6),
.O5(CLBLL_L_X4Y111_SLICE_X5Y111_DO5),
.O6(CLBLL_L_X4Y111_SLICE_X5Y111_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h6699060906090000)
  ) CLBLL_L_X4Y111_SLICE_X5Y111_CLUT (
.I0(CLBLM_L_X8Y112_SLICE_X10Y112_DO6),
.I1(CLBLL_L_X4Y114_SLICE_X4Y114_AO6),
.I2(CLBLM_R_X7Y112_SLICE_X9Y112_DO6),
.I3(CLBLM_R_X7Y112_SLICE_X9Y112_BO6),
.I4(CLBLL_L_X4Y110_SLICE_X5Y110_BO5),
.I5(CLBLM_R_X5Y109_SLICE_X7Y109_BO6),
.O5(CLBLL_L_X4Y111_SLICE_X5Y111_CO5),
.O6(CLBLL_L_X4Y111_SLICE_X5Y111_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h8eff08ef08ef008e)
  ) CLBLL_L_X4Y111_SLICE_X5Y111_BLUT (
.I0(CLBLM_R_X7Y112_SLICE_X8Y112_CO6),
.I1(CLBLL_L_X4Y111_SLICE_X4Y111_DO6),
.I2(CLBLL_L_X4Y109_SLICE_X5Y109_AO5),
.I3(CLBLM_R_X5Y112_SLICE_X6Y112_BO6),
.I4(CLBLL_L_X4Y112_SLICE_X4Y112_CO6),
.I5(CLBLL_L_X4Y111_SLICE_X5Y111_AO5),
.O5(CLBLL_L_X4Y111_SLICE_X5Y111_BO5),
.O6(CLBLL_L_X4Y111_SLICE_X5Y111_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0aafaaff0f0fffff)
  ) CLBLL_L_X4Y111_SLICE_X5Y111_ALUT (
.I0(CLBLM_R_X7Y112_SLICE_X8Y112_CO6),
.I1(1'b1),
.I2(RIOB33_X105Y101_IOB_X1Y101_I),
.I3(CLBLL_L_X4Y109_SLICE_X5Y109_AO5),
.I4(LIOB33_X0Y115_IOB_X0Y115_I),
.I5(1'b1),
.O5(CLBLL_L_X4Y111_SLICE_X5Y111_AO5),
.O6(CLBLL_L_X4Y111_SLICE_X5Y111_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h599aa665a665599a)
  ) CLBLL_L_X4Y112_SLICE_X4Y112_DLUT (
.I0(CLBLL_L_X4Y114_SLICE_X4Y114_AO6),
.I1(CLBLM_R_X7Y112_SLICE_X9Y112_DO6),
.I2(CLBLL_L_X4Y110_SLICE_X5Y110_BO5),
.I3(CLBLM_R_X5Y109_SLICE_X7Y109_BO6),
.I4(CLBLM_L_X8Y112_SLICE_X10Y112_DO6),
.I5(CLBLM_R_X7Y112_SLICE_X9Y112_BO6),
.O5(CLBLL_L_X4Y112_SLICE_X4Y112_DO5),
.O6(CLBLL_L_X4Y112_SLICE_X4Y112_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h71f5d450f3fffcf0)
  ) CLBLL_L_X4Y112_SLICE_X4Y112_CLUT (
.I0(LIOB33_X0Y115_IOB_X0Y115_I),
.I1(RIOB33_X105Y101_IOB_X1Y101_I),
.I2(CLBLM_R_X7Y112_SLICE_X9Y112_CO6),
.I3(LIOB33_X0Y113_IOB_X0Y113_I),
.I4(CLBLM_R_X7Y112_SLICE_X8Y112_AO5),
.I5(LIOB33_X0Y117_IOB_X0Y117_I),
.O5(CLBLL_L_X4Y112_SLICE_X4Y112_CO5),
.O6(CLBLL_L_X4Y112_SLICE_X4Y112_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h6996a55a996655aa)
  ) CLBLL_L_X4Y112_SLICE_X4Y112_BLUT (
.I0(CLBLM_R_X7Y112_SLICE_X8Y112_AO5),
.I1(LIOB33_X0Y117_IOB_X0Y117_I),
.I2(RIOB33_X105Y101_IOB_X1Y101_I),
.I3(CLBLM_R_X7Y112_SLICE_X9Y112_CO6),
.I4(LIOB33_X0Y115_IOB_X0Y115_I),
.I5(LIOB33_X0Y113_IOB_X0Y113_I),
.O5(CLBLL_L_X4Y112_SLICE_X4Y112_BO5),
.O6(CLBLL_L_X4Y112_SLICE_X4Y112_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h999966668778e11e)
  ) CLBLL_L_X4Y112_SLICE_X4Y112_ALUT (
.I0(CLBLL_L_X4Y111_SLICE_X4Y111_DO6),
.I1(CLBLL_L_X4Y112_SLICE_X4Y112_CO6),
.I2(CLBLM_R_X5Y112_SLICE_X6Y112_BO6),
.I3(CLBLL_L_X4Y111_SLICE_X5Y111_AO6),
.I4(CLBLM_R_X5Y111_SLICE_X6Y111_AO6),
.I5(1'b1),
.O5(CLBLL_L_X4Y112_SLICE_X4Y112_AO5),
.O6(CLBLL_L_X4Y112_SLICE_X4Y112_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h9999999966666666)
  ) CLBLL_L_X4Y112_SLICE_X5Y112_DLUT (
.I0(CLBLL_L_X4Y112_SLICE_X5Y112_AO6),
.I1(CLBLL_L_X4Y113_SLICE_X5Y113_AO6),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(CLBLL_L_X4Y111_SLICE_X5Y111_BO6),
.O5(CLBLL_L_X4Y112_SLICE_X5Y112_DO5),
.O6(CLBLL_L_X4Y112_SLICE_X5Y112_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000b2bb000022b2)
  ) CLBLL_L_X4Y112_SLICE_X5Y112_CLUT (
.I0(CLBLL_L_X4Y112_SLICE_X5Y112_AO6),
.I1(CLBLL_L_X4Y113_SLICE_X5Y113_AO6),
.I2(CLBLL_L_X4Y111_SLICE_X5Y111_DO6),
.I3(CLBLM_R_X5Y112_SLICE_X6Y112_BO6),
.I4(CLBLL_L_X4Y113_SLICE_X5Y113_BO6),
.I5(CLBLL_L_X4Y111_SLICE_X5Y111_AO6),
.O5(CLBLL_L_X4Y112_SLICE_X5Y112_CO5),
.O6(CLBLL_L_X4Y112_SLICE_X5Y112_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hbf3b3b233b232302)
  ) CLBLL_L_X4Y112_SLICE_X5Y112_BLUT (
.I0(CLBLM_R_X5Y110_SLICE_X7Y110_DO6),
.I1(CLBLL_L_X4Y113_SLICE_X5Y113_AO6),
.I2(CLBLM_R_X5Y112_SLICE_X6Y112_AO6),
.I3(CLBLM_R_X5Y112_SLICE_X7Y112_AO5),
.I4(CLBLL_L_X4Y111_SLICE_X5Y111_AO6),
.I5(CLBLL_L_X4Y111_SLICE_X5Y111_DO6),
.O5(CLBLL_L_X4Y112_SLICE_X5Y112_BO5),
.O6(CLBLL_L_X4Y112_SLICE_X5Y112_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h2abfbf2abfbf2a2a)
  ) CLBLL_L_X4Y112_SLICE_X5Y112_ALUT (
.I0(CLBLM_R_X5Y110_SLICE_X7Y110_DO6),
.I1(LIOB33_X0Y115_IOB_X0Y115_I),
.I2(RIOB33_X105Y101_IOB_X1Y102_I),
.I3(RIOB33_X105Y103_IOB_X1Y103_I),
.I4(CLBLM_R_X5Y111_SLICE_X6Y111_DO6),
.I5(LIOB33_X0Y113_IOB_X0Y113_I),
.O5(CLBLL_L_X4Y112_SLICE_X5Y112_AO5),
.O6(CLBLL_L_X4Y112_SLICE_X5Y112_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h55555555ffffffff)
  ) CLBLL_L_X4Y113_SLICE_X4Y113_DLUT (
.I0(LIOB33_X0Y115_IOB_X0Y115_I),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(RIOB33_X105Y107_IOB_X1Y108_I),
.O5(CLBLL_L_X4Y113_SLICE_X4Y113_DO5),
.O6(CLBLL_L_X4Y113_SLICE_X4Y113_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hef000e00ffefff0e)
  ) CLBLL_L_X4Y113_SLICE_X4Y113_CLUT (
.I0(CLBLL_L_X4Y112_SLICE_X5Y112_CO6),
.I1(CLBLL_L_X4Y113_SLICE_X5Y113_CO6),
.I2(CLBLM_R_X7Y114_SLICE_X8Y114_CO6),
.I3(CLBLM_R_X7Y114_SLICE_X8Y114_DO6),
.I4(CLBLL_L_X4Y114_SLICE_X4Y114_BO6),
.I5(CLBLM_R_X7Y113_SLICE_X8Y113_CO6),
.O5(CLBLL_L_X4Y113_SLICE_X4Y113_CO5),
.O6(CLBLL_L_X4Y113_SLICE_X4Y113_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfbbf32b3b33b2032)
  ) CLBLL_L_X4Y113_SLICE_X4Y113_BLUT (
.I0(CLBLM_R_X7Y113_SLICE_X8Y113_DO6),
.I1(CLBLM_R_X5Y113_SLICE_X7Y113_BO6),
.I2(CLBLL_L_X4Y113_SLICE_X4Y113_DO6),
.I3(CLBLM_R_X5Y110_SLICE_X6Y110_CO6),
.I4(CLBLM_R_X5Y112_SLICE_X6Y112_DO6),
.I5(CLBLL_L_X4Y113_SLICE_X4Y113_CO6),
.O5(CLBLL_L_X4Y113_SLICE_X4Y113_BO5),
.O6(CLBLL_L_X4Y113_SLICE_X4Y113_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'ha05fa05f3333cc93)
  ) CLBLL_L_X4Y113_SLICE_X4Y113_ALUT (
.I0(RIOB33_X105Y107_IOB_X1Y108_I),
.I1(CLBLM_R_X5Y113_SLICE_X7Y113_BO6),
.I2(LIOB33_X0Y115_IOB_X0Y115_I),
.I3(CLBLM_R_X5Y110_SLICE_X6Y110_CO6),
.I4(CLBLM_R_X5Y112_SLICE_X6Y112_DO6),
.I5(1'b1),
.O5(CLBLL_L_X4Y113_SLICE_X4Y113_AO5),
.O6(CLBLL_L_X4Y113_SLICE_X4Y113_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X4Y113_SLICE_X5Y113_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y113_SLICE_X5Y113_DO5),
.O6(CLBLL_L_X4Y113_SLICE_X5Y113_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h44006c006c446c6c)
  ) CLBLL_L_X4Y113_SLICE_X5Y113_CLUT (
.I0(LIOB33_X0Y115_IOB_X0Y115_I),
.I1(CLBLM_R_X7Y114_SLICE_X8Y114_BO6),
.I2(RIOB33_X105Y103_IOB_X1Y104_I),
.I3(CLBLM_R_X5Y111_SLICE_X6Y111_BO6),
.I4(RIOB33_X105Y103_IOB_X1Y103_I),
.I5(CLBLM_R_X5Y113_SLICE_X7Y113_AO6),
.O5(CLBLL_L_X4Y113_SLICE_X5Y113_CO5),
.O6(CLBLL_L_X4Y113_SLICE_X5Y113_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h9666cccc999633cc)
  ) CLBLL_L_X4Y113_SLICE_X5Y113_BLUT (
.I0(RIOB33_X105Y103_IOB_X1Y104_I),
.I1(CLBLM_R_X7Y114_SLICE_X8Y114_BO6),
.I2(RIOB33_X105Y103_IOB_X1Y103_I),
.I3(CLBLM_R_X5Y113_SLICE_X7Y113_AO6),
.I4(LIOB33_X0Y115_IOB_X0Y115_I),
.I5(CLBLM_R_X5Y111_SLICE_X6Y111_BO6),
.O5(CLBLL_L_X4Y113_SLICE_X5Y113_BO5),
.O6(CLBLL_L_X4Y113_SLICE_X5Y113_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h3cc3cc330ccfccff)
  ) CLBLL_L_X4Y113_SLICE_X5Y113_ALUT (
.I0(1'b1),
.I1(CLBLM_R_X5Y111_SLICE_X6Y111_BO6),
.I2(RIOB33_X105Y103_IOB_X1Y103_I),
.I3(CLBLM_R_X5Y113_SLICE_X7Y113_AO6),
.I4(LIOB33_X0Y115_IOB_X0Y115_I),
.I5(1'b1),
.O5(CLBLL_L_X4Y113_SLICE_X5Y113_AO5),
.O6(CLBLL_L_X4Y113_SLICE_X5Y113_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h55555555aaaaaaaa)
  ) CLBLL_L_X4Y114_SLICE_X4Y114_DLUT (
.I0(CLBLL_L_X4Y113_SLICE_X5Y113_BO6),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(CLBLL_L_X4Y112_SLICE_X5Y112_BO6),
.O5(CLBLL_L_X4Y114_SLICE_X4Y114_DO5),
.O6(CLBLL_L_X4Y114_SLICE_X4Y114_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hdf5d5d455d454504)
  ) CLBLL_L_X4Y114_SLICE_X4Y114_CLUT (
.I0(CLBLM_R_X7Y114_SLICE_X8Y114_CO6),
.I1(CLBLL_L_X4Y113_SLICE_X5Y113_AO5),
.I2(CLBLM_R_X7Y114_SLICE_X8Y114_AO5),
.I3(CLBLL_L_X4Y114_SLICE_X4Y114_AO5),
.I4(CLBLL_L_X4Y112_SLICE_X5Y112_BO6),
.I5(CLBLM_R_X5Y113_SLICE_X7Y113_AO5),
.O5(CLBLL_L_X4Y114_SLICE_X4Y114_CO5),
.O6(CLBLL_L_X4Y114_SLICE_X4Y114_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h5f05ff55c3c33333)
  ) CLBLL_L_X4Y114_SLICE_X4Y114_BLUT (
.I0(CLBLM_R_X7Y114_SLICE_X8Y114_AO5),
.I1(CLBLM_R_X7Y114_SLICE_X8Y114_BO6),
.I2(LIOB33_X0Y115_IOB_X0Y115_I),
.I3(CLBLM_R_X5Y113_SLICE_X7Y113_AO5),
.I4(RIOB33_X105Y103_IOB_X1Y104_I),
.I5(1'b1),
.O5(CLBLL_L_X4Y114_SLICE_X4Y114_BO5),
.O6(CLBLL_L_X4Y114_SLICE_X4Y114_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h3f3f3f3f0f0fffff)
  ) CLBLL_L_X4Y114_SLICE_X4Y114_ALUT (
.I0(1'b1),
.I1(LIOB33_X0Y115_IOB_X0Y116_I),
.I2(LIOB33_X0Y115_IOB_X0Y115_I),
.I3(1'b1),
.I4(RIOB33_X105Y103_IOB_X1Y104_I),
.I5(1'b1),
.O5(CLBLL_L_X4Y114_SLICE_X4Y114_AO5),
.O6(CLBLL_L_X4Y114_SLICE_X4Y114_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X4Y114_SLICE_X5Y114_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y114_SLICE_X5Y114_DO5),
.O6(CLBLL_L_X4Y114_SLICE_X5Y114_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X4Y114_SLICE_X5Y114_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y114_SLICE_X5Y114_CO5),
.O6(CLBLL_L_X4Y114_SLICE_X5Y114_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X4Y114_SLICE_X5Y114_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y114_SLICE_X5Y114_BO5),
.O6(CLBLL_L_X4Y114_SLICE_X5Y114_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X4Y114_SLICE_X5Y114_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y114_SLICE_X5Y114_AO5),
.O6(CLBLL_L_X4Y114_SLICE_X5Y114_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h963c963cc396c396)
  ) CLBLL_L_X4Y115_SLICE_X4Y115_DLUT (
.I0(CLBLL_L_X4Y112_SLICE_X5Y112_BO6),
.I1(CLBLM_R_X7Y114_SLICE_X8Y114_CO6),
.I2(CLBLL_L_X4Y114_SLICE_X4Y114_BO6),
.I3(CLBLL_L_X4Y113_SLICE_X5Y113_AO5),
.I4(1'b1),
.I5(CLBLL_L_X4Y114_SLICE_X4Y114_BO5),
.O5(CLBLL_L_X4Y115_SLICE_X4Y115_DO5),
.O6(CLBLL_L_X4Y115_SLICE_X4Y115_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h00ffaa558a75ef10)
  ) CLBLL_L_X4Y115_SLICE_X4Y115_CLUT (
.I0(CLBLL_L_X4Y113_SLICE_X4Y113_AO6),
.I1(CLBLM_R_X7Y113_SLICE_X8Y113_CO6),
.I2(CLBLM_R_X7Y114_SLICE_X8Y114_DO6),
.I3(CLBLL_L_X4Y113_SLICE_X4Y113_AO5),
.I4(CLBLM_R_X7Y113_SLICE_X8Y113_DO6),
.I5(CLBLL_L_X4Y115_SLICE_X4Y115_BO6),
.O5(CLBLL_L_X4Y115_SLICE_X4Y115_CO5),
.O6(CLBLL_L_X4Y115_SLICE_X4Y115_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h00008ecf00000c8e)
  ) CLBLL_L_X4Y115_SLICE_X4Y115_BLUT (
.I0(CLBLL_L_X4Y112_SLICE_X5Y112_BO6),
.I1(CLBLL_L_X4Y114_SLICE_X4Y114_BO6),
.I2(CLBLM_R_X7Y114_SLICE_X8Y114_CO6),
.I3(CLBLL_L_X4Y114_SLICE_X4Y114_BO5),
.I4(CLBLL_L_X4Y115_SLICE_X4Y115_AO6),
.I5(CLBLL_L_X4Y113_SLICE_X5Y113_AO5),
.O5(CLBLL_L_X4Y115_SLICE_X4Y115_BO5),
.O6(CLBLL_L_X4Y115_SLICE_X4Y115_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h3333cccca55aa596)
  ) CLBLL_L_X4Y115_SLICE_X4Y115_ALUT (
.I0(CLBLM_R_X7Y113_SLICE_X8Y113_DO6),
.I1(CLBLM_R_X7Y114_SLICE_X8Y114_DO6),
.I2(CLBLL_L_X4Y113_SLICE_X4Y113_AO6),
.I3(CLBLL_L_X4Y115_SLICE_X4Y115_BO6),
.I4(CLBLM_R_X7Y113_SLICE_X8Y113_CO6),
.I5(1'b1),
.O5(CLBLL_L_X4Y115_SLICE_X4Y115_AO5),
.O6(CLBLL_L_X4Y115_SLICE_X4Y115_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X4Y115_SLICE_X5Y115_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y115_SLICE_X5Y115_DO5),
.O6(CLBLL_L_X4Y115_SLICE_X5Y115_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X4Y115_SLICE_X5Y115_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y115_SLICE_X5Y115_CO5),
.O6(CLBLL_L_X4Y115_SLICE_X5Y115_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X4Y115_SLICE_X5Y115_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y115_SLICE_X5Y115_BO5),
.O6(CLBLL_L_X4Y115_SLICE_X5Y115_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X4Y115_SLICE_X5Y115_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y115_SLICE_X5Y115_AO5),
.O6(CLBLL_L_X4Y115_SLICE_X5Y115_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X4Y116_SLICE_X4Y116_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y116_SLICE_X4Y116_DO5),
.O6(CLBLL_L_X4Y116_SLICE_X4Y116_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X4Y116_SLICE_X4Y116_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y116_SLICE_X4Y116_CO5),
.O6(CLBLL_L_X4Y116_SLICE_X4Y116_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X4Y116_SLICE_X4Y116_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y116_SLICE_X4Y116_BO5),
.O6(CLBLL_L_X4Y116_SLICE_X4Y116_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0f0f0f0ff0f0f0f0)
  ) CLBLL_L_X4Y116_SLICE_X4Y116_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(CLBLL_L_X4Y115_SLICE_X4Y115_AO6),
.I3(1'b1),
.I4(1'b1),
.I5(CLBLL_L_X4Y114_SLICE_X4Y114_CO6),
.O5(CLBLL_L_X4Y116_SLICE_X4Y116_AO5),
.O6(CLBLL_L_X4Y116_SLICE_X4Y116_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X4Y116_SLICE_X5Y116_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y116_SLICE_X5Y116_DO5),
.O6(CLBLL_L_X4Y116_SLICE_X5Y116_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X4Y116_SLICE_X5Y116_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y116_SLICE_X5Y116_CO5),
.O6(CLBLL_L_X4Y116_SLICE_X5Y116_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X4Y116_SLICE_X5Y116_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y116_SLICE_X5Y116_BO5),
.O6(CLBLL_L_X4Y116_SLICE_X5Y116_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X4Y116_SLICE_X5Y116_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y116_SLICE_X5Y116_AO5),
.O6(CLBLL_L_X4Y116_SLICE_X5Y116_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X8Y103_SLICE_X10Y103_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X8Y103_SLICE_X10Y103_DO5),
.O6(CLBLM_L_X8Y103_SLICE_X10Y103_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X8Y103_SLICE_X10Y103_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X8Y103_SLICE_X10Y103_CO5),
.O6(CLBLM_L_X8Y103_SLICE_X10Y103_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h47080b0844084408)
  ) CLBLM_L_X8Y103_SLICE_X10Y103_BLUT (
.I0(LIOB33_SING_X0Y100_IOB_X0Y100_I),
.I1(RIOB33_X105Y101_IOB_X1Y102_I),
.I2(RIOB33_X105Y101_IOB_X1Y101_I),
.I3(RIOB33_X105Y113_IOB_X1Y113_I),
.I4(RIOB33_X105Y111_IOB_X1Y112_I),
.I5(RIOB33_X105Y103_IOB_X1Y103_I),
.O5(CLBLM_L_X8Y103_SLICE_X10Y103_BO5),
.O6(CLBLM_L_X8Y103_SLICE_X10Y103_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'ha0a05f5fff00ff5f)
  ) CLBLM_L_X8Y103_SLICE_X10Y103_ALUT (
.I0(LIOB33_X0Y101_IOB_X0Y101_I),
.I1(1'b1),
.I2(RIOB33_X105Y101_IOB_X1Y101_I),
.I3(CLBLM_L_X8Y103_SLICE_X10Y103_BO6),
.I4(CLBLM_R_X7Y103_SLICE_X8Y103_BO6),
.I5(1'b1),
.O5(CLBLM_L_X8Y103_SLICE_X10Y103_AO5),
.O6(CLBLM_L_X8Y103_SLICE_X10Y103_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X8Y103_SLICE_X11Y103_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X8Y103_SLICE_X11Y103_DO5),
.O6(CLBLM_L_X8Y103_SLICE_X11Y103_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X8Y103_SLICE_X11Y103_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X8Y103_SLICE_X11Y103_CO5),
.O6(CLBLM_L_X8Y103_SLICE_X11Y103_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hbc703bf7438fc408)
  ) CLBLM_L_X8Y103_SLICE_X11Y103_BLUT (
.I0(RIOB33_X105Y101_IOB_X1Y101_I),
.I1(LIOB33_X0Y101_IOB_X0Y102_I),
.I2(CLBLM_L_X8Y103_SLICE_X10Y103_AO5),
.I3(RIOB33_X105Y101_IOB_X1Y102_I),
.I4(CLBLM_L_X10Y103_SLICE_X12Y103_AO6),
.I5(CLBLM_L_X10Y103_SLICE_X12Y103_CO6),
.O5(CLBLM_L_X8Y103_SLICE_X11Y103_BO5),
.O6(CLBLM_L_X8Y103_SLICE_X11Y103_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h7887878787787878)
  ) CLBLM_L_X8Y103_SLICE_X11Y103_ALUT (
.I0(RIOB33_X105Y101_IOB_X1Y101_I),
.I1(LIOB33_X0Y103_IOB_X0Y104_I),
.I2(CLBLM_L_X8Y104_SLICE_X10Y104_CO6),
.I3(LIOB33_X0Y101_IOB_X0Y102_I),
.I4(RIOB33_X105Y101_IOB_X1Y102_I),
.I5(CLBLM_L_X10Y103_SLICE_X12Y103_CO6),
.O5(CLBLM_L_X8Y103_SLICE_X11Y103_AO5),
.O6(CLBLM_L_X8Y103_SLICE_X11Y103_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h3fc03fc0c53a956a)
  ) CLBLM_L_X8Y104_SLICE_X10Y104_DLUT (
.I0(CLBLM_R_X7Y103_SLICE_X8Y103_BO6),
.I1(RIOB33_X105Y101_IOB_X1Y102_I),
.I2(LIOB33_X0Y101_IOB_X0Y101_I),
.I3(CLBLM_L_X10Y104_SLICE_X12Y104_AO6),
.I4(RIOB33_X105Y101_IOB_X1Y101_I),
.I5(CLBLM_L_X8Y103_SLICE_X10Y103_BO6),
.O5(CLBLM_L_X8Y104_SLICE_X10Y104_DO5),
.O6(CLBLM_L_X8Y104_SLICE_X10Y104_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hffc3ffc3d741c300)
  ) CLBLM_L_X8Y104_SLICE_X10Y104_CLUT (
.I0(CLBLM_R_X7Y103_SLICE_X8Y103_BO6),
.I1(CLBLM_L_X10Y102_SLICE_X12Y102_AO6),
.I2(CLBLM_L_X10Y104_SLICE_X12Y104_AO6),
.I3(CLBLM_L_X8Y104_SLICE_X10Y104_AO5),
.I4(CLBLM_L_X8Y104_SLICE_X10Y104_AO6),
.I5(CLBLM_L_X8Y103_SLICE_X10Y103_BO6),
.O5(CLBLM_L_X8Y104_SLICE_X10Y104_CO5),
.O6(CLBLM_L_X8Y104_SLICE_X10Y104_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h639c66999c639966)
  ) CLBLM_L_X8Y104_SLICE_X10Y104_BLUT (
.I0(CLBLM_L_X8Y103_SLICE_X10Y103_BO6),
.I1(CLBLM_L_X10Y104_SLICE_X12Y104_AO6),
.I2(CLBLM_R_X7Y103_SLICE_X8Y103_BO6),
.I3(CLBLM_L_X10Y102_SLICE_X12Y102_AO6),
.I4(CLBLM_L_X8Y104_SLICE_X10Y104_AO6),
.I5(CLBLM_L_X8Y104_SLICE_X10Y104_AO5),
.O5(CLBLM_L_X8Y104_SLICE_X10Y104_BO5),
.O6(CLBLM_L_X8Y104_SLICE_X10Y104_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h5f5f5f5f0f0fffff)
  ) CLBLM_L_X8Y104_SLICE_X10Y104_ALUT (
.I0(LIOB33_X0Y101_IOB_X0Y101_I),
.I1(1'b1),
.I2(RIOB33_X105Y101_IOB_X1Y101_I),
.I3(1'b1),
.I4(LIOB33_X0Y101_IOB_X0Y102_I),
.I5(1'b1),
.O5(CLBLM_L_X8Y104_SLICE_X10Y104_AO5),
.O6(CLBLM_L_X8Y104_SLICE_X10Y104_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hfdc4f731dc407310)
  ) CLBLM_L_X8Y104_SLICE_X11Y104_DLUT (
.I0(CLBLM_L_X8Y103_SLICE_X11Y103_AO6),
.I1(CLBLM_L_X8Y105_SLICE_X11Y105_AO5),
.I2(CLBLM_R_X7Y104_SLICE_X9Y104_AO5),
.I3(CLBLM_R_X7Y105_SLICE_X8Y105_AO6),
.I4(CLBLM_L_X10Y104_SLICE_X12Y104_CO6),
.I5(CLBLM_L_X8Y104_SLICE_X11Y104_BO6),
.O5(CLBLM_L_X8Y104_SLICE_X11Y104_DO5),
.O6(CLBLM_L_X8Y104_SLICE_X11Y104_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h7fffbf3f153f2a00)
  ) CLBLM_L_X8Y104_SLICE_X11Y104_CLUT (
.I0(RIOB33_X105Y101_IOB_X1Y101_I),
.I1(LIOB33_X0Y117_IOB_X0Y117_I),
.I2(LIOB33_X0Y105_IOB_X0Y105_I),
.I3(LIOB33_X0Y103_IOB_X0Y104_I),
.I4(CLBLM_L_X8Y103_SLICE_X11Y103_BO6),
.I5(CLBLM_L_X8Y104_SLICE_X11Y104_BO6),
.O5(CLBLM_L_X8Y104_SLICE_X11Y104_CO5),
.O6(CLBLM_L_X8Y104_SLICE_X11Y104_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h7f13b320ff5fffa0)
  ) CLBLM_L_X8Y104_SLICE_X11Y104_BLUT (
.I0(RIOB33_X105Y101_IOB_X1Y101_I),
.I1(LIOB33_X0Y117_IOB_X0Y117_I),
.I2(LIOB33_X0Y101_IOB_X0Y102_I),
.I3(CLBLM_R_X7Y104_SLICE_X8Y104_DO6),
.I4(CLBLM_L_X8Y104_SLICE_X10Y104_DO6),
.I5(LIOB33_X0Y103_IOB_X0Y104_I),
.O5(CLBLM_L_X8Y104_SLICE_X11Y104_BO5),
.O6(CLBLM_L_X8Y104_SLICE_X11Y104_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h69a55a69965aa596)
  ) CLBLM_L_X8Y104_SLICE_X11Y104_ALUT (
.I0(CLBLM_R_X7Y105_SLICE_X8Y105_AO6),
.I1(CLBLM_R_X7Y104_SLICE_X9Y104_AO5),
.I2(CLBLM_L_X10Y104_SLICE_X12Y104_CO6),
.I3(CLBLM_L_X8Y104_SLICE_X11Y104_BO6),
.I4(CLBLM_L_X8Y103_SLICE_X11Y103_AO6),
.I5(CLBLM_L_X8Y105_SLICE_X11Y105_AO5),
.O5(CLBLM_L_X8Y104_SLICE_X11Y104_AO5),
.O6(CLBLM_L_X8Y104_SLICE_X11Y104_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X8Y105_SLICE_X10Y105_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X8Y105_SLICE_X10Y105_DO5),
.O6(CLBLM_L_X8Y105_SLICE_X10Y105_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X8Y105_SLICE_X10Y105_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X8Y105_SLICE_X10Y105_CO5),
.O6(CLBLM_L_X8Y105_SLICE_X10Y105_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h6fff06669fff0999)
  ) CLBLM_L_X8Y105_SLICE_X10Y105_BLUT (
.I0(CLBLM_R_X7Y105_SLICE_X8Y105_AO6),
.I1(CLBLM_L_X8Y104_SLICE_X11Y104_CO6),
.I2(LIOB33_X0Y115_IOB_X0Y116_I),
.I3(LIOB33_X0Y107_IOB_X0Y107_I),
.I4(CLBLM_R_X7Y105_SLICE_X9Y105_BO6),
.I5(CLBLM_L_X8Y106_SLICE_X11Y106_AO6),
.O5(CLBLM_L_X8Y105_SLICE_X10Y105_BO5),
.O6(CLBLM_L_X8Y105_SLICE_X10Y105_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0fff0fff55ff55ff)
  ) CLBLM_L_X8Y105_SLICE_X10Y105_ALUT (
.I0(RIOB33_X105Y101_IOB_X1Y101_I),
.I1(1'b1),
.I2(LIOB33_X0Y115_IOB_X0Y116_I),
.I3(LIOB33_X0Y105_IOB_X0Y106_I),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X8Y105_SLICE_X10Y105_AO5),
.O6(CLBLM_L_X8Y105_SLICE_X10Y105_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h96996696cc33cccc)
  ) CLBLM_L_X8Y105_SLICE_X11Y105_DLUT (
.I0(RIOB33_X105Y101_IOB_X1Y102_I),
.I1(CLBLM_L_X10Y105_SLICE_X13Y105_BO6),
.I2(RIOB33_X105Y101_IOB_X1Y101_I),
.I3(CLBLM_L_X10Y103_SLICE_X12Y103_DO6),
.I4(CLBLM_L_X10Y105_SLICE_X12Y105_CO6),
.I5(LIOB33_X0Y105_IOB_X0Y105_I),
.O5(CLBLM_L_X8Y105_SLICE_X11Y105_DO5),
.O6(CLBLM_L_X8Y105_SLICE_X11Y105_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hf9ff99f990990090)
  ) CLBLM_L_X8Y105_SLICE_X11Y105_CLUT (
.I0(CLBLM_L_X10Y105_SLICE_X13Y105_AO5),
.I1(CLBLM_L_X10Y105_SLICE_X13Y105_BO6),
.I2(CLBLM_L_X8Y105_SLICE_X11Y105_AO5),
.I3(CLBLM_L_X10Y105_SLICE_X12Y105_CO6),
.I4(CLBLM_L_X10Y103_SLICE_X12Y103_DO6),
.I5(CLBLM_L_X8Y105_SLICE_X10Y105_AO5),
.O5(CLBLM_L_X8Y105_SLICE_X11Y105_CO5),
.O6(CLBLM_L_X8Y105_SLICE_X11Y105_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h3c96c36996c3693c)
  ) CLBLM_L_X8Y105_SLICE_X11Y105_BLUT (
.I0(CLBLM_L_X10Y105_SLICE_X12Y105_CO6),
.I1(CLBLM_L_X10Y105_SLICE_X13Y105_BO6),
.I2(CLBLM_L_X8Y105_SLICE_X10Y105_AO5),
.I3(CLBLM_L_X10Y103_SLICE_X12Y103_DO6),
.I4(CLBLM_L_X10Y105_SLICE_X13Y105_AO5),
.I5(CLBLM_L_X8Y105_SLICE_X11Y105_AO5),
.O5(CLBLM_L_X8Y105_SLICE_X11Y105_BO5),
.O6(CLBLM_L_X8Y105_SLICE_X11Y105_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h33ff33ff0fff0fff)
  ) CLBLM_L_X8Y105_SLICE_X11Y105_ALUT (
.I0(1'b1),
.I1(LIOB33_X0Y103_IOB_X0Y104_I),
.I2(LIOB33_X0Y105_IOB_X0Y105_I),
.I3(RIOB33_X105Y101_IOB_X1Y101_I),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X8Y105_SLICE_X11Y105_AO5),
.O6(CLBLM_L_X8Y105_SLICE_X11Y105_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h2dd2b44bd22d4bb4)
  ) CLBLM_L_X8Y106_SLICE_X10Y106_DLUT (
.I0(CLBLM_L_X8Y104_SLICE_X11Y104_AO6),
.I1(CLBLM_L_X8Y106_SLICE_X10Y106_AO6),
.I2(CLBLM_L_X8Y104_SLICE_X11Y104_DO6),
.I3(CLBLM_L_X8Y106_SLICE_X10Y106_AO5),
.I4(CLBLM_R_X7Y105_SLICE_X9Y105_BO6),
.I5(CLBLM_L_X8Y105_SLICE_X11Y105_BO6),
.O5(CLBLM_L_X8Y106_SLICE_X10Y106_DO5),
.O6(CLBLM_L_X8Y106_SLICE_X10Y106_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h002b2bffafffafff)
  ) CLBLM_L_X8Y106_SLICE_X10Y106_CLUT (
.I0(CLBLM_L_X8Y104_SLICE_X11Y104_CO6),
.I1(LIOB33_X0Y105_IOB_X0Y106_I),
.I2(CLBLM_L_X8Y106_SLICE_X11Y106_AO6),
.I3(CLBLM_L_X8Y105_SLICE_X11Y105_BO6),
.I4(LIOB33_X0Y107_IOB_X0Y107_I),
.I5(LIOB33_X0Y117_IOB_X0Y117_I),
.O5(CLBLM_L_X8Y106_SLICE_X10Y106_CO5),
.O6(CLBLM_L_X8Y106_SLICE_X10Y106_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hb7488b7477888778)
  ) CLBLM_L_X8Y106_SLICE_X10Y106_BLUT (
.I0(LIOB33_X0Y107_IOB_X0Y107_I),
.I1(LIOB33_X0Y117_IOB_X0Y117_I),
.I2(CLBLM_L_X8Y106_SLICE_X11Y106_AO6),
.I3(CLBLM_L_X8Y105_SLICE_X11Y105_BO6),
.I4(CLBLM_L_X8Y104_SLICE_X11Y104_CO6),
.I5(LIOB33_X0Y105_IOB_X0Y106_I),
.O5(CLBLM_L_X8Y106_SLICE_X10Y106_BO5),
.O6(CLBLM_L_X8Y106_SLICE_X10Y106_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h3f3f3f3f33ff33ff)
  ) CLBLM_L_X8Y106_SLICE_X10Y106_ALUT (
.I0(1'b1),
.I1(LIOB33_X0Y107_IOB_X0Y107_I),
.I2(LIOB33_X0Y115_IOB_X0Y116_I),
.I3(LIOB33_X0Y117_IOB_X0Y117_I),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X8Y106_SLICE_X10Y106_AO5),
.O6(CLBLM_L_X8Y106_SLICE_X10Y106_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hefbf8c23ce3b0802)
  ) CLBLM_L_X8Y106_SLICE_X11Y106_DLUT (
.I0(CLBLM_R_X7Y106_SLICE_X8Y106_AO6),
.I1(CLBLM_L_X8Y107_SLICE_X11Y107_AO6),
.I2(CLBLM_L_X8Y106_SLICE_X10Y106_BO6),
.I3(CLBLM_L_X8Y106_SLICE_X11Y106_CO6),
.I4(CLBLM_L_X8Y107_SLICE_X11Y107_BO5),
.I5(CLBLM_L_X8Y105_SLICE_X10Y105_BO6),
.O5(CLBLM_L_X8Y106_SLICE_X11Y106_DO5),
.O6(CLBLM_L_X8Y106_SLICE_X11Y106_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h6996a55a5aa56996)
  ) CLBLM_L_X8Y106_SLICE_X11Y106_CLUT (
.I0(CLBLM_L_X10Y108_SLICE_X13Y108_BO6),
.I1(CLBLM_L_X8Y106_SLICE_X10Y106_AO5),
.I2(CLBLM_L_X10Y106_SLICE_X13Y106_DO6),
.I3(CLBLM_L_X8Y105_SLICE_X11Y105_CO6),
.I4(CLBLM_L_X8Y104_SLICE_X11Y104_DO6),
.I5(CLBLM_L_X8Y105_SLICE_X11Y105_BO6),
.O5(CLBLM_L_X8Y106_SLICE_X11Y106_CO5),
.O6(CLBLM_L_X8Y106_SLICE_X11Y106_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h6999666996669996)
  ) CLBLM_L_X8Y106_SLICE_X11Y106_BLUT (
.I0(CLBLM_L_X8Y107_SLICE_X11Y107_BO5),
.I1(CLBLM_L_X8Y107_SLICE_X11Y107_AO6),
.I2(CLBLM_R_X7Y106_SLICE_X8Y106_AO6),
.I3(CLBLM_L_X8Y105_SLICE_X10Y105_BO6),
.I4(CLBLM_L_X8Y106_SLICE_X10Y106_BO6),
.I5(CLBLM_L_X8Y106_SLICE_X11Y106_CO6),
.O5(CLBLM_L_X8Y106_SLICE_X11Y106_BO5),
.O6(CLBLM_L_X8Y106_SLICE_X11Y106_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h69999666c3333ccc)
  ) CLBLM_L_X8Y106_SLICE_X11Y106_ALUT (
.I0(LIOB33_X0Y105_IOB_X0Y105_I),
.I1(CLBLM_L_X10Y103_SLICE_X12Y103_DO6),
.I2(RIOB33_X105Y101_IOB_X1Y102_I),
.I3(LIOB33_X0Y103_IOB_X0Y104_I),
.I4(CLBLM_L_X10Y105_SLICE_X12Y105_BO6),
.I5(RIOB33_X105Y101_IOB_X1Y101_I),
.O5(CLBLM_L_X8Y106_SLICE_X11Y106_AO5),
.O6(CLBLM_L_X8Y106_SLICE_X11Y106_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h82c3283c00820028)
  ) CLBLM_L_X8Y107_SLICE_X10Y107_DLUT (
.I0(CLBLM_L_X8Y105_SLICE_X10Y105_BO6),
.I1(CLBLM_L_X8Y107_SLICE_X11Y107_AO6),
.I2(CLBLM_L_X10Y106_SLICE_X12Y106_AO6),
.I3(CLBLM_L_X8Y106_SLICE_X10Y106_BO6),
.I4(CLBLM_L_X8Y106_SLICE_X10Y106_CO6),
.I5(CLBLM_R_X7Y106_SLICE_X8Y106_AO6),
.O5(CLBLM_L_X8Y107_SLICE_X10Y107_DO5),
.O6(CLBLM_L_X8Y107_SLICE_X10Y107_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hc639af50639caf50)
  ) CLBLM_L_X8Y107_SLICE_X10Y107_CLUT (
.I0(CLBLM_L_X8Y106_SLICE_X10Y106_CO6),
.I1(RIOB33_X105Y101_IOB_X1Y101_I),
.I2(CLBLM_L_X10Y106_SLICE_X12Y106_AO6),
.I3(CLBLM_L_X10Y107_SLICE_X12Y107_AO6),
.I4(LIOB33_X0Y107_IOB_X0Y108_I),
.I5(LIOB33_X0Y117_IOB_X0Y117_I),
.O5(CLBLM_L_X8Y107_SLICE_X10Y107_CO5),
.O6(CLBLM_L_X8Y107_SLICE_X10Y107_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h69c33c69963cc396)
  ) CLBLM_L_X8Y107_SLICE_X10Y107_BLUT (
.I0(CLBLM_R_X7Y106_SLICE_X9Y106_DO6),
.I1(CLBLM_L_X8Y106_SLICE_X11Y106_DO6),
.I2(CLBLM_L_X8Y107_SLICE_X11Y107_CO6),
.I3(CLBLM_R_X5Y107_SLICE_X7Y107_AO5),
.I4(CLBLM_L_X8Y106_SLICE_X11Y106_BO6),
.I5(CLBLM_L_X8Y108_SLICE_X10Y108_AO5),
.O5(CLBLM_L_X8Y107_SLICE_X10Y107_BO5),
.O6(CLBLM_L_X8Y107_SLICE_X10Y107_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h9669696996969669)
  ) CLBLM_L_X8Y107_SLICE_X10Y107_ALUT (
.I0(CLBLM_L_X8Y106_SLICE_X10Y106_CO6),
.I1(CLBLM_L_X10Y106_SLICE_X12Y106_AO6),
.I2(CLBLM_L_X8Y107_SLICE_X11Y107_AO6),
.I3(CLBLM_R_X7Y106_SLICE_X8Y106_AO6),
.I4(CLBLM_L_X8Y105_SLICE_X10Y105_BO6),
.I5(CLBLM_L_X8Y106_SLICE_X10Y106_BO6),
.O5(CLBLM_L_X8Y107_SLICE_X10Y107_AO5),
.O6(CLBLM_L_X8Y107_SLICE_X10Y107_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hfbbff22fb00b2002)
  ) CLBLM_L_X8Y107_SLICE_X11Y107_DLUT (
.I0(CLBLM_L_X8Y106_SLICE_X10Y106_CO6),
.I1(CLBLM_L_X10Y106_SLICE_X12Y106_AO6),
.I2(CLBLM_L_X10Y107_SLICE_X12Y107_AO6),
.I3(CLBLM_L_X8Y107_SLICE_X11Y107_AO5),
.I4(CLBLM_L_X8Y107_SLICE_X11Y107_AO6),
.I5(CLBLM_L_X8Y107_SLICE_X11Y107_BO6),
.O5(CLBLM_L_X8Y107_SLICE_X11Y107_DO5),
.O6(CLBLM_L_X8Y107_SLICE_X11Y107_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h39c69c63c639639c)
  ) CLBLM_L_X8Y107_SLICE_X11Y107_CLUT (
.I0(CLBLM_L_X10Y106_SLICE_X12Y106_AO6),
.I1(CLBLM_L_X10Y107_SLICE_X12Y107_AO6),
.I2(CLBLM_L_X8Y106_SLICE_X10Y106_CO6),
.I3(CLBLM_L_X8Y107_SLICE_X11Y107_AO5),
.I4(CLBLM_L_X8Y107_SLICE_X11Y107_AO6),
.I5(CLBLM_L_X8Y107_SLICE_X11Y107_BO6),
.O5(CLBLM_L_X8Y107_SLICE_X11Y107_CO5),
.O6(CLBLM_L_X8Y107_SLICE_X11Y107_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h33ff33ff77777777)
  ) CLBLM_L_X8Y107_SLICE_X11Y107_BLUT (
.I0(LIOB33_X0Y115_IOB_X0Y116_I),
.I1(LIOB33_X0Y109_IOB_X0Y109_I),
.I2(1'b1),
.I3(LIOB33_X0Y117_IOB_X0Y117_I),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X8Y107_SLICE_X11Y107_BO5),
.O6(CLBLM_L_X8Y107_SLICE_X11Y107_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h33ff33ff55ff55ff)
  ) CLBLM_L_X8Y107_SLICE_X11Y107_ALUT (
.I0(RIOB33_X105Y101_IOB_X1Y101_I),
.I1(LIOB33_X0Y117_IOB_X0Y117_I),
.I2(1'b1),
.I3(LIOB33_X0Y107_IOB_X0Y108_I),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X8Y107_SLICE_X11Y107_AO5),
.O6(CLBLM_L_X8Y107_SLICE_X11Y107_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h693c96c3c3693c96)
  ) CLBLM_L_X8Y108_SLICE_X10Y108_DLUT (
.I0(CLBLM_L_X8Y108_SLICE_X10Y108_AO6),
.I1(CLBLM_R_X11Y109_SLICE_X14Y109_BO6),
.I2(CLBLM_L_X10Y110_SLICE_X13Y110_AO6),
.I3(CLBLM_L_X10Y108_SLICE_X12Y108_AO6),
.I4(CLBLM_L_X10Y108_SLICE_X12Y108_DO6),
.I5(CLBLM_L_X8Y107_SLICE_X11Y107_DO6),
.O5(CLBLM_L_X8Y108_SLICE_X10Y108_DO5),
.O6(CLBLM_L_X8Y108_SLICE_X10Y108_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h5a9696a5a569695a)
  ) CLBLM_L_X8Y108_SLICE_X10Y108_CLUT (
.I0(CLBLM_L_X8Y108_SLICE_X10Y108_AO6),
.I1(CLBLM_L_X8Y107_SLICE_X11Y107_CO6),
.I2(CLBLM_L_X10Y108_SLICE_X12Y108_AO6),
.I3(CLBLM_L_X8Y108_SLICE_X10Y108_AO5),
.I4(CLBLM_L_X8Y106_SLICE_X11Y106_DO6),
.I5(CLBLM_L_X8Y107_SLICE_X11Y107_DO6),
.O5(CLBLM_L_X8Y108_SLICE_X10Y108_CO5),
.O6(CLBLM_L_X8Y108_SLICE_X10Y108_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h69c3963ca50f5af0)
  ) CLBLM_L_X8Y108_SLICE_X10Y108_BLUT (
.I0(LIOB33_X0Y107_IOB_X0Y108_I),
.I1(LIOB33_X0Y107_IOB_X0Y107_I),
.I2(CLBLM_L_X10Y106_SLICE_X12Y106_BO6),
.I3(LIOB33_X0Y117_IOB_X0Y117_I),
.I4(CLBLM_L_X8Y106_SLICE_X10Y106_CO6),
.I5(RIOB33_X105Y101_IOB_X1Y101_I),
.O5(CLBLM_L_X8Y108_SLICE_X10Y108_BO5),
.O6(CLBLM_L_X8Y108_SLICE_X10Y108_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h33ff33ff55ff55ff)
  ) CLBLM_L_X8Y108_SLICE_X10Y108_ALUT (
.I0(LIOB33_X0Y115_IOB_X0Y116_I),
.I1(LIOB33_X0Y117_IOB_X0Y117_I),
.I2(1'b1),
.I3(LIOB33_X0Y109_IOB_X0Y110_I),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X8Y108_SLICE_X10Y108_AO5),
.O6(CLBLM_L_X8Y108_SLICE_X10Y108_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h7fbf152abfbf2a2a)
  ) CLBLM_L_X8Y108_SLICE_X11Y108_DLUT (
.I0(CLBLM_L_X10Y106_SLICE_X12Y106_BO6),
.I1(LIOB33_X0Y117_IOB_X0Y117_I),
.I2(LIOB33_X0Y107_IOB_X0Y108_I),
.I3(LIOB33_X0Y107_IOB_X0Y107_I),
.I4(CLBLM_L_X8Y106_SLICE_X10Y106_CO6),
.I5(RIOB33_X105Y101_IOB_X1Y101_I),
.O5(CLBLM_L_X8Y108_SLICE_X11Y108_DO5),
.O6(CLBLM_L_X8Y108_SLICE_X11Y108_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hc6669c966ccc363c)
  ) CLBLM_L_X8Y108_SLICE_X11Y108_CLUT (
.I0(LIOB33_X0Y109_IOB_X0Y109_I),
.I1(CLBLM_L_X10Y108_SLICE_X12Y108_BO6),
.I2(CLBLM_L_X10Y109_SLICE_X12Y109_BO6),
.I3(LIOB33_X0Y117_IOB_X0Y117_I),
.I4(CLBLM_L_X8Y108_SLICE_X11Y108_DO6),
.I5(RIOB33_X105Y101_IOB_X1Y101_I),
.O5(CLBLM_L_X8Y108_SLICE_X11Y108_CO5),
.O6(CLBLM_L_X8Y108_SLICE_X11Y108_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hc639639caa55ff00)
  ) CLBLM_L_X8Y108_SLICE_X11Y108_BLUT (
.I0(CLBLM_L_X8Y108_SLICE_X11Y108_DO6),
.I1(LIOB33_X0Y109_IOB_X0Y110_I),
.I2(LIOB33_X0Y109_IOB_X0Y109_I),
.I3(CLBLM_L_X10Y108_SLICE_X12Y108_AO6),
.I4(CLBLM_L_X10Y109_SLICE_X12Y109_BO6),
.I5(LIOB33_X0Y117_IOB_X0Y117_I),
.O5(CLBLM_L_X8Y108_SLICE_X11Y108_BO5),
.O6(CLBLM_L_X8Y108_SLICE_X11Y108_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h02233bbfaaffffff)
  ) CLBLM_L_X8Y108_SLICE_X11Y108_ALUT (
.I0(CLBLM_L_X8Y108_SLICE_X11Y108_DO6),
.I1(LIOB33_X0Y109_IOB_X0Y110_I),
.I2(LIOB33_X0Y109_IOB_X0Y109_I),
.I3(CLBLM_L_X10Y109_SLICE_X12Y109_BO6),
.I4(CLBLM_L_X10Y108_SLICE_X12Y108_AO6),
.I5(LIOB33_X0Y117_IOB_X0Y117_I),
.O5(CLBLM_L_X8Y108_SLICE_X11Y108_AO5),
.O6(CLBLM_L_X8Y108_SLICE_X11Y108_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h9fa0a350a0a06ca0)
  ) CLBLM_L_X8Y109_SLICE_X10Y109_DLUT (
.I0(LIOB33_X0Y107_IOB_X0Y108_I),
.I1(LIOB33_X0Y105_IOB_X0Y106_I),
.I2(RIOB33_X105Y109_IOB_X1Y110_I),
.I3(RIOB33_X105Y111_IOB_X1Y111_I),
.I4(CLBLM_L_X10Y109_SLICE_X12Y109_DO6),
.I5(LIOB33_X0Y107_IOB_X0Y107_I),
.O5(CLBLM_L_X8Y109_SLICE_X10Y109_DO5),
.O6(CLBLM_L_X8Y109_SLICE_X10Y109_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h95ff6a00a93356cc)
  ) CLBLM_L_X8Y109_SLICE_X10Y109_CLUT (
.I0(LIOB33_X0Y109_IOB_X0Y109_I),
.I1(CLBLM_R_X7Y109_SLICE_X9Y109_AO6),
.I2(LIOB33_X0Y107_IOB_X0Y108_I),
.I3(RIOB33_X105Y109_IOB_X1Y109_I),
.I4(CLBLM_L_X8Y109_SLICE_X10Y109_DO6),
.I5(CLBLM_R_X11Y106_SLICE_X15Y106_AO5),
.O5(CLBLM_L_X8Y109_SLICE_X10Y109_CO5),
.O6(CLBLM_L_X8Y109_SLICE_X10Y109_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h69a5c30f965a3cf0)
  ) CLBLM_L_X8Y109_SLICE_X10Y109_BLUT (
.I0(RIOB33_X105Y109_IOB_X1Y110_I),
.I1(LIOB33_X0Y107_IOB_X0Y108_I),
.I2(CLBLM_L_X10Y109_SLICE_X12Y109_CO6),
.I3(RIOB33_X105Y109_IOB_X1Y109_I),
.I4(LIOB33_X0Y107_IOB_X0Y107_I),
.I5(CLBLM_R_X11Y106_SLICE_X15Y106_AO5),
.O5(CLBLM_L_X8Y109_SLICE_X10Y109_BO5),
.O6(CLBLM_L_X8Y109_SLICE_X10Y109_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h1f5f7fff051f557f)
  ) CLBLM_L_X8Y109_SLICE_X10Y109_ALUT (
.I0(CLBLM_L_X8Y109_SLICE_X10Y109_DO6),
.I1(LIOB33_X0Y107_IOB_X0Y108_I),
.I2(RIOB33_X105Y109_IOB_X1Y109_I),
.I3(CLBLM_R_X7Y109_SLICE_X9Y109_AO6),
.I4(LIOB33_X0Y109_IOB_X0Y109_I),
.I5(CLBLM_R_X11Y106_SLICE_X15Y106_AO5),
.O5(CLBLM_L_X8Y109_SLICE_X10Y109_AO5),
.O6(CLBLM_L_X8Y109_SLICE_X10Y109_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X8Y109_SLICE_X11Y109_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X8Y109_SLICE_X11Y109_DO5),
.O6(CLBLM_L_X8Y109_SLICE_X11Y109_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X8Y109_SLICE_X11Y109_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X8Y109_SLICE_X11Y109_CO5),
.O6(CLBLM_L_X8Y109_SLICE_X11Y109_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X8Y109_SLICE_X11Y109_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X8Y109_SLICE_X11Y109_BO5),
.O6(CLBLM_L_X8Y109_SLICE_X11Y109_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X8Y109_SLICE_X11Y109_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X8Y109_SLICE_X11Y109_AO5),
.O6(CLBLM_L_X8Y109_SLICE_X11Y109_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X8Y110_SLICE_X10Y110_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X8Y110_SLICE_X10Y110_DO5),
.O6(CLBLM_L_X8Y110_SLICE_X10Y110_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h238c8c2302080802)
  ) CLBLM_L_X8Y110_SLICE_X10Y110_CLUT (
.I0(CLBLM_L_X8Y108_SLICE_X11Y108_AO6),
.I1(CLBLM_L_X8Y110_SLICE_X11Y110_CO6),
.I2(CLBLM_L_X8Y110_SLICE_X11Y110_BO6),
.I3(CLBLM_L_X10Y112_SLICE_X12Y112_AO6),
.I4(CLBLM_L_X8Y110_SLICE_X11Y110_AO5),
.I5(CLBLM_L_X8Y110_SLICE_X11Y110_AO6),
.O5(CLBLM_L_X8Y110_SLICE_X10Y110_CO5),
.O6(CLBLM_L_X8Y110_SLICE_X10Y110_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h59a69a65a659659a)
  ) CLBLM_L_X8Y110_SLICE_X10Y110_BLUT (
.I0(CLBLM_L_X8Y110_SLICE_X11Y110_AO5),
.I1(CLBLM_L_X8Y110_SLICE_X11Y110_BO6),
.I2(CLBLM_L_X8Y110_SLICE_X11Y110_AO6),
.I3(CLBLM_L_X8Y112_SLICE_X10Y112_AO6),
.I4(CLBLM_L_X8Y108_SLICE_X11Y108_AO6),
.I5(CLBLM_L_X10Y110_SLICE_X13Y110_BO6),
.O5(CLBLM_L_X8Y110_SLICE_X10Y110_BO5),
.O6(CLBLM_L_X8Y110_SLICE_X10Y110_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h59a69a65a659659a)
  ) CLBLM_L_X8Y110_SLICE_X10Y110_ALUT (
.I0(CLBLM_L_X8Y110_SLICE_X11Y110_AO5),
.I1(CLBLM_L_X8Y110_SLICE_X11Y110_BO6),
.I2(CLBLM_L_X8Y110_SLICE_X11Y110_AO6),
.I3(CLBLM_L_X8Y110_SLICE_X11Y110_CO6),
.I4(CLBLM_L_X8Y108_SLICE_X11Y108_AO6),
.I5(CLBLM_L_X10Y112_SLICE_X12Y112_AO6),
.O5(CLBLM_L_X8Y110_SLICE_X10Y110_AO5),
.O6(CLBLM_L_X8Y110_SLICE_X10Y110_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X8Y110_SLICE_X11Y110_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X8Y110_SLICE_X11Y110_DO5),
.O6(CLBLM_L_X8Y110_SLICE_X11Y110_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h10f775f751f7f7f7)
  ) CLBLM_L_X8Y110_SLICE_X11Y110_CLUT (
.I0(CLBLM_R_X11Y109_SLICE_X14Y109_BO6),
.I1(CLBLM_L_X10Y110_SLICE_X12Y110_AO6),
.I2(CLBLM_L_X10Y109_SLICE_X12Y109_AO6),
.I3(RIOB33_X105Y101_IOB_X1Y101_I),
.I4(LIOB33_X0Y109_IOB_X0Y110_I),
.I5(LIOB33_X0Y109_IOB_X0Y109_I),
.O5(CLBLM_L_X8Y110_SLICE_X11Y110_CO5),
.O6(CLBLM_L_X8Y110_SLICE_X11Y110_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hd2aa2d554bffb400)
  ) CLBLM_L_X8Y110_SLICE_X11Y110_BLUT (
.I0(CLBLM_L_X10Y109_SLICE_X12Y109_AO6),
.I1(LIOB33_X0Y109_IOB_X0Y109_I),
.I2(LIOB33_X0Y109_IOB_X0Y110_I),
.I3(RIOB33_X105Y101_IOB_X1Y101_I),
.I4(CLBLM_R_X11Y109_SLICE_X14Y109_BO6),
.I5(CLBLM_L_X10Y110_SLICE_X12Y110_AO6),
.O5(CLBLM_L_X8Y110_SLICE_X11Y110_BO5),
.O6(CLBLM_L_X8Y110_SLICE_X11Y110_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h33ff33ff3f3f3f3f)
  ) CLBLM_L_X8Y110_SLICE_X11Y110_ALUT (
.I0(1'b1),
.I1(LIOB33_X0Y111_IOB_X0Y111_I),
.I2(RIOB33_X105Y101_IOB_X1Y101_I),
.I3(LIOB33_X0Y117_IOB_X0Y117_I),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X8Y110_SLICE_X11Y110_AO5),
.O6(CLBLM_L_X8Y110_SLICE_X11Y110_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X8Y111_SLICE_X10Y111_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X8Y111_SLICE_X10Y111_DO5),
.O6(CLBLM_L_X8Y111_SLICE_X10Y111_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h2b8ebbeeaf0affaa)
  ) CLBLM_L_X8Y111_SLICE_X10Y111_CLUT (
.I0(CLBLM_L_X8Y108_SLICE_X11Y108_AO6),
.I1(RIOB33_X105Y101_IOB_X1Y101_I),
.I2(LIOB33_X0Y111_IOB_X0Y111_I),
.I3(CLBLM_L_X10Y110_SLICE_X12Y110_BO6),
.I4(LIOB33_X0Y117_IOB_X0Y117_I),
.I5(LIOB33_X0Y109_IOB_X0Y110_I),
.O5(CLBLM_L_X8Y111_SLICE_X10Y111_CO5),
.O6(CLBLM_L_X8Y111_SLICE_X10Y111_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h7887877887788778)
  ) CLBLM_L_X8Y111_SLICE_X10Y111_BLUT (
.I0(LIOB33_X0Y111_IOB_X0Y111_I),
.I1(LIOB33_X0Y117_IOB_X0Y117_I),
.I2(CLBLM_L_X8Y108_SLICE_X11Y108_AO6),
.I3(CLBLM_L_X10Y110_SLICE_X12Y110_BO6),
.I4(LIOB33_X0Y109_IOB_X0Y110_I),
.I5(RIOB33_X105Y101_IOB_X1Y101_I),
.O5(CLBLM_L_X8Y111_SLICE_X10Y111_BO5),
.O6(CLBLM_L_X8Y111_SLICE_X10Y111_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h3fc0c03f956a6a95)
  ) CLBLM_L_X8Y111_SLICE_X10Y111_ALUT (
.I0(CLBLM_L_X10Y111_SLICE_X12Y111_CO6),
.I1(RIOB33_X105Y103_IOB_X1Y104_I),
.I2(LIOB33_X0Y109_IOB_X0Y110_I),
.I3(CLBLM_R_X11Y111_SLICE_X14Y111_AO5),
.I4(CLBLM_L_X10Y111_SLICE_X12Y111_BO6),
.I5(1'b1),
.O5(CLBLM_L_X8Y111_SLICE_X10Y111_AO5),
.O6(CLBLM_L_X8Y111_SLICE_X10Y111_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h33333333ffffffff)
  ) CLBLM_L_X8Y111_SLICE_X11Y111_DLUT (
.I0(1'b1),
.I1(LIOB33_X0Y109_IOB_X0Y110_I),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(RIOB33_X105Y103_IOB_X1Y104_I),
.O5(CLBLM_L_X8Y111_SLICE_X11Y111_DO5),
.O6(CLBLM_L_X8Y111_SLICE_X11Y111_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h1f5f7fff07175777)
  ) CLBLM_L_X8Y111_SLICE_X11Y111_CLUT (
.I0(CLBLM_L_X8Y111_SLICE_X11Y111_AO6),
.I1(CLBLM_L_X10Y111_SLICE_X12Y111_BO6),
.I2(RIOB33_X105Y103_IOB_X1Y104_I),
.I3(LIOB33_X0Y109_IOB_X0Y110_I),
.I4(LIOB33_X0Y111_IOB_X0Y111_I),
.I5(CLBLM_R_X11Y111_SLICE_X14Y111_AO5),
.O5(CLBLM_L_X8Y111_SLICE_X11Y111_CO5),
.O6(CLBLM_L_X8Y111_SLICE_X11Y111_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h4bd2b42db42d4bd2)
  ) CLBLM_L_X8Y111_SLICE_X11Y111_BLUT (
.I0(CLBLM_L_X8Y111_SLICE_X11Y111_DO6),
.I1(CLBLM_L_X10Y111_SLICE_X12Y111_BO6),
.I2(CLBLM_L_X10Y111_SLICE_X13Y111_AO5),
.I3(CLBLM_R_X11Y111_SLICE_X14Y111_AO5),
.I4(CLBLM_L_X10Y111_SLICE_X12Y111_DO6),
.I5(CLBLM_L_X10Y112_SLICE_X13Y112_CO6),
.O5(CLBLM_L_X8Y111_SLICE_X11Y111_BO5),
.O6(CLBLM_L_X8Y111_SLICE_X11Y111_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h66aa995577ff1155)
  ) CLBLM_L_X8Y111_SLICE_X11Y111_ALUT (
.I0(CLBLM_L_X10Y112_SLICE_X13Y112_CO6),
.I1(LIOB33_X0Y109_IOB_X0Y110_I),
.I2(1'b1),
.I3(RIOB33_X105Y105_IOB_X1Y105_I),
.I4(CLBLM_L_X10Y111_SLICE_X12Y111_DO6),
.I5(1'b1),
.O5(CLBLM_L_X8Y111_SLICE_X11Y111_AO5),
.O6(CLBLM_L_X8Y111_SLICE_X11Y111_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hb24dcf304db2cf30)
  ) CLBLM_L_X8Y112_SLICE_X10Y112_DLUT (
.I0(LIOB33_X0Y111_IOB_X0Y112_I),
.I1(CLBLM_L_X8Y111_SLICE_X10Y111_CO6),
.I2(CLBLM_L_X8Y112_SLICE_X11Y112_AO6),
.I3(CLBLM_L_X8Y112_SLICE_X10Y112_CO6),
.I4(LIOB33_X0Y117_IOB_X0Y117_I),
.I5(LIOB33_X0Y113_IOB_X0Y113_I),
.O5(CLBLM_L_X8Y112_SLICE_X10Y112_DO5),
.O6(CLBLM_L_X8Y112_SLICE_X10Y112_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h4bd2b42db42d4bd2)
  ) CLBLM_L_X8Y112_SLICE_X10Y112_CLUT (
.I0(CLBLM_L_X8Y110_SLICE_X11Y110_AO5),
.I1(CLBLM_L_X10Y112_SLICE_X12Y112_AO6),
.I2(CLBLM_L_X10Y110_SLICE_X13Y110_CO6),
.I3(CLBLM_L_X8Y110_SLICE_X11Y110_CO6),
.I4(CLBLM_R_X7Y112_SLICE_X8Y112_AO6),
.I5(CLBLM_R_X5Y112_SLICE_X7Y112_AO6),
.O5(CLBLM_L_X8Y112_SLICE_X10Y112_CO5),
.O6(CLBLM_L_X8Y112_SLICE_X10Y112_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h639cc6399c6339c6)
  ) CLBLM_L_X8Y112_SLICE_X10Y112_BLUT (
.I0(CLBLM_L_X8Y110_SLICE_X11Y110_CO6),
.I1(CLBLM_L_X10Y111_SLICE_X12Y111_AO6),
.I2(CLBLM_L_X10Y112_SLICE_X12Y112_AO6),
.I3(CLBLM_R_X5Y112_SLICE_X7Y112_AO6),
.I4(CLBLM_L_X8Y110_SLICE_X11Y110_AO5),
.I5(CLBLM_L_X10Y112_SLICE_X12Y112_BO6),
.O5(CLBLM_L_X8Y112_SLICE_X10Y112_BO5),
.O6(CLBLM_L_X8Y112_SLICE_X10Y112_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h00ffffff0aafafaf)
  ) CLBLM_L_X8Y112_SLICE_X10Y112_ALUT (
.I0(CLBLM_L_X8Y111_SLICE_X10Y111_CO6),
.I1(1'b1),
.I2(CLBLM_L_X8Y112_SLICE_X11Y112_AO6),
.I3(LIOB33_X0Y117_IOB_X0Y117_I),
.I4(LIOB33_X0Y111_IOB_X0Y112_I),
.I5(1'b1),
.O5(CLBLM_L_X8Y112_SLICE_X10Y112_AO5),
.O6(CLBLM_L_X8Y112_SLICE_X10Y112_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h4ddd8eeecfff0ccc)
  ) CLBLM_L_X8Y112_SLICE_X11Y112_DLUT (
.I0(LIOB33_X0Y109_IOB_X0Y110_I),
.I1(CLBLM_L_X10Y112_SLICE_X12Y112_BO6),
.I2(LIOB33_X0Y111_IOB_X0Y111_I),
.I3(RIOB33_X105Y101_IOB_X1Y102_I),
.I4(CLBLM_L_X10Y111_SLICE_X13Y111_CO6),
.I5(RIOB33_X105Y103_IOB_X1Y103_I),
.O5(CLBLM_L_X8Y112_SLICE_X11Y112_DO5),
.O6(CLBLM_L_X8Y112_SLICE_X11Y112_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h4dcf8e0cddffeecc)
  ) CLBLM_L_X8Y112_SLICE_X11Y112_CLUT (
.I0(LIOB33_X0Y109_IOB_X0Y110_I),
.I1(CLBLM_L_X8Y110_SLICE_X11Y110_CO6),
.I2(LIOB33_X0Y111_IOB_X0Y111_I),
.I3(RIOB33_X105Y101_IOB_X1Y102_I),
.I4(CLBLM_L_X10Y110_SLICE_X12Y110_DO6),
.I5(RIOB33_X105Y101_IOB_X1Y101_I),
.O5(CLBLM_L_X8Y112_SLICE_X11Y112_CO5),
.O6(CLBLM_L_X8Y112_SLICE_X11Y112_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h69999666c3333ccc)
  ) CLBLM_L_X8Y112_SLICE_X11Y112_BLUT (
.I0(LIOB33_X0Y111_IOB_X0Y111_I),
.I1(CLBLM_L_X10Y112_SLICE_X12Y112_BO6),
.I2(LIOB33_X0Y109_IOB_X0Y110_I),
.I3(RIOB33_X105Y103_IOB_X1Y103_I),
.I4(CLBLM_L_X10Y111_SLICE_X13Y111_CO6),
.I5(RIOB33_X105Y101_IOB_X1Y102_I),
.O5(CLBLM_L_X8Y112_SLICE_X11Y112_BO5),
.O6(CLBLM_L_X8Y112_SLICE_X11Y112_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h69a5c30f965a3cf0)
  ) CLBLM_L_X8Y112_SLICE_X11Y112_ALUT (
.I0(RIOB33_X105Y101_IOB_X1Y102_I),
.I1(LIOB33_X0Y111_IOB_X0Y111_I),
.I2(CLBLM_L_X10Y110_SLICE_X12Y110_DO6),
.I3(RIOB33_X105Y101_IOB_X1Y101_I),
.I4(LIOB33_X0Y109_IOB_X0Y110_I),
.I5(CLBLM_L_X8Y110_SLICE_X11Y110_CO6),
.O5(CLBLM_L_X8Y112_SLICE_X11Y112_AO5),
.O6(CLBLM_L_X8Y112_SLICE_X11Y112_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X8Y113_SLICE_X10Y113_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X8Y113_SLICE_X10Y113_DO5),
.O6(CLBLM_L_X8Y113_SLICE_X10Y113_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h7d14ff3cdd44ffcc)
  ) CLBLM_L_X8Y113_SLICE_X10Y113_CLUT (
.I0(LIOB33_X0Y111_IOB_X0Y112_I),
.I1(CLBLM_L_X8Y113_SLICE_X10Y113_AO6),
.I2(RIOB33_X105Y105_IOB_X1Y105_I),
.I3(CLBLM_L_X8Y111_SLICE_X11Y111_CO6),
.I4(RIOB33_X105Y103_IOB_X1Y104_I),
.I5(LIOB33_X0Y111_IOB_X0Y111_I),
.O5(CLBLM_L_X8Y113_SLICE_X10Y113_CO5),
.O6(CLBLM_L_X8Y113_SLICE_X10Y113_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h6ac0953f953f6ac0)
  ) CLBLM_L_X8Y113_SLICE_X10Y113_BLUT (
.I0(RIOB33_X105Y105_IOB_X1Y105_I),
.I1(RIOB33_X105Y103_IOB_X1Y104_I),
.I2(LIOB33_X0Y111_IOB_X0Y112_I),
.I3(LIOB33_X0Y111_IOB_X0Y111_I),
.I4(CLBLM_L_X8Y113_SLICE_X10Y113_AO6),
.I5(CLBLM_L_X8Y111_SLICE_X11Y111_CO6),
.O5(CLBLM_L_X8Y113_SLICE_X10Y113_BO5),
.O6(CLBLM_L_X8Y113_SLICE_X10Y113_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h96693cc36969c3c3)
  ) CLBLM_L_X8Y113_SLICE_X10Y113_ALUT (
.I0(RIOB33_X105Y107_IOB_X1Y107_I),
.I1(CLBLM_R_X7Y110_SLICE_X9Y110_BO5),
.I2(CLBLM_L_X10Y112_SLICE_X13Y112_BO6),
.I3(CLBLM_L_X8Y111_SLICE_X11Y111_AO5),
.I4(LIOB33_X0Y109_IOB_X0Y110_I),
.I5(1'b1),
.O5(CLBLM_L_X8Y113_SLICE_X10Y113_AO5),
.O6(CLBLM_L_X8Y113_SLICE_X10Y113_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X8Y113_SLICE_X11Y113_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X8Y113_SLICE_X11Y113_DO5),
.O6(CLBLM_L_X8Y113_SLICE_X11Y113_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X8Y113_SLICE_X11Y113_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X8Y113_SLICE_X11Y113_CO5),
.O6(CLBLM_L_X8Y113_SLICE_X11Y113_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X8Y113_SLICE_X11Y113_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X8Y113_SLICE_X11Y113_BO5),
.O6(CLBLM_L_X8Y113_SLICE_X11Y113_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X8Y113_SLICE_X11Y113_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X8Y113_SLICE_X11Y113_AO5),
.O6(CLBLM_L_X8Y113_SLICE_X11Y113_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X10Y102_SLICE_X12Y102_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X10Y102_SLICE_X12Y102_DO5),
.O6(CLBLM_L_X10Y102_SLICE_X12Y102_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hffaaff55ae085d04)
  ) CLBLM_L_X10Y102_SLICE_X12Y102_CLUT (
.I0(CLBLM_L_X10Y104_SLICE_X13Y104_AO6),
.I1(CLBLM_L_X10Y102_SLICE_X12Y102_AO6),
.I2(CLBLM_L_X10Y104_SLICE_X12Y104_AO6),
.I3(CLBLM_L_X10Y102_SLICE_X12Y102_AO5),
.I4(CLBLM_L_X10Y104_SLICE_X12Y104_BO6),
.I5(CLBLM_L_X10Y103_SLICE_X12Y103_BO6),
.O5(CLBLM_L_X10Y102_SLICE_X12Y102_CO5),
.O6(CLBLM_L_X10Y102_SLICE_X12Y102_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h6696669999699966)
  ) CLBLM_L_X10Y102_SLICE_X12Y102_BLUT (
.I0(CLBLM_L_X10Y104_SLICE_X12Y104_BO6),
.I1(CLBLM_L_X10Y104_SLICE_X13Y104_AO6),
.I2(CLBLM_L_X10Y104_SLICE_X12Y104_AO6),
.I3(CLBLM_L_X10Y103_SLICE_X12Y103_BO6),
.I4(CLBLM_L_X10Y102_SLICE_X12Y102_AO6),
.I5(CLBLM_L_X10Y102_SLICE_X12Y102_AO5),
.O5(CLBLM_L_X10Y102_SLICE_X12Y102_BO5),
.O6(CLBLM_L_X10Y102_SLICE_X12Y102_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h7777777733ff33ff)
  ) CLBLM_L_X10Y102_SLICE_X12Y102_ALUT (
.I0(LIOB33_X0Y101_IOB_X0Y101_I),
.I1(RIOB33_X105Y101_IOB_X1Y102_I),
.I2(1'b1),
.I3(LIOB33_X0Y101_IOB_X0Y102_I),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X10Y102_SLICE_X12Y102_AO5),
.O6(CLBLM_L_X10Y102_SLICE_X12Y102_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X10Y102_SLICE_X13Y102_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X10Y102_SLICE_X13Y102_DO5),
.O6(CLBLM_L_X10Y102_SLICE_X13Y102_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X10Y102_SLICE_X13Y102_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X10Y102_SLICE_X13Y102_CO5),
.O6(CLBLM_L_X10Y102_SLICE_X13Y102_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X10Y102_SLICE_X13Y102_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X10Y102_SLICE_X13Y102_BO5),
.O6(CLBLM_L_X10Y102_SLICE_X13Y102_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X10Y102_SLICE_X13Y102_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X10Y102_SLICE_X13Y102_AO5),
.O6(CLBLM_L_X10Y102_SLICE_X13Y102_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h4dd4dd44cffcffcc)
  ) CLBLM_L_X10Y103_SLICE_X12Y103_DLUT (
.I0(RIOB33_X105Y101_IOB_X1Y101_I),
.I1(CLBLM_L_X8Y104_SLICE_X10Y104_CO6),
.I2(RIOB33_X105Y101_IOB_X1Y102_I),
.I3(CLBLM_L_X10Y103_SLICE_X12Y103_CO6),
.I4(LIOB33_X0Y101_IOB_X0Y102_I),
.I5(LIOB33_X0Y103_IOB_X0Y104_I),
.O5(CLBLM_L_X10Y103_SLICE_X12Y103_DO5),
.O6(CLBLM_L_X10Y103_SLICE_X12Y103_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h6c6c6c6c939c936c)
  ) CLBLM_L_X10Y103_SLICE_X12Y103_CLUT (
.I0(RIOB33_X105Y103_IOB_X1Y103_I),
.I1(CLBLM_L_X10Y104_SLICE_X12Y104_BO6),
.I2(LIOB33_X0Y101_IOB_X0Y101_I),
.I3(CLBLM_L_X10Y104_SLICE_X12Y104_AO6),
.I4(RIOB33_X105Y101_IOB_X1Y102_I),
.I5(CLBLM_L_X10Y103_SLICE_X12Y103_BO6),
.O5(CLBLM_L_X10Y103_SLICE_X12Y103_CO5),
.O6(CLBLM_L_X10Y103_SLICE_X12Y103_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h1500d1cc44440000)
  ) CLBLM_L_X10Y103_SLICE_X12Y103_BLUT (
.I0(RIOB33_X105Y101_IOB_X1Y102_I),
.I1(RIOB33_X105Y103_IOB_X1Y103_I),
.I2(RIOB33_X105Y111_IOB_X1Y112_I),
.I3(RIOB33_X105Y103_IOB_X1Y104_I),
.I4(LIOB33_SING_X0Y100_IOB_X0Y100_I),
.I5(RIOB33_X105Y113_IOB_X1Y113_I),
.O5(CLBLM_L_X10Y103_SLICE_X12Y103_BO5),
.O6(CLBLM_L_X10Y103_SLICE_X12Y103_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'ha5a50f0fff05ff0f)
  ) CLBLM_L_X10Y103_SLICE_X12Y103_ALUT (
.I0(LIOB33_X0Y101_IOB_X0Y101_I),
.I1(1'b1),
.I2(CLBLM_L_X10Y104_SLICE_X12Y104_AO6),
.I3(CLBLM_L_X10Y103_SLICE_X12Y103_BO6),
.I4(RIOB33_X105Y101_IOB_X1Y102_I),
.I5(1'b1),
.O5(CLBLM_L_X10Y103_SLICE_X12Y103_AO5),
.O6(CLBLM_L_X10Y103_SLICE_X12Y103_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X10Y103_SLICE_X13Y103_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X10Y103_SLICE_X13Y103_DO5),
.O6(CLBLM_L_X10Y103_SLICE_X13Y103_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X10Y103_SLICE_X13Y103_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X10Y103_SLICE_X13Y103_CO5),
.O6(CLBLM_L_X10Y103_SLICE_X13Y103_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X10Y103_SLICE_X13Y103_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X10Y103_SLICE_X13Y103_BO5),
.O6(CLBLM_L_X10Y103_SLICE_X13Y103_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X10Y103_SLICE_X13Y103_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X10Y103_SLICE_X13Y103_AO5),
.O6(CLBLM_L_X10Y103_SLICE_X13Y103_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h260c0a0a26260000)
  ) CLBLM_L_X10Y104_SLICE_X12Y104_DLUT (
.I0(RIOB33_X105Y113_IOB_X1Y113_I),
.I1(LIOB33_SING_X0Y100_IOB_X0Y100_I),
.I2(RIOB33_X105Y103_IOB_X1Y103_I),
.I3(RIOB33_X105Y111_IOB_X1Y112_I),
.I4(RIOB33_X105Y103_IOB_X1Y104_I),
.I5(RIOB33_X105Y105_IOB_X1Y105_I),
.O5(CLBLM_L_X10Y104_SLICE_X12Y104_DO5),
.O6(CLBLM_L_X10Y104_SLICE_X12Y104_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h659a9a65a65959a6)
  ) CLBLM_L_X10Y104_SLICE_X12Y104_CLUT (
.I0(CLBLM_L_X10Y105_SLICE_X13Y105_AO6),
.I1(CLBLM_L_X8Y104_SLICE_X10Y104_CO6),
.I2(CLBLM_L_X10Y102_SLICE_X12Y102_BO6),
.I3(CLBLM_L_X10Y102_SLICE_X12Y102_CO6),
.I4(CLBLM_L_X10Y104_SLICE_X13Y104_BO6),
.I5(CLBLM_L_X8Y105_SLICE_X11Y105_AO6),
.O5(CLBLM_L_X10Y104_SLICE_X12Y104_CO5),
.O6(CLBLM_L_X10Y104_SLICE_X12Y104_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h134c6666b1ee0000)
  ) CLBLM_L_X10Y104_SLICE_X12Y104_BLUT (
.I0(RIOB33_X105Y103_IOB_X1Y104_I),
.I1(RIOB33_X105Y103_IOB_X1Y103_I),
.I2(RIOB33_X105Y111_IOB_X1Y112_I),
.I3(RIOB33_X105Y105_IOB_X1Y105_I),
.I4(RIOB33_X105Y113_IOB_X1Y113_I),
.I5(LIOB33_SING_X0Y100_IOB_X0Y100_I),
.O5(CLBLM_L_X10Y104_SLICE_X12Y104_BO5),
.O6(CLBLM_L_X10Y104_SLICE_X12Y104_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h15255aaac0f050a0)
  ) CLBLM_L_X10Y104_SLICE_X12Y104_ALUT (
.I0(RIOB33_X105Y101_IOB_X1Y102_I),
.I1(RIOB33_X105Y111_IOB_X1Y112_I),
.I2(RIOB33_X105Y113_IOB_X1Y113_I),
.I3(RIOB33_X105Y103_IOB_X1Y104_I),
.I4(RIOB33_X105Y103_IOB_X1Y103_I),
.I5(LIOB33_SING_X0Y100_IOB_X0Y100_I),
.O5(CLBLM_L_X10Y104_SLICE_X12Y104_AO5),
.O6(CLBLM_L_X10Y104_SLICE_X12Y104_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hff99ff999f099900)
  ) CLBLM_L_X10Y104_SLICE_X13Y104_DLUT (
.I0(CLBLM_R_X11Y104_SLICE_X14Y104_AO6),
.I1(CLBLM_R_X11Y104_SLICE_X15Y104_BO6),
.I2(CLBLM_L_X10Y104_SLICE_X12Y104_BO6),
.I3(CLBLM_L_X10Y104_SLICE_X13Y104_AO5),
.I4(CLBLM_L_X10Y104_SLICE_X13Y104_AO6),
.I5(CLBLM_L_X10Y104_SLICE_X12Y104_DO6),
.O5(CLBLM_L_X10Y104_SLICE_X13Y104_DO5),
.O6(CLBLM_L_X10Y104_SLICE_X13Y104_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h55aaff00a9560ff0)
  ) CLBLM_L_X10Y104_SLICE_X13Y104_CLUT (
.I0(RIOB33_X105Y103_IOB_X1Y104_I),
.I1(RIOB33_X105Y103_IOB_X1Y103_I),
.I2(CLBLM_L_X10Y104_SLICE_X12Y104_BO6),
.I3(CLBLM_R_X11Y104_SLICE_X15Y104_BO6),
.I4(LIOB33_X0Y101_IOB_X0Y101_I),
.I5(CLBLM_L_X10Y104_SLICE_X12Y104_DO6),
.O5(CLBLM_L_X10Y104_SLICE_X13Y104_CO5),
.O6(CLBLM_L_X10Y104_SLICE_X13Y104_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h559aaa65aa65559a)
  ) CLBLM_L_X10Y104_SLICE_X13Y104_BLUT (
.I0(CLBLM_R_X11Y104_SLICE_X15Y104_BO6),
.I1(CLBLM_L_X10Y104_SLICE_X12Y104_BO6),
.I2(CLBLM_L_X10Y104_SLICE_X13Y104_AO6),
.I3(CLBLM_L_X10Y104_SLICE_X12Y104_DO6),
.I4(CLBLM_R_X11Y104_SLICE_X14Y104_AO6),
.I5(CLBLM_L_X10Y104_SLICE_X13Y104_AO5),
.O5(CLBLM_L_X10Y104_SLICE_X13Y104_BO5),
.O6(CLBLM_L_X10Y104_SLICE_X13Y104_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h55ff55ff0fff0fff)
  ) CLBLM_L_X10Y104_SLICE_X13Y104_ALUT (
.I0(LIOB33_X0Y101_IOB_X0Y101_I),
.I1(1'b1),
.I2(LIOB33_X0Y101_IOB_X0Y102_I),
.I3(RIOB33_X105Y103_IOB_X1Y103_I),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X10Y104_SLICE_X13Y104_AO5),
.O6(CLBLM_L_X10Y104_SLICE_X13Y104_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h96c3f05a3c96f05a)
  ) CLBLM_L_X10Y105_SLICE_X12Y105_DLUT (
.I0(CLBLM_R_X11Y104_SLICE_X15Y104_AO6),
.I1(RIOB33_X105Y103_IOB_X1Y104_I),
.I2(CLBLM_R_X11Y104_SLICE_X14Y104_DO6),
.I3(CLBLM_L_X10Y105_SLICE_X12Y105_AO5),
.I4(LIOB33_X0Y101_IOB_X0Y102_I),
.I5(RIOB33_X105Y103_IOB_X1Y103_I),
.O5(CLBLM_L_X10Y105_SLICE_X12Y105_DO5),
.O6(CLBLM_L_X10Y105_SLICE_X12Y105_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h6c93a05f936c5fa0)
  ) CLBLM_L_X10Y105_SLICE_X12Y105_CLUT (
.I0(LIOB33_X0Y103_IOB_X0Y104_I),
.I1(RIOB33_X105Y103_IOB_X1Y103_I),
.I2(RIOB33_X105Y101_IOB_X1Y102_I),
.I3(CLBLM_L_X10Y102_SLICE_X12Y102_CO6),
.I4(LIOB33_X0Y101_IOB_X0Y102_I),
.I5(CLBLM_L_X10Y104_SLICE_X13Y104_CO6),
.O5(CLBLM_L_X10Y105_SLICE_X12Y105_CO5),
.O6(CLBLM_L_X10Y105_SLICE_X12Y105_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hb4783cf0c30fb478)
  ) CLBLM_L_X10Y105_SLICE_X12Y105_BLUT (
.I0(RIOB33_X105Y101_IOB_X1Y102_I),
.I1(LIOB33_X0Y101_IOB_X0Y102_I),
.I2(CLBLM_L_X10Y104_SLICE_X13Y104_CO6),
.I3(RIOB33_X105Y103_IOB_X1Y103_I),
.I4(CLBLM_L_X10Y105_SLICE_X12Y105_AO6),
.I5(CLBLM_L_X10Y103_SLICE_X12Y103_AO5),
.O5(CLBLM_L_X10Y105_SLICE_X12Y105_BO5),
.O6(CLBLM_L_X10Y105_SLICE_X12Y105_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h93939393ff13ff13)
  ) CLBLM_L_X10Y105_SLICE_X12Y105_ALUT (
.I0(RIOB33_X105Y103_IOB_X1Y103_I),
.I1(CLBLM_L_X10Y104_SLICE_X12Y104_BO6),
.I2(LIOB33_X0Y101_IOB_X0Y101_I),
.I3(CLBLM_L_X10Y104_SLICE_X12Y104_DO6),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X10Y105_SLICE_X12Y105_AO5),
.O6(CLBLM_L_X10Y105_SLICE_X12Y105_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h7b12ff5af330fff0)
  ) CLBLM_L_X10Y105_SLICE_X13Y105_DLUT (
.I0(LIOB33_X0Y103_IOB_X0Y104_I),
.I1(LIOB33_X0Y105_IOB_X0Y105_I),
.I2(CLBLM_L_X10Y105_SLICE_X12Y105_DO6),
.I3(CLBLM_L_X10Y105_SLICE_X13Y105_CO6),
.I4(RIOB33_X105Y101_IOB_X1Y102_I),
.I5(RIOB33_X105Y103_IOB_X1Y103_I),
.O5(CLBLM_L_X10Y105_SLICE_X13Y105_DO5),
.O6(CLBLM_L_X10Y105_SLICE_X13Y105_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h4dd4cffcdd44ffcc)
  ) CLBLM_L_X10Y105_SLICE_X13Y105_CLUT (
.I0(LIOB33_X0Y103_IOB_X0Y104_I),
.I1(CLBLM_L_X10Y102_SLICE_X12Y102_CO6),
.I2(RIOB33_X105Y103_IOB_X1Y103_I),
.I3(CLBLM_L_X10Y104_SLICE_X13Y104_CO6),
.I4(RIOB33_X105Y101_IOB_X1Y102_I),
.I5(LIOB33_X0Y101_IOB_X0Y102_I),
.O5(CLBLM_L_X10Y105_SLICE_X13Y105_CO5),
.O6(CLBLM_L_X10Y105_SLICE_X13Y105_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h6699966996699966)
  ) CLBLM_L_X10Y105_SLICE_X13Y105_BLUT (
.I0(CLBLM_L_X10Y104_SLICE_X13Y104_DO6),
.I1(CLBLM_R_X11Y105_SLICE_X14Y105_AO6),
.I2(CLBLM_L_X10Y104_SLICE_X13Y104_BO6),
.I3(CLBLM_R_X11Y104_SLICE_X14Y104_BO6),
.I4(CLBLM_L_X10Y105_SLICE_X13Y105_AO6),
.I5(CLBLM_L_X10Y102_SLICE_X12Y102_CO6),
.O5(CLBLM_L_X10Y105_SLICE_X13Y105_BO5),
.O6(CLBLM_L_X10Y105_SLICE_X13Y105_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h55ff55ff77777777)
  ) CLBLM_L_X10Y105_SLICE_X13Y105_ALUT (
.I0(RIOB33_X105Y101_IOB_X1Y102_I),
.I1(LIOB33_X0Y105_IOB_X0Y105_I),
.I2(1'b1),
.I3(LIOB33_X0Y103_IOB_X0Y104_I),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X10Y105_SLICE_X13Y105_AO5),
.O6(CLBLM_L_X10Y105_SLICE_X13Y105_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h6f06ff66cf0cffcc)
  ) CLBLM_L_X10Y106_SLICE_X12Y106_DLUT (
.I0(RIOB33_X105Y101_IOB_X1Y102_I),
.I1(CLBLM_L_X10Y106_SLICE_X13Y106_AO6),
.I2(LIOB33_X0Y107_IOB_X0Y107_I),
.I3(CLBLM_L_X8Y105_SLICE_X11Y105_CO6),
.I4(RIOB33_X105Y101_IOB_X1Y101_I),
.I5(LIOB33_X0Y105_IOB_X0Y106_I),
.O5(CLBLM_L_X10Y106_SLICE_X12Y106_DO5),
.O6(CLBLM_L_X10Y106_SLICE_X12Y106_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h7f07ff778f08ff88)
  ) CLBLM_L_X10Y106_SLICE_X12Y106_CLUT (
.I0(RIOB33_X105Y101_IOB_X1Y102_I),
.I1(LIOB33_X0Y103_IOB_X0Y104_I),
.I2(LIOB33_X0Y105_IOB_X0Y105_I),
.I3(CLBLM_L_X10Y103_SLICE_X12Y103_DO6),
.I4(RIOB33_X105Y101_IOB_X1Y101_I),
.I5(CLBLM_L_X10Y105_SLICE_X12Y105_BO6),
.O5(CLBLM_L_X10Y106_SLICE_X12Y106_CO5),
.O6(CLBLM_L_X10Y106_SLICE_X12Y106_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h87f078f0e13c1e3c)
  ) CLBLM_L_X10Y106_SLICE_X12Y106_BLUT (
.I0(RIOB33_X105Y101_IOB_X1Y101_I),
.I1(CLBLM_L_X10Y106_SLICE_X13Y106_BO6),
.I2(CLBLM_L_X10Y106_SLICE_X13Y106_AO6),
.I3(LIOB33_X0Y105_IOB_X0Y106_I),
.I4(RIOB33_X105Y101_IOB_X1Y102_I),
.I5(CLBLM_L_X10Y106_SLICE_X12Y106_CO6),
.O5(CLBLM_L_X10Y106_SLICE_X12Y106_BO5),
.O6(CLBLM_L_X10Y106_SLICE_X12Y106_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h7887878787787878)
  ) CLBLM_L_X10Y106_SLICE_X12Y106_ALUT (
.I0(RIOB33_X105Y101_IOB_X1Y101_I),
.I1(LIOB33_X0Y107_IOB_X0Y107_I),
.I2(CLBLM_L_X10Y106_SLICE_X13Y106_AO6),
.I3(LIOB33_X0Y105_IOB_X0Y106_I),
.I4(RIOB33_X105Y101_IOB_X1Y102_I),
.I5(CLBLM_L_X8Y105_SLICE_X11Y105_CO6),
.O5(CLBLM_L_X10Y106_SLICE_X12Y106_AO5),
.O6(CLBLM_L_X10Y106_SLICE_X12Y106_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h59a6a6599a65659a)
  ) CLBLM_L_X10Y106_SLICE_X13Y106_DLUT (
.I0(CLBLM_R_X11Y105_SLICE_X14Y105_BO6),
.I1(CLBLM_R_X11Y105_SLICE_X14Y105_CO6),
.I2(CLBLM_L_X10Y105_SLICE_X13Y105_AO5),
.I3(CLBLM_L_X10Y108_SLICE_X13Y108_AO5),
.I4(CLBLM_R_X11Y105_SLICE_X14Y105_AO5),
.I5(CLBLM_L_X10Y105_SLICE_X13Y105_CO6),
.O5(CLBLM_L_X10Y106_SLICE_X13Y106_DO5),
.O6(CLBLM_L_X10Y106_SLICE_X13Y106_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hffa5b721b721a500)
  ) CLBLM_L_X10Y106_SLICE_X13Y106_CLUT (
.I0(CLBLM_R_X11Y105_SLICE_X14Y105_BO6),
.I1(CLBLM_R_X11Y105_SLICE_X14Y105_CO6),
.I2(CLBLM_R_X11Y105_SLICE_X14Y105_AO5),
.I3(CLBLM_L_X10Y108_SLICE_X13Y108_AO5),
.I4(CLBLM_L_X10Y105_SLICE_X13Y105_AO5),
.I5(CLBLM_L_X10Y105_SLICE_X13Y105_CO6),
.O5(CLBLM_L_X10Y106_SLICE_X13Y106_CO5),
.O6(CLBLM_L_X10Y106_SLICE_X13Y106_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h69969966c33c33cc)
  ) CLBLM_L_X10Y106_SLICE_X13Y106_BLUT (
.I0(RIOB33_X105Y103_IOB_X1Y103_I),
.I1(CLBLM_L_X10Y105_SLICE_X12Y105_DO6),
.I2(RIOB33_X105Y101_IOB_X1Y102_I),
.I3(CLBLM_L_X10Y105_SLICE_X13Y105_CO6),
.I4(LIOB33_X0Y105_IOB_X0Y105_I),
.I5(LIOB33_X0Y103_IOB_X0Y104_I),
.O5(CLBLM_L_X10Y106_SLICE_X13Y106_BO5),
.O6(CLBLM_L_X10Y106_SLICE_X13Y106_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hd52ab9467f8013ec)
  ) CLBLM_L_X10Y106_SLICE_X13Y106_ALUT (
.I0(LIOB33_X0Y105_IOB_X0Y105_I),
.I1(CLBLM_R_X11Y105_SLICE_X14Y105_CO6),
.I2(RIOB33_X105Y101_IOB_X1Y102_I),
.I3(CLBLM_R_X11Y105_SLICE_X14Y105_BO6),
.I4(CLBLM_L_X10Y105_SLICE_X13Y105_CO6),
.I5(RIOB33_X105Y103_IOB_X1Y103_I),
.O5(CLBLM_L_X10Y106_SLICE_X13Y106_AO5),
.O6(CLBLM_L_X10Y106_SLICE_X13Y106_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X10Y107_SLICE_X12Y107_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X10Y107_SLICE_X12Y107_DO5),
.O6(CLBLM_L_X10Y107_SLICE_X12Y107_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h777f7fff377f7fff)
  ) CLBLM_L_X10Y107_SLICE_X12Y107_CLUT (
.I0(LIOB33_SING_X0Y100_IOB_X0Y100_I),
.I1(RIOB33_X105Y109_IOB_X1Y110_I),
.I2(RIOB33_X105Y111_IOB_X1Y111_I),
.I3(RIOB33_X105Y113_IOB_X1Y113_I),
.I4(LIOB33_X0Y101_IOB_X0Y101_I),
.I5(RIOB33_X105Y111_IOB_X1Y112_I),
.O5(CLBLM_L_X10Y107_SLICE_X12Y107_CO5),
.O6(CLBLM_L_X10Y107_SLICE_X12Y107_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h5fff7fff175f1fff)
  ) CLBLM_L_X10Y107_SLICE_X12Y107_BLUT (
.I0(RIOB33_X105Y109_IOB_X1Y110_I),
.I1(LIOB33_X0Y101_IOB_X0Y101_I),
.I2(LIOB33_X0Y101_IOB_X0Y102_I),
.I3(RIOB33_X105Y111_IOB_X1Y111_I),
.I4(LIOB33_X0Y103_IOB_X0Y104_I),
.I5(CLBLM_L_X10Y107_SLICE_X12Y107_CO6),
.O5(CLBLM_L_X10Y107_SLICE_X12Y107_BO5),
.O6(CLBLM_L_X10Y107_SLICE_X12Y107_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h2dd2d22db44b4bb4)
  ) CLBLM_L_X10Y107_SLICE_X12Y107_ALUT (
.I0(CLBLM_L_X10Y106_SLICE_X13Y106_DO6),
.I1(CLBLM_L_X10Y108_SLICE_X13Y108_BO6),
.I2(CLBLM_L_X10Y106_SLICE_X13Y106_CO6),
.I3(CLBLM_L_X10Y108_SLICE_X13Y108_AO6),
.I4(CLBLM_R_X11Y106_SLICE_X14Y106_AO6),
.I5(CLBLM_L_X8Y105_SLICE_X11Y105_CO6),
.O5(CLBLM_L_X10Y107_SLICE_X12Y107_AO5),
.O6(CLBLM_L_X10Y107_SLICE_X12Y107_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hb75f5f5fb75fdf5f)
  ) CLBLM_L_X10Y107_SLICE_X13Y107_DLUT (
.I0(LIOB33_X0Y101_IOB_X0Y101_I),
.I1(RIOB33_X105Y113_IOB_X1Y113_I),
.I2(RIOB33_X105Y111_IOB_X1Y111_I),
.I3(RIOB33_X105Y109_IOB_X1Y110_I),
.I4(LIOB33_SING_X0Y100_IOB_X0Y100_I),
.I5(RIOB33_X105Y111_IOB_X1Y112_I),
.O5(CLBLM_L_X10Y107_SLICE_X13Y107_DO5),
.O6(CLBLM_L_X10Y107_SLICE_X13Y107_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hb2df5dffa0dfdfff)
  ) CLBLM_L_X10Y107_SLICE_X13Y107_CLUT (
.I0(LIOB33_X0Y101_IOB_X0Y102_I),
.I1(CLBLM_L_X10Y107_SLICE_X12Y107_CO6),
.I2(RIOB33_X105Y109_IOB_X1Y110_I),
.I3(RIOB33_X105Y111_IOB_X1Y111_I),
.I4(LIOB33_X0Y103_IOB_X0Y104_I),
.I5(LIOB33_X0Y101_IOB_X0Y101_I),
.O5(CLBLM_L_X10Y107_SLICE_X13Y107_CO5),
.O6(CLBLM_L_X10Y107_SLICE_X13Y107_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'ha599699969aa5aaa)
  ) CLBLM_L_X10Y107_SLICE_X13Y107_BLUT (
.I0(CLBLM_L_X10Y108_SLICE_X13Y108_DO6),
.I1(CLBLM_R_X11Y107_SLICE_X15Y107_AO5),
.I2(LIOB33_X0Y107_IOB_X0Y107_I),
.I3(RIOB33_X105Y109_IOB_X1Y109_I),
.I4(LIOB33_X0Y105_IOB_X0Y106_I),
.I5(CLBLM_R_X11Y107_SLICE_X14Y107_BO6),
.O5(CLBLM_L_X10Y107_SLICE_X13Y107_BO5),
.O6(CLBLM_L_X10Y107_SLICE_X13Y107_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h6999c33396663ccc)
  ) CLBLM_L_X10Y107_SLICE_X13Y107_ALUT (
.I0(LIOB33_X0Y105_IOB_X0Y105_I),
.I1(CLBLM_R_X11Y107_SLICE_X15Y107_AO5),
.I2(RIOB33_X105Y109_IOB_X1Y109_I),
.I3(LIOB33_X0Y105_IOB_X0Y106_I),
.I4(RIOB33_X105Y109_IOB_X1Y110_I),
.I5(CLBLM_L_X10Y107_SLICE_X13Y107_CO6),
.O5(CLBLM_L_X10Y107_SLICE_X13Y107_AO5),
.O6(CLBLM_L_X10Y107_SLICE_X13Y107_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hecfe80c8b3fb2032)
  ) CLBLM_L_X10Y108_SLICE_X12Y108_DLUT (
.I0(CLBLM_L_X10Y106_SLICE_X12Y106_DO6),
.I1(CLBLM_L_X10Y108_SLICE_X13Y108_CO6),
.I2(CLBLM_L_X8Y107_SLICE_X11Y107_AO5),
.I3(CLBLM_L_X10Y108_SLICE_X12Y108_CO6),
.I4(CLBLM_L_X10Y109_SLICE_X13Y109_AO5),
.I5(CLBLM_R_X11Y110_SLICE_X15Y110_AO6),
.O5(CLBLM_L_X10Y108_SLICE_X12Y108_DO5),
.O6(CLBLM_L_X10Y108_SLICE_X12Y108_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h6996c33c996633cc)
  ) CLBLM_L_X10Y108_SLICE_X12Y108_CLUT (
.I0(LIOB33_X0Y105_IOB_X0Y106_I),
.I1(CLBLM_R_X11Y106_SLICE_X14Y106_DO6),
.I2(RIOB33_X105Y101_IOB_X1Y102_I),
.I3(CLBLM_L_X10Y106_SLICE_X13Y106_CO6),
.I4(RIOB33_X105Y103_IOB_X1Y103_I),
.I5(LIOB33_X0Y107_IOB_X0Y107_I),
.O5(CLBLM_L_X10Y108_SLICE_X12Y108_CO5),
.O6(CLBLM_L_X10Y108_SLICE_X12Y108_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hd278a50f5af0d278)
  ) CLBLM_L_X10Y108_SLICE_X12Y108_BLUT (
.I0(LIOB33_X0Y107_IOB_X0Y108_I),
.I1(RIOB33_X105Y101_IOB_X1Y101_I),
.I2(CLBLM_L_X10Y108_SLICE_X13Y108_CO6),
.I3(RIOB33_X105Y101_IOB_X1Y102_I),
.I4(CLBLM_L_X10Y106_SLICE_X12Y106_DO6),
.I5(CLBLM_L_X10Y108_SLICE_X12Y108_CO6),
.O5(CLBLM_L_X10Y108_SLICE_X12Y108_BO5),
.O6(CLBLM_L_X10Y108_SLICE_X12Y108_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h6996a55a5aa56996)
  ) CLBLM_L_X10Y108_SLICE_X12Y108_ALUT (
.I0(CLBLM_L_X10Y109_SLICE_X13Y109_AO5),
.I1(CLBLM_L_X8Y107_SLICE_X11Y107_AO5),
.I2(CLBLM_L_X10Y108_SLICE_X13Y108_CO6),
.I3(CLBLM_R_X11Y110_SLICE_X15Y110_AO6),
.I4(CLBLM_L_X10Y106_SLICE_X12Y106_DO6),
.I5(CLBLM_L_X10Y108_SLICE_X12Y108_CO6),
.O5(CLBLM_L_X10Y108_SLICE_X12Y108_AO5),
.O6(CLBLM_L_X10Y108_SLICE_X12Y108_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hb878888884b47888)
  ) CLBLM_L_X10Y108_SLICE_X13Y108_DLUT (
.I0(LIOB33_X0Y105_IOB_X0Y106_I),
.I1(RIOB33_X105Y109_IOB_X1Y110_I),
.I2(RIOB33_X105Y111_IOB_X1Y111_I),
.I3(LIOB33_X0Y103_IOB_X0Y104_I),
.I4(LIOB33_X0Y105_IOB_X0Y105_I),
.I5(CLBLM_L_X10Y107_SLICE_X12Y107_BO6),
.O5(CLBLM_L_X10Y108_SLICE_X13Y108_DO5),
.O6(CLBLM_L_X10Y108_SLICE_X13Y108_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h63c69c399c3963c6)
  ) CLBLM_L_X10Y108_SLICE_X13Y108_CLUT (
.I0(CLBLM_L_X10Y108_SLICE_X13Y108_AO6),
.I1(CLBLM_R_X11Y108_SLICE_X15Y108_BO6),
.I2(CLBLM_R_X11Y106_SLICE_X14Y106_AO6),
.I3(CLBLM_L_X10Y106_SLICE_X13Y106_CO6),
.I4(CLBLM_L_X10Y108_SLICE_X13Y108_BO5),
.I5(CLBLM_R_X11Y106_SLICE_X14Y106_CO6),
.O5(CLBLM_L_X10Y108_SLICE_X13Y108_CO5),
.O6(CLBLM_L_X10Y108_SLICE_X13Y108_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h3333ffff33ff33ff)
  ) CLBLM_L_X10Y108_SLICE_X13Y108_BLUT (
.I0(1'b1),
.I1(LIOB33_X0Y107_IOB_X0Y107_I),
.I2(1'b1),
.I3(RIOB33_X105Y103_IOB_X1Y103_I),
.I4(RIOB33_X105Y101_IOB_X1Y101_I),
.I5(1'b1),
.O5(CLBLM_L_X10Y108_SLICE_X13Y108_BO5),
.O6(CLBLM_L_X10Y108_SLICE_X13Y108_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h00ffffff0f0fffff)
  ) CLBLM_L_X10Y108_SLICE_X13Y108_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(LIOB33_X0Y105_IOB_X0Y106_I),
.I3(LIOB33_X0Y107_IOB_X0Y107_I),
.I4(RIOB33_X105Y101_IOB_X1Y102_I),
.I5(1'b1),
.O5(CLBLM_L_X10Y108_SLICE_X13Y108_AO5),
.O6(CLBLM_L_X10Y108_SLICE_X13Y108_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h2b2fbfff3fbfbfff)
  ) CLBLM_L_X10Y109_SLICE_X12Y109_DLUT (
.I0(CLBLM_L_X10Y107_SLICE_X12Y107_BO6),
.I1(RIOB33_X105Y109_IOB_X1Y110_I),
.I2(LIOB33_X0Y105_IOB_X0Y105_I),
.I3(LIOB33_X0Y105_IOB_X0Y106_I),
.I4(RIOB33_X105Y111_IOB_X1Y111_I),
.I5(LIOB33_X0Y103_IOB_X0Y104_I),
.O5(CLBLM_L_X10Y109_SLICE_X12Y109_DO5),
.O6(CLBLM_L_X10Y109_SLICE_X12Y109_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hc7bf63ffe3bf33ff)
  ) CLBLM_L_X10Y109_SLICE_X12Y109_CLUT (
.I0(CLBLM_L_X10Y107_SLICE_X12Y107_BO6),
.I1(LIOB33_X0Y105_IOB_X0Y106_I),
.I2(LIOB33_X0Y105_IOB_X0Y105_I),
.I3(RIOB33_X105Y111_IOB_X1Y111_I),
.I4(RIOB33_X105Y109_IOB_X1Y110_I),
.I5(LIOB33_X0Y103_IOB_X0Y104_I),
.O5(CLBLM_L_X10Y109_SLICE_X12Y109_CO5),
.O6(CLBLM_L_X10Y109_SLICE_X12Y109_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h6996c33c996633cc)
  ) CLBLM_L_X10Y109_SLICE_X12Y109_BLUT (
.I0(LIOB33_X0Y107_IOB_X0Y108_I),
.I1(CLBLM_L_X10Y106_SLICE_X12Y106_DO6),
.I2(RIOB33_X105Y101_IOB_X1Y102_I),
.I3(CLBLM_L_X10Y109_SLICE_X13Y109_CO6),
.I4(RIOB33_X105Y101_IOB_X1Y101_I),
.I5(LIOB33_X0Y107_IOB_X0Y107_I),
.O5(CLBLM_L_X10Y109_SLICE_X12Y109_BO5),
.O6(CLBLM_L_X10Y109_SLICE_X12Y109_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h4dd4cffcdd44ffcc)
  ) CLBLM_L_X10Y109_SLICE_X12Y109_ALUT (
.I0(LIOB33_X0Y107_IOB_X0Y108_I),
.I1(CLBLM_L_X10Y106_SLICE_X12Y106_DO6),
.I2(RIOB33_X105Y101_IOB_X1Y102_I),
.I3(CLBLM_L_X10Y109_SLICE_X13Y109_CO6),
.I4(RIOB33_X105Y101_IOB_X1Y101_I),
.I5(LIOB33_X0Y107_IOB_X0Y107_I),
.O5(CLBLM_L_X10Y109_SLICE_X12Y109_AO5),
.O6(CLBLM_L_X10Y109_SLICE_X12Y109_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h9a6a6a6a959a956a)
  ) CLBLM_L_X10Y109_SLICE_X13Y109_DLUT (
.I0(CLBLM_R_X11Y109_SLICE_X15Y109_AO6),
.I1(RIOB33_X105Y103_IOB_X1Y103_I),
.I2(LIOB33_X0Y107_IOB_X0Y108_I),
.I3(CLBLM_R_X11Y109_SLICE_X14Y109_CO6),
.I4(RIOB33_X105Y101_IOB_X1Y102_I),
.I5(CLBLM_L_X10Y109_SLICE_X13Y109_BO6),
.O5(CLBLM_L_X10Y109_SLICE_X13Y109_DO5),
.O6(CLBLM_L_X10Y109_SLICE_X13Y109_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h9cc339cc63c3c6cc)
  ) CLBLM_L_X10Y109_SLICE_X13Y109_CLUT (
.I0(RIOB33_X105Y101_IOB_X1Y102_I),
.I1(CLBLM_R_X11Y106_SLICE_X14Y106_DO6),
.I2(CLBLM_L_X10Y105_SLICE_X13Y105_DO6),
.I3(LIOB33_X0Y105_IOB_X0Y106_I),
.I4(CLBLM_R_X11Y108_SLICE_X14Y108_DO6),
.I5(RIOB33_X105Y103_IOB_X1Y103_I),
.O5(CLBLM_L_X10Y109_SLICE_X13Y109_CO5),
.O6(CLBLM_L_X10Y109_SLICE_X13Y109_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h7dff143cddff44cc)
  ) CLBLM_L_X10Y109_SLICE_X13Y109_BLUT (
.I0(RIOB33_X105Y101_IOB_X1Y102_I),
.I1(CLBLM_R_X11Y106_SLICE_X14Y106_DO6),
.I2(RIOB33_X105Y103_IOB_X1Y103_I),
.I3(LIOB33_X0Y107_IOB_X0Y107_I),
.I4(CLBLM_L_X10Y106_SLICE_X13Y106_CO6),
.I5(LIOB33_X0Y105_IOB_X0Y106_I),
.O5(CLBLM_L_X10Y109_SLICE_X13Y109_BO5),
.O6(CLBLM_L_X10Y109_SLICE_X13Y109_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h00ffffff0fff0fff)
  ) CLBLM_L_X10Y109_SLICE_X13Y109_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(RIOB33_X105Y101_IOB_X1Y101_I),
.I3(LIOB33_X0Y109_IOB_X0Y109_I),
.I4(RIOB33_X105Y101_IOB_X1Y102_I),
.I5(1'b1),
.O5(CLBLM_L_X10Y109_SLICE_X13Y109_AO5),
.O6(CLBLM_L_X10Y109_SLICE_X13Y109_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hb4c3780f3cb4f078)
  ) CLBLM_L_X10Y110_SLICE_X12Y110_DLUT (
.I0(RIOB33_X105Y101_IOB_X1Y102_I),
.I1(LIOB33_X0Y109_IOB_X0Y109_I),
.I2(CLBLM_R_X11Y110_SLICE_X14Y110_CO6),
.I3(CLBLM_L_X10Y110_SLICE_X12Y110_CO6),
.I4(RIOB33_X105Y103_IOB_X1Y103_I),
.I5(CLBLM_L_X12Y110_SLICE_X16Y110_BO6),
.O5(CLBLM_L_X10Y110_SLICE_X12Y110_DO5),
.O6(CLBLM_L_X10Y110_SLICE_X12Y110_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h7fdfff5f134c5f00)
  ) CLBLM_L_X10Y110_SLICE_X12Y110_CLUT (
.I0(RIOB33_X105Y101_IOB_X1Y102_I),
.I1(LIOB33_X0Y107_IOB_X0Y107_I),
.I2(LIOB33_X0Y107_IOB_X0Y108_I),
.I3(CLBLM_R_X11Y108_SLICE_X14Y108_AO6),
.I4(RIOB33_X105Y103_IOB_X1Y103_I),
.I5(CLBLM_L_X10Y109_SLICE_X13Y109_BO6),
.O5(CLBLM_L_X10Y110_SLICE_X12Y110_CO5),
.O6(CLBLM_L_X10Y110_SLICE_X12Y110_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hb4cc2dff4b33d200)
  ) CLBLM_L_X10Y110_SLICE_X12Y110_BLUT (
.I0(RIOB33_X105Y101_IOB_X1Y101_I),
.I1(CLBLM_L_X10Y109_SLICE_X12Y109_AO6),
.I2(RIOB33_X105Y101_IOB_X1Y102_I),
.I3(LIOB33_X0Y109_IOB_X0Y109_I),
.I4(CLBLM_L_X10Y110_SLICE_X12Y110_AO6),
.I5(CLBLM_L_X10Y109_SLICE_X13Y109_DO6),
.O5(CLBLM_L_X10Y110_SLICE_X12Y110_BO5),
.O6(CLBLM_L_X10Y110_SLICE_X12Y110_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h6996c33c996633cc)
  ) CLBLM_L_X10Y110_SLICE_X12Y110_ALUT (
.I0(LIOB33_X0Y107_IOB_X0Y108_I),
.I1(CLBLM_R_X11Y108_SLICE_X14Y108_AO6),
.I2(RIOB33_X105Y103_IOB_X1Y103_I),
.I3(CLBLM_L_X10Y109_SLICE_X13Y109_BO6),
.I4(RIOB33_X105Y101_IOB_X1Y102_I),
.I5(LIOB33_X0Y107_IOB_X0Y107_I),
.O5(CLBLM_L_X10Y110_SLICE_X12Y110_AO5),
.O6(CLBLM_L_X10Y110_SLICE_X12Y110_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h020baaff2fbfffff)
  ) CLBLM_L_X10Y110_SLICE_X13Y110_DLUT (
.I0(CLBLM_L_X12Y108_SLICE_X16Y108_BO6),
.I1(LIOB33_X0Y107_IOB_X0Y107_I),
.I2(LIOB33_X0Y107_IOB_X0Y108_I),
.I3(CLBLM_L_X10Y107_SLICE_X13Y107_AO6),
.I4(RIOB33_X105Y107_IOB_X1Y108_I),
.I5(CLBLM_L_X10Y107_SLICE_X13Y107_BO6),
.O5(CLBLM_L_X10Y110_SLICE_X13Y110_DO5),
.O6(CLBLM_L_X10Y110_SLICE_X13Y110_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h3c9696c3c369693c)
  ) CLBLM_L_X10Y110_SLICE_X13Y110_CLUT (
.I0(CLBLM_R_X11Y110_SLICE_X14Y110_BO6),
.I1(CLBLM_R_X11Y110_SLICE_X14Y110_AO5),
.I2(CLBLM_L_X10Y111_SLICE_X13Y111_BO6),
.I3(CLBLM_L_X10Y110_SLICE_X13Y110_AO5),
.I4(CLBLM_R_X11Y109_SLICE_X14Y109_DO6),
.I5(CLBLM_R_X11Y110_SLICE_X14Y110_DO6),
.O5(CLBLM_L_X10Y110_SLICE_X13Y110_CO5),
.O6(CLBLM_L_X10Y110_SLICE_X13Y110_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h693cc36996c33c96)
  ) CLBLM_L_X10Y110_SLICE_X13Y110_BLUT (
.I0(CLBLM_L_X10Y108_SLICE_X12Y108_DO6),
.I1(CLBLM_R_X11Y110_SLICE_X14Y110_BO6),
.I2(CLBLM_R_X11Y109_SLICE_X14Y109_DO6),
.I3(CLBLM_R_X11Y109_SLICE_X14Y109_BO6),
.I4(CLBLM_L_X10Y110_SLICE_X13Y110_AO6),
.I5(CLBLM_L_X10Y110_SLICE_X13Y110_AO5),
.O5(CLBLM_L_X10Y110_SLICE_X13Y110_BO5),
.O6(CLBLM_L_X10Y110_SLICE_X13Y110_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h55ff55ff5555ffff)
  ) CLBLM_L_X10Y110_SLICE_X13Y110_ALUT (
.I0(LIOB33_X0Y109_IOB_X0Y110_I),
.I1(1'b1),
.I2(1'b1),
.I3(RIOB33_X105Y101_IOB_X1Y101_I),
.I4(RIOB33_X105Y101_IOB_X1Y102_I),
.I5(1'b1),
.O5(CLBLM_L_X10Y110_SLICE_X13Y110_AO5),
.O6(CLBLM_L_X10Y110_SLICE_X13Y110_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h2bb2bb22affaffaa)
  ) CLBLM_L_X10Y111_SLICE_X12Y111_DLUT (
.I0(CLBLM_R_X11Y111_SLICE_X14Y111_BO6),
.I1(RIOB33_X105Y105_IOB_X1Y105_I),
.I2(RIOB33_X105Y107_IOB_X1Y107_I),
.I3(CLBLM_L_X10Y112_SLICE_X13Y112_AO5),
.I4(LIOB33_X0Y107_IOB_X0Y108_I),
.I5(LIOB33_X0Y109_IOB_X0Y109_I),
.O5(CLBLM_L_X10Y111_SLICE_X12Y111_DO5),
.O6(CLBLM_L_X10Y111_SLICE_X12Y111_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h37077f077f377f7f)
  ) CLBLM_L_X10Y111_SLICE_X12Y111_CLUT (
.I0(LIOB33_X0Y109_IOB_X0Y110_I),
.I1(RIOB33_X105Y103_IOB_X1Y103_I),
.I2(CLBLM_L_X10Y111_SLICE_X13Y111_BO6),
.I3(CLBLM_L_X12Y110_SLICE_X16Y110_CO6),
.I4(LIOB33_X0Y109_IOB_X0Y109_I),
.I5(CLBLM_R_X11Y111_SLICE_X14Y111_CO6),
.O5(CLBLM_L_X10Y111_SLICE_X12Y111_CO5),
.O6(CLBLM_L_X10Y111_SLICE_X12Y111_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h7887878787787878)
  ) CLBLM_L_X10Y111_SLICE_X12Y111_BLUT (
.I0(RIOB33_X105Y105_IOB_X1Y105_I),
.I1(LIOB33_X0Y109_IOB_X0Y109_I),
.I2(CLBLM_R_X11Y111_SLICE_X14Y111_BO6),
.I3(LIOB33_X0Y107_IOB_X0Y108_I),
.I4(RIOB33_X105Y107_IOB_X1Y107_I),
.I5(CLBLM_L_X10Y112_SLICE_X13Y112_AO5),
.O5(CLBLM_L_X10Y111_SLICE_X12Y111_BO5),
.O6(CLBLM_L_X10Y111_SLICE_X12Y111_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h963cccccc39633cc)
  ) CLBLM_L_X10Y111_SLICE_X12Y111_ALUT (
.I0(LIOB33_X0Y109_IOB_X0Y109_I),
.I1(CLBLM_L_X10Y111_SLICE_X13Y111_BO6),
.I2(LIOB33_X0Y109_IOB_X0Y110_I),
.I3(CLBLM_R_X11Y111_SLICE_X14Y111_CO6),
.I4(RIOB33_X105Y103_IOB_X1Y103_I),
.I5(CLBLM_L_X12Y110_SLICE_X16Y110_CO6),
.O5(CLBLM_L_X10Y111_SLICE_X12Y111_AO5),
.O6(CLBLM_L_X10Y111_SLICE_X12Y111_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hd7b1284e5f93a06c)
  ) CLBLM_L_X10Y111_SLICE_X13Y111_DLUT (
.I0(LIOB33_X0Y107_IOB_X0Y108_I),
.I1(CLBLM_R_X11Y109_SLICE_X15Y109_CO6),
.I2(RIOB33_X105Y105_IOB_X1Y105_I),
.I3(CLBLM_R_X11Y111_SLICE_X15Y111_DO6),
.I4(CLBLM_L_X12Y110_SLICE_X16Y110_DO6),
.I5(RIOB33_X105Y103_IOB_X1Y104_I),
.O5(CLBLM_L_X10Y111_SLICE_X13Y111_DO5),
.O6(CLBLM_L_X10Y111_SLICE_X13Y111_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h9fa0605f5f9fa060)
  ) CLBLM_L_X10Y111_SLICE_X13Y111_CLUT (
.I0(RIOB33_X105Y103_IOB_X1Y104_I),
.I1(RIOB33_X105Y103_IOB_X1Y103_I),
.I2(LIOB33_X0Y109_IOB_X0Y109_I),
.I3(CLBLM_L_X12Y110_SLICE_X16Y110_CO6),
.I4(CLBLM_L_X10Y111_SLICE_X13Y111_DO6),
.I5(CLBLM_R_X11Y111_SLICE_X14Y111_CO6),
.O5(CLBLM_L_X10Y111_SLICE_X13Y111_CO5),
.O6(CLBLM_L_X10Y111_SLICE_X13Y111_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h718e8e718e71718e)
  ) CLBLM_L_X10Y111_SLICE_X13Y111_BLUT (
.I0(CLBLM_R_X11Y111_SLICE_X15Y111_DO6),
.I1(CLBLM_R_X11Y110_SLICE_X15Y110_AO5),
.I2(CLBLM_R_X11Y109_SLICE_X15Y109_CO6),
.I3(CLBLM_R_X11Y111_SLICE_X14Y111_AO6),
.I4(CLBLM_L_X10Y111_SLICE_X13Y111_AO6),
.I5(CLBLM_L_X12Y110_SLICE_X16Y110_DO6),
.O5(CLBLM_L_X10Y111_SLICE_X13Y111_BO5),
.O6(CLBLM_L_X10Y111_SLICE_X13Y111_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h777777775f5f5f5f)
  ) CLBLM_L_X10Y111_SLICE_X13Y111_ALUT (
.I0(RIOB33_X105Y105_IOB_X1Y105_I),
.I1(LIOB33_X0Y107_IOB_X0Y108_I),
.I2(LIOB33_X0Y109_IOB_X0Y110_I),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X10Y111_SLICE_X13Y111_AO5),
.O6(CLBLM_L_X10Y111_SLICE_X13Y111_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X10Y112_SLICE_X12Y112_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X10Y112_SLICE_X12Y112_DO5),
.O6(CLBLM_L_X10Y112_SLICE_X12Y112_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X10Y112_SLICE_X12Y112_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X10Y112_SLICE_X12Y112_CO5),
.O6(CLBLM_L_X10Y112_SLICE_X12Y112_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h1f077f575f17ff77)
  ) CLBLM_L_X10Y112_SLICE_X12Y112_BLUT (
.I0(CLBLM_R_X11Y110_SLICE_X14Y110_BO6),
.I1(CLBLM_L_X12Y110_SLICE_X16Y110_BO6),
.I2(RIOB33_X105Y101_IOB_X1Y102_I),
.I3(CLBLM_L_X10Y110_SLICE_X12Y110_CO6),
.I4(LIOB33_X0Y109_IOB_X0Y110_I),
.I5(LIOB33_X0Y109_IOB_X0Y109_I),
.O5(CLBLM_L_X10Y112_SLICE_X12Y112_BO5),
.O6(CLBLM_L_X10Y112_SLICE_X12Y112_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h9a5a6aaaa59a556a)
  ) CLBLM_L_X10Y112_SLICE_X12Y112_ALUT (
.I0(CLBLM_R_X11Y110_SLICE_X14Y110_BO6),
.I1(LIOB33_X0Y109_IOB_X0Y109_I),
.I2(RIOB33_X105Y101_IOB_X1Y102_I),
.I3(CLBLM_L_X12Y110_SLICE_X16Y110_BO6),
.I4(LIOB33_X0Y109_IOB_X0Y110_I),
.I5(CLBLM_L_X10Y110_SLICE_X12Y110_CO6),
.O5(CLBLM_L_X10Y112_SLICE_X12Y112_AO5),
.O6(CLBLM_L_X10Y112_SLICE_X12Y112_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hd24bbbbb2db44444)
  ) CLBLM_L_X10Y112_SLICE_X13Y112_DLUT (
.I0(CLBLM_L_X12Y108_SLICE_X16Y108_BO6),
.I1(CLBLM_L_X10Y107_SLICE_X13Y107_AO6),
.I2(LIOB33_X0Y107_IOB_X0Y108_I),
.I3(LIOB33_X0Y107_IOB_X0Y107_I),
.I4(RIOB33_X105Y107_IOB_X1Y108_I),
.I5(CLBLM_L_X10Y107_SLICE_X13Y107_BO6),
.O5(CLBLM_L_X10Y112_SLICE_X13Y112_DO5),
.O6(CLBLM_L_X10Y112_SLICE_X13Y112_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hbd3942c671f58e0a)
  ) CLBLM_L_X10Y112_SLICE_X13Y112_CLUT (
.I0(CLBLM_L_X10Y112_SLICE_X13Y112_AO6),
.I1(RIOB33_X105Y107_IOB_X1Y107_I),
.I2(CLBLM_R_X11Y110_SLICE_X15Y110_CO6),
.I3(LIOB33_X0Y107_IOB_X0Y108_I),
.I4(CLBLM_L_X10Y112_SLICE_X13Y112_DO6),
.I5(LIOB33_X0Y109_IOB_X0Y109_I),
.O5(CLBLM_L_X10Y112_SLICE_X13Y112_CO5),
.O6(CLBLM_L_X10Y112_SLICE_X13Y112_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h377f7f7f1515377f)
  ) CLBLM_L_X10Y112_SLICE_X13Y112_BLUT (
.I0(CLBLM_L_X10Y112_SLICE_X13Y112_DO6),
.I1(RIOB33_X105Y107_IOB_X1Y107_I),
.I2(LIOB33_X0Y109_IOB_X0Y109_I),
.I3(LIOB33_X0Y107_IOB_X0Y108_I),
.I4(CLBLM_L_X10Y112_SLICE_X13Y112_AO6),
.I5(CLBLM_R_X11Y110_SLICE_X15Y110_CO6),
.O5(CLBLM_L_X10Y112_SLICE_X13Y112_BO5),
.O6(CLBLM_L_X10Y112_SLICE_X13Y112_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h3cc3cc3396696699)
  ) CLBLM_L_X10Y112_SLICE_X13Y112_ALUT (
.I0(CLBLM_R_X11Y110_SLICE_X15Y110_CO6),
.I1(CLBLM_L_X10Y107_SLICE_X13Y107_AO6),
.I2(RIOB33_X105Y107_IOB_X1Y108_I),
.I3(CLBLM_L_X12Y108_SLICE_X16Y108_BO6),
.I4(LIOB33_X0Y107_IOB_X0Y107_I),
.I5(1'b1),
.O5(CLBLM_L_X10Y112_SLICE_X13Y112_AO5),
.O6(CLBLM_L_X10Y112_SLICE_X13Y112_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hfaa0fea8f550fd54)
  ) CLBLM_L_X12Y104_SLICE_X16Y104_DLUT (
.I0(CLBLM_L_X12Y106_SLICE_X17Y106_AO6),
.I1(CLBLM_L_X12Y104_SLICE_X16Y104_AO6),
.I2(CLBLM_L_X12Y104_SLICE_X16Y104_CO6),
.I3(CLBLM_L_X12Y104_SLICE_X16Y104_AO5),
.I4(CLBLM_R_X11Y104_SLICE_X15Y104_CO6),
.I5(CLBLM_L_X12Y105_SLICE_X16Y105_BO6),
.O5(CLBLM_L_X12Y104_SLICE_X16Y104_DO5),
.O6(CLBLM_L_X12Y104_SLICE_X16Y104_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h206c00aa22660000)
  ) CLBLM_L_X12Y104_SLICE_X16Y104_CLUT (
.I0(RIOB33_X105Y113_IOB_X1Y113_I),
.I1(LIOB33_SING_X0Y100_IOB_X0Y100_I),
.I2(RIOB33_X105Y111_IOB_X1Y112_I),
.I3(RIOB33_X105Y105_IOB_X1Y105_I),
.I4(RIOB33_X105Y107_IOB_X1Y107_I),
.I5(RIOB33_X105Y107_IOB_X1Y108_I),
.O5(CLBLM_L_X12Y104_SLICE_X16Y104_CO5),
.O6(CLBLM_L_X12Y104_SLICE_X16Y104_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h3c963cc3c369c33c)
  ) CLBLM_L_X12Y104_SLICE_X16Y104_BLUT (
.I0(CLBLM_R_X11Y104_SLICE_X15Y104_CO6),
.I1(CLBLM_L_X12Y106_SLICE_X17Y106_AO6),
.I2(CLBLM_L_X12Y105_SLICE_X16Y105_BO6),
.I3(CLBLM_L_X12Y104_SLICE_X16Y104_CO6),
.I4(CLBLM_L_X12Y104_SLICE_X16Y104_AO6),
.I5(CLBLM_L_X12Y104_SLICE_X16Y104_AO5),
.O5(CLBLM_L_X12Y104_SLICE_X16Y104_BO5),
.O6(CLBLM_L_X12Y104_SLICE_X16Y104_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h33ff33ff3f3f3f3f)
  ) CLBLM_L_X12Y104_SLICE_X16Y104_ALUT (
.I0(1'b1),
.I1(RIOB33_X105Y105_IOB_X1Y105_I),
.I2(LIOB33_X0Y101_IOB_X0Y102_I),
.I3(LIOB33_X0Y101_IOB_X0Y101_I),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X12Y104_SLICE_X16Y104_AO5),
.O6(CLBLM_L_X12Y104_SLICE_X16Y104_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X12Y104_SLICE_X17Y104_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X12Y104_SLICE_X17Y104_DO5),
.O6(CLBLM_L_X12Y104_SLICE_X17Y104_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X12Y104_SLICE_X17Y104_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X12Y104_SLICE_X17Y104_CO5),
.O6(CLBLM_L_X12Y104_SLICE_X17Y104_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X12Y104_SLICE_X17Y104_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X12Y104_SLICE_X17Y104_BO5),
.O6(CLBLM_L_X12Y104_SLICE_X17Y104_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X12Y104_SLICE_X17Y104_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X12Y104_SLICE_X17Y104_AO5),
.O6(CLBLM_L_X12Y104_SLICE_X17Y104_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h078805aa0a0a0000)
  ) CLBLM_L_X12Y105_SLICE_X16Y105_DLUT (
.I0(RIOB33_X105Y113_IOB_X1Y113_I),
.I1(RIOB33_X105Y111_IOB_X1Y112_I),
.I2(RIOB33_X105Y107_IOB_X1Y107_I),
.I3(LIOB33_SING_X0Y100_IOB_X0Y100_I),
.I4(RIOB33_X105Y109_IOB_X1Y109_I),
.I5(RIOB33_X105Y107_IOB_X1Y108_I),
.O5(CLBLM_L_X12Y105_SLICE_X16Y105_DO5),
.O6(CLBLM_L_X12Y105_SLICE_X16Y105_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h6663afaf999c5050)
  ) CLBLM_L_X12Y105_SLICE_X16Y105_CLUT (
.I0(CLBLM_L_X12Y104_SLICE_X16Y104_CO6),
.I1(RIOB33_X105Y107_IOB_X1Y107_I),
.I2(CLBLM_R_X11Y104_SLICE_X15Y104_CO6),
.I3(RIOB33_X105Y105_IOB_X1Y105_I),
.I4(LIOB33_X0Y101_IOB_X0Y101_I),
.I5(CLBLM_L_X12Y105_SLICE_X16Y105_BO6),
.O5(CLBLM_L_X12Y105_SLICE_X16Y105_CO5),
.O6(CLBLM_L_X12Y105_SLICE_X16Y105_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h06f533006666cc00)
  ) CLBLM_L_X12Y105_SLICE_X16Y105_BLUT (
.I0(RIOB33_X105Y109_IOB_X1Y109_I),
.I1(RIOB33_X105Y107_IOB_X1Y107_I),
.I2(RIOB33_X105Y111_IOB_X1Y112_I),
.I3(LIOB33_SING_X0Y100_IOB_X0Y100_I),
.I4(RIOB33_X105Y113_IOB_X1Y113_I),
.I5(RIOB33_X105Y107_IOB_X1Y108_I),
.O5(CLBLM_L_X12Y105_SLICE_X16Y105_BO5),
.O6(CLBLM_L_X12Y105_SLICE_X16Y105_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f0f3ffcc0033ff)
  ) CLBLM_L_X12Y105_SLICE_X16Y105_ALUT (
.I0(1'b1),
.I1(RIOB33_X105Y105_IOB_X1Y105_I),
.I2(CLBLM_L_X12Y104_SLICE_X16Y104_CO6),
.I3(LIOB33_X0Y101_IOB_X0Y101_I),
.I4(CLBLM_R_X11Y104_SLICE_X15Y104_CO6),
.I5(1'b1),
.O5(CLBLM_L_X12Y105_SLICE_X16Y105_AO5),
.O6(CLBLM_L_X12Y105_SLICE_X16Y105_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h9931111199395f5f)
  ) CLBLM_L_X12Y105_SLICE_X17Y105_DLUT (
.I0(RIOB33_X105Y113_IOB_X1Y113_I),
.I1(LIOB33_SING_X0Y100_IOB_X0Y100_I),
.I2(RIOB33_X105Y111_IOB_X1Y111_I),
.I3(RIOB33_X105Y111_IOB_X1Y112_I),
.I4(RIOB33_X105Y109_IOB_X1Y110_I),
.I5(RIOB33_X105Y109_IOB_X1Y109_I),
.O5(CLBLM_L_X12Y105_SLICE_X17Y105_DO5),
.O6(CLBLM_L_X12Y105_SLICE_X17Y105_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hafd050f05f20a000)
  ) CLBLM_L_X12Y105_SLICE_X17Y105_CLUT (
.I0(RIOB33_X105Y113_IOB_X1Y113_I),
.I1(RIOB33_X105Y111_IOB_X1Y112_I),
.I2(RIOB33_X105Y109_IOB_X1Y110_I),
.I3(LIOB33_SING_X0Y100_IOB_X0Y100_I),
.I4(RIOB33_X105Y111_IOB_X1Y111_I),
.I5(LIOB33_X0Y101_IOB_X0Y101_I),
.O5(CLBLM_L_X12Y105_SLICE_X17Y105_CO5),
.O6(CLBLM_L_X12Y105_SLICE_X17Y105_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h5aaa4bffa555b400)
  ) CLBLM_L_X12Y105_SLICE_X17Y105_BLUT (
.I0(CLBLM_L_X12Y105_SLICE_X17Y105_DO6),
.I1(LIOB33_X0Y101_IOB_X0Y101_I),
.I2(LIOB33_X0Y101_IOB_X0Y102_I),
.I3(RIOB33_X105Y109_IOB_X1Y109_I),
.I4(CLBLM_R_X13Y105_SLICE_X18Y105_AO6),
.I5(CLBLM_L_X12Y105_SLICE_X17Y105_CO6),
.O5(CLBLM_L_X12Y105_SLICE_X17Y105_BO5),
.O6(CLBLM_L_X12Y105_SLICE_X17Y105_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0a0bbbbbafbfffff)
  ) CLBLM_L_X12Y105_SLICE_X17Y105_ALUT (
.I0(CLBLM_L_X12Y105_SLICE_X17Y105_DO6),
.I1(CLBLM_R_X13Y105_SLICE_X18Y105_AO6),
.I2(LIOB33_X0Y101_IOB_X0Y102_I),
.I3(LIOB33_X0Y101_IOB_X0Y101_I),
.I4(RIOB33_X105Y109_IOB_X1Y109_I),
.I5(CLBLM_L_X12Y105_SLICE_X17Y105_CO6),
.O5(CLBLM_L_X12Y105_SLICE_X17Y105_AO5),
.O6(CLBLM_L_X12Y105_SLICE_X17Y105_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h787887877878b478)
  ) CLBLM_L_X12Y106_SLICE_X16Y106_DLUT (
.I0(RIOB33_X105Y107_IOB_X1Y108_I),
.I1(LIOB33_X0Y101_IOB_X0Y101_I),
.I2(CLBLM_R_X13Y106_SLICE_X19Y106_CO6),
.I3(RIOB33_X105Y107_IOB_X1Y107_I),
.I4(CLBLM_L_X12Y105_SLICE_X16Y105_DO6),
.I5(CLBLM_L_X12Y105_SLICE_X16Y105_BO6),
.O5(CLBLM_L_X12Y106_SLICE_X16Y106_DO5),
.O6(CLBLM_L_X12Y106_SLICE_X16Y106_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hda2a25d54fbfb040)
  ) CLBLM_L_X12Y106_SLICE_X16Y106_CLUT (
.I0(CLBLM_L_X12Y105_SLICE_X16Y105_AO6),
.I1(RIOB33_X105Y105_IOB_X1Y105_I),
.I2(LIOB33_X0Y101_IOB_X0Y102_I),
.I3(RIOB33_X105Y107_IOB_X1Y107_I),
.I4(CLBLM_L_X12Y106_SLICE_X16Y106_DO6),
.I5(CLBLM_L_X12Y106_SLICE_X16Y106_BO6),
.O5(CLBLM_L_X12Y106_SLICE_X16Y106_CO5),
.O6(CLBLM_L_X12Y106_SLICE_X16Y106_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hcc333333aabbbbbb)
  ) CLBLM_L_X12Y106_SLICE_X16Y106_BLUT (
.I0(CLBLM_L_X12Y105_SLICE_X16Y105_DO6),
.I1(CLBLM_L_X12Y105_SLICE_X16Y105_BO6),
.I2(1'b1),
.I3(RIOB33_X105Y107_IOB_X1Y107_I),
.I4(LIOB33_X0Y101_IOB_X0Y101_I),
.I5(1'b1),
.O5(CLBLM_L_X12Y106_SLICE_X16Y106_BO5),
.O6(CLBLM_L_X12Y106_SLICE_X16Y106_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h3333ffff3f3f3f3f)
  ) CLBLM_L_X12Y106_SLICE_X16Y106_ALUT (
.I0(1'b1),
.I1(RIOB33_X105Y107_IOB_X1Y108_I),
.I2(LIOB33_X0Y103_IOB_X0Y104_I),
.I3(1'b1),
.I4(LIOB33_X0Y101_IOB_X0Y101_I),
.I5(1'b1),
.O5(CLBLM_L_X12Y106_SLICE_X16Y106_AO5),
.O6(CLBLM_L_X12Y106_SLICE_X16Y106_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hfcc0f330fec8fb32)
  ) CLBLM_L_X12Y106_SLICE_X17Y106_DLUT (
.I0(CLBLM_L_X12Y106_SLICE_X17Y106_AO6),
.I1(CLBLM_L_X12Y106_SLICE_X16Y106_AO6),
.I2(CLBLM_L_X12Y105_SLICE_X16Y105_DO6),
.I3(CLBLM_L_X12Y106_SLICE_X17Y106_AO5),
.I4(CLBLM_R_X13Y106_SLICE_X19Y106_CO6),
.I5(CLBLM_L_X12Y105_SLICE_X16Y105_BO6),
.O5(CLBLM_L_X12Y106_SLICE_X17Y106_DO5),
.O6(CLBLM_L_X12Y106_SLICE_X17Y106_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h9a65f00f59a6ff00)
  ) CLBLM_L_X12Y106_SLICE_X17Y106_CLUT (
.I0(RIOB33_X105Y107_IOB_X1Y108_I),
.I1(RIOB33_X105Y107_IOB_X1Y107_I),
.I2(CLBLM_L_X12Y106_SLICE_X16Y106_BO5),
.I3(CLBLM_R_X13Y106_SLICE_X18Y106_DO6),
.I4(LIOB33_X0Y101_IOB_X0Y102_I),
.I5(CLBLM_R_X13Y106_SLICE_X19Y106_AO6),
.O5(CLBLM_L_X12Y106_SLICE_X17Y106_CO5),
.O6(CLBLM_L_X12Y106_SLICE_X17Y106_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h695a696996a59696)
  ) CLBLM_L_X12Y106_SLICE_X17Y106_BLUT (
.I0(CLBLM_R_X13Y106_SLICE_X19Y106_CO6),
.I1(CLBLM_L_X12Y105_SLICE_X16Y105_DO6),
.I2(CLBLM_L_X12Y106_SLICE_X16Y106_AO6),
.I3(CLBLM_L_X12Y105_SLICE_X16Y105_BO6),
.I4(CLBLM_L_X12Y106_SLICE_X17Y106_AO6),
.I5(CLBLM_L_X12Y106_SLICE_X17Y106_AO5),
.O5(CLBLM_L_X12Y106_SLICE_X17Y106_BO5),
.O6(CLBLM_L_X12Y106_SLICE_X17Y106_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h3f3f3f3f77777777)
  ) CLBLM_L_X12Y106_SLICE_X17Y106_ALUT (
.I0(LIOB33_X0Y101_IOB_X0Y102_I),
.I1(RIOB33_X105Y107_IOB_X1Y107_I),
.I2(LIOB33_X0Y101_IOB_X0Y101_I),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X12Y106_SLICE_X17Y106_AO5),
.O6(CLBLM_L_X12Y106_SLICE_X17Y106_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h599aa665a665599a)
  ) CLBLM_L_X12Y107_SLICE_X16Y107_DLUT (
.I0(CLBLM_L_X12Y105_SLICE_X17Y105_AO6),
.I1(CLBLM_L_X12Y105_SLICE_X17Y105_BO6),
.I2(CLBLM_R_X13Y106_SLICE_X18Y106_BO6),
.I3(CLBLM_L_X12Y106_SLICE_X16Y106_AO5),
.I4(CLBLM_R_X11Y107_SLICE_X15Y107_AO6),
.I5(CLBLM_R_X11Y107_SLICE_X14Y107_BO5),
.O5(CLBLM_L_X12Y107_SLICE_X16Y107_DO5),
.O6(CLBLM_L_X12Y107_SLICE_X16Y107_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h2dd2d22db44b4bb4)
  ) CLBLM_L_X12Y107_SLICE_X16Y107_CLUT (
.I0(CLBLM_L_X12Y106_SLICE_X17Y106_BO6),
.I1(CLBLM_R_X11Y107_SLICE_X14Y107_AO6),
.I2(CLBLM_R_X13Y106_SLICE_X18Y106_CO6),
.I3(CLBLM_L_X12Y106_SLICE_X17Y106_DO6),
.I4(CLBLM_L_X12Y108_SLICE_X16Y108_AO5),
.I5(CLBLM_L_X12Y104_SLICE_X16Y104_DO6),
.O5(CLBLM_L_X12Y107_SLICE_X16Y107_CO5),
.O6(CLBLM_L_X12Y107_SLICE_X16Y107_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h7fbfbfbf152a2a2a)
  ) CLBLM_L_X12Y107_SLICE_X16Y107_BLUT (
.I0(CLBLM_L_X12Y106_SLICE_X16Y106_DO6),
.I1(RIOB33_X105Y105_IOB_X1Y105_I),
.I2(LIOB33_X0Y103_IOB_X0Y104_I),
.I3(RIOB33_X105Y107_IOB_X1Y107_I),
.I4(LIOB33_X0Y101_IOB_X0Y102_I),
.I5(CLBLM_L_X12Y104_SLICE_X16Y104_DO6),
.O5(CLBLM_L_X12Y107_SLICE_X16Y107_BO5),
.O6(CLBLM_L_X12Y107_SLICE_X16Y107_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h399cc663c663399c)
  ) CLBLM_L_X12Y107_SLICE_X16Y107_ALUT (
.I0(CLBLM_R_X13Y106_SLICE_X18Y106_CO6),
.I1(CLBLM_L_X12Y105_SLICE_X17Y105_BO6),
.I2(CLBLM_L_X12Y108_SLICE_X16Y108_AO5),
.I3(CLBLM_L_X12Y106_SLICE_X17Y106_DO6),
.I4(CLBLM_R_X13Y106_SLICE_X18Y106_BO6),
.I5(CLBLM_L_X12Y106_SLICE_X16Y106_AO5),
.O5(CLBLM_L_X12Y107_SLICE_X16Y107_AO5),
.O6(CLBLM_L_X12Y107_SLICE_X16Y107_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h4cdfdf4cdf4cdf4c)
  ) CLBLM_L_X12Y107_SLICE_X17Y107_DLUT (
.I0(LIOB33_X0Y103_IOB_X0Y104_I),
.I1(CLBLM_L_X12Y106_SLICE_X17Y106_DO6),
.I2(RIOB33_X105Y107_IOB_X1Y107_I),
.I3(CLBLM_R_X13Y106_SLICE_X18Y106_DO6),
.I4(RIOB33_X105Y107_IOB_X1Y108_I),
.I5(LIOB33_X0Y101_IOB_X0Y102_I),
.O5(CLBLM_L_X12Y107_SLICE_X17Y107_DO5),
.O6(CLBLM_L_X12Y107_SLICE_X17Y107_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0c5f4fdf4cdf5fff)
  ) CLBLM_L_X12Y107_SLICE_X17Y107_CLUT (
.I0(LIOB33_X0Y103_IOB_X0Y104_I),
.I1(CLBLM_R_X13Y106_SLICE_X19Y106_AO5),
.I2(RIOB33_X105Y107_IOB_X1Y108_I),
.I3(CLBLM_L_X12Y105_SLICE_X17Y105_BO6),
.I4(CLBLM_R_X13Y106_SLICE_X18Y106_AO6),
.I5(LIOB33_X0Y101_IOB_X0Y102_I),
.O5(CLBLM_L_X12Y107_SLICE_X17Y107_CO5),
.O6(CLBLM_L_X12Y107_SLICE_X17Y107_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hb44b2dd2dd22dd22)
  ) CLBLM_L_X12Y107_SLICE_X17Y107_BLUT (
.I0(CLBLM_R_X13Y106_SLICE_X18Y106_AO6),
.I1(CLBLM_R_X13Y106_SLICE_X19Y106_AO5),
.I2(LIOB33_X0Y103_IOB_X0Y104_I),
.I3(CLBLM_L_X12Y105_SLICE_X17Y105_BO6),
.I4(LIOB33_X0Y101_IOB_X0Y102_I),
.I5(RIOB33_X105Y107_IOB_X1Y108_I),
.O5(CLBLM_L_X12Y107_SLICE_X17Y107_BO5),
.O6(CLBLM_L_X12Y107_SLICE_X17Y107_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h5555ffffb24d30cf)
  ) CLBLM_L_X12Y107_SLICE_X17Y107_ALUT (
.I0(RIOB33_X105Y107_IOB_X1Y108_I),
.I1(CLBLM_R_X13Y106_SLICE_X19Y106_AO5),
.I2(CLBLM_R_X13Y106_SLICE_X18Y106_AO6),
.I3(CLBLM_L_X12Y105_SLICE_X17Y105_BO6),
.I4(LIOB33_X0Y101_IOB_X0Y102_I),
.I5(1'b1),
.O5(CLBLM_L_X12Y107_SLICE_X17Y107_AO5),
.O6(CLBLM_L_X12Y107_SLICE_X17Y107_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h7fdf134cdfdf4c4c)
  ) CLBLM_L_X12Y108_SLICE_X16Y108_DLUT (
.I0(LIOB33_X0Y105_IOB_X0Y105_I),
.I1(CLBLM_L_X12Y107_SLICE_X17Y107_AO5),
.I2(RIOB33_X105Y107_IOB_X1Y107_I),
.I3(RIOB33_X105Y107_IOB_X1Y108_I),
.I4(CLBLM_L_X12Y107_SLICE_X17Y107_DO6),
.I5(LIOB33_X0Y103_IOB_X0Y104_I),
.O5(CLBLM_L_X12Y108_SLICE_X16Y108_DO5),
.O6(CLBLM_L_X12Y108_SLICE_X16Y108_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h9aa66a565a96aa66)
  ) CLBLM_L_X12Y108_SLICE_X16Y108_CLUT (
.I0(CLBLM_R_X11Y107_SLICE_X15Y107_DO6),
.I1(CLBLM_R_X11Y106_SLICE_X15Y106_BO6),
.I2(RIOB33_X105Y107_IOB_X1Y108_I),
.I3(CLBLM_L_X12Y107_SLICE_X17Y107_CO6),
.I4(LIOB33_X0Y105_IOB_X0Y106_I),
.I5(LIOB33_X0Y105_IOB_X0Y105_I),
.O5(CLBLM_L_X12Y108_SLICE_X16Y108_CO5),
.O6(CLBLM_L_X12Y108_SLICE_X16Y108_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h1f5f7fff03135f7f)
  ) CLBLM_L_X12Y108_SLICE_X16Y108_BLUT (
.I0(LIOB33_X0Y105_IOB_X0Y106_I),
.I1(CLBLM_R_X11Y106_SLICE_X15Y106_BO6),
.I2(RIOB33_X105Y107_IOB_X1Y108_I),
.I3(LIOB33_X0Y105_IOB_X0Y105_I),
.I4(CLBLM_R_X11Y107_SLICE_X15Y107_DO6),
.I5(CLBLM_L_X12Y107_SLICE_X17Y107_CO6),
.O5(CLBLM_L_X12Y108_SLICE_X16Y108_BO5),
.O6(CLBLM_L_X12Y108_SLICE_X16Y108_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h3333ffff00ffffff)
  ) CLBLM_L_X12Y108_SLICE_X16Y108_ALUT (
.I0(1'b1),
.I1(LIOB33_X0Y105_IOB_X0Y105_I),
.I2(1'b1),
.I3(LIOB33_X0Y103_IOB_X0Y104_I),
.I4(RIOB33_X105Y107_IOB_X1Y107_I),
.I5(1'b1),
.O5(CLBLM_L_X12Y108_SLICE_X16Y108_AO5),
.O6(CLBLM_L_X12Y108_SLICE_X16Y108_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h7dddffff14443ccc)
  ) CLBLM_L_X12Y108_SLICE_X17Y108_DLUT (
.I0(LIOB33_X0Y105_IOB_X0Y105_I),
.I1(CLBLM_L_X12Y106_SLICE_X17Y106_CO6),
.I2(LIOB33_X0Y103_IOB_X0Y104_I),
.I3(RIOB33_X105Y107_IOB_X1Y107_I),
.I4(RIOB33_X105Y105_IOB_X1Y105_I),
.I5(CLBLM_L_X12Y107_SLICE_X16Y107_BO6),
.O5(CLBLM_L_X12Y108_SLICE_X17Y108_DO5),
.O6(CLBLM_L_X12Y108_SLICE_X17Y108_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h7ddd1444ffff3ccc)
  ) CLBLM_L_X12Y108_SLICE_X17Y108_CLUT (
.I0(RIOB33_X105Y103_IOB_X1Y104_I),
.I1(CLBLM_L_X12Y106_SLICE_X16Y106_CO6),
.I2(LIOB33_X0Y103_IOB_X0Y104_I),
.I3(RIOB33_X105Y105_IOB_X1Y105_I),
.I4(CLBLM_R_X11Y105_SLICE_X15Y105_CO6),
.I5(LIOB33_X0Y105_IOB_X0Y105_I),
.O5(CLBLM_L_X12Y108_SLICE_X17Y108_CO5),
.O6(CLBLM_L_X12Y108_SLICE_X17Y108_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h6c93a05f936c5fa0)
  ) CLBLM_L_X12Y108_SLICE_X17Y108_BLUT (
.I0(RIOB33_X105Y105_IOB_X1Y105_I),
.I1(LIOB33_X0Y103_IOB_X0Y104_I),
.I2(LIOB33_X0Y105_IOB_X0Y105_I),
.I3(CLBLM_L_X12Y107_SLICE_X16Y107_BO6),
.I4(RIOB33_X105Y107_IOB_X1Y107_I),
.I5(CLBLM_L_X12Y106_SLICE_X17Y106_CO6),
.O5(CLBLM_L_X12Y108_SLICE_X17Y108_BO5),
.O6(CLBLM_L_X12Y108_SLICE_X17Y108_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'ha6cf593065cf9a30)
  ) CLBLM_L_X12Y108_SLICE_X17Y108_ALUT (
.I0(RIOB33_X105Y107_IOB_X1Y107_I),
.I1(CLBLM_L_X12Y107_SLICE_X16Y107_BO6),
.I2(CLBLM_R_X13Y107_SLICE_X18Y107_AO6),
.I3(LIOB33_X0Y105_IOB_X0Y105_I),
.I4(CLBLM_L_X12Y107_SLICE_X16Y107_AO6),
.I5(RIOB33_X105Y105_IOB_X1Y105_I),
.O5(CLBLM_L_X12Y108_SLICE_X17Y108_AO5),
.O6(CLBLM_L_X12Y108_SLICE_X17Y108_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hff999f099f099900)
  ) CLBLM_L_X12Y109_SLICE_X16Y109_DLUT (
.I0(CLBLM_L_X12Y109_SLICE_X16Y109_AO6),
.I1(CLBLM_L_X12Y107_SLICE_X16Y107_DO6),
.I2(CLBLM_L_X12Y107_SLICE_X17Y107_BO6),
.I3(CLBLM_L_X12Y110_SLICE_X16Y110_AO6),
.I4(CLBLM_L_X12Y108_SLICE_X16Y108_AO6),
.I5(CLBLM_L_X12Y107_SLICE_X17Y107_DO6),
.O5(CLBLM_L_X12Y109_SLICE_X16Y109_DO5),
.O6(CLBLM_L_X12Y109_SLICE_X16Y109_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h87f078f0e13c1e3c)
  ) CLBLM_L_X12Y109_SLICE_X16Y109_CLUT (
.I0(RIOB33_X105Y105_IOB_X1Y105_I),
.I1(CLBLM_R_X11Y108_SLICE_X15Y108_DO6),
.I2(CLBLM_L_X12Y109_SLICE_X17Y109_BO6),
.I3(LIOB33_X0Y105_IOB_X0Y106_I),
.I4(RIOB33_X105Y107_IOB_X1Y107_I),
.I5(CLBLM_L_X12Y108_SLICE_X17Y108_DO6),
.O5(CLBLM_L_X12Y109_SLICE_X16Y109_CO5),
.O6(CLBLM_L_X12Y109_SLICE_X16Y109_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h59a6a6599a65659a)
  ) CLBLM_L_X12Y109_SLICE_X16Y109_BLUT (
.I0(CLBLM_L_X12Y107_SLICE_X16Y107_DO6),
.I1(CLBLM_L_X12Y107_SLICE_X17Y107_BO6),
.I2(CLBLM_L_X12Y108_SLICE_X16Y108_AO6),
.I3(CLBLM_L_X12Y110_SLICE_X16Y110_AO6),
.I4(CLBLM_L_X12Y109_SLICE_X16Y109_AO6),
.I5(CLBLM_L_X12Y107_SLICE_X17Y107_DO6),
.O5(CLBLM_L_X12Y109_SLICE_X16Y109_BO5),
.O6(CLBLM_L_X12Y109_SLICE_X16Y109_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h7777777778877887)
  ) CLBLM_L_X12Y109_SLICE_X16Y109_ALUT (
.I0(LIOB33_X0Y105_IOB_X0Y105_I),
.I1(RIOB33_X105Y107_IOB_X1Y108_I),
.I2(CLBLM_L_X12Y107_SLICE_X17Y107_CO6),
.I3(CLBLM_R_X11Y106_SLICE_X15Y106_BO6),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X12Y109_SLICE_X16Y109_AO5),
.O6(CLBLM_L_X12Y109_SLICE_X16Y109_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X12Y109_SLICE_X17Y109_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X12Y109_SLICE_X17Y109_DO5),
.O6(CLBLM_L_X12Y109_SLICE_X17Y109_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X12Y109_SLICE_X17Y109_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X12Y109_SLICE_X17Y109_CO5),
.O6(CLBLM_L_X12Y109_SLICE_X17Y109_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'ha66a66aa9955a66a)
  ) CLBLM_L_X12Y109_SLICE_X17Y109_BLUT (
.I0(CLBLM_L_X12Y107_SLICE_X16Y107_DO6),
.I1(LIOB33_X0Y105_IOB_X0Y105_I),
.I2(RIOB33_X105Y107_IOB_X1Y107_I),
.I3(RIOB33_X105Y107_IOB_X1Y108_I),
.I4(CLBLM_L_X12Y107_SLICE_X17Y107_BO6),
.I5(CLBLM_L_X12Y107_SLICE_X17Y107_DO6),
.O5(CLBLM_L_X12Y109_SLICE_X17Y109_BO5),
.O6(CLBLM_L_X12Y109_SLICE_X17Y109_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hc663399c9c9c9c9c)
  ) CLBLM_L_X12Y109_SLICE_X17Y109_ALUT (
.I0(CLBLM_L_X12Y108_SLICE_X17Y108_CO6),
.I1(CLBLM_L_X12Y108_SLICE_X17Y108_AO6),
.I2(CLBLM_L_X12Y108_SLICE_X17Y108_BO6),
.I3(RIOB33_X105Y103_IOB_X1Y104_I),
.I4(RIOB33_X105Y105_IOB_X1Y105_I),
.I5(LIOB33_X0Y105_IOB_X0Y106_I),
.O5(CLBLM_L_X12Y109_SLICE_X17Y109_AO5),
.O6(CLBLM_L_X12Y109_SLICE_X17Y109_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h6996c33c3cc36996)
  ) CLBLM_L_X12Y110_SLICE_X16Y110_DLUT (
.I0(CLBLM_R_X11Y107_SLICE_X15Y107_CO6),
.I1(CLBLM_L_X12Y108_SLICE_X16Y108_CO6),
.I2(CLBLM_L_X12Y109_SLICE_X16Y109_DO6),
.I3(CLBLM_L_X12Y110_SLICE_X16Y110_AO5),
.I4(CLBLM_R_X11Y111_SLICE_X15Y111_BO5),
.I5(CLBLM_L_X12Y109_SLICE_X16Y109_BO6),
.O5(CLBLM_L_X12Y110_SLICE_X16Y110_DO5),
.O6(CLBLM_L_X12Y110_SLICE_X16Y110_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h6fafffff060a66aa)
  ) CLBLM_L_X12Y110_SLICE_X16Y110_CLUT (
.I0(CLBLM_L_X12Y109_SLICE_X17Y109_AO6),
.I1(LIOB33_X0Y107_IOB_X0Y107_I),
.I2(RIOB33_X105Y103_IOB_X1Y103_I),
.I3(RIOB33_X105Y103_IOB_X1Y104_I),
.I4(LIOB33_X0Y107_IOB_X0Y108_I),
.I5(CLBLM_R_X11Y109_SLICE_X15Y109_BO6),
.O5(CLBLM_L_X12Y110_SLICE_X16Y110_CO5),
.O6(CLBLM_L_X12Y110_SLICE_X16Y110_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h69999666c3333ccc)
  ) CLBLM_L_X12Y110_SLICE_X16Y110_BLUT (
.I0(LIOB33_X0Y107_IOB_X0Y108_I),
.I1(CLBLM_R_X11Y109_SLICE_X15Y109_BO6),
.I2(LIOB33_X0Y107_IOB_X0Y107_I),
.I3(RIOB33_X105Y103_IOB_X1Y104_I),
.I4(CLBLM_L_X12Y109_SLICE_X17Y109_AO6),
.I5(RIOB33_X105Y103_IOB_X1Y103_I),
.O5(CLBLM_L_X12Y110_SLICE_X16Y110_BO5),
.O6(CLBLM_L_X12Y110_SLICE_X16Y110_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h33ff33ff0fff0fff)
  ) CLBLM_L_X12Y110_SLICE_X16Y110_ALUT (
.I0(1'b1),
.I1(LIOB33_X0Y105_IOB_X0Y106_I),
.I2(LIOB33_X0Y107_IOB_X0Y107_I),
.I3(RIOB33_X105Y107_IOB_X1Y107_I),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X12Y110_SLICE_X16Y110_AO5),
.O6(CLBLM_L_X12Y110_SLICE_X16Y110_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X12Y110_SLICE_X17Y110_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X12Y110_SLICE_X17Y110_DO5),
.O6(CLBLM_L_X12Y110_SLICE_X17Y110_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X12Y110_SLICE_X17Y110_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X12Y110_SLICE_X17Y110_CO5),
.O6(CLBLM_L_X12Y110_SLICE_X17Y110_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X12Y110_SLICE_X17Y110_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X12Y110_SLICE_X17Y110_BO5),
.O6(CLBLM_L_X12Y110_SLICE_X17Y110_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X12Y110_SLICE_X17Y110_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X12Y110_SLICE_X17Y110_AO5),
.O6(CLBLM_L_X12Y110_SLICE_X17Y110_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y103_SLICE_X2Y103_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y103_SLICE_X2Y103_DO5),
.O6(CLBLM_R_X3Y103_SLICE_X2Y103_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y103_SLICE_X2Y103_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y103_SLICE_X2Y103_CO5),
.O6(CLBLM_R_X3Y103_SLICE_X2Y103_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h939f939f539f539f)
  ) CLBLM_R_X3Y103_SLICE_X2Y103_BLUT (
.I0(LIOB33_SING_X0Y100_IOB_X0Y100_I),
.I1(RIOB33_X105Y113_IOB_X1Y113_I),
.I2(LIOB33_X0Y115_IOB_X0Y116_I),
.I3(LIOB33_X0Y117_IOB_X0Y117_I),
.I4(1'b1),
.I5(RIOB33_X105Y111_IOB_X1Y112_I),
.O5(CLBLM_R_X3Y103_SLICE_X2Y103_BO5),
.O6(CLBLM_R_X3Y103_SLICE_X2Y103_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h4278724802b8f248)
  ) CLBLM_R_X3Y103_SLICE_X2Y103_ALUT (
.I0(LIOB33_SING_X0Y100_IOB_X0Y100_I),
.I1(LIOB33_X0Y115_IOB_X0Y116_I),
.I2(RIOB33_X105Y113_IOB_X1Y113_I),
.I3(LIOB33_X0Y113_IOB_X0Y114_I),
.I4(LIOB33_X0Y117_IOB_X0Y117_I),
.I5(RIOB33_X105Y111_IOB_X1Y112_I),
.O5(CLBLM_R_X3Y103_SLICE_X2Y103_AO5),
.O6(CLBLM_R_X3Y103_SLICE_X2Y103_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y103_SLICE_X3Y103_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y103_SLICE_X3Y103_DO5),
.O6(CLBLM_R_X3Y103_SLICE_X3Y103_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y103_SLICE_X3Y103_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y103_SLICE_X3Y103_CO5),
.O6(CLBLM_R_X3Y103_SLICE_X3Y103_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0ff55ff50ff55ff)
  ) CLBLM_R_X3Y103_SLICE_X3Y103_BLUT (
.I0(LIOB33_SING_X0Y100_IOB_X0Y100_I),
.I1(1'b1),
.I2(LIOB33_X0Y115_IOB_X0Y116_I),
.I3(LIOB33_X0Y113_IOB_X0Y114_I),
.I4(RIOB33_X105Y113_IOB_X1Y113_I),
.I5(RIOB33_X105Y111_IOB_X1Y112_I),
.O5(CLBLM_R_X3Y103_SLICE_X3Y103_BO5),
.O6(CLBLM_R_X3Y103_SLICE_X3Y103_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'ha5a50f0f7711ff33)
  ) CLBLM_R_X3Y103_SLICE_X3Y103_ALUT (
.I0(LIOB33_X0Y113_IOB_X0Y114_I),
.I1(CLBLM_R_X3Y103_SLICE_X2Y103_BO6),
.I2(CLBLM_R_X3Y103_SLICE_X2Y103_AO6),
.I3(CLBLM_R_X3Y103_SLICE_X3Y103_BO6),
.I4(LIOB33_X0Y101_IOB_X0Y101_I),
.I5(1'b1),
.O5(CLBLM_R_X3Y103_SLICE_X3Y103_AO5),
.O6(CLBLM_R_X3Y103_SLICE_X3Y103_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h8fe5701a7f1580ea)
  ) CLBLM_R_X3Y104_SLICE_X2Y104_DLUT (
.I0(CLBLM_R_X3Y103_SLICE_X3Y103_AO6),
.I1(LIOB33_X0Y103_IOB_X0Y103_I),
.I2(LIOB33_X0Y101_IOB_X0Y102_I),
.I3(CLBLM_R_X3Y104_SLICE_X2Y104_AO5),
.I4(CLBLL_L_X4Y103_SLICE_X4Y103_BO6),
.I5(LIOB33_X0Y113_IOB_X0Y114_I),
.O5(CLBLM_R_X3Y104_SLICE_X2Y104_DO5),
.O6(CLBLM_R_X3Y104_SLICE_X2Y104_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h1c441c0050441c00)
  ) CLBLM_R_X3Y104_SLICE_X2Y104_CLUT (
.I0(LIOB33_X0Y103_IOB_X0Y103_I),
.I1(RIOB33_X105Y113_IOB_X1Y113_I),
.I2(LIOB33_SING_X0Y100_IOB_X0Y100_I),
.I3(LIOB33_X0Y113_IOB_X0Y114_I),
.I4(LIOB33_X0Y115_IOB_X0Y116_I),
.I5(RIOB33_X105Y111_IOB_X1Y112_I),
.O5(CLBLM_R_X3Y104_SLICE_X2Y104_CO5),
.O6(CLBLM_R_X3Y104_SLICE_X2Y104_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h3ccc3cccc3339c6c)
  ) CLBLM_R_X3Y104_SLICE_X2Y104_BLUT (
.I0(LIOB33_X0Y103_IOB_X0Y103_I),
.I1(CLBLM_R_X3Y103_SLICE_X2Y103_AO6),
.I2(LIOB33_X0Y101_IOB_X0Y101_I),
.I3(LIOB33_X0Y113_IOB_X0Y114_I),
.I4(CLBLM_R_X3Y105_SLICE_X2Y105_AO6),
.I5(CLBLM_R_X3Y104_SLICE_X2Y104_CO6),
.O5(CLBLM_R_X3Y104_SLICE_X2Y104_BO5),
.O6(CLBLM_R_X3Y104_SLICE_X2Y104_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'ha5a50f0fcdcdcfcf)
  ) CLBLM_R_X3Y104_SLICE_X2Y104_ALUT (
.I0(LIOB33_X0Y103_IOB_X0Y103_I),
.I1(CLBLM_R_X3Y104_SLICE_X2Y104_CO6),
.I2(CLBLM_R_X3Y105_SLICE_X2Y105_AO6),
.I3(1'b1),
.I4(LIOB33_X0Y101_IOB_X0Y101_I),
.I5(1'b1),
.O5(CLBLM_R_X3Y104_SLICE_X2Y104_AO5),
.O6(CLBLM_R_X3Y104_SLICE_X2Y104_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'he8fae8e88eaf8e8e)
  ) CLBLM_R_X3Y104_SLICE_X3Y104_DLUT (
.I0(CLBLM_R_X3Y104_SLICE_X3Y104_AO6),
.I1(CLBLM_R_X3Y104_SLICE_X2Y104_CO6),
.I2(CLBLM_R_X3Y106_SLICE_X2Y106_BO5),
.I3(CLBLM_R_X3Y105_SLICE_X2Y105_AO6),
.I4(CLBLL_L_X4Y103_SLICE_X4Y103_AO6),
.I5(CLBLM_R_X3Y103_SLICE_X2Y103_AO6),
.O5(CLBLM_R_X3Y104_SLICE_X3Y104_DO5),
.O6(CLBLM_R_X3Y104_SLICE_X3Y104_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hfba2f751faa0f550)
  ) CLBLM_R_X3Y104_SLICE_X3Y104_CLUT (
.I0(CLBLM_R_X3Y105_SLICE_X2Y105_AO6),
.I1(CLBLL_L_X2Y104_SLICE_X0Y104_BO6),
.I2(CLBLL_L_X2Y104_SLICE_X0Y104_CO6),
.I3(CLBLM_R_X3Y104_SLICE_X3Y104_AO5),
.I4(CLBLL_L_X4Y103_SLICE_X4Y103_AO6),
.I5(CLBLM_R_X13Y106_SLICE_X18Y106_AO5),
.O5(CLBLM_R_X3Y104_SLICE_X3Y104_CO5),
.O6(CLBLM_R_X3Y104_SLICE_X3Y104_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h6cffffff006c6c6c)
  ) CLBLM_R_X3Y104_SLICE_X3Y104_BLUT (
.I0(LIOB33_X0Y101_IOB_X0Y102_I),
.I1(CLBLM_R_X3Y104_SLICE_X2Y104_BO6),
.I2(LIOB33_X0Y103_IOB_X0Y103_I),
.I3(RIOB33_X105Y105_IOB_X1Y106_I),
.I4(LIOB33_X0Y103_IOB_X0Y104_I),
.I5(CLBLM_R_X3Y104_SLICE_X3Y104_CO6),
.O5(CLBLM_R_X3Y104_SLICE_X3Y104_BO5),
.O6(CLBLM_R_X3Y104_SLICE_X3Y104_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0f0fffff3f3f3f3f)
  ) CLBLM_R_X3Y104_SLICE_X3Y104_ALUT (
.I0(1'b1),
.I1(RIOB33_X105Y105_IOB_X1Y106_I),
.I2(LIOB33_X0Y101_IOB_X0Y102_I),
.I3(1'b1),
.I4(LIOB33_X0Y103_IOB_X0Y103_I),
.I5(1'b1),
.O5(CLBLM_R_X3Y104_SLICE_X3Y104_AO5),
.O6(CLBLM_R_X3Y104_SLICE_X3Y104_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y105_SLICE_X2Y105_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y105_SLICE_X2Y105_DO5),
.O6(CLBLM_R_X3Y105_SLICE_X2Y105_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h7fb31320ffff5fa0)
  ) CLBLM_R_X3Y105_SLICE_X2Y105_CLUT (
.I0(LIOB33_X0Y103_IOB_X0Y103_I),
.I1(RIOB33_X105Y105_IOB_X1Y106_I),
.I2(LIOB33_X0Y103_IOB_X0Y104_I),
.I3(CLBLM_R_X3Y104_SLICE_X2Y104_DO6),
.I4(CLBLM_R_X3Y104_SLICE_X3Y104_BO6),
.I5(LIOB33_X0Y105_IOB_X0Y105_I),
.O5(CLBLM_R_X3Y105_SLICE_X2Y105_CO5),
.O6(CLBLM_R_X3Y105_SLICE_X2Y105_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h6a95956ac03f3fc0)
  ) CLBLM_R_X3Y105_SLICE_X2Y105_BLUT (
.I0(RIOB33_X105Y105_IOB_X1Y106_I),
.I1(LIOB33_X0Y103_IOB_X0Y104_I),
.I2(LIOB33_X0Y103_IOB_X0Y103_I),
.I3(CLBLM_R_X3Y104_SLICE_X2Y104_DO6),
.I4(CLBLM_R_X3Y104_SLICE_X3Y104_BO6),
.I5(LIOB33_X0Y105_IOB_X0Y105_I),
.O5(CLBLM_R_X3Y105_SLICE_X2Y105_BO5),
.O6(CLBLM_R_X3Y105_SLICE_X2Y105_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h472874280b28f428)
  ) CLBLM_R_X3Y105_SLICE_X2Y105_ALUT (
.I0(LIOB33_SING_X0Y100_IOB_X0Y100_I),
.I1(LIOB33_X0Y113_IOB_X0Y114_I),
.I2(LIOB33_X0Y103_IOB_X0Y103_I),
.I3(RIOB33_X105Y113_IOB_X1Y113_I),
.I4(LIOB33_X0Y115_IOB_X0Y116_I),
.I5(RIOB33_X105Y111_IOB_X1Y112_I),
.O5(CLBLM_R_X3Y105_SLICE_X2Y105_AO5),
.O6(CLBLM_R_X3Y105_SLICE_X2Y105_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y105_SLICE_X3Y105_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y105_SLICE_X3Y105_DO5),
.O6(CLBLM_R_X3Y105_SLICE_X3Y105_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y105_SLICE_X3Y105_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y105_SLICE_X3Y105_CO5),
.O6(CLBLM_R_X3Y105_SLICE_X3Y105_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y105_SLICE_X3Y105_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y105_SLICE_X3Y105_BO5),
.O6(CLBLM_R_X3Y105_SLICE_X3Y105_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y105_SLICE_X3Y105_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y105_SLICE_X3Y105_AO5),
.O6(CLBLM_R_X3Y105_SLICE_X3Y105_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h96669996cccc3c3c)
  ) CLBLM_R_X3Y106_SLICE_X2Y106_DLUT (
.I0(LIOB33_X0Y103_IOB_X0Y103_I),
.I1(CLBLL_L_X4Y104_SLICE_X4Y104_AO6),
.I2(CLBLL_L_X4Y104_SLICE_X4Y104_BO6),
.I3(RIOB33_X105Y105_IOB_X1Y106_I),
.I4(CLBLM_R_X3Y104_SLICE_X3Y104_BO6),
.I5(LIOB33_X0Y105_IOB_X0Y105_I),
.O5(CLBLM_R_X3Y106_SLICE_X2Y106_DO5),
.O6(CLBLM_R_X3Y106_SLICE_X2Y106_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0c043cb400008888)
  ) CLBLM_R_X3Y106_SLICE_X2Y106_CLUT (
.I0(LIOB33_X0Y103_IOB_X0Y103_I),
.I1(RIOB33_X105Y113_IOB_X1Y113_I),
.I2(LIOB33_SING_X0Y100_IOB_X0Y100_I),
.I3(RIOB33_X105Y111_IOB_X1Y112_I),
.I4(RIOB33_SING_X105Y100_IOB_X1Y100_I),
.I5(RIOB33_X105Y105_IOB_X1Y106_I),
.O5(CLBLM_R_X3Y106_SLICE_X2Y106_CO5),
.O6(CLBLM_R_X3Y106_SLICE_X2Y106_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h20a020a03333ffff)
  ) CLBLM_R_X3Y106_SLICE_X2Y106_BLUT (
.I0(RIOB33_X105Y113_IOB_X1Y113_I),
.I1(LIOB33_X0Y113_IOB_X0Y114_I),
.I2(LIOB33_X0Y103_IOB_X0Y103_I),
.I3(RIOB33_X105Y111_IOB_X1Y112_I),
.I4(LIOB33_X0Y101_IOB_X0Y101_I),
.I5(1'b1),
.O5(CLBLM_R_X3Y106_SLICE_X2Y106_BO5),
.O6(CLBLM_R_X3Y106_SLICE_X2Y106_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h2000000099993333)
  ) CLBLM_R_X3Y106_SLICE_X2Y106_ALUT (
.I0(RIOB33_SING_X105Y100_IOB_X1Y100_I),
.I1(CLBLL_L_X2Y106_SLICE_X1Y106_BO6),
.I2(CLBLM_R_X3Y103_SLICE_X2Y103_BO6),
.I3(CLBLM_R_X3Y106_SLICE_X2Y106_BO6),
.I4(LIOB33_X0Y101_IOB_X0Y101_I),
.I5(1'b1),
.O5(CLBLM_R_X3Y106_SLICE_X2Y106_AO5),
.O6(CLBLM_R_X3Y106_SLICE_X2Y106_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hfab2f571b2a07150)
  ) CLBLM_R_X3Y106_SLICE_X3Y106_DLUT (
.I0(CLBLM_R_X3Y106_SLICE_X3Y106_AO6),
.I1(CLBLL_L_X4Y104_SLICE_X4Y104_BO6),
.I2(CLBLM_R_X3Y107_SLICE_X2Y107_AO5),
.I3(CLBLM_R_X3Y106_SLICE_X3Y106_AO5),
.I4(CLBLL_L_X4Y104_SLICE_X4Y104_AO6),
.I5(CLBLM_R_X3Y104_SLICE_X3Y104_BO6),
.O5(CLBLM_R_X3Y106_SLICE_X3Y106_DO5),
.O6(CLBLM_R_X3Y106_SLICE_X3Y106_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h5a96a56996a5695a)
  ) CLBLM_R_X3Y106_SLICE_X3Y106_CLUT (
.I0(CLBLM_R_X3Y106_SLICE_X3Y106_AO6),
.I1(CLBLL_L_X4Y104_SLICE_X4Y104_BO6),
.I2(CLBLM_R_X3Y107_SLICE_X2Y107_AO5),
.I3(CLBLM_R_X3Y106_SLICE_X3Y106_AO5),
.I4(CLBLL_L_X4Y104_SLICE_X4Y104_AO6),
.I5(CLBLM_R_X3Y104_SLICE_X3Y104_BO6),
.O5(CLBLM_R_X3Y106_SLICE_X3Y106_CO5),
.O6(CLBLM_R_X3Y106_SLICE_X3Y106_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'ha66a6a6a95a6956a)
  ) CLBLM_R_X3Y106_SLICE_X3Y106_BLUT (
.I0(CLBLL_L_X4Y105_SLICE_X4Y105_AO6),
.I1(LIOB33_X0Y105_IOB_X0Y106_I),
.I2(LIOB33_X0Y103_IOB_X0Y103_I),
.I3(CLBLL_L_X4Y106_SLICE_X4Y106_AO6),
.I4(RIOB33_X105Y105_IOB_X1Y106_I),
.I5(CLBLM_R_X3Y105_SLICE_X2Y105_CO6),
.O5(CLBLM_R_X3Y106_SLICE_X3Y106_BO5),
.O6(CLBLM_R_X3Y106_SLICE_X3Y106_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0fff0fff33ff33ff)
  ) CLBLM_R_X3Y106_SLICE_X3Y106_ALUT (
.I0(1'b1),
.I1(RIOB33_X105Y105_IOB_X1Y106_I),
.I2(LIOB33_X0Y103_IOB_X0Y103_I),
.I3(LIOB33_X0Y105_IOB_X0Y105_I),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y106_SLICE_X3Y106_AO5),
.O6(CLBLM_R_X3Y106_SLICE_X3Y106_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0b2f2b3f3bbfbbff)
  ) CLBLM_R_X3Y107_SLICE_X2Y107_DLUT (
.I0(CLBLL_L_X2Y107_SLICE_X0Y107_BO6),
.I1(CLBLM_R_X3Y106_SLICE_X3Y106_CO6),
.I2(RIOB33_SING_X105Y100_IOB_X1Y100_I),
.I3(CLBLM_R_X3Y105_SLICE_X2Y105_BO6),
.I4(LIOB33_X0Y105_IOB_X0Y106_I),
.I5(LIOB33_X0Y107_IOB_X0Y107_I),
.O5(CLBLM_R_X3Y107_SLICE_X2Y107_DO5),
.O6(CLBLM_R_X3Y107_SLICE_X2Y107_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h6a95956ac03f3fc0)
  ) CLBLM_R_X3Y107_SLICE_X2Y107_CLUT (
.I0(RIOB33_X105Y105_IOB_X1Y106_I),
.I1(RIOB33_SING_X105Y100_IOB_X1Y100_I),
.I2(LIOB33_X0Y107_IOB_X0Y108_I),
.I3(CLBLM_R_X3Y106_SLICE_X3Y106_BO6),
.I4(CLBLM_R_X3Y107_SLICE_X2Y107_DO6),
.I5(LIOB33_X0Y107_IOB_X0Y107_I),
.O5(CLBLM_R_X3Y107_SLICE_X2Y107_CO5),
.O6(CLBLM_R_X3Y107_SLICE_X2Y107_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h8ef371f3710c8e0c)
  ) CLBLM_R_X3Y107_SLICE_X2Y107_BLUT (
.I0(RIOB33_SING_X105Y100_IOB_X1Y100_I),
.I1(CLBLM_R_X3Y105_SLICE_X2Y105_BO6),
.I2(CLBLL_L_X2Y107_SLICE_X0Y107_BO6),
.I3(LIOB33_X0Y105_IOB_X0Y106_I),
.I4(RIOB33_X105Y105_IOB_X1Y106_I),
.I5(CLBLM_R_X3Y106_SLICE_X2Y106_DO6),
.O5(CLBLM_R_X3Y107_SLICE_X2Y107_BO5),
.O6(CLBLM_R_X3Y107_SLICE_X2Y107_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h6969c3c355ff55ff)
  ) CLBLM_R_X3Y107_SLICE_X2Y107_ALUT (
.I0(LIOB33_X0Y105_IOB_X0Y106_I),
.I1(CLBLM_R_X3Y105_SLICE_X2Y105_BO6),
.I2(CLBLL_L_X2Y107_SLICE_X0Y107_BO6),
.I3(RIOB33_X105Y105_IOB_X1Y106_I),
.I4(RIOB33_SING_X105Y100_IOB_X1Y100_I),
.I5(1'b1),
.O5(CLBLM_R_X3Y107_SLICE_X2Y107_AO5),
.O6(CLBLM_R_X3Y107_SLICE_X2Y107_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hc6936c936cc66c6c)
  ) CLBLM_R_X3Y107_SLICE_X3Y107_DLUT (
.I0(LIOB33_X0Y109_IOB_X0Y109_I),
.I1(CLBLL_L_X4Y107_SLICE_X5Y107_BO6),
.I2(RIOB33_X105Y105_IOB_X1Y106_I),
.I3(CLBLM_R_X3Y107_SLICE_X3Y107_CO6),
.I4(RIOB33_SING_X105Y100_IOB_X1Y100_I),
.I5(CLBLL_L_X4Y107_SLICE_X4Y107_AO6),
.O5(CLBLM_R_X3Y107_SLICE_X3Y107_DO5),
.O6(CLBLM_R_X3Y107_SLICE_X3Y107_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h70f7f7f780f8f8f8)
  ) CLBLM_R_X3Y107_SLICE_X3Y107_CLUT (
.I0(RIOB33_X105Y105_IOB_X1Y106_I),
.I1(LIOB33_X0Y107_IOB_X0Y107_I),
.I2(CLBLM_R_X3Y107_SLICE_X2Y107_DO6),
.I3(RIOB33_SING_X105Y100_IOB_X1Y100_I),
.I4(LIOB33_X0Y107_IOB_X0Y108_I),
.I5(CLBLM_R_X3Y106_SLICE_X3Y106_BO6),
.O5(CLBLM_R_X3Y107_SLICE_X3Y107_CO5),
.O6(CLBLM_R_X3Y107_SLICE_X3Y107_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'ha5a555553333ffff)
  ) CLBLM_R_X3Y107_SLICE_X3Y107_BLUT (
.I0(CLBLM_R_X3Y107_SLICE_X3Y107_DO6),
.I1(RIOB33_X105Y105_IOB_X1Y106_I),
.I2(RIOB33_SING_X105Y100_IOB_X1Y100_I),
.I3(1'b1),
.I4(LIOB33_X0Y109_IOB_X0Y110_I),
.I5(1'b1),
.O5(CLBLM_R_X3Y107_SLICE_X3Y107_BO5),
.O6(CLBLM_R_X3Y107_SLICE_X3Y107_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h66cc99330fff0fff)
  ) CLBLM_R_X3Y107_SLICE_X3Y107_ALUT (
.I0(RIOB33_SING_X105Y100_IOB_X1Y100_I),
.I1(CLBLL_L_X4Y107_SLICE_X4Y107_AO6),
.I2(RIOB33_X105Y105_IOB_X1Y106_I),
.I3(LIOB33_X0Y109_IOB_X0Y109_I),
.I4(CLBLM_R_X3Y107_SLICE_X3Y107_CO6),
.I5(1'b1),
.O5(CLBLM_R_X3Y107_SLICE_X3Y107_AO5),
.O6(CLBLM_R_X3Y107_SLICE_X3Y107_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y108_SLICE_X2Y108_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y108_SLICE_X2Y108_DO5),
.O6(CLBLM_R_X3Y108_SLICE_X2Y108_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y108_SLICE_X2Y108_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y108_SLICE_X2Y108_CO5),
.O6(CLBLM_R_X3Y108_SLICE_X2Y108_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y108_SLICE_X2Y108_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y108_SLICE_X2Y108_BO5),
.O6(CLBLM_R_X3Y108_SLICE_X2Y108_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y108_SLICE_X2Y108_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y108_SLICE_X2Y108_AO5),
.O6(CLBLM_R_X3Y108_SLICE_X2Y108_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y108_SLICE_X3Y108_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y108_SLICE_X3Y108_DO5),
.O6(CLBLM_R_X3Y108_SLICE_X3Y108_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y108_SLICE_X3Y108_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y108_SLICE_X3Y108_CO5),
.O6(CLBLM_R_X3Y108_SLICE_X3Y108_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y108_SLICE_X3Y108_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y108_SLICE_X3Y108_BO5),
.O6(CLBLM_R_X3Y108_SLICE_X3Y108_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h6999c33396663ccc)
  ) CLBLM_R_X3Y108_SLICE_X3Y108_ALUT (
.I0(LIOB33_X0Y111_IOB_X0Y111_I),
.I1(CLBLM_R_X5Y107_SLICE_X6Y107_AO6),
.I2(RIOB33_X105Y105_IOB_X1Y106_I),
.I3(LIOB33_X0Y109_IOB_X0Y110_I),
.I4(RIOB33_SING_X105Y100_IOB_X1Y100_I),
.I5(CLBLL_L_X4Y107_SLICE_X4Y107_BO6),
.O5(CLBLM_R_X3Y108_SLICE_X3Y108_AO5),
.O6(CLBLM_R_X3Y108_SLICE_X3Y108_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y109_SLICE_X2Y109_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y109_SLICE_X2Y109_DO5),
.O6(CLBLM_R_X3Y109_SLICE_X2Y109_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y109_SLICE_X2Y109_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y109_SLICE_X2Y109_CO5),
.O6(CLBLM_R_X3Y109_SLICE_X2Y109_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y109_SLICE_X2Y109_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y109_SLICE_X2Y109_BO5),
.O6(CLBLM_R_X3Y109_SLICE_X2Y109_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y109_SLICE_X2Y109_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y109_SLICE_X2Y109_AO5),
.O6(CLBLM_R_X3Y109_SLICE_X2Y109_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y109_SLICE_X3Y109_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y109_SLICE_X3Y109_DO5),
.O6(CLBLM_R_X3Y109_SLICE_X3Y109_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y109_SLICE_X3Y109_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y109_SLICE_X3Y109_CO5),
.O6(CLBLM_R_X3Y109_SLICE_X3Y109_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y109_SLICE_X3Y109_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y109_SLICE_X3Y109_BO5),
.O6(CLBLM_R_X3Y109_SLICE_X3Y109_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h69c3963ca50f5af0)
  ) CLBLM_R_X3Y109_SLICE_X3Y109_ALUT (
.I0(LIOB33_X0Y113_IOB_X0Y113_I),
.I1(LIOB33_X0Y115_IOB_X0Y115_I),
.I2(CLBLL_L_X4Y108_SLICE_X5Y108_AO6),
.I3(RIOB33_X105Y105_IOB_X1Y106_I),
.I4(CLBLL_L_X4Y108_SLICE_X4Y108_DO6),
.I5(RIOB33_SING_X105Y100_IOB_X1Y100_I),
.O5(CLBLM_R_X3Y109_SLICE_X3Y109_AO5),
.O6(CLBLM_R_X3Y109_SLICE_X3Y109_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h3933363c9c3c6ccc)
  ) CLBLM_R_X3Y112_SLICE_X2Y112_DLUT (
.I0(RIOB33_X105Y109_IOB_X1Y110_I),
.I1(CLBLM_R_X3Y112_SLICE_X3Y112_AO6),
.I2(CLBLM_R_X5Y113_SLICE_X7Y113_CO6),
.I3(LIOB33_X0Y115_IOB_X0Y115_I),
.I4(CLBLM_R_X3Y112_SLICE_X2Y112_BO6),
.I5(CLBLL_L_X4Y113_SLICE_X4Y113_BO6),
.O5(CLBLM_R_X3Y112_SLICE_X2Y112_DO5),
.O6(CLBLM_R_X3Y112_SLICE_X2Y112_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h3b020202bf232323)
  ) CLBLM_R_X3Y112_SLICE_X2Y112_CLUT (
.I0(CLBLM_R_X3Y112_SLICE_X2Y112_AO6),
.I1(CLBLM_R_X3Y112_SLICE_X3Y112_AO5),
.I2(CLBLM_R_X5Y113_SLICE_X7Y113_CO6),
.I3(RIOB33_X105Y111_IOB_X1Y111_I),
.I4(LIOB33_X0Y115_IOB_X0Y115_I),
.I5(CLBLL_L_X4Y113_SLICE_X4Y113_BO6),
.O5(CLBLM_R_X3Y112_SLICE_X2Y112_CO5),
.O6(CLBLM_R_X3Y112_SLICE_X2Y112_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'ha79f97dfdf5f5f5f)
  ) CLBLM_R_X3Y112_SLICE_X2Y112_BLUT (
.I0(LIOB33_X0Y113_IOB_X0Y113_I),
.I1(RIOB33_X105Y109_IOB_X1Y110_I),
.I2(RIOB33_X105Y111_IOB_X1Y111_I),
.I3(CLBLM_R_X5Y112_SLICE_X7Y112_DO6),
.I4(LIOB33_X0Y111_IOB_X0Y111_I),
.I5(LIOB33_X0Y111_IOB_X0Y112_I),
.O5(CLBLM_R_X3Y112_SLICE_X2Y112_BO5),
.O6(CLBLM_R_X3Y112_SLICE_X2Y112_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'ha5a5555596696699)
  ) CLBLM_R_X3Y112_SLICE_X2Y112_ALUT (
.I0(CLBLM_R_X3Y112_SLICE_X2Y112_BO6),
.I1(CLBLM_R_X5Y113_SLICE_X7Y113_CO6),
.I2(LIOB33_X0Y115_IOB_X0Y115_I),
.I3(CLBLL_L_X4Y113_SLICE_X4Y113_BO6),
.I4(RIOB33_X105Y109_IOB_X1Y110_I),
.I5(1'b1),
.O5(CLBLM_R_X3Y112_SLICE_X2Y112_AO5),
.O6(CLBLM_R_X3Y112_SLICE_X2Y112_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y112_SLICE_X3Y112_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y112_SLICE_X3Y112_DO5),
.O6(CLBLM_R_X3Y112_SLICE_X3Y112_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y112_SLICE_X3Y112_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y112_SLICE_X3Y112_CO5),
.O6(CLBLM_R_X3Y112_SLICE_X3Y112_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h133f77ff37ffffff)
  ) CLBLM_R_X3Y112_SLICE_X3Y112_BLUT (
.I0(LIOB33_X0Y113_IOB_X0Y113_I),
.I1(LIOB33_X0Y111_IOB_X0Y112_I),
.I2(LIOB33_X0Y111_IOB_X0Y111_I),
.I3(RIOB33_X105Y109_IOB_X1Y110_I),
.I4(RIOB33_X105Y111_IOB_X1Y111_I),
.I5(CLBLM_R_X5Y112_SLICE_X7Y112_DO6),
.O5(CLBLM_R_X3Y112_SLICE_X3Y112_BO5),
.O6(CLBLM_R_X3Y112_SLICE_X3Y112_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hbfd33f9f7f13ff5f)
  ) CLBLM_R_X3Y112_SLICE_X3Y112_ALUT (
.I0(LIOB33_X0Y113_IOB_X0Y113_I),
.I1(LIOB33_X0Y115_IOB_X0Y115_I),
.I2(RIOB33_X105Y111_IOB_X1Y111_I),
.I3(CLBLM_R_X3Y112_SLICE_X3Y112_BO6),
.I4(RIOB33_X105Y109_IOB_X1Y110_I),
.I5(1'b1),
.O5(CLBLM_R_X3Y112_SLICE_X3Y112_AO5),
.O6(CLBLM_R_X3Y112_SLICE_X3Y112_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h9a5965a6a5aaa5aa)
  ) CLBLM_R_X5Y104_SLICE_X6Y104_DLUT (
.I0(CLBLM_R_X7Y103_SLICE_X8Y103_DO6),
.I1(LIOB33_X0Y115_IOB_X0Y116_I),
.I2(CLBLL_L_X4Y104_SLICE_X5Y104_AO5),
.I3(CLBLM_R_X7Y104_SLICE_X8Y104_BO6),
.I4(LIOB33_X0Y117_IOB_X0Y117_I),
.I5(LIOB33_X0Y101_IOB_X0Y102_I),
.O5(CLBLM_R_X5Y104_SLICE_X6Y104_DO5),
.O6(CLBLM_R_X5Y104_SLICE_X6Y104_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h6a95956a956a956a)
  ) CLBLM_R_X5Y104_SLICE_X6Y104_CLUT (
.I0(CLBLM_R_X7Y103_SLICE_X8Y103_DO6),
.I1(LIOB33_X0Y115_IOB_X0Y116_I),
.I2(LIOB33_X0Y103_IOB_X0Y104_I),
.I3(CLBLL_L_X4Y103_SLICE_X5Y103_CO6),
.I4(LIOB33_X0Y117_IOB_X0Y117_I),
.I5(LIOB33_X0Y101_IOB_X0Y102_I),
.O5(CLBLM_R_X5Y104_SLICE_X6Y104_CO5),
.O6(CLBLM_R_X5Y104_SLICE_X6Y104_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h406f00a0505000a0)
  ) CLBLM_R_X5Y104_SLICE_X6Y104_BLUT (
.I0(LIOB33_SING_X0Y100_IOB_X0Y100_I),
.I1(RIOB33_X105Y111_IOB_X1Y112_I),
.I2(LIOB33_X0Y117_IOB_X0Y117_I),
.I3(LIOB33_X0Y115_IOB_X0Y116_I),
.I4(RIOB33_X105Y113_IOB_X1Y113_I),
.I5(RIOB33_X105Y101_IOB_X1Y101_I),
.O5(CLBLM_R_X5Y104_SLICE_X6Y104_BO5),
.O6(CLBLM_R_X5Y104_SLICE_X6Y104_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h00ffffff0fff0fff)
  ) CLBLM_R_X5Y104_SLICE_X6Y104_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(LIOB33_X0Y115_IOB_X0Y116_I),
.I3(LIOB33_X0Y103_IOB_X0Y104_I),
.I4(LIOB33_X0Y113_IOB_X0Y114_I),
.I5(1'b1),
.O5(CLBLM_R_X5Y104_SLICE_X6Y104_AO5),
.O6(CLBLM_R_X5Y104_SLICE_X6Y104_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X5Y104_SLICE_X7Y104_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y104_SLICE_X7Y104_DO5),
.O6(CLBLM_R_X5Y104_SLICE_X7Y104_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X5Y104_SLICE_X7Y104_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y104_SLICE_X7Y104_CO5),
.O6(CLBLM_R_X5Y104_SLICE_X7Y104_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h7ff7f7f707707070)
  ) CLBLM_R_X5Y104_SLICE_X7Y104_BLUT (
.I0(LIOB33_X0Y115_IOB_X0Y116_I),
.I1(LIOB33_X0Y103_IOB_X0Y104_I),
.I2(CLBLM_R_X7Y103_SLICE_X8Y103_DO6),
.I3(LIOB33_X0Y101_IOB_X0Y102_I),
.I4(LIOB33_X0Y117_IOB_X0Y117_I),
.I5(CLBLL_L_X4Y103_SLICE_X5Y103_CO6),
.O5(CLBLM_R_X5Y104_SLICE_X7Y104_BO5),
.O6(CLBLM_R_X5Y104_SLICE_X7Y104_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h39c6c6399c63639c)
  ) CLBLM_R_X5Y104_SLICE_X7Y104_ALUT (
.I0(CLBLM_R_X7Y104_SLICE_X8Y104_CO6),
.I1(CLBLM_L_X8Y104_SLICE_X10Y104_BO6),
.I2(CLBLM_R_X5Y104_SLICE_X6Y104_AO5),
.I3(CLBLM_R_X7Y104_SLICE_X9Y104_AO6),
.I4(CLBLM_R_X7Y104_SLICE_X8Y104_DO6),
.I5(CLBLL_L_X4Y103_SLICE_X5Y103_CO6),
.O5(CLBLM_R_X5Y104_SLICE_X7Y104_AO5),
.O6(CLBLM_R_X5Y104_SLICE_X7Y104_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h7fbfff3f152a3f00)
  ) CLBLM_R_X5Y105_SLICE_X6Y105_DLUT (
.I0(LIOB33_X0Y103_IOB_X0Y104_I),
.I1(LIOB33_X0Y113_IOB_X0Y114_I),
.I2(LIOB33_X0Y105_IOB_X0Y105_I),
.I3(CLBLM_R_X5Y104_SLICE_X6Y104_DO6),
.I4(LIOB33_X0Y115_IOB_X0Y116_I),
.I5(CLBLL_L_X4Y105_SLICE_X5Y105_AO6),
.O5(CLBLM_R_X5Y105_SLICE_X6Y105_DO5),
.O6(CLBLM_R_X5Y105_SLICE_X6Y105_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hb43cc3b478f00f78)
  ) CLBLM_R_X5Y105_SLICE_X6Y105_CLUT (
.I0(LIOB33_X0Y113_IOB_X0Y114_I),
.I1(LIOB33_X0Y105_IOB_X0Y106_I),
.I2(CLBLM_R_X7Y105_SLICE_X9Y105_CO6),
.I3(CLBLM_R_X7Y105_SLICE_X9Y105_DO6),
.I4(CLBLM_R_X5Y105_SLICE_X6Y105_DO6),
.I5(LIOB33_X0Y115_IOB_X0Y116_I),
.O5(CLBLM_R_X5Y105_SLICE_X6Y105_CO5),
.O6(CLBLM_R_X5Y105_SLICE_X6Y105_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h6a95c03f956a3fc0)
  ) CLBLM_R_X5Y105_SLICE_X6Y105_BLUT (
.I0(LIOB33_X0Y105_IOB_X0Y105_I),
.I1(LIOB33_X0Y115_IOB_X0Y116_I),
.I2(LIOB33_X0Y103_IOB_X0Y104_I),
.I3(CLBLM_R_X5Y104_SLICE_X6Y104_DO6),
.I4(LIOB33_X0Y113_IOB_X0Y114_I),
.I5(CLBLL_L_X4Y105_SLICE_X5Y105_AO6),
.O5(CLBLM_R_X5Y105_SLICE_X6Y105_BO5),
.O6(CLBLM_R_X5Y105_SLICE_X6Y105_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hd2785af0b41e963c)
  ) CLBLM_R_X5Y105_SLICE_X6Y105_ALUT (
.I0(LIOB33_X0Y105_IOB_X0Y105_I),
.I1(CLBLM_R_X5Y104_SLICE_X6Y104_CO6),
.I2(CLBLM_R_X5Y104_SLICE_X7Y104_AO6),
.I3(LIOB33_X0Y115_IOB_X0Y116_I),
.I4(LIOB33_X0Y113_IOB_X0Y114_I),
.I5(CLBLL_L_X4Y105_SLICE_X5Y105_AO6),
.O5(CLBLM_R_X5Y105_SLICE_X6Y105_AO5),
.O6(CLBLM_R_X5Y105_SLICE_X6Y105_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X5Y105_SLICE_X7Y105_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y105_SLICE_X7Y105_DO5),
.O6(CLBLM_R_X5Y105_SLICE_X7Y105_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'he8b2eebb8822e8b2)
  ) CLBLM_R_X5Y105_SLICE_X7Y105_CLUT (
.I0(CLBLM_R_X5Y105_SLICE_X7Y105_AO6),
.I1(CLBLM_R_X5Y106_SLICE_X7Y106_AO6),
.I2(CLBLM_R_X5Y106_SLICE_X7Y106_AO5),
.I3(CLBLM_R_X5Y104_SLICE_X7Y104_AO6),
.I4(CLBLM_R_X5Y104_SLICE_X6Y104_CO6),
.I5(CLBLL_L_X4Y105_SLICE_X5Y105_AO6),
.O5(CLBLM_R_X5Y105_SLICE_X7Y105_CO5),
.O6(CLBLM_R_X5Y105_SLICE_X7Y105_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h3c96c36996c3693c)
  ) CLBLM_R_X5Y105_SLICE_X7Y105_BLUT (
.I0(CLBLM_R_X5Y104_SLICE_X6Y104_CO6),
.I1(CLBLM_R_X5Y106_SLICE_X7Y106_AO6),
.I2(CLBLM_R_X5Y104_SLICE_X7Y104_AO6),
.I3(CLBLL_L_X4Y105_SLICE_X5Y105_AO6),
.I4(CLBLM_R_X5Y105_SLICE_X7Y105_AO6),
.I5(CLBLM_R_X5Y106_SLICE_X7Y106_AO5),
.O5(CLBLM_R_X5Y105_SLICE_X7Y105_BO5),
.O6(CLBLM_R_X5Y105_SLICE_X7Y105_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h5f5f5f5f0f0fffff)
  ) CLBLM_R_X5Y105_SLICE_X7Y105_ALUT (
.I0(LIOB33_X0Y113_IOB_X0Y114_I),
.I1(1'b1),
.I2(LIOB33_X0Y105_IOB_X0Y106_I),
.I3(1'b1),
.I4(LIOB33_X0Y103_IOB_X0Y103_I),
.I5(1'b1),
.O5(CLBLM_R_X5Y105_SLICE_X7Y105_AO5),
.O6(CLBLM_R_X5Y105_SLICE_X7Y105_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hefae8a088a08efae)
  ) CLBLM_R_X5Y106_SLICE_X6Y106_DLUT (
.I0(CLBLM_R_X5Y106_SLICE_X6Y106_AO6),
.I1(CLBLL_L_X4Y107_SLICE_X5Y107_AO6),
.I2(CLBLM_R_X5Y106_SLICE_X7Y106_DO6),
.I3(CLBLL_L_X4Y106_SLICE_X5Y106_BO6),
.I4(CLBLM_R_X7Y106_SLICE_X8Y106_AO5),
.I5(CLBLM_R_X7Y106_SLICE_X8Y106_BO6),
.O5(CLBLM_R_X5Y106_SLICE_X6Y106_DO5),
.O6(CLBLM_R_X5Y106_SLICE_X6Y106_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h65a69a599a5965a6)
  ) CLBLM_R_X5Y106_SLICE_X6Y106_CLUT (
.I0(CLBLM_R_X5Y106_SLICE_X6Y106_AO6),
.I1(CLBLL_L_X4Y107_SLICE_X5Y107_AO6),
.I2(CLBLM_R_X5Y106_SLICE_X7Y106_DO6),
.I3(CLBLL_L_X4Y106_SLICE_X5Y106_BO6),
.I4(CLBLM_R_X7Y106_SLICE_X8Y106_AO5),
.I5(CLBLM_R_X7Y106_SLICE_X8Y106_BO6),
.O5(CLBLM_R_X5Y106_SLICE_X6Y106_CO5),
.O6(CLBLM_R_X5Y106_SLICE_X6Y106_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hd728b14e5fa0936c)
  ) CLBLM_R_X5Y106_SLICE_X6Y106_BLUT (
.I0(LIOB33_X0Y107_IOB_X0Y108_I),
.I1(CLBLM_R_X5Y106_SLICE_X7Y106_DO6),
.I2(LIOB33_X0Y113_IOB_X0Y114_I),
.I3(CLBLM_R_X7Y106_SLICE_X8Y106_BO6),
.I4(CLBLL_L_X4Y106_SLICE_X5Y106_BO6),
.I5(LIOB33_X0Y103_IOB_X0Y103_I),
.O5(CLBLM_R_X5Y106_SLICE_X6Y106_BO5),
.O6(CLBLM_R_X5Y106_SLICE_X6Y106_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h00ffffff0fff0fff)
  ) CLBLM_R_X5Y106_SLICE_X6Y106_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(LIOB33_X0Y113_IOB_X0Y114_I),
.I3(LIOB33_X0Y109_IOB_X0Y109_I),
.I4(LIOB33_X0Y103_IOB_X0Y103_I),
.I5(1'b1),
.O5(CLBLM_R_X5Y106_SLICE_X6Y106_AO5),
.O6(CLBLM_R_X5Y106_SLICE_X6Y106_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h6c93936c936c936c)
  ) CLBLM_R_X5Y106_SLICE_X7Y106_DLUT (
.I0(LIOB33_X0Y107_IOB_X0Y107_I),
.I1(CLBLM_R_X7Y105_SLICE_X9Y105_CO6),
.I2(LIOB33_X0Y113_IOB_X0Y114_I),
.I3(CLBLM_R_X5Y105_SLICE_X7Y105_CO6),
.I4(LIOB33_X0Y115_IOB_X0Y116_I),
.I5(LIOB33_X0Y105_IOB_X0Y106_I),
.O5(CLBLM_R_X5Y106_SLICE_X7Y106_DO5),
.O6(CLBLM_R_X5Y106_SLICE_X7Y106_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h639cc6399c6339c6)
  ) CLBLM_R_X5Y106_SLICE_X7Y106_CLUT (
.I0(CLBLL_L_X4Y105_SLICE_X5Y105_BO6),
.I1(CLBLM_R_X7Y105_SLICE_X9Y105_AO6),
.I2(CLBLM_R_X5Y105_SLICE_X7Y105_BO6),
.I3(CLBLM_R_X5Y105_SLICE_X7Y105_CO6),
.I4(CLBLM_R_X5Y106_SLICE_X7Y106_BO5),
.I5(CLBLM_R_X5Y106_SLICE_X7Y106_BO6),
.O5(CLBLM_R_X5Y106_SLICE_X7Y106_CO5),
.O6(CLBLM_R_X5Y106_SLICE_X7Y106_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h5555ffff0f0fffff)
  ) CLBLM_R_X5Y106_SLICE_X7Y106_BLUT (
.I0(LIOB33_X0Y113_IOB_X0Y114_I),
.I1(1'b1),
.I2(LIOB33_X0Y103_IOB_X0Y103_I),
.I3(1'b1),
.I4(LIOB33_X0Y107_IOB_X0Y107_I),
.I5(1'b1),
.O5(CLBLM_R_X5Y106_SLICE_X7Y106_BO5),
.O6(CLBLM_R_X5Y106_SLICE_X7Y106_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0fff0fff5f5f5f5f)
  ) CLBLM_R_X5Y106_SLICE_X7Y106_ALUT (
.I0(LIOB33_X0Y113_IOB_X0Y114_I),
.I1(1'b1),
.I2(LIOB33_X0Y105_IOB_X0Y105_I),
.I3(LIOB33_X0Y115_IOB_X0Y116_I),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y106_SLICE_X7Y106_AO5),
.O6(CLBLM_R_X5Y106_SLICE_X7Y106_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hac536c936f905fa0)
  ) CLBLM_R_X5Y107_SLICE_X6Y107_DLUT (
.I0(LIOB33_X0Y109_IOB_X0Y110_I),
.I1(CLBLL_L_X4Y107_SLICE_X4Y107_CO6),
.I2(RIOB33_X105Y105_IOB_X1Y106_I),
.I3(CLBLM_R_X5Y106_SLICE_X6Y106_CO6),
.I4(LIOB33_X0Y109_IOB_X0Y109_I),
.I5(CLBLL_L_X4Y106_SLICE_X5Y106_CO6),
.O5(CLBLM_R_X5Y107_SLICE_X6Y107_DO5),
.O6(CLBLM_R_X5Y107_SLICE_X6Y107_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h6969966996699696)
  ) CLBLM_R_X5Y107_SLICE_X6Y107_CLUT (
.I0(CLBLM_R_X7Y106_SLICE_X9Y106_BO6),
.I1(CLBLM_R_X5Y107_SLICE_X7Y107_AO6),
.I2(CLBLM_R_X5Y106_SLICE_X6Y106_DO6),
.I3(CLBLM_R_X5Y106_SLICE_X6Y106_CO6),
.I4(CLBLM_R_X3Y107_SLICE_X3Y107_BO5),
.I5(CLBLL_L_X4Y107_SLICE_X5Y107_DO6),
.O5(CLBLM_R_X5Y107_SLICE_X6Y107_CO5),
.O6(CLBLM_R_X5Y107_SLICE_X6Y107_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h445d4c5f5fdfdfff)
  ) CLBLM_R_X5Y107_SLICE_X6Y107_BLUT (
.I0(RIOB33_X105Y105_IOB_X1Y106_I),
.I1(CLBLL_L_X4Y107_SLICE_X4Y107_CO6),
.I2(LIOB33_X0Y109_IOB_X0Y110_I),
.I3(CLBLL_L_X4Y106_SLICE_X5Y106_CO6),
.I4(LIOB33_X0Y109_IOB_X0Y109_I),
.I5(CLBLM_R_X5Y106_SLICE_X6Y106_CO6),
.O5(CLBLM_R_X5Y107_SLICE_X6Y107_BO5),
.O6(CLBLM_R_X5Y107_SLICE_X6Y107_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h9cc36c333c9ccc6c)
  ) CLBLM_R_X5Y107_SLICE_X6Y107_ALUT (
.I0(RIOB33_X105Y105_IOB_X1Y106_I),
.I1(CLBLM_R_X5Y106_SLICE_X6Y106_BO6),
.I2(LIOB33_X0Y109_IOB_X0Y109_I),
.I3(CLBLL_L_X4Y107_SLICE_X4Y107_CO6),
.I4(LIOB33_X0Y103_IOB_X0Y103_I),
.I5(CLBLL_L_X4Y106_SLICE_X5Y106_CO6),
.O5(CLBLM_R_X5Y107_SLICE_X6Y107_AO5),
.O6(CLBLM_R_X5Y107_SLICE_X6Y107_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X5Y107_SLICE_X7Y107_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y107_SLICE_X7Y107_DO5),
.O6(CLBLM_R_X5Y107_SLICE_X7Y107_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0b2b0bbb2fffbfff)
  ) CLBLM_R_X5Y107_SLICE_X7Y107_CLUT (
.I0(CLBLL_L_X4Y106_SLICE_X5Y106_DO6),
.I1(CLBLM_R_X7Y105_SLICE_X8Y105_CO6),
.I2(LIOB33_X0Y103_IOB_X0Y103_I),
.I3(LIOB33_X0Y109_IOB_X0Y110_I),
.I4(LIOB33_X0Y109_IOB_X0Y109_I),
.I5(CLBLM_R_X7Y106_SLICE_X9Y106_BO6),
.O5(CLBLM_R_X5Y107_SLICE_X7Y107_CO5),
.O6(CLBLM_R_X5Y107_SLICE_X7Y107_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h8f70e31c7f8013ec)
  ) CLBLM_R_X5Y107_SLICE_X7Y107_BLUT (
.I0(LIOB33_X0Y103_IOB_X0Y103_I),
.I1(CLBLM_R_X7Y105_SLICE_X8Y105_CO6),
.I2(LIOB33_X0Y109_IOB_X0Y109_I),
.I3(CLBLM_R_X7Y106_SLICE_X9Y106_AO6),
.I4(CLBLL_L_X4Y106_SLICE_X5Y106_DO6),
.I5(LIOB33_X0Y113_IOB_X0Y114_I),
.O5(CLBLM_R_X5Y107_SLICE_X7Y107_BO5),
.O6(CLBLM_R_X5Y107_SLICE_X7Y107_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h5555ffff5f5f5f5f)
  ) CLBLM_R_X5Y107_SLICE_X7Y107_ALUT (
.I0(LIOB33_X0Y109_IOB_X0Y110_I),
.I1(1'b1),
.I2(LIOB33_X0Y113_IOB_X0Y114_I),
.I3(1'b1),
.I4(LIOB33_X0Y103_IOB_X0Y103_I),
.I5(1'b1),
.O5(CLBLM_R_X5Y107_SLICE_X7Y107_AO5),
.O6(CLBLM_R_X5Y107_SLICE_X7Y107_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X5Y108_SLICE_X6Y108_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y108_SLICE_X6Y108_DO5),
.O6(CLBLM_R_X5Y108_SLICE_X6Y108_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hebc38200ffebc382)
  ) CLBLM_R_X5Y108_SLICE_X6Y108_CLUT (
.I0(CLBLL_L_X4Y107_SLICE_X4Y107_BO6),
.I1(CLBLM_R_X5Y107_SLICE_X6Y107_CO6),
.I2(CLBLM_R_X5Y108_SLICE_X7Y108_AO6),
.I3(CLBLM_R_X5Y110_SLICE_X6Y110_AO6),
.I4(CLBLM_R_X5Y110_SLICE_X7Y110_AO6),
.I5(CLBLM_R_X5Y107_SLICE_X6Y107_DO6),
.O5(CLBLM_R_X5Y108_SLICE_X6Y108_CO5),
.O6(CLBLM_R_X5Y108_SLICE_X6Y108_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h4dddd444cffffccc)
  ) CLBLM_R_X5Y108_SLICE_X6Y108_BLUT (
.I0(RIOB33_X105Y105_IOB_X1Y106_I),
.I1(CLBLM_R_X5Y107_SLICE_X6Y107_BO6),
.I2(LIOB33_X0Y109_IOB_X0Y110_I),
.I3(LIOB33_X0Y103_IOB_X0Y103_I),
.I4(CLBLM_R_X5Y107_SLICE_X7Y107_BO6),
.I5(LIOB33_X0Y111_IOB_X0Y111_I),
.O5(CLBLM_R_X5Y108_SLICE_X6Y108_BO5),
.O6(CLBLM_R_X5Y108_SLICE_X6Y108_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h7887877888777788)
  ) CLBLM_R_X5Y108_SLICE_X6Y108_ALUT (
.I0(RIOB33_X105Y105_IOB_X1Y106_I),
.I1(LIOB33_X0Y111_IOB_X0Y111_I),
.I2(LIOB33_X0Y109_IOB_X0Y110_I),
.I3(CLBLM_R_X5Y107_SLICE_X6Y107_BO6),
.I4(CLBLM_R_X5Y107_SLICE_X7Y107_BO6),
.I5(LIOB33_X0Y103_IOB_X0Y103_I),
.O5(CLBLM_R_X5Y108_SLICE_X6Y108_AO5),
.O6(CLBLM_R_X5Y108_SLICE_X6Y108_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X5Y108_SLICE_X7Y108_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y108_SLICE_X7Y108_DO5),
.O6(CLBLM_R_X5Y108_SLICE_X7Y108_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h69a5c30f965a3cf0)
  ) CLBLM_R_X5Y108_SLICE_X7Y108_CLUT (
.I0(LIOB33_X0Y109_IOB_X0Y110_I),
.I1(LIOB33_X0Y111_IOB_X0Y111_I),
.I2(CLBLM_R_X7Y108_SLICE_X9Y108_DO6),
.I3(LIOB33_X0Y113_IOB_X0Y114_I),
.I4(LIOB33_X0Y115_IOB_X0Y116_I),
.I5(CLBLM_R_X7Y107_SLICE_X9Y107_DO6),
.O5(CLBLM_R_X5Y108_SLICE_X7Y108_CO5),
.O6(CLBLM_R_X5Y108_SLICE_X7Y108_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h4dd4dd44cffcffcc)
  ) CLBLM_R_X5Y108_SLICE_X7Y108_BLUT (
.I0(LIOB33_X0Y111_IOB_X0Y111_I),
.I1(CLBLM_R_X7Y107_SLICE_X9Y107_DO6),
.I2(LIOB33_X0Y109_IOB_X0Y110_I),
.I3(CLBLM_R_X7Y108_SLICE_X9Y108_DO6),
.I4(LIOB33_X0Y115_IOB_X0Y116_I),
.I5(LIOB33_X0Y113_IOB_X0Y114_I),
.O5(CLBLM_R_X5Y108_SLICE_X7Y108_BO5),
.O6(CLBLM_R_X5Y108_SLICE_X7Y108_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h55ff55ff00ffffff)
  ) CLBLM_R_X5Y108_SLICE_X7Y108_ALUT (
.I0(RIOB33_X105Y105_IOB_X1Y106_I),
.I1(1'b1),
.I2(1'b1),
.I3(LIOB33_X0Y111_IOB_X0Y111_I),
.I4(LIOB33_X0Y103_IOB_X0Y103_I),
.I5(1'b1),
.O5(CLBLM_R_X5Y108_SLICE_X7Y108_AO5),
.O6(CLBLM_R_X5Y108_SLICE_X7Y108_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X5Y109_SLICE_X6Y109_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y109_SLICE_X6Y109_DO5),
.O6(CLBLM_R_X5Y109_SLICE_X6Y109_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X5Y109_SLICE_X6Y109_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y109_SLICE_X6Y109_CO5),
.O6(CLBLM_R_X5Y109_SLICE_X6Y109_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X5Y109_SLICE_X6Y109_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y109_SLICE_X6Y109_BO5),
.O6(CLBLM_R_X5Y109_SLICE_X6Y109_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X5Y109_SLICE_X6Y109_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y109_SLICE_X6Y109_AO5),
.O6(CLBLM_R_X5Y109_SLICE_X6Y109_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X5Y109_SLICE_X7Y109_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y109_SLICE_X7Y109_DO5),
.O6(CLBLM_R_X5Y109_SLICE_X7Y109_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X5Y109_SLICE_X7Y109_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y109_SLICE_X7Y109_CO5),
.O6(CLBLM_R_X5Y109_SLICE_X7Y109_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0d4f0ddf4dffddff)
  ) CLBLM_R_X5Y109_SLICE_X7Y109_BLUT (
.I0(CLBLM_R_X7Y109_SLICE_X8Y109_CO6),
.I1(CLBLM_R_X5Y108_SLICE_X7Y108_BO6),
.I2(LIOB33_X0Y113_IOB_X0Y114_I),
.I3(CLBLM_R_X7Y109_SLICE_X8Y109_DO6),
.I4(LIOB33_X0Y111_IOB_X0Y112_I),
.I5(LIOB33_X0Y113_IOB_X0Y113_I),
.O5(CLBLM_R_X5Y109_SLICE_X7Y109_BO5),
.O6(CLBLM_R_X5Y109_SLICE_X7Y109_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h96c3cc663c96cc66)
  ) CLBLM_R_X5Y109_SLICE_X7Y109_ALUT (
.I0(CLBLM_R_X7Y109_SLICE_X8Y109_CO6),
.I1(CLBLM_R_X7Y109_SLICE_X8Y109_BO6),
.I2(LIOB33_X0Y115_IOB_X0Y116_I),
.I3(CLBLM_R_X5Y108_SLICE_X7Y108_BO6),
.I4(LIOB33_X0Y111_IOB_X0Y112_I),
.I5(LIOB33_X0Y113_IOB_X0Y114_I),
.O5(CLBLM_R_X5Y109_SLICE_X7Y109_AO5),
.O6(CLBLM_R_X5Y109_SLICE_X7Y109_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h00000000f0f0f0f0)
  ) CLBLM_R_X5Y110_SLICE_X6Y110_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(CLBLM_R_X5Y108_SLICE_X6Y108_BO6),
.I3(1'b1),
.I4(1'b1),
.I5(CLBLM_R_X7Y107_SLICE_X8Y107_AO6),
.O5(CLBLM_R_X5Y110_SLICE_X6Y110_DO5),
.O6(CLBLM_R_X5Y110_SLICE_X6Y110_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0ff00ff00ff08ff0)
  ) CLBLM_R_X5Y110_SLICE_X6Y110_CLUT (
.I0(CLBLM_L_X8Y110_SLICE_X10Y110_CO6),
.I1(CLBLM_R_X7Y110_SLICE_X8Y110_CO6),
.I2(CLBLM_R_X5Y112_SLICE_X6Y112_AO5),
.I3(CLBLM_R_X5Y111_SLICE_X6Y111_CO6),
.I4(CLBLM_R_X5Y110_SLICE_X6Y110_DO6),
.I5(CLBLM_R_X5Y110_SLICE_X6Y110_BO6),
.O5(CLBLM_R_X5Y110_SLICE_X6Y110_CO5),
.O6(CLBLM_R_X5Y110_SLICE_X6Y110_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h05055555965a66aa)
  ) CLBLM_R_X5Y110_SLICE_X6Y110_BLUT (
.I0(CLBLM_R_X5Y112_SLICE_X7Y112_DO6),
.I1(RIOB33_X105Y109_IOB_X1Y110_I),
.I2(LIOB33_X0Y111_IOB_X0Y111_I),
.I3(LIOB33_X0Y111_IOB_X0Y112_I),
.I4(RIOB33_X105Y111_IOB_X1Y111_I),
.I5(1'b1),
.O5(CLBLM_R_X5Y110_SLICE_X6Y110_BO5),
.O6(CLBLM_R_X5Y110_SLICE_X6Y110_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h3333ffffa5a55555)
  ) CLBLM_R_X5Y110_SLICE_X6Y110_ALUT (
.I0(CLBLM_L_X8Y111_SLICE_X11Y111_BO6),
.I1(RIOB33_SING_X105Y100_IOB_X1Y100_I),
.I2(RIOB33_X105Y103_IOB_X1Y104_I),
.I3(1'b1),
.I4(LIOB33_X0Y111_IOB_X0Y111_I),
.I5(1'b1),
.O5(CLBLM_R_X5Y110_SLICE_X6Y110_AO5),
.O6(CLBLM_R_X5Y110_SLICE_X6Y110_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h517175ff51f3f7ff)
  ) CLBLM_R_X5Y110_SLICE_X7Y110_DLUT (
.I0(RIOB33_X105Y101_IOB_X1Y102_I),
.I1(CLBLM_R_X7Y111_SLICE_X8Y111_AO6),
.I2(CLBLM_L_X8Y112_SLICE_X11Y112_DO6),
.I3(LIOB33_X0Y113_IOB_X0Y113_I),
.I4(CLBLM_R_X5Y110_SLICE_X7Y110_BO5),
.I5(LIOB33_X0Y111_IOB_X0Y112_I),
.O5(CLBLM_R_X5Y110_SLICE_X7Y110_DO5),
.O6(CLBLM_R_X5Y110_SLICE_X7Y110_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'ha96a696665a6a5aa)
  ) CLBLM_R_X5Y110_SLICE_X7Y110_CLUT (
.I0(CLBLM_R_X7Y111_SLICE_X8Y111_BO6),
.I1(LIOB33_X0Y111_IOB_X0Y112_I),
.I2(CLBLM_L_X8Y112_SLICE_X11Y112_DO6),
.I3(CLBLM_R_X7Y111_SLICE_X8Y111_AO6),
.I4(RIOB33_X105Y101_IOB_X1Y102_I),
.I5(RIOB33_X105Y103_IOB_X1Y103_I),
.O5(CLBLM_R_X5Y110_SLICE_X7Y110_CO5),
.O6(CLBLM_R_X5Y110_SLICE_X7Y110_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0fff0fffcc0033ff)
  ) CLBLM_R_X5Y110_SLICE_X7Y110_BLUT (
.I0(1'b1),
.I1(RIOB33_X105Y103_IOB_X1Y103_I),
.I2(LIOB33_X0Y103_IOB_X0Y103_I),
.I3(LIOB33_X0Y111_IOB_X0Y112_I),
.I4(CLBLM_R_X7Y111_SLICE_X8Y111_BO6),
.I5(1'b1),
.O5(CLBLM_R_X5Y110_SLICE_X7Y110_BO5),
.O6(CLBLM_R_X5Y110_SLICE_X7Y110_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0fff0fff69699999)
  ) CLBLM_R_X5Y110_SLICE_X7Y110_ALUT (
.I0(CLBLM_R_X7Y110_SLICE_X9Y110_AO5),
.I1(CLBLM_R_X7Y111_SLICE_X9Y111_AO6),
.I2(LIOB33_X0Y111_IOB_X0Y112_I),
.I3(RIOB33_SING_X105Y100_IOB_X1Y100_I),
.I4(RIOB33_X105Y107_IOB_X1Y108_I),
.I5(1'b1),
.O5(CLBLM_R_X5Y110_SLICE_X7Y110_AO5),
.O6(CLBLM_R_X5Y110_SLICE_X7Y110_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'haf0a0f0050f5f0ff)
  ) CLBLM_R_X5Y111_SLICE_X6Y111_DLUT (
.I0(LIOB33_X0Y111_IOB_X0Y112_I),
.I1(1'b1),
.I2(CLBLM_R_X7Y111_SLICE_X8Y111_AO5),
.I3(CLBLM_R_X5Y110_SLICE_X6Y110_AO5),
.I4(RIOB33_X105Y103_IOB_X1Y103_I),
.I5(CLBLM_L_X8Y113_SLICE_X10Y113_BO6),
.O5(CLBLM_R_X5Y111_SLICE_X6Y111_DO5),
.O6(CLBLM_R_X5Y111_SLICE_X6Y111_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h57157f1f5f17ff3f)
  ) CLBLM_R_X5Y111_SLICE_X6Y111_CLUT (
.I0(RIOB33_X105Y107_IOB_X1Y108_I),
.I1(CLBLM_R_X7Y111_SLICE_X9Y111_AO6),
.I2(CLBLM_R_X5Y111_SLICE_X7Y111_AO6),
.I3(CLBLM_R_X7Y110_SLICE_X9Y110_AO5),
.I4(LIOB33_X0Y113_IOB_X0Y113_I),
.I5(LIOB33_X0Y111_IOB_X0Y112_I),
.O5(CLBLM_R_X5Y111_SLICE_X6Y111_CO5),
.O6(CLBLM_R_X5Y111_SLICE_X6Y111_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h307770f773f777ff)
  ) CLBLM_R_X5Y111_SLICE_X6Y111_BLUT (
.I0(LIOB33_X0Y113_IOB_X0Y113_I),
.I1(RIOB33_X105Y103_IOB_X1Y103_I),
.I2(CLBLM_R_X7Y111_SLICE_X8Y111_AO5),
.I3(CLBLM_L_X8Y113_SLICE_X10Y113_BO6),
.I4(LIOB33_X0Y111_IOB_X0Y112_I),
.I5(CLBLM_R_X5Y110_SLICE_X6Y110_AO5),
.O5(CLBLM_R_X5Y111_SLICE_X6Y111_BO5),
.O6(CLBLM_R_X5Y111_SLICE_X6Y111_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h69c3a50f963c5af0)
  ) CLBLM_R_X5Y111_SLICE_X6Y111_ALUT (
.I0(LIOB33_X0Y113_IOB_X0Y113_I),
.I1(RIOB33_X105Y101_IOB_X1Y101_I),
.I2(CLBLM_R_X5Y110_SLICE_X7Y110_CO6),
.I3(RIOB33_X105Y101_IOB_X1Y102_I),
.I4(LIOB33_X0Y115_IOB_X0Y115_I),
.I5(CLBLM_R_X7Y112_SLICE_X8Y112_CO6),
.O5(CLBLM_R_X5Y111_SLICE_X6Y111_AO5),
.O6(CLBLM_R_X5Y111_SLICE_X6Y111_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h2a80bfeabfeabfea)
  ) CLBLM_R_X5Y111_SLICE_X7Y111_DLUT (
.I0(CLBLM_R_X7Y111_SLICE_X9Y111_AO5),
.I1(LIOB33_X0Y111_IOB_X0Y111_I),
.I2(RIOB33_X105Y109_IOB_X1Y110_I),
.I3(CLBLM_R_X5Y111_SLICE_X7Y111_CO6),
.I4(RIOB33_X105Y109_IOB_X1Y109_I),
.I5(LIOB33_X0Y111_IOB_X0Y112_I),
.O5(CLBLM_R_X5Y111_SLICE_X7Y111_DO5),
.O6(CLBLM_R_X5Y111_SLICE_X7Y111_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hb5ad2d0fdfdfffff)
  ) CLBLM_R_X5Y111_SLICE_X7Y111_CLUT (
.I0(LIOB33_X0Y109_IOB_X0Y109_I),
.I1(CLBLM_R_X7Y111_SLICE_X9Y111_CO6),
.I2(LIOB33_X0Y109_IOB_X0Y110_I),
.I3(LIOB33_X0Y107_IOB_X0Y108_I),
.I4(RIOB33_X105Y109_IOB_X1Y110_I),
.I5(RIOB33_X105Y111_IOB_X1Y111_I),
.O5(CLBLM_R_X5Y111_SLICE_X7Y111_CO5),
.O6(CLBLM_R_X5Y111_SLICE_X7Y111_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hac6c6f5f539390a0)
  ) CLBLM_R_X5Y111_SLICE_X7Y111_BLUT (
.I0(LIOB33_X0Y113_IOB_X0Y113_I),
.I1(CLBLM_R_X7Y110_SLICE_X9Y110_AO5),
.I2(RIOB33_X105Y107_IOB_X1Y108_I),
.I3(LIOB33_X0Y111_IOB_X0Y112_I),
.I4(CLBLM_R_X7Y111_SLICE_X9Y111_AO6),
.I5(CLBLM_R_X5Y111_SLICE_X7Y111_AO6),
.O5(CLBLM_R_X5Y111_SLICE_X7Y111_BO5),
.O6(CLBLM_R_X5Y111_SLICE_X7Y111_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h6a95c03f956a3fc0)
  ) CLBLM_R_X5Y111_SLICE_X7Y111_ALUT (
.I0(RIOB33_X105Y109_IOB_X1Y109_I),
.I1(RIOB33_X105Y109_IOB_X1Y110_I),
.I2(LIOB33_X0Y111_IOB_X0Y111_I),
.I3(CLBLM_R_X7Y111_SLICE_X9Y111_AO5),
.I4(LIOB33_X0Y111_IOB_X0Y112_I),
.I5(CLBLM_R_X5Y111_SLICE_X7Y111_CO6),
.O5(CLBLM_R_X5Y111_SLICE_X7Y111_AO5),
.O6(CLBLM_R_X5Y111_SLICE_X7Y111_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h00cc00cc00cc00cc)
  ) CLBLM_R_X5Y112_SLICE_X6Y112_DLUT (
.I0(1'b1),
.I1(CLBLM_R_X5Y111_SLICE_X6Y111_CO6),
.I2(1'b1),
.I3(CLBLM_R_X5Y112_SLICE_X6Y112_AO5),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y112_SLICE_X6Y112_DO5),
.O6(CLBLM_R_X5Y112_SLICE_X6Y112_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h7887877887788778)
  ) CLBLM_R_X5Y112_SLICE_X6Y112_CLUT (
.I0(LIOB33_X0Y111_IOB_X0Y111_I),
.I1(RIOB33_X105Y111_IOB_X1Y111_I),
.I2(CLBLM_R_X5Y112_SLICE_X7Y112_DO6),
.I3(CLBLM_R_X5Y111_SLICE_X7Y111_DO6),
.I4(RIOB33_X105Y109_IOB_X1Y110_I),
.I5(LIOB33_X0Y111_IOB_X0Y112_I),
.O5(CLBLM_R_X5Y112_SLICE_X6Y112_CO5),
.O6(CLBLM_R_X5Y112_SLICE_X6Y112_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h6999a55596665aaa)
  ) CLBLM_R_X5Y112_SLICE_X6Y112_BLUT (
.I0(CLBLM_R_X5Y111_SLICE_X6Y111_DO6),
.I1(LIOB33_X0Y113_IOB_X0Y113_I),
.I2(RIOB33_X105Y101_IOB_X1Y102_I),
.I3(LIOB33_X0Y115_IOB_X0Y115_I),
.I4(RIOB33_X105Y103_IOB_X1Y103_I),
.I5(CLBLM_R_X5Y110_SLICE_X7Y110_DO6),
.O5(CLBLM_R_X5Y112_SLICE_X6Y112_BO5),
.O6(CLBLM_R_X5Y112_SLICE_X6Y112_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h99559955f0000fff)
  ) CLBLM_R_X5Y112_SLICE_X6Y112_ALUT (
.I0(CLBLM_R_X5Y111_SLICE_X6Y111_DO6),
.I1(RIOB33_X105Y103_IOB_X1Y103_I),
.I2(RIOB33_X105Y109_IOB_X1Y109_I),
.I3(LIOB33_X0Y113_IOB_X0Y113_I),
.I4(CLBLM_R_X5Y112_SLICE_X6Y112_CO6),
.I5(1'b1),
.O5(CLBLM_R_X5Y112_SLICE_X6Y112_AO5),
.O6(CLBLM_R_X5Y112_SLICE_X6Y112_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h88000000eeccaa00)
  ) CLBLM_R_X5Y112_SLICE_X7Y112_DLUT (
.I0(LIOB33_X0Y111_IOB_X0Y111_I),
.I1(LIOB33_X0Y109_IOB_X0Y110_I),
.I2(1'b1),
.I3(RIOB33_X105Y109_IOB_X1Y110_I),
.I4(RIOB33_X105Y111_IOB_X1Y111_I),
.I5(CLBLM_R_X5Y112_SLICE_X7Y112_BO6),
.O5(CLBLM_R_X5Y112_SLICE_X7Y112_DO5),
.O6(CLBLM_R_X5Y112_SLICE_X7Y112_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hd10cb7c06ac0c0c0)
  ) CLBLM_R_X5Y112_SLICE_X7Y112_CLUT (
.I0(LIOB33_X0Y111_IOB_X0Y111_I),
.I1(RIOB33_X105Y109_IOB_X1Y110_I),
.I2(LIOB33_X0Y113_IOB_X0Y113_I),
.I3(RIOB33_X105Y111_IOB_X1Y111_I),
.I4(CLBLM_R_X5Y112_SLICE_X7Y112_DO6),
.I5(LIOB33_X0Y111_IOB_X0Y112_I),
.O5(CLBLM_R_X5Y112_SLICE_X7Y112_CO5),
.O6(CLBLM_R_X5Y112_SLICE_X7Y112_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h77ff137f7fff777f)
  ) CLBLM_R_X5Y112_SLICE_X7Y112_BLUT (
.I0(RIOB33_X105Y111_IOB_X1Y111_I),
.I1(LIOB33_X0Y109_IOB_X0Y109_I),
.I2(LIOB33_X0Y107_IOB_X0Y108_I),
.I3(RIOB33_X105Y109_IOB_X1Y110_I),
.I4(CLBLM_R_X7Y111_SLICE_X9Y111_CO6),
.I5(LIOB33_X0Y109_IOB_X0Y110_I),
.O5(CLBLM_R_X5Y112_SLICE_X7Y112_BO5),
.O6(CLBLM_R_X5Y112_SLICE_X7Y112_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0fff0fff33ff33ff)
  ) CLBLM_R_X5Y112_SLICE_X7Y112_ALUT (
.I0(1'b1),
.I1(LIOB33_X0Y115_IOB_X0Y115_I),
.I2(LIOB33_X0Y111_IOB_X0Y111_I),
.I3(RIOB33_X105Y101_IOB_X1Y102_I),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y112_SLICE_X7Y112_AO5),
.O6(CLBLM_R_X5Y112_SLICE_X7Y112_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X5Y113_SLICE_X6Y113_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y113_SLICE_X6Y113_DO5),
.O6(CLBLM_R_X5Y113_SLICE_X6Y113_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X5Y113_SLICE_X6Y113_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y113_SLICE_X6Y113_CO5),
.O6(CLBLM_R_X5Y113_SLICE_X6Y113_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X5Y113_SLICE_X6Y113_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y113_SLICE_X6Y113_BO5),
.O6(CLBLM_R_X5Y113_SLICE_X6Y113_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X5Y113_SLICE_X6Y113_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y113_SLICE_X6Y113_AO5),
.O6(CLBLM_R_X5Y113_SLICE_X6Y113_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X5Y113_SLICE_X7Y113_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y113_SLICE_X7Y113_DO5),
.O6(CLBLM_R_X5Y113_SLICE_X7Y113_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h570577077f77ff7f)
  ) CLBLM_R_X5Y113_SLICE_X7Y113_CLUT (
.I0(RIOB33_X105Y109_IOB_X1Y109_I),
.I1(LIOB33_X0Y115_IOB_X0Y115_I),
.I2(CLBLM_R_X5Y110_SLICE_X6Y110_BO5),
.I3(CLBLM_R_X5Y111_SLICE_X7Y111_DO6),
.I4(LIOB33_X0Y113_IOB_X0Y113_I),
.I5(CLBLM_R_X5Y112_SLICE_X7Y112_CO6),
.O5(CLBLM_R_X5Y113_SLICE_X7Y113_CO5),
.O6(CLBLM_R_X5Y113_SLICE_X7Y113_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h936cff00c93655aa)
  ) CLBLM_R_X5Y113_SLICE_X7Y113_BLUT (
.I0(CLBLM_R_X5Y110_SLICE_X6Y110_BO5),
.I1(LIOB33_X0Y115_IOB_X0Y115_I),
.I2(LIOB33_X0Y113_IOB_X0Y113_I),
.I3(CLBLM_R_X5Y112_SLICE_X7Y112_CO6),
.I4(RIOB33_X105Y109_IOB_X1Y109_I),
.I5(CLBLM_R_X5Y111_SLICE_X7Y111_DO6),
.O5(CLBLM_R_X5Y113_SLICE_X7Y113_BO5),
.O6(CLBLM_R_X5Y113_SLICE_X7Y113_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h5fa0a05f5fff005f)
  ) CLBLM_R_X5Y113_SLICE_X7Y113_ALUT (
.I0(RIOB33_X105Y103_IOB_X1Y104_I),
.I1(1'b1),
.I2(LIOB33_X0Y113_IOB_X0Y113_I),
.I3(CLBLM_R_X7Y113_SLICE_X9Y113_AO6),
.I4(CLBLM_L_X8Y113_SLICE_X10Y113_CO6),
.I5(1'b1),
.O5(CLBLM_R_X5Y113_SLICE_X7Y113_AO5),
.O6(CLBLM_R_X5Y113_SLICE_X7Y113_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h33d9ff15cc2600ea)
  ) CLBLM_R_X7Y103_SLICE_X8Y103_DLUT (
.I0(CLBLM_R_X7Y103_SLICE_X8Y103_AO6),
.I1(LIOB33_X0Y101_IOB_X0Y101_I),
.I2(LIOB33_X0Y117_IOB_X0Y117_I),
.I3(CLBLM_R_X7Y103_SLICE_X8Y103_CO6),
.I4(RIOB33_X105Y101_IOB_X1Y101_I),
.I5(CLBLM_R_X7Y103_SLICE_X8Y103_BO6),
.O5(CLBLM_R_X7Y103_SLICE_X8Y103_DO5),
.O6(CLBLM_R_X7Y103_SLICE_X8Y103_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h226600a002c600a0)
  ) CLBLM_R_X7Y103_SLICE_X8Y103_CLUT (
.I0(RIOB33_X105Y113_IOB_X1Y113_I),
.I1(LIOB33_SING_X0Y100_IOB_X0Y100_I),
.I2(RIOB33_X105Y101_IOB_X1Y102_I),
.I3(LIOB33_X0Y117_IOB_X0Y117_I),
.I4(RIOB33_X105Y101_IOB_X1Y101_I),
.I5(RIOB33_X105Y111_IOB_X1Y112_I),
.O5(CLBLM_R_X7Y103_SLICE_X8Y103_CO5),
.O6(CLBLM_R_X7Y103_SLICE_X8Y103_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h165626a6d010e0e0)
  ) CLBLM_R_X7Y103_SLICE_X8Y103_BLUT (
.I0(RIOB33_X105Y101_IOB_X1Y101_I),
.I1(RIOB33_X105Y101_IOB_X1Y102_I),
.I2(RIOB33_X105Y113_IOB_X1Y113_I),
.I3(RIOB33_X105Y111_IOB_X1Y112_I),
.I4(RIOB33_X105Y103_IOB_X1Y103_I),
.I5(LIOB33_SING_X0Y100_IOB_X0Y100_I),
.O5(CLBLM_R_X7Y103_SLICE_X8Y103_BO5),
.O6(CLBLM_R_X7Y103_SLICE_X8Y103_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h154a35cab0e03060)
  ) CLBLM_R_X7Y103_SLICE_X8Y103_ALUT (
.I0(RIOB33_X105Y101_IOB_X1Y101_I),
.I1(RIOB33_X105Y101_IOB_X1Y102_I),
.I2(RIOB33_X105Y113_IOB_X1Y113_I),
.I3(LIOB33_X0Y117_IOB_X0Y117_I),
.I4(RIOB33_X105Y111_IOB_X1Y112_I),
.I5(LIOB33_SING_X0Y100_IOB_X0Y100_I),
.O5(CLBLM_R_X7Y103_SLICE_X8Y103_AO5),
.O6(CLBLM_R_X7Y103_SLICE_X8Y103_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X7Y103_SLICE_X9Y103_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y103_SLICE_X9Y103_DO5),
.O6(CLBLM_R_X7Y103_SLICE_X9Y103_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X7Y103_SLICE_X9Y103_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y103_SLICE_X9Y103_CO5),
.O6(CLBLM_R_X7Y103_SLICE_X9Y103_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X7Y103_SLICE_X9Y103_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y103_SLICE_X9Y103_BO5),
.O6(CLBLM_R_X7Y103_SLICE_X9Y103_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X7Y103_SLICE_X9Y103_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y103_SLICE_X9Y103_AO5),
.O6(CLBLM_R_X7Y103_SLICE_X9Y103_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hffcece00ce00ffce)
  ) CLBLM_R_X7Y104_SLICE_X8Y104_DLUT (
.I0(CLBLM_R_X7Y104_SLICE_X8Y104_AO6),
.I1(CLBLM_R_X7Y103_SLICE_X8Y103_CO6),
.I2(CLBLM_R_X7Y103_SLICE_X8Y103_AO6),
.I3(CLBLM_R_X7Y104_SLICE_X8Y104_AO5),
.I4(CLBLM_L_X8Y104_SLICE_X10Y104_AO6),
.I5(CLBLM_R_X7Y103_SLICE_X8Y103_BO6),
.O5(CLBLM_R_X7Y104_SLICE_X8Y104_DO5),
.O6(CLBLM_R_X7Y104_SLICE_X8Y104_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h31cece31ce3131ce)
  ) CLBLM_R_X7Y104_SLICE_X8Y104_CLUT (
.I0(CLBLM_R_X7Y104_SLICE_X8Y104_AO6),
.I1(CLBLM_R_X7Y103_SLICE_X8Y103_CO6),
.I2(CLBLM_R_X7Y103_SLICE_X8Y103_AO6),
.I3(CLBLM_R_X7Y104_SLICE_X8Y104_AO5),
.I4(CLBLM_L_X8Y104_SLICE_X10Y104_AO6),
.I5(CLBLM_R_X7Y103_SLICE_X8Y103_BO6),
.O5(CLBLM_R_X7Y104_SLICE_X8Y104_CO5),
.O6(CLBLM_R_X7Y104_SLICE_X8Y104_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf00f0f0fcccfcfcf)
  ) CLBLM_R_X7Y104_SLICE_X8Y104_BLUT (
.I0(1'b1),
.I1(CLBLM_R_X7Y103_SLICE_X8Y103_CO6),
.I2(CLBLM_R_X7Y103_SLICE_X8Y103_AO6),
.I3(LIOB33_X0Y117_IOB_X0Y117_I),
.I4(LIOB33_X0Y101_IOB_X0Y101_I),
.I5(1'b1),
.O5(CLBLM_R_X7Y104_SLICE_X8Y104_BO5),
.O6(CLBLM_R_X7Y104_SLICE_X8Y104_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h3f3f3f3f33ff33ff)
  ) CLBLM_R_X7Y104_SLICE_X8Y104_ALUT (
.I0(1'b1),
.I1(LIOB33_X0Y117_IOB_X0Y117_I),
.I2(LIOB33_X0Y101_IOB_X0Y101_I),
.I3(LIOB33_X0Y101_IOB_X0Y102_I),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y104_SLICE_X8Y104_AO5),
.O6(CLBLM_R_X7Y104_SLICE_X8Y104_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h9c3963c6c3ccc3cc)
  ) CLBLM_R_X7Y104_SLICE_X9Y104_DLUT (
.I0(LIOB33_X0Y117_IOB_X0Y117_I),
.I1(CLBLM_L_X8Y104_SLICE_X10Y104_DO6),
.I2(CLBLM_R_X7Y104_SLICE_X8Y104_BO5),
.I3(CLBLM_L_X8Y103_SLICE_X10Y103_AO6),
.I4(RIOB33_X105Y101_IOB_X1Y101_I),
.I5(LIOB33_X0Y101_IOB_X0Y102_I),
.O5(CLBLM_R_X7Y104_SLICE_X9Y104_DO5),
.O6(CLBLM_R_X7Y104_SLICE_X9Y104_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h7887877887788778)
  ) CLBLM_R_X7Y104_SLICE_X9Y104_CLUT (
.I0(LIOB33_X0Y117_IOB_X0Y117_I),
.I1(LIOB33_X0Y103_IOB_X0Y104_I),
.I2(CLBLM_R_X7Y104_SLICE_X8Y104_DO6),
.I3(CLBLM_L_X8Y104_SLICE_X10Y104_DO6),
.I4(RIOB33_X105Y101_IOB_X1Y101_I),
.I5(LIOB33_X0Y101_IOB_X0Y102_I),
.O5(CLBLM_R_X7Y104_SLICE_X9Y104_CO5),
.O6(CLBLM_R_X7Y104_SLICE_X9Y104_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h6996969669696996)
  ) CLBLM_R_X7Y104_SLICE_X9Y104_BLUT (
.I0(CLBLM_L_X8Y104_SLICE_X10Y104_CO6),
.I1(CLBLM_L_X10Y102_SLICE_X12Y102_BO6),
.I2(CLBLM_L_X8Y105_SLICE_X11Y105_AO6),
.I3(CLBLM_R_X7Y104_SLICE_X8Y104_DO6),
.I4(CLBLM_R_X7Y104_SLICE_X9Y104_AO6),
.I5(CLBLM_L_X8Y104_SLICE_X10Y104_BO6),
.O5(CLBLM_R_X7Y104_SLICE_X9Y104_BO5),
.O6(CLBLM_R_X7Y104_SLICE_X9Y104_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h33ff33ff55ff55ff)
  ) CLBLM_R_X7Y104_SLICE_X9Y104_ALUT (
.I0(LIOB33_X0Y105_IOB_X0Y105_I),
.I1(LIOB33_X0Y103_IOB_X0Y104_I),
.I2(1'b1),
.I3(LIOB33_X0Y117_IOB_X0Y117_I),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y104_SLICE_X9Y104_AO5),
.O6(CLBLM_R_X7Y104_SLICE_X9Y104_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h7fbfff3f152a3f00)
  ) CLBLM_R_X7Y105_SLICE_X8Y105_DLUT (
.I0(LIOB33_X0Y115_IOB_X0Y116_I),
.I1(LIOB33_X0Y113_IOB_X0Y114_I),
.I2(LIOB33_X0Y107_IOB_X0Y108_I),
.I3(CLBLM_R_X7Y105_SLICE_X8Y105_AO5),
.I4(LIOB33_X0Y107_IOB_X0Y107_I),
.I5(CLBLM_R_X7Y105_SLICE_X8Y105_BO6),
.O5(CLBLM_R_X7Y105_SLICE_X8Y105_DO5),
.O6(CLBLM_R_X7Y105_SLICE_X8Y105_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h6a95c03f956a3fc0)
  ) CLBLM_R_X7Y105_SLICE_X8Y105_CLUT (
.I0(LIOB33_X0Y115_IOB_X0Y116_I),
.I1(LIOB33_X0Y113_IOB_X0Y114_I),
.I2(LIOB33_X0Y107_IOB_X0Y108_I),
.I3(CLBLM_R_X7Y105_SLICE_X8Y105_AO5),
.I4(LIOB33_X0Y107_IOB_X0Y107_I),
.I5(CLBLM_R_X7Y105_SLICE_X8Y105_BO6),
.O5(CLBLM_R_X7Y105_SLICE_X8Y105_CO5),
.O6(CLBLM_R_X7Y105_SLICE_X8Y105_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h7b12bb22ff5affaa)
  ) CLBLM_R_X7Y105_SLICE_X8Y105_BLUT (
.I0(CLBLM_R_X7Y105_SLICE_X9Y105_CO6),
.I1(LIOB33_X0Y107_IOB_X0Y107_I),
.I2(LIOB33_X0Y105_IOB_X0Y106_I),
.I3(CLBLM_R_X5Y105_SLICE_X7Y105_CO6),
.I4(LIOB33_X0Y115_IOB_X0Y116_I),
.I5(LIOB33_X0Y113_IOB_X0Y114_I),
.O5(CLBLM_R_X7Y105_SLICE_X8Y105_BO5),
.O6(CLBLM_R_X7Y105_SLICE_X8Y105_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h5555ffff96693cc3)
  ) CLBLM_R_X7Y105_SLICE_X8Y105_ALUT (
.I0(LIOB33_X0Y117_IOB_X0Y117_I),
.I1(CLBLM_R_X7Y105_SLICE_X9Y105_BO6),
.I2(CLBLM_L_X8Y106_SLICE_X11Y106_AO6),
.I3(CLBLM_L_X8Y104_SLICE_X11Y104_CO6),
.I4(LIOB33_X0Y105_IOB_X0Y106_I),
.I5(1'b1),
.O5(CLBLM_R_X7Y105_SLICE_X8Y105_AO5),
.O6(CLBLM_R_X7Y105_SLICE_X8Y105_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h6c93936ca05f5fa0)
  ) CLBLM_R_X7Y105_SLICE_X9Y105_DLUT (
.I0(LIOB33_X0Y115_IOB_X0Y116_I),
.I1(LIOB33_X0Y103_IOB_X0Y104_I),
.I2(LIOB33_X0Y105_IOB_X0Y105_I),
.I3(CLBLM_R_X5Y104_SLICE_X7Y104_BO6),
.I4(CLBLM_R_X7Y104_SLICE_X9Y104_DO6),
.I5(LIOB33_X0Y117_IOB_X0Y117_I),
.O5(CLBLM_R_X7Y105_SLICE_X9Y105_DO5),
.O6(CLBLM_R_X7Y105_SLICE_X9Y105_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h9f60c03f3fc09f60)
  ) CLBLM_R_X7Y105_SLICE_X9Y105_CLUT (
.I0(LIOB33_X0Y115_IOB_X0Y116_I),
.I1(LIOB33_X0Y117_IOB_X0Y117_I),
.I2(LIOB33_X0Y105_IOB_X0Y105_I),
.I3(CLBLM_R_X7Y104_SLICE_X9Y104_BO6),
.I4(CLBLM_R_X5Y104_SLICE_X7Y104_BO6),
.I5(CLBLM_R_X7Y104_SLICE_X9Y104_CO6),
.O5(CLBLM_R_X7Y105_SLICE_X9Y105_CO5),
.O6(CLBLM_R_X7Y105_SLICE_X9Y105_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'he8c0fce88e0ccf8e)
  ) CLBLM_R_X7Y105_SLICE_X9Y105_BLUT (
.I0(CLBLM_R_X5Y104_SLICE_X7Y104_BO6),
.I1(CLBLM_L_X8Y105_SLICE_X10Y105_AO6),
.I2(CLBLM_R_X7Y104_SLICE_X9Y104_BO6),
.I3(CLBLM_R_X5Y106_SLICE_X7Y106_AO6),
.I4(CLBLM_R_X7Y104_SLICE_X9Y104_CO6),
.I5(CLBLM_R_X7Y104_SLICE_X9Y104_AO5),
.O5(CLBLM_R_X7Y105_SLICE_X9Y105_BO5),
.O6(CLBLM_R_X7Y105_SLICE_X9Y105_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h78871ee18778e11e)
  ) CLBLM_R_X7Y105_SLICE_X9Y105_ALUT (
.I0(CLBLM_R_X5Y104_SLICE_X7Y104_BO6),
.I1(CLBLM_R_X5Y106_SLICE_X7Y106_AO6),
.I2(CLBLM_R_X7Y104_SLICE_X9Y104_BO6),
.I3(CLBLM_L_X8Y105_SLICE_X10Y105_AO6),
.I4(CLBLM_R_X7Y104_SLICE_X9Y104_CO6),
.I5(CLBLM_R_X7Y104_SLICE_X9Y104_AO5),
.O5(CLBLM_R_X7Y105_SLICE_X9Y105_AO5),
.O6(CLBLM_R_X7Y105_SLICE_X9Y105_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000002000)
  ) CLBLM_R_X7Y106_SLICE_X8Y106_DLUT (
.I0(CLBLM_R_X3Y106_SLICE_X2Y106_AO6),
.I1(CLBLM_L_X8Y104_SLICE_X11Y104_CO6),
.I2(RIOB33_X105Y107_IOB_X1Y108_I),
.I3(LIOB33_X0Y103_IOB_X0Y104_I),
.I4(CLBLM_L_X8Y106_SLICE_X11Y106_AO6),
.I5(CLBLM_L_X12Y107_SLICE_X17Y107_AO5),
.O5(CLBLM_R_X7Y106_SLICE_X8Y106_DO5),
.O6(CLBLM_R_X7Y106_SLICE_X8Y106_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h6999966696666999)
  ) CLBLM_R_X7Y106_SLICE_X8Y106_CLUT (
.I0(CLBLM_R_X7Y105_SLICE_X9Y105_BO6),
.I1(CLBLM_L_X8Y104_SLICE_X11Y104_CO6),
.I2(LIOB33_X0Y105_IOB_X0Y106_I),
.I3(LIOB33_X0Y117_IOB_X0Y117_I),
.I4(CLBLM_L_X8Y106_SLICE_X10Y106_AO6),
.I5(CLBLM_L_X8Y106_SLICE_X11Y106_AO6),
.O5(CLBLM_R_X7Y106_SLICE_X8Y106_CO5),
.O6(CLBLM_R_X7Y106_SLICE_X8Y106_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h6696996996996966)
  ) CLBLM_R_X7Y106_SLICE_X8Y106_BLUT (
.I0(CLBLM_L_X8Y106_SLICE_X10Y106_AO6),
.I1(CLBLM_L_X8Y104_SLICE_X11Y104_AO6),
.I2(CLBLM_R_X7Y105_SLICE_X9Y105_AO6),
.I3(CLBLM_R_X5Y106_SLICE_X7Y106_BO6),
.I4(CLBLM_R_X7Y105_SLICE_X9Y105_BO6),
.I5(CLBLM_R_X5Y105_SLICE_X7Y105_CO6),
.O5(CLBLM_R_X7Y106_SLICE_X8Y106_BO5),
.O6(CLBLM_R_X7Y106_SLICE_X8Y106_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h5555ffff5f5f5f5f)
  ) CLBLM_R_X7Y106_SLICE_X8Y106_ALUT (
.I0(LIOB33_X0Y107_IOB_X0Y108_I),
.I1(1'b1),
.I2(LIOB33_X0Y113_IOB_X0Y114_I),
.I3(1'b1),
.I4(LIOB33_X0Y115_IOB_X0Y116_I),
.I5(1'b1),
.O5(CLBLM_R_X7Y106_SLICE_X8Y106_AO5),
.O6(CLBLM_R_X7Y106_SLICE_X8Y106_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hfbb0bf0bf2202f02)
  ) CLBLM_R_X7Y106_SLICE_X9Y106_DLUT (
.I0(CLBLM_R_X7Y105_SLICE_X8Y105_BO6),
.I1(CLBLM_R_X7Y106_SLICE_X8Y106_CO6),
.I2(CLBLM_L_X8Y106_SLICE_X10Y106_DO6),
.I3(CLBLM_R_X5Y106_SLICE_X6Y106_AO5),
.I4(CLBLM_R_X7Y106_SLICE_X8Y106_AO6),
.I5(CLBLM_R_X7Y106_SLICE_X8Y106_AO5),
.O5(CLBLM_R_X7Y106_SLICE_X9Y106_DO5),
.O6(CLBLM_R_X7Y106_SLICE_X9Y106_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h8fe3701c7f1380ec)
  ) CLBLM_R_X7Y106_SLICE_X9Y106_CLUT (
.I0(LIOB33_X0Y117_IOB_X0Y117_I),
.I1(CLBLM_L_X8Y106_SLICE_X11Y106_AO6),
.I2(LIOB33_X0Y105_IOB_X0Y106_I),
.I3(CLBLM_L_X8Y104_SLICE_X11Y104_CO6),
.I4(CLBLM_L_X8Y105_SLICE_X11Y105_DO6),
.I5(RIOB33_X105Y101_IOB_X1Y101_I),
.O5(CLBLM_R_X7Y106_SLICE_X9Y106_CO5),
.O6(CLBLM_R_X7Y106_SLICE_X9Y106_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h65a69a599a5965a6)
  ) CLBLM_R_X7Y106_SLICE_X9Y106_BLUT (
.I0(CLBLM_R_X7Y106_SLICE_X8Y106_AO6),
.I1(CLBLM_R_X7Y105_SLICE_X8Y105_BO6),
.I2(CLBLM_R_X7Y106_SLICE_X8Y106_CO6),
.I3(CLBLM_R_X7Y106_SLICE_X8Y106_AO5),
.I4(CLBLM_L_X8Y106_SLICE_X10Y106_DO6),
.I5(CLBLM_R_X5Y106_SLICE_X6Y106_AO5),
.O5(CLBLM_R_X7Y106_SLICE_X9Y106_BO5),
.O6(CLBLM_R_X7Y106_SLICE_X9Y106_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h65a69a599a5965a6)
  ) CLBLM_R_X7Y106_SLICE_X9Y106_ALUT (
.I0(CLBLM_R_X7Y106_SLICE_X8Y106_AO6),
.I1(CLBLM_R_X7Y105_SLICE_X8Y105_BO6),
.I2(CLBLM_R_X7Y106_SLICE_X8Y106_CO6),
.I3(CLBLM_R_X7Y106_SLICE_X8Y106_AO5),
.I4(CLBLM_L_X8Y105_SLICE_X10Y105_BO6),
.I5(CLBLM_L_X8Y106_SLICE_X10Y106_BO6),
.O5(CLBLM_R_X7Y106_SLICE_X9Y106_AO5),
.O6(CLBLM_R_X7Y106_SLICE_X9Y106_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h5a96a56996a5695a)
  ) CLBLM_R_X7Y107_SLICE_X8Y107_DLUT (
.I0(CLBLM_L_X8Y107_SLICE_X10Y107_BO6),
.I1(CLBLM_R_X7Y107_SLICE_X9Y107_CO6),
.I2(CLBLM_R_X5Y110_SLICE_X7Y110_BO6),
.I3(CLBLM_R_X5Y107_SLICE_X7Y107_CO6),
.I4(CLBLM_R_X7Y108_SLICE_X8Y108_AO6),
.I5(CLBLM_R_X5Y108_SLICE_X7Y108_AO5),
.O5(CLBLM_R_X7Y107_SLICE_X8Y107_DO5),
.O6(CLBLM_R_X7Y107_SLICE_X8Y107_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h7800ff78ff78ff78)
  ) CLBLM_R_X7Y107_SLICE_X8Y107_CLUT (
.I0(LIOB33_X0Y113_IOB_X0Y114_I),
.I1(LIOB33_X0Y109_IOB_X0Y110_I),
.I2(CLBLM_R_X7Y107_SLICE_X9Y107_BO6),
.I3(CLBLM_R_X5Y107_SLICE_X7Y107_CO6),
.I4(LIOB33_X0Y103_IOB_X0Y103_I),
.I5(LIOB33_X0Y111_IOB_X0Y111_I),
.O5(CLBLM_R_X7Y107_SLICE_X8Y107_CO5),
.O6(CLBLM_R_X7Y107_SLICE_X8Y107_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h659a9a65a65959a6)
  ) CLBLM_R_X7Y107_SLICE_X8Y107_BLUT (
.I0(CLBLM_R_X7Y108_SLICE_X9Y108_BO6),
.I1(CLBLM_R_X5Y108_SLICE_X7Y108_AO5),
.I2(CLBLM_R_X7Y107_SLICE_X9Y107_CO6),
.I3(CLBLM_R_X7Y108_SLICE_X8Y108_AO6),
.I4(CLBLM_R_X7Y107_SLICE_X9Y107_DO6),
.I5(CLBLM_R_X5Y107_SLICE_X7Y107_CO6),
.O5(CLBLM_R_X7Y107_SLICE_X8Y107_BO5),
.O6(CLBLM_R_X7Y107_SLICE_X8Y107_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h69c39933963c66cc)
  ) CLBLM_R_X7Y107_SLICE_X8Y107_ALUT (
.I0(LIOB33_X0Y103_IOB_X0Y103_I),
.I1(CLBLM_R_X7Y107_SLICE_X9Y107_BO6),
.I2(LIOB33_X0Y113_IOB_X0Y114_I),
.I3(LIOB33_X0Y111_IOB_X0Y111_I),
.I4(LIOB33_X0Y109_IOB_X0Y110_I),
.I5(CLBLM_R_X5Y107_SLICE_X7Y107_CO6),
.O5(CLBLM_R_X7Y107_SLICE_X8Y107_AO5),
.O6(CLBLM_R_X7Y107_SLICE_X8Y107_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0701ff557f1fffff)
  ) CLBLM_R_X7Y107_SLICE_X9Y107_DLUT (
.I0(CLBLM_R_X7Y107_SLICE_X9Y107_AO6),
.I1(LIOB33_X0Y109_IOB_X0Y109_I),
.I2(LIOB33_X0Y109_IOB_X0Y110_I),
.I3(CLBLM_R_X7Y105_SLICE_X8Y105_DO6),
.I4(LIOB33_X0Y113_IOB_X0Y114_I),
.I5(CLBLM_L_X8Y106_SLICE_X11Y106_BO6),
.O5(CLBLM_R_X7Y107_SLICE_X9Y107_DO5),
.O6(CLBLM_R_X7Y107_SLICE_X9Y107_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h9c39f5f563c60a0a)
  ) CLBLM_R_X7Y107_SLICE_X9Y107_CLUT (
.I0(CLBLM_R_X7Y107_SLICE_X9Y107_AO6),
.I1(LIOB33_X0Y109_IOB_X0Y110_I),
.I2(CLBLM_R_X7Y105_SLICE_X8Y105_DO6),
.I3(LIOB33_X0Y109_IOB_X0Y109_I),
.I4(LIOB33_X0Y113_IOB_X0Y114_I),
.I5(CLBLM_L_X8Y106_SLICE_X11Y106_BO6),
.O5(CLBLM_R_X7Y107_SLICE_X9Y107_CO5),
.O6(CLBLM_R_X7Y107_SLICE_X9Y107_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h39c69c6355aa00ff)
  ) CLBLM_R_X7Y107_SLICE_X9Y107_BLUT (
.I0(CLBLM_R_X7Y105_SLICE_X8Y105_DO6),
.I1(LIOB33_X0Y115_IOB_X0Y116_I),
.I2(LIOB33_X0Y113_IOB_X0Y114_I),
.I3(CLBLM_L_X8Y107_SLICE_X10Y107_AO6),
.I4(CLBLM_R_X7Y107_SLICE_X9Y107_AO6),
.I5(LIOB33_X0Y109_IOB_X0Y109_I),
.O5(CLBLM_R_X7Y107_SLICE_X9Y107_BO5),
.O6(CLBLM_R_X7Y107_SLICE_X9Y107_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h6a95c03f956a3fc0)
  ) CLBLM_R_X7Y107_SLICE_X9Y107_ALUT (
.I0(LIOB33_X0Y107_IOB_X0Y108_I),
.I1(LIOB33_X0Y107_IOB_X0Y107_I),
.I2(LIOB33_X0Y117_IOB_X0Y117_I),
.I3(CLBLM_L_X8Y105_SLICE_X10Y105_BO6),
.I4(LIOB33_X0Y115_IOB_X0Y116_I),
.I5(CLBLM_R_X7Y106_SLICE_X9Y106_CO6),
.O5(CLBLM_R_X7Y107_SLICE_X9Y107_AO5),
.O6(CLBLM_R_X7Y107_SLICE_X9Y107_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X7Y108_SLICE_X8Y108_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y108_SLICE_X8Y108_DO5),
.O6(CLBLM_R_X7Y108_SLICE_X8Y108_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h639c9c63c63939c6)
  ) CLBLM_R_X7Y108_SLICE_X8Y108_CLUT (
.I0(CLBLM_R_X7Y108_SLICE_X8Y108_AO6),
.I1(CLBLM_R_X7Y108_SLICE_X9Y108_CO6),
.I2(CLBLM_R_X7Y108_SLICE_X9Y108_BO6),
.I3(CLBLM_R_X7Y108_SLICE_X8Y108_AO5),
.I4(CLBLM_L_X8Y108_SLICE_X11Y108_BO6),
.I5(CLBLM_R_X7Y107_SLICE_X9Y107_DO6),
.O5(CLBLM_R_X7Y108_SLICE_X8Y108_CO5),
.O6(CLBLM_R_X7Y108_SLICE_X8Y108_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h4bb4d22db44b2dd2)
  ) CLBLM_R_X7Y108_SLICE_X8Y108_BLUT (
.I0(CLBLM_R_X7Y107_SLICE_X9Y107_DO6),
.I1(CLBLM_R_X7Y108_SLICE_X9Y108_BO6),
.I2(CLBLM_R_X7Y109_SLICE_X8Y109_AO6),
.I3(CLBLM_L_X8Y108_SLICE_X10Y108_CO6),
.I4(CLBLM_R_X7Y108_SLICE_X8Y108_AO6),
.I5(CLBLM_R_X7Y108_SLICE_X8Y108_AO5),
.O5(CLBLM_R_X7Y108_SLICE_X8Y108_BO5),
.O6(CLBLM_R_X7Y108_SLICE_X8Y108_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h00ffffff0fff0fff)
  ) CLBLM_R_X7Y108_SLICE_X8Y108_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(LIOB33_X0Y115_IOB_X0Y116_I),
.I3(LIOB33_X0Y111_IOB_X0Y111_I),
.I4(LIOB33_X0Y113_IOB_X0Y114_I),
.I5(1'b1),
.O5(CLBLM_R_X7Y108_SLICE_X8Y108_AO5),
.O6(CLBLM_R_X7Y108_SLICE_X8Y108_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h93ccc9666ccc3666)
  ) CLBLM_R_X7Y108_SLICE_X9Y108_DLUT (
.I0(CLBLM_L_X8Y108_SLICE_X10Y108_BO6),
.I1(CLBLM_L_X8Y107_SLICE_X10Y107_CO6),
.I2(LIOB33_X0Y115_IOB_X0Y116_I),
.I3(LIOB33_X0Y109_IOB_X0Y109_I),
.I4(CLBLM_R_X7Y108_SLICE_X9Y108_AO6),
.I5(LIOB33_X0Y117_IOB_X0Y117_I),
.O5(CLBLM_R_X7Y108_SLICE_X9Y108_DO5),
.O6(CLBLM_R_X7Y108_SLICE_X9Y108_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h077f011fffff5f5f)
  ) CLBLM_R_X7Y108_SLICE_X9Y108_CLUT (
.I0(CLBLM_L_X8Y108_SLICE_X10Y108_BO6),
.I1(LIOB33_X0Y109_IOB_X0Y109_I),
.I2(CLBLM_L_X8Y107_SLICE_X11Y107_CO6),
.I3(LIOB33_X0Y109_IOB_X0Y110_I),
.I4(CLBLM_R_X7Y108_SLICE_X9Y108_AO6),
.I5(LIOB33_X0Y115_IOB_X0Y116_I),
.O5(CLBLM_R_X7Y108_SLICE_X9Y108_CO5),
.O6(CLBLM_R_X7Y108_SLICE_X9Y108_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hc39969cc69993ccc)
  ) CLBLM_R_X7Y108_SLICE_X9Y108_BLUT (
.I0(CLBLM_R_X7Y108_SLICE_X9Y108_AO6),
.I1(CLBLM_L_X8Y107_SLICE_X11Y107_CO6),
.I2(LIOB33_X0Y109_IOB_X0Y110_I),
.I3(LIOB33_X0Y115_IOB_X0Y116_I),
.I4(CLBLM_L_X8Y108_SLICE_X10Y108_BO6),
.I5(LIOB33_X0Y109_IOB_X0Y109_I),
.O5(CLBLM_R_X7Y108_SLICE_X9Y108_BO5),
.O6(CLBLM_R_X7Y108_SLICE_X9Y108_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h71d4f3fcf550fff0)
  ) CLBLM_R_X7Y108_SLICE_X9Y108_ALUT (
.I0(LIOB33_X0Y107_IOB_X0Y108_I),
.I1(LIOB33_X0Y117_IOB_X0Y117_I),
.I2(CLBLM_L_X8Y105_SLICE_X10Y105_BO6),
.I3(CLBLM_R_X7Y106_SLICE_X9Y106_CO6),
.I4(LIOB33_X0Y115_IOB_X0Y116_I),
.I5(LIOB33_X0Y107_IOB_X0Y107_I),
.O5(CLBLM_R_X7Y108_SLICE_X9Y108_AO5),
.O6(CLBLM_R_X7Y108_SLICE_X9Y108_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h6a95956a56a9a956)
  ) CLBLM_R_X7Y109_SLICE_X8Y109_DLUT (
.I0(CLBLM_L_X8Y108_SLICE_X10Y108_DO6),
.I1(CLBLM_R_X7Y108_SLICE_X8Y108_AO5),
.I2(CLBLM_R_X7Y108_SLICE_X9Y108_CO6),
.I3(CLBLM_R_X7Y109_SLICE_X8Y109_AO5),
.I4(CLBLM_L_X8Y110_SLICE_X11Y110_AO6),
.I5(CLBLM_L_X8Y108_SLICE_X11Y108_BO6),
.O5(CLBLM_R_X7Y109_SLICE_X8Y109_DO5),
.O6(CLBLM_R_X7Y109_SLICE_X8Y109_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h7887877887788778)
  ) CLBLM_R_X7Y109_SLICE_X8Y109_CLUT (
.I0(LIOB33_X0Y111_IOB_X0Y111_I),
.I1(LIOB33_X0Y115_IOB_X0Y116_I),
.I2(CLBLM_R_X7Y108_SLICE_X9Y108_CO6),
.I3(CLBLM_L_X8Y108_SLICE_X11Y108_CO6),
.I4(LIOB33_X0Y109_IOB_X0Y110_I),
.I5(LIOB33_X0Y117_IOB_X0Y117_I),
.O5(CLBLM_R_X7Y109_SLICE_X8Y109_CO5),
.O6(CLBLM_R_X7Y109_SLICE_X8Y109_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h5a96a56996a5695a)
  ) CLBLM_R_X7Y109_SLICE_X8Y109_BLUT (
.I0(CLBLM_L_X8Y110_SLICE_X11Y110_BO6),
.I1(CLBLM_L_X8Y108_SLICE_X11Y108_BO6),
.I2(CLBLM_L_X8Y110_SLICE_X11Y110_AO6),
.I3(CLBLM_R_X7Y108_SLICE_X9Y108_CO6),
.I4(CLBLM_L_X8Y108_SLICE_X11Y108_AO6),
.I5(CLBLM_R_X7Y108_SLICE_X8Y108_AO5),
.O5(CLBLM_R_X7Y109_SLICE_X8Y109_BO5),
.O6(CLBLM_R_X7Y109_SLICE_X8Y109_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h00ffffff0fff0fff)
  ) CLBLM_R_X7Y109_SLICE_X8Y109_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(LIOB33_X0Y115_IOB_X0Y116_I),
.I3(LIOB33_X0Y111_IOB_X0Y112_I),
.I4(LIOB33_X0Y113_IOB_X0Y114_I),
.I5(1'b1),
.O5(CLBLM_R_X7Y109_SLICE_X8Y109_AO5),
.O6(CLBLM_R_X7Y109_SLICE_X8Y109_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h7ff70770ff777700)
  ) CLBLM_R_X7Y109_SLICE_X9Y109_DLUT (
.I0(LIOB33_X0Y109_IOB_X0Y110_I),
.I1(RIOB33_X105Y109_IOB_X1Y109_I),
.I2(LIOB33_X0Y109_IOB_X0Y109_I),
.I3(CLBLM_R_X7Y109_SLICE_X9Y109_CO6),
.I4(CLBLM_L_X8Y109_SLICE_X10Y109_AO6),
.I5(RIOB33_X105Y109_IOB_X1Y110_I),
.O5(CLBLM_R_X7Y109_SLICE_X9Y109_DO5),
.O6(CLBLM_R_X7Y109_SLICE_X9Y109_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hdf9977f777d77777)
  ) CLBLM_R_X7Y109_SLICE_X9Y109_CLUT (
.I0(RIOB33_X105Y111_IOB_X1Y111_I),
.I1(LIOB33_X0Y107_IOB_X0Y108_I),
.I2(LIOB33_X0Y105_IOB_X0Y106_I),
.I3(CLBLM_L_X10Y109_SLICE_X12Y109_DO6),
.I4(LIOB33_X0Y107_IOB_X0Y107_I),
.I5(RIOB33_X105Y109_IOB_X1Y110_I),
.O5(CLBLM_R_X7Y109_SLICE_X9Y109_CO5),
.O6(CLBLM_R_X7Y109_SLICE_X9Y109_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h69a59955965a66aa)
  ) CLBLM_R_X7Y109_SLICE_X9Y109_BLUT (
.I0(CLBLM_L_X8Y109_SLICE_X10Y109_AO6),
.I1(RIOB33_X105Y109_IOB_X1Y110_I),
.I2(LIOB33_X0Y109_IOB_X0Y110_I),
.I3(LIOB33_X0Y109_IOB_X0Y109_I),
.I4(RIOB33_X105Y109_IOB_X1Y109_I),
.I5(CLBLM_R_X7Y109_SLICE_X9Y109_CO6),
.O5(CLBLM_R_X7Y109_SLICE_X9Y109_BO5),
.O6(CLBLM_R_X7Y109_SLICE_X9Y109_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h99993333a05fa05f)
  ) CLBLM_R_X7Y109_SLICE_X9Y109_ALUT (
.I0(LIOB33_X0Y107_IOB_X0Y107_I),
.I1(CLBLM_L_X10Y109_SLICE_X12Y109_CO6),
.I2(RIOB33_SING_X105Y100_IOB_X1Y100_I),
.I3(CLBLM_R_X3Y107_SLICE_X2Y107_BO6),
.I4(RIOB33_X105Y109_IOB_X1Y110_I),
.I5(1'b1),
.O5(CLBLM_R_X7Y109_SLICE_X9Y109_AO5),
.O6(CLBLM_R_X7Y109_SLICE_X9Y109_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X7Y110_SLICE_X8Y110_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y110_SLICE_X8Y110_DO5),
.O6(CLBLM_R_X7Y110_SLICE_X8Y110_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000200000000)
  ) CLBLM_R_X7Y110_SLICE_X8Y110_CLUT (
.I0(CLBLM_L_X8Y107_SLICE_X10Y107_DO6),
.I1(CLBLM_R_X7Y107_SLICE_X8Y107_AO6),
.I2(CLBLM_R_X7Y110_SLICE_X9Y110_BO6),
.I3(CLBLM_L_X8Y109_SLICE_X10Y109_CO6),
.I4(CLBLM_R_X5Y112_SLICE_X7Y112_DO6),
.I5(CLBLM_R_X7Y106_SLICE_X8Y106_DO6),
.O5(CLBLM_R_X7Y110_SLICE_X8Y110_CO5),
.O6(CLBLM_R_X7Y110_SLICE_X8Y110_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h7bf3ffff12305af0)
  ) CLBLM_R_X7Y110_SLICE_X8Y110_BLUT (
.I0(LIOB33_X0Y117_IOB_X0Y117_I),
.I1(LIOB33_X0Y115_IOB_X0Y116_I),
.I2(CLBLM_L_X8Y108_SLICE_X11Y108_CO6),
.I3(LIOB33_X0Y109_IOB_X0Y110_I),
.I4(LIOB33_X0Y111_IOB_X0Y111_I),
.I5(CLBLM_R_X7Y108_SLICE_X9Y108_CO6),
.O5(CLBLM_R_X7Y110_SLICE_X8Y110_BO5),
.O6(CLBLM_R_X7Y110_SLICE_X8Y110_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hc3699999693ccccc)
  ) CLBLM_R_X7Y110_SLICE_X8Y110_ALUT (
.I0(CLBLM_R_X7Y110_SLICE_X8Y110_BO6),
.I1(CLBLM_L_X8Y110_SLICE_X10Y110_AO6),
.I2(LIOB33_X0Y117_IOB_X0Y117_I),
.I3(LIOB33_X0Y115_IOB_X0Y116_I),
.I4(LIOB33_X0Y111_IOB_X0Y112_I),
.I5(CLBLM_L_X8Y111_SLICE_X10Y111_BO6),
.O5(CLBLM_R_X7Y110_SLICE_X8Y110_AO5),
.O6(CLBLM_R_X7Y110_SLICE_X8Y110_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h9c936c936c9c6c6c)
  ) CLBLM_R_X7Y110_SLICE_X9Y110_DLUT (
.I0(LIOB33_X0Y109_IOB_X0Y110_I),
.I1(CLBLM_L_X8Y109_SLICE_X10Y109_CO6),
.I2(RIOB33_X105Y107_IOB_X1Y108_I),
.I3(CLBLM_L_X10Y110_SLICE_X13Y110_DO6),
.I4(LIOB33_X0Y109_IOB_X0Y109_I),
.I5(CLBLM_L_X8Y109_SLICE_X10Y109_BO6),
.O5(CLBLM_R_X7Y110_SLICE_X9Y110_DO5),
.O6(CLBLM_R_X7Y110_SLICE_X9Y110_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h1f7f13137f7f1f7f)
  ) CLBLM_R_X7Y110_SLICE_X9Y110_CLUT (
.I0(LIOB33_X0Y109_IOB_X0Y110_I),
.I1(CLBLM_L_X8Y109_SLICE_X10Y109_CO6),
.I2(RIOB33_X105Y107_IOB_X1Y108_I),
.I3(LIOB33_X0Y109_IOB_X0Y109_I),
.I4(CLBLM_L_X10Y110_SLICE_X13Y110_DO6),
.I5(CLBLM_L_X8Y109_SLICE_X10Y109_BO6),
.O5(CLBLM_R_X7Y110_SLICE_X9Y110_CO5),
.O6(CLBLM_R_X7Y110_SLICE_X9Y110_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h022223335aaaa555)
  ) CLBLM_R_X7Y110_SLICE_X9Y110_BLUT (
.I0(CLBLM_L_X10Y110_SLICE_X13Y110_DO6),
.I1(CLBLM_L_X8Y109_SLICE_X10Y109_CO6),
.I2(LIOB33_X0Y109_IOB_X0Y109_I),
.I3(RIOB33_X105Y107_IOB_X1Y108_I),
.I4(CLBLM_L_X8Y109_SLICE_X10Y109_BO6),
.I5(1'b1),
.O5(CLBLM_R_X7Y110_SLICE_X9Y110_BO5),
.O6(CLBLM_R_X7Y110_SLICE_X9Y110_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h3cccc3333fff0333)
  ) CLBLM_R_X7Y110_SLICE_X9Y110_ALUT (
.I0(1'b1),
.I1(CLBLM_R_X7Y109_SLICE_X9Y109_BO6),
.I2(LIOB33_X0Y111_IOB_X0Y111_I),
.I3(RIOB33_X105Y107_IOB_X1Y108_I),
.I4(CLBLM_R_X7Y110_SLICE_X9Y110_CO6),
.I5(1'b1),
.O5(CLBLM_R_X7Y110_SLICE_X9Y110_AO5),
.O6(CLBLM_R_X7Y110_SLICE_X9Y110_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X7Y111_SLICE_X8Y111_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y111_SLICE_X8Y111_DO5),
.O6(CLBLM_R_X7Y111_SLICE_X8Y111_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X7Y111_SLICE_X8Y111_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y111_SLICE_X8Y111_CO5),
.O6(CLBLM_R_X7Y111_SLICE_X8Y111_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h8fe37f13701c80ec)
  ) CLBLM_R_X7Y111_SLICE_X8Y111_BLUT (
.I0(RIOB33_X105Y103_IOB_X1Y103_I),
.I1(CLBLM_L_X8Y111_SLICE_X10Y111_AO6),
.I2(LIOB33_X0Y111_IOB_X0Y111_I),
.I3(CLBLM_L_X10Y111_SLICE_X12Y111_CO6),
.I4(RIOB33_X105Y103_IOB_X1Y104_I),
.I5(CLBLM_L_X8Y111_SLICE_X11Y111_BO6),
.O5(CLBLM_R_X7Y111_SLICE_X8Y111_BO5),
.O6(CLBLM_R_X7Y111_SLICE_X8Y111_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'ha5a555553f03ff33)
  ) CLBLM_R_X7Y111_SLICE_X8Y111_ALUT (
.I0(CLBLM_L_X8Y111_SLICE_X10Y111_AO5),
.I1(CLBLM_L_X8Y111_SLICE_X10Y111_AO6),
.I2(RIOB33_X105Y103_IOB_X1Y103_I),
.I3(CLBLM_L_X10Y111_SLICE_X12Y111_CO6),
.I4(LIOB33_X0Y111_IOB_X0Y111_I),
.I5(1'b1),
.O5(CLBLM_R_X7Y111_SLICE_X8Y111_AO5),
.O6(CLBLM_R_X7Y111_SLICE_X8Y111_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X7Y111_SLICE_X9Y111_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y111_SLICE_X9Y111_DO5),
.O6(CLBLM_R_X7Y111_SLICE_X9Y111_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h10f5f3fff7ffffff)
  ) CLBLM_R_X7Y111_SLICE_X9Y111_CLUT (
.I0(LIOB33_X0Y105_IOB_X0Y106_I),
.I1(LIOB33_X0Y107_IOB_X0Y108_I),
.I2(CLBLM_L_X10Y109_SLICE_X12Y109_DO6),
.I3(RIOB33_X105Y109_IOB_X1Y110_I),
.I4(RIOB33_X105Y111_IOB_X1Y111_I),
.I5(LIOB33_X0Y107_IOB_X0Y107_I),
.O5(CLBLM_R_X7Y111_SLICE_X9Y111_CO5),
.O6(CLBLM_R_X7Y111_SLICE_X9Y111_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'he26ac0c084a66ac0)
  ) CLBLM_R_X7Y111_SLICE_X9Y111_BLUT (
.I0(RIOB33_X105Y111_IOB_X1Y111_I),
.I1(RIOB33_X105Y109_IOB_X1Y110_I),
.I2(LIOB33_X0Y109_IOB_X0Y110_I),
.I3(LIOB33_X0Y107_IOB_X0Y108_I),
.I4(LIOB33_X0Y109_IOB_X0Y109_I),
.I5(CLBLM_R_X7Y111_SLICE_X9Y111_CO6),
.O5(CLBLM_R_X7Y111_SLICE_X9Y111_BO5),
.O6(CLBLM_R_X7Y111_SLICE_X9Y111_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h3fc0c03f3fff003f)
  ) CLBLM_R_X7Y111_SLICE_X9Y111_ALUT (
.I0(1'b1),
.I1(RIOB33_X105Y109_IOB_X1Y109_I),
.I2(LIOB33_X0Y111_IOB_X0Y111_I),
.I3(CLBLM_R_X7Y111_SLICE_X9Y111_BO6),
.I4(CLBLM_R_X7Y109_SLICE_X9Y109_DO6),
.I5(1'b1),
.O5(CLBLM_R_X7Y111_SLICE_X9Y111_AO5),
.O6(CLBLM_R_X7Y111_SLICE_X9Y111_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X7Y112_SLICE_X8Y112_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y112_SLICE_X8Y112_DO5),
.O6(CLBLM_R_X7Y112_SLICE_X8Y112_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h505570f775f7ffff)
  ) CLBLM_R_X7Y112_SLICE_X8Y112_CLUT (
.I0(RIOB33_X105Y101_IOB_X1Y101_I),
.I1(LIOB33_X0Y111_IOB_X0Y112_I),
.I2(CLBLM_L_X8Y112_SLICE_X11Y112_CO6),
.I3(CLBLM_L_X8Y112_SLICE_X11Y112_BO6),
.I4(LIOB33_X0Y113_IOB_X0Y113_I),
.I5(CLBLM_R_X7Y112_SLICE_X8Y112_BO6),
.O5(CLBLM_R_X7Y112_SLICE_X8Y112_CO5),
.O6(CLBLM_R_X7Y112_SLICE_X8Y112_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h69c39933963c66cc)
  ) CLBLM_R_X7Y112_SLICE_X8Y112_BLUT (
.I0(RIOB33_X105Y101_IOB_X1Y102_I),
.I1(CLBLM_L_X8Y112_SLICE_X11Y112_DO6),
.I2(LIOB33_X0Y111_IOB_X0Y111_I),
.I3(LIOB33_X0Y111_IOB_X0Y112_I),
.I4(RIOB33_X105Y103_IOB_X1Y103_I),
.I5(CLBLM_L_X8Y111_SLICE_X10Y111_AO5),
.O5(CLBLM_R_X7Y112_SLICE_X8Y112_BO5),
.O6(CLBLM_R_X7Y112_SLICE_X8Y112_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h3f3f3f3fd52a40bf)
  ) CLBLM_R_X7Y112_SLICE_X8Y112_ALUT (
.I0(CLBLM_L_X8Y112_SLICE_X11Y112_CO6),
.I1(LIOB33_X0Y111_IOB_X0Y112_I),
.I2(RIOB33_X105Y101_IOB_X1Y101_I),
.I3(CLBLM_R_X7Y112_SLICE_X8Y112_BO6),
.I4(CLBLM_L_X8Y112_SLICE_X11Y112_BO6),
.I5(1'b1),
.O5(CLBLM_R_X7Y112_SLICE_X8Y112_AO5),
.O6(CLBLM_R_X7Y112_SLICE_X8Y112_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'he27b1d846a3f95c0)
  ) CLBLM_R_X7Y112_SLICE_X9Y112_DLUT (
.I0(CLBLM_R_X7Y110_SLICE_X8Y110_BO6),
.I1(LIOB33_X0Y115_IOB_X0Y116_I),
.I2(LIOB33_X0Y113_IOB_X0Y113_I),
.I3(CLBLM_L_X8Y111_SLICE_X10Y111_BO6),
.I4(CLBLM_L_X8Y110_SLICE_X10Y110_BO6),
.I5(LIOB33_X0Y111_IOB_X0Y112_I),
.O5(CLBLM_R_X7Y112_SLICE_X9Y112_DO5),
.O6(CLBLM_R_X7Y112_SLICE_X9Y112_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h48dedede88eeeeee)
  ) CLBLM_R_X7Y112_SLICE_X9Y112_CLUT (
.I0(CLBLM_L_X8Y112_SLICE_X10Y112_BO6),
.I1(CLBLM_L_X8Y112_SLICE_X10Y112_AO5),
.I2(LIOB33_X0Y111_IOB_X0Y112_I),
.I3(LIOB33_X0Y117_IOB_X0Y117_I),
.I4(LIOB33_X0Y113_IOB_X0Y113_I),
.I5(RIOB33_X105Y101_IOB_X1Y101_I),
.O5(CLBLM_R_X7Y112_SLICE_X9Y112_CO5),
.O6(CLBLM_R_X7Y112_SLICE_X9Y112_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h377f07377f7f077f)
  ) CLBLM_R_X7Y112_SLICE_X9Y112_BLUT (
.I0(LIOB33_X0Y113_IOB_X0Y113_I),
.I1(LIOB33_X0Y115_IOB_X0Y116_I),
.I2(CLBLM_L_X8Y110_SLICE_X10Y110_BO6),
.I3(CLBLM_L_X8Y111_SLICE_X10Y111_BO6),
.I4(CLBLM_R_X7Y110_SLICE_X8Y110_BO6),
.I5(LIOB33_X0Y111_IOB_X0Y112_I),
.O5(CLBLM_R_X7Y112_SLICE_X9Y112_BO5),
.O6(CLBLM_R_X7Y112_SLICE_X9Y112_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h87ff7800e1331ecc)
  ) CLBLM_R_X7Y112_SLICE_X9Y112_ALUT (
.I0(LIOB33_X0Y117_IOB_X0Y117_I),
.I1(CLBLM_L_X8Y112_SLICE_X11Y112_AO6),
.I2(RIOB33_X105Y101_IOB_X1Y101_I),
.I3(LIOB33_X0Y111_IOB_X0Y112_I),
.I4(CLBLM_L_X8Y112_SLICE_X10Y112_BO6),
.I5(CLBLM_L_X8Y111_SLICE_X10Y111_CO6),
.O5(CLBLM_R_X7Y112_SLICE_X9Y112_AO5),
.O6(CLBLM_R_X7Y112_SLICE_X9Y112_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h15ff01777fff5777)
  ) CLBLM_R_X7Y113_SLICE_X8Y113_DLUT (
.I0(CLBLM_R_X5Y111_SLICE_X7Y111_BO6),
.I1(CLBLM_R_X5Y110_SLICE_X7Y110_AO5),
.I2(LIOB33_X0Y113_IOB_X0Y113_I),
.I3(RIOB33_X105Y107_IOB_X1Y107_I),
.I4(CLBLM_R_X7Y113_SLICE_X8Y113_BO5),
.I5(LIOB33_X0Y115_IOB_X0Y115_I),
.O5(CLBLM_R_X7Y113_SLICE_X8Y113_DO5),
.O6(CLBLM_R_X7Y113_SLICE_X8Y113_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h95aaa9666aaa5666)
  ) CLBLM_R_X7Y113_SLICE_X8Y113_CLUT (
.I0(CLBLM_R_X5Y111_SLICE_X7Y111_BO6),
.I1(CLBLM_R_X5Y110_SLICE_X7Y110_AO5),
.I2(LIOB33_X0Y113_IOB_X0Y113_I),
.I3(RIOB33_X105Y107_IOB_X1Y107_I),
.I4(CLBLM_R_X7Y113_SLICE_X8Y113_BO5),
.I5(LIOB33_X0Y115_IOB_X0Y115_I),
.O5(CLBLM_R_X7Y113_SLICE_X8Y113_CO5),
.O6(CLBLM_R_X7Y113_SLICE_X8Y113_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h3cc3c3c30ccfcfcf)
  ) CLBLM_R_X7Y113_SLICE_X8Y113_BLUT (
.I0(1'b1),
.I1(CLBLM_R_X7Y113_SLICE_X9Y113_BO6),
.I2(CLBLM_R_X7Y110_SLICE_X9Y110_AO6),
.I3(RIOB33_X105Y107_IOB_X1Y107_I),
.I4(LIOB33_X0Y111_IOB_X0Y112_I),
.I5(1'b1),
.O5(CLBLM_R_X7Y113_SLICE_X8Y113_BO5),
.O6(CLBLM_R_X7Y113_SLICE_X8Y113_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h5f5f5f5f66cc9933)
  ) CLBLM_R_X7Y113_SLICE_X8Y113_ALUT (
.I0(LIOB33_X0Y113_IOB_X0Y113_I),
.I1(CLBLM_R_X7Y113_SLICE_X8Y113_BO5),
.I2(RIOB33_X105Y103_IOB_X1Y104_I),
.I3(RIOB33_X105Y107_IOB_X1Y107_I),
.I4(CLBLM_R_X5Y110_SLICE_X7Y110_AO5),
.I5(1'b1),
.O5(CLBLM_R_X7Y113_SLICE_X8Y113_AO5),
.O6(CLBLM_R_X7Y113_SLICE_X8Y113_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h1f7f005f5fff1f7f)
  ) CLBLM_R_X7Y113_SLICE_X9Y113_DLUT (
.I0(LIOB33_X0Y111_IOB_X0Y112_I),
.I1(LIOB33_X0Y111_IOB_X0Y111_I),
.I2(RIOB33_X105Y105_IOB_X1Y105_I),
.I3(CLBLM_R_X7Y113_SLICE_X9Y113_CO6),
.I4(CLBLM_L_X8Y111_SLICE_X11Y111_AO5),
.I5(CLBLM_L_X8Y113_SLICE_X10Y113_AO5),
.O5(CLBLM_R_X7Y113_SLICE_X9Y113_DO5),
.O6(CLBLM_R_X7Y113_SLICE_X9Y113_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hd2b4781e5a96f03c)
  ) CLBLM_R_X7Y113_SLICE_X9Y113_CLUT (
.I0(RIOB33_X105Y107_IOB_X1Y107_I),
.I1(CLBLM_R_X7Y110_SLICE_X9Y110_BO5),
.I2(CLBLM_R_X7Y110_SLICE_X9Y110_DO6),
.I3(CLBLM_L_X10Y112_SLICE_X13Y112_BO6),
.I4(LIOB33_X0Y111_IOB_X0Y111_I),
.I5(LIOB33_X0Y109_IOB_X0Y110_I),
.O5(CLBLM_R_X7Y113_SLICE_X9Y113_CO5),
.O6(CLBLM_R_X7Y113_SLICE_X9Y113_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h1f7f5fff07571777)
  ) CLBLM_R_X7Y113_SLICE_X9Y113_BLUT (
.I0(CLBLM_R_X7Y110_SLICE_X9Y110_DO6),
.I1(CLBLM_R_X7Y110_SLICE_X9Y110_BO5),
.I2(RIOB33_X105Y107_IOB_X1Y107_I),
.I3(LIOB33_X0Y111_IOB_X0Y111_I),
.I4(LIOB33_X0Y109_IOB_X0Y110_I),
.I5(CLBLM_L_X10Y112_SLICE_X13Y112_BO6),
.O5(CLBLM_R_X7Y113_SLICE_X9Y113_BO5),
.O6(CLBLM_R_X7Y113_SLICE_X9Y113_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hd24bbbbb2db44444)
  ) CLBLM_R_X7Y113_SLICE_X9Y113_ALUT (
.I0(CLBLM_L_X8Y111_SLICE_X11Y111_AO5),
.I1(CLBLM_L_X8Y113_SLICE_X10Y113_AO5),
.I2(LIOB33_X0Y111_IOB_X0Y112_I),
.I3(LIOB33_X0Y111_IOB_X0Y111_I),
.I4(RIOB33_X105Y105_IOB_X1Y105_I),
.I5(CLBLM_R_X7Y113_SLICE_X9Y113_CO6),
.O5(CLBLM_R_X7Y113_SLICE_X9Y113_AO5),
.O6(CLBLM_R_X7Y113_SLICE_X9Y113_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h13017f37ff77ff77)
  ) CLBLM_R_X7Y114_SLICE_X8Y114_DLUT (
.I0(CLBLM_R_X7Y113_SLICE_X8Y113_BO6),
.I1(CLBLM_R_X7Y113_SLICE_X8Y113_AO5),
.I2(LIOB33_X0Y113_IOB_X0Y113_I),
.I3(CLBLM_R_X7Y113_SLICE_X9Y113_DO6),
.I4(LIOB33_X0Y115_IOB_X0Y115_I),
.I5(RIOB33_X105Y105_IOB_X1Y105_I),
.O5(CLBLM_R_X7Y114_SLICE_X8Y114_DO5),
.O6(CLBLM_R_X7Y114_SLICE_X8Y114_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h93c96c36cc66cc66)
  ) CLBLM_R_X7Y114_SLICE_X8Y114_CLUT (
.I0(CLBLM_R_X7Y113_SLICE_X8Y113_BO6),
.I1(CLBLM_R_X7Y113_SLICE_X8Y113_AO5),
.I2(LIOB33_X0Y113_IOB_X0Y113_I),
.I3(CLBLM_R_X7Y113_SLICE_X9Y113_DO6),
.I4(LIOB33_X0Y115_IOB_X0Y115_I),
.I5(RIOB33_X105Y105_IOB_X1Y105_I),
.O5(CLBLM_R_X7Y114_SLICE_X8Y114_CO5),
.O6(CLBLM_R_X7Y114_SLICE_X8Y114_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h599aa665a665599a)
  ) CLBLM_R_X7Y114_SLICE_X8Y114_BLUT (
.I0(CLBLM_R_X7Y113_SLICE_X8Y113_BO6),
.I1(CLBLM_R_X7Y113_SLICE_X9Y113_AO6),
.I2(CLBLM_R_X7Y113_SLICE_X8Y113_AO6),
.I3(CLBLM_L_X8Y113_SLICE_X10Y113_CO6),
.I4(CLBLM_R_X7Y114_SLICE_X8Y114_AO6),
.I5(CLBLM_R_X7Y113_SLICE_X9Y113_DO6),
.O5(CLBLM_R_X7Y114_SLICE_X8Y114_BO5),
.O6(CLBLM_R_X7Y114_SLICE_X8Y114_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h5f5f5f5f5fa0a05f)
  ) CLBLM_R_X7Y114_SLICE_X8Y114_ALUT (
.I0(LIOB33_X0Y113_IOB_X0Y113_I),
.I1(1'b1),
.I2(RIOB33_X105Y105_IOB_X1Y105_I),
.I3(CLBLM_R_X7Y113_SLICE_X9Y113_DO6),
.I4(CLBLM_R_X7Y113_SLICE_X8Y113_BO6),
.I5(1'b1),
.O5(CLBLM_R_X7Y114_SLICE_X8Y114_AO5),
.O6(CLBLM_R_X7Y114_SLICE_X8Y114_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X7Y114_SLICE_X9Y114_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y114_SLICE_X9Y114_DO5),
.O6(CLBLM_R_X7Y114_SLICE_X9Y114_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X7Y114_SLICE_X9Y114_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y114_SLICE_X9Y114_CO5),
.O6(CLBLM_R_X7Y114_SLICE_X9Y114_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X7Y114_SLICE_X9Y114_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y114_SLICE_X9Y114_BO5),
.O6(CLBLM_R_X7Y114_SLICE_X9Y114_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X7Y114_SLICE_X9Y114_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y114_SLICE_X9Y114_AO5),
.O6(CLBLM_R_X7Y114_SLICE_X9Y114_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h69696966c3ccc3cc)
  ) CLBLM_R_X11Y104_SLICE_X14Y104_DLUT (
.I0(RIOB33_X105Y105_IOB_X1Y105_I),
.I1(CLBLM_R_X11Y104_SLICE_X15Y104_CO6),
.I2(CLBLM_R_X11Y104_SLICE_X15Y104_DO6),
.I3(CLBLM_R_X11Y104_SLICE_X15Y104_BO6),
.I4(RIOB33_X105Y103_IOB_X1Y104_I),
.I5(LIOB33_X0Y101_IOB_X0Y101_I),
.O5(CLBLM_R_X11Y104_SLICE_X14Y104_DO5),
.O6(CLBLM_R_X11Y104_SLICE_X14Y104_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hfcc0fec8f330fb32)
  ) CLBLM_R_X11Y104_SLICE_X14Y104_CLUT (
.I0(CLBLM_R_X11Y104_SLICE_X14Y104_AO6),
.I1(CLBLM_R_X11Y104_SLICE_X15Y104_CO6),
.I2(CLBLM_R_X11Y104_SLICE_X15Y104_DO6),
.I3(CLBLM_R_X11Y104_SLICE_X14Y104_AO5),
.I4(CLBLM_R_X11Y104_SLICE_X15Y104_BO6),
.I5(CLBLM_L_X12Y104_SLICE_X16Y104_AO6),
.O5(CLBLM_R_X11Y104_SLICE_X14Y104_CO5),
.O6(CLBLM_R_X11Y104_SLICE_X14Y104_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h59a65aa5a659a55a)
  ) CLBLM_R_X11Y104_SLICE_X14Y104_BLUT (
.I0(CLBLM_R_X11Y104_SLICE_X15Y104_CO6),
.I1(CLBLM_R_X11Y104_SLICE_X15Y104_BO6),
.I2(CLBLM_R_X11Y104_SLICE_X15Y104_DO6),
.I3(CLBLM_L_X12Y104_SLICE_X16Y104_AO6),
.I4(CLBLM_R_X11Y104_SLICE_X14Y104_AO6),
.I5(CLBLM_R_X11Y104_SLICE_X14Y104_AO5),
.O5(CLBLM_R_X11Y104_SLICE_X14Y104_BO5),
.O6(CLBLM_R_X11Y104_SLICE_X14Y104_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h3333ffff00ffffff)
  ) CLBLM_R_X11Y104_SLICE_X14Y104_ALUT (
.I0(1'b1),
.I1(LIOB33_X0Y101_IOB_X0Y101_I),
.I2(1'b1),
.I3(LIOB33_X0Y101_IOB_X0Y102_I),
.I4(RIOB33_X105Y103_IOB_X1Y104_I),
.I5(1'b1),
.O5(CLBLM_R_X11Y104_SLICE_X14Y104_AO5),
.O6(CLBLM_R_X11Y104_SLICE_X14Y104_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h20206a600020ca60)
  ) CLBLM_R_X11Y104_SLICE_X15Y104_DLUT (
.I0(RIOB33_X105Y113_IOB_X1Y113_I),
.I1(LIOB33_SING_X0Y100_IOB_X0Y100_I),
.I2(RIOB33_X105Y105_IOB_X1Y105_I),
.I3(RIOB33_X105Y107_IOB_X1Y107_I),
.I4(RIOB33_X105Y103_IOB_X1Y104_I),
.I5(RIOB33_X105Y111_IOB_X1Y112_I),
.O5(CLBLM_R_X11Y104_SLICE_X15Y104_DO5),
.O6(CLBLM_R_X11Y104_SLICE_X15Y104_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h462c0a2c46e0c6e0)
  ) CLBLM_R_X11Y104_SLICE_X15Y104_CLUT (
.I0(LIOB33_SING_X0Y100_IOB_X0Y100_I),
.I1(RIOB33_X105Y113_IOB_X1Y113_I),
.I2(RIOB33_X105Y105_IOB_X1Y105_I),
.I3(RIOB33_X105Y107_IOB_X1Y107_I),
.I4(RIOB33_X105Y111_IOB_X1Y112_I),
.I5(RIOB33_X105Y107_IOB_X1Y108_I),
.O5(CLBLM_R_X11Y104_SLICE_X15Y104_CO5),
.O6(CLBLM_R_X11Y104_SLICE_X15Y104_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h125a0ff0dd5a0000)
  ) CLBLM_R_X11Y104_SLICE_X15Y104_BLUT (
.I0(RIOB33_X105Y107_IOB_X1Y107_I),
.I1(RIOB33_X105Y111_IOB_X1Y112_I),
.I2(RIOB33_X105Y103_IOB_X1Y104_I),
.I3(RIOB33_X105Y105_IOB_X1Y105_I),
.I4(RIOB33_X105Y113_IOB_X1Y113_I),
.I5(LIOB33_SING_X0Y100_IOB_X0Y100_I),
.O5(CLBLM_R_X11Y104_SLICE_X15Y104_BO5),
.O6(CLBLM_R_X11Y104_SLICE_X15Y104_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'ha05fa05fffff005f)
  ) CLBLM_R_X11Y104_SLICE_X15Y104_ALUT (
.I0(RIOB33_X105Y103_IOB_X1Y104_I),
.I1(1'b1),
.I2(LIOB33_X0Y101_IOB_X0Y101_I),
.I3(CLBLM_R_X11Y104_SLICE_X15Y104_BO6),
.I4(CLBLM_R_X11Y104_SLICE_X15Y104_DO6),
.I5(1'b1),
.O5(CLBLM_R_X11Y104_SLICE_X15Y104_AO5),
.O6(CLBLM_R_X11Y104_SLICE_X15Y104_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h7dfff5ff143c50f0)
  ) CLBLM_R_X11Y105_SLICE_X14Y105_DLUT (
.I0(RIOB33_X105Y103_IOB_X1Y103_I),
.I1(LIOB33_X0Y101_IOB_X0Y102_I),
.I2(CLBLM_R_X11Y104_SLICE_X14Y104_DO6),
.I3(LIOB33_X0Y103_IOB_X0Y104_I),
.I4(RIOB33_X105Y103_IOB_X1Y104_I),
.I5(CLBLM_L_X10Y104_SLICE_X13Y104_DO6),
.O5(CLBLM_R_X11Y105_SLICE_X14Y105_DO5),
.O6(CLBLM_R_X11Y105_SLICE_X14Y105_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h69c3a50f963c5af0)
  ) CLBLM_R_X11Y105_SLICE_X14Y105_CLUT (
.I0(RIOB33_X105Y103_IOB_X1Y103_I),
.I1(LIOB33_X0Y101_IOB_X0Y102_I),
.I2(CLBLM_R_X11Y104_SLICE_X14Y104_DO6),
.I3(LIOB33_X0Y103_IOB_X0Y104_I),
.I4(RIOB33_X105Y103_IOB_X1Y104_I),
.I5(CLBLM_L_X10Y104_SLICE_X13Y104_DO6),
.O5(CLBLM_R_X11Y105_SLICE_X14Y105_CO5),
.O6(CLBLM_R_X11Y105_SLICE_X14Y105_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h6969966996699696)
  ) CLBLM_R_X11Y105_SLICE_X14Y105_BLUT (
.I0(CLBLM_L_X12Y104_SLICE_X16Y104_BO6),
.I1(CLBLM_R_X11Y104_SLICE_X14Y104_CO6),
.I2(CLBLM_R_X11Y105_SLICE_X15Y105_AO6),
.I3(CLBLM_R_X11Y104_SLICE_X14Y104_BO6),
.I4(CLBLM_R_X11Y105_SLICE_X14Y105_AO6),
.I5(CLBLM_L_X10Y104_SLICE_X13Y104_DO6),
.O5(CLBLM_R_X11Y105_SLICE_X14Y105_BO5),
.O6(CLBLM_R_X11Y105_SLICE_X14Y105_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h3f3f3f3f33ff33ff)
  ) CLBLM_R_X11Y105_SLICE_X14Y105_ALUT (
.I0(1'b1),
.I1(RIOB33_X105Y103_IOB_X1Y103_I),
.I2(LIOB33_X0Y103_IOB_X0Y104_I),
.I3(LIOB33_X0Y105_IOB_X0Y105_I),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X11Y105_SLICE_X14Y105_AO5),
.O6(CLBLM_R_X11Y105_SLICE_X14Y105_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hbc2f4cdf43d0b320)
  ) CLBLM_R_X11Y105_SLICE_X15Y105_DLUT (
.I0(RIOB33_X105Y103_IOB_X1Y104_I),
.I1(CLBLM_R_X11Y104_SLICE_X15Y104_AO5),
.I2(LIOB33_X0Y101_IOB_X0Y102_I),
.I3(CLBLM_L_X12Y105_SLICE_X16Y105_AO5),
.I4(RIOB33_X105Y105_IOB_X1Y105_I),
.I5(CLBLM_L_X12Y105_SLICE_X16Y105_CO6),
.O5(CLBLM_R_X11Y105_SLICE_X15Y105_DO5),
.O6(CLBLM_R_X11Y105_SLICE_X15Y105_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h2abfbfbfbf2a2a2a)
  ) CLBLM_R_X11Y105_SLICE_X15Y105_CLUT (
.I0(CLBLM_R_X11Y104_SLICE_X14Y104_CO6),
.I1(LIOB33_X0Y103_IOB_X0Y104_I),
.I2(RIOB33_X105Y103_IOB_X1Y104_I),
.I3(LIOB33_X0Y101_IOB_X0Y102_I),
.I4(RIOB33_X105Y105_IOB_X1Y105_I),
.I5(CLBLM_L_X12Y105_SLICE_X16Y105_CO6),
.O5(CLBLM_R_X11Y105_SLICE_X15Y105_CO5),
.O6(CLBLM_R_X11Y105_SLICE_X15Y105_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h69999666c3333ccc)
  ) CLBLM_R_X11Y105_SLICE_X15Y105_BLUT (
.I0(RIOB33_X105Y105_IOB_X1Y105_I),
.I1(CLBLM_L_X12Y105_SLICE_X16Y105_CO6),
.I2(LIOB33_X0Y103_IOB_X0Y104_I),
.I3(RIOB33_X105Y103_IOB_X1Y104_I),
.I4(CLBLM_R_X11Y104_SLICE_X14Y104_CO6),
.I5(LIOB33_X0Y101_IOB_X0Y102_I),
.O5(CLBLM_R_X11Y105_SLICE_X15Y105_BO5),
.O6(CLBLM_R_X11Y105_SLICE_X15Y105_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h3f3f3f3f33ff33ff)
  ) CLBLM_R_X11Y105_SLICE_X15Y105_ALUT (
.I0(1'b1),
.I1(RIOB33_X105Y103_IOB_X1Y104_I),
.I2(LIOB33_X0Y103_IOB_X0Y104_I),
.I3(LIOB33_X0Y105_IOB_X0Y105_I),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X11Y105_SLICE_X15Y105_AO5),
.O6(CLBLM_R_X11Y105_SLICE_X15Y105_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h87e1ff55781e00aa)
  ) CLBLM_R_X11Y106_SLICE_X14Y106_DLUT (
.I0(CLBLM_R_X11Y105_SLICE_X15Y105_BO6),
.I1(RIOB33_X105Y103_IOB_X1Y103_I),
.I2(RIOB33_X105Y103_IOB_X1Y104_I),
.I3(CLBLM_R_X11Y105_SLICE_X14Y105_DO6),
.I4(LIOB33_X0Y105_IOB_X0Y105_I),
.I5(CLBLM_R_X11Y106_SLICE_X14Y106_BO6),
.O5(CLBLM_R_X11Y106_SLICE_X14Y106_DO5),
.O6(CLBLM_R_X11Y106_SLICE_X14Y106_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'he8a0fae88e0aaf8e)
  ) CLBLM_R_X11Y106_SLICE_X14Y106_CLUT (
.I0(CLBLM_R_X11Y109_SLICE_X14Y109_AO6),
.I1(CLBLM_R_X11Y105_SLICE_X14Y105_AO5),
.I2(CLBLM_R_X11Y105_SLICE_X15Y105_AO5),
.I3(CLBLM_R_X11Y105_SLICE_X14Y105_DO6),
.I4(CLBLM_R_X11Y105_SLICE_X15Y105_BO6),
.I5(CLBLM_R_X11Y106_SLICE_X14Y106_BO6),
.O5(CLBLM_R_X11Y106_SLICE_X14Y106_CO5),
.O6(CLBLM_R_X11Y106_SLICE_X14Y106_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h639cc6399c6339c6)
  ) CLBLM_R_X11Y106_SLICE_X14Y106_BLUT (
.I0(CLBLM_R_X11Y105_SLICE_X15Y105_AO6),
.I1(CLBLM_L_X12Y106_SLICE_X17Y106_BO6),
.I2(CLBLM_L_X12Y104_SLICE_X16Y104_BO6),
.I3(CLBLM_R_X11Y107_SLICE_X14Y107_AO6),
.I4(CLBLM_R_X11Y104_SLICE_X14Y104_CO6),
.I5(CLBLM_L_X12Y104_SLICE_X16Y104_DO6),
.O5(CLBLM_R_X11Y106_SLICE_X14Y106_BO5),
.O6(CLBLM_R_X11Y106_SLICE_X14Y106_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h6996696996966996)
  ) CLBLM_R_X11Y106_SLICE_X14Y106_ALUT (
.I0(CLBLM_R_X11Y106_SLICE_X14Y106_BO6),
.I1(CLBLM_R_X11Y105_SLICE_X15Y105_AO5),
.I2(CLBLM_R_X11Y109_SLICE_X14Y109_AO6),
.I3(CLBLM_R_X11Y105_SLICE_X14Y105_DO6),
.I4(CLBLM_R_X11Y105_SLICE_X15Y105_BO6),
.I5(CLBLM_R_X11Y105_SLICE_X14Y105_AO5),
.O5(CLBLM_R_X11Y106_SLICE_X14Y106_AO5),
.O6(CLBLM_R_X11Y106_SLICE_X14Y106_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h71f5f3ffd450fcf0)
  ) CLBLM_R_X11Y106_SLICE_X15Y106_DLUT (
.I0(RIOB33_X105Y109_IOB_X1Y109_I),
.I1(LIOB33_X0Y105_IOB_X0Y105_I),
.I2(CLBLM_R_X11Y107_SLICE_X15Y107_AO5),
.I3(RIOB33_X105Y109_IOB_X1Y110_I),
.I4(LIOB33_X0Y105_IOB_X0Y106_I),
.I5(CLBLM_L_X10Y107_SLICE_X13Y107_CO6),
.O5(CLBLM_R_X11Y106_SLICE_X15Y106_DO5),
.O6(CLBLM_R_X11Y106_SLICE_X15Y106_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h4dd4dd44cffcffcc)
  ) CLBLM_R_X11Y106_SLICE_X15Y106_CLUT (
.I0(RIOB33_X105Y109_IOB_X1Y109_I),
.I1(CLBLM_L_X12Y105_SLICE_X17Y105_AO6),
.I2(LIOB33_X0Y101_IOB_X0Y102_I),
.I3(CLBLM_L_X10Y107_SLICE_X13Y107_DO6),
.I4(RIOB33_X105Y109_IOB_X1Y110_I),
.I5(LIOB33_X0Y103_IOB_X0Y104_I),
.O5(CLBLM_R_X11Y106_SLICE_X15Y106_CO5),
.O6(CLBLM_R_X11Y106_SLICE_X15Y106_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h69a5c30f965a3cf0)
  ) CLBLM_R_X11Y106_SLICE_X15Y106_BLUT (
.I0(RIOB33_X105Y109_IOB_X1Y110_I),
.I1(LIOB33_X0Y103_IOB_X0Y104_I),
.I2(CLBLM_L_X12Y105_SLICE_X17Y105_AO6),
.I3(RIOB33_X105Y109_IOB_X1Y109_I),
.I4(LIOB33_X0Y101_IOB_X0Y102_I),
.I5(CLBLM_L_X10Y107_SLICE_X13Y107_DO6),
.O5(CLBLM_R_X11Y106_SLICE_X15Y106_BO5),
.O6(CLBLM_R_X11Y106_SLICE_X15Y106_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h3333ffff2abf2abf)
  ) CLBLM_R_X11Y106_SLICE_X15Y106_ALUT (
.I0(CLBLM_R_X11Y106_SLICE_X15Y106_DO6),
.I1(RIOB33_X105Y109_IOB_X1Y109_I),
.I2(LIOB33_X0Y107_IOB_X0Y107_I),
.I3(CLBLM_L_X10Y108_SLICE_X13Y108_DO6),
.I4(LIOB33_X0Y101_IOB_X0Y101_I),
.I5(1'b1),
.O5(CLBLM_R_X11Y106_SLICE_X15Y106_AO5),
.O6(CLBLM_R_X11Y106_SLICE_X15Y106_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h9cc6c3ccf50a0000)
  ) CLBLM_R_X11Y107_SLICE_X14Y107_DLUT (
.I0(LIOB33_X0Y101_IOB_X0Y101_I),
.I1(LIOB33_X0Y103_IOB_X0Y104_I),
.I2(CLBLM_L_X10Y107_SLICE_X12Y107_CO6),
.I3(LIOB33_X0Y101_IOB_X0Y102_I),
.I4(RIOB33_X105Y111_IOB_X1Y111_I),
.I5(RIOB33_X105Y109_IOB_X1Y110_I),
.O5(CLBLM_R_X11Y107_SLICE_X14Y107_DO5),
.O6(CLBLM_R_X11Y107_SLICE_X14Y107_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h69c3963c963c963c)
  ) CLBLM_R_X11Y107_SLICE_X14Y107_CLUT (
.I0(LIOB33_X0Y101_IOB_X0Y102_I),
.I1(CLBLM_L_X12Y104_SLICE_X16Y104_DO6),
.I2(CLBLM_L_X12Y106_SLICE_X16Y106_DO6),
.I3(RIOB33_X105Y107_IOB_X1Y107_I),
.I4(LIOB33_X0Y103_IOB_X0Y104_I),
.I5(RIOB33_X105Y105_IOB_X1Y105_I),
.O5(CLBLM_R_X11Y107_SLICE_X14Y107_CO5),
.O6(CLBLM_R_X11Y107_SLICE_X14Y107_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h93939393f00f00ff)
  ) CLBLM_R_X11Y107_SLICE_X14Y107_BLUT (
.I0(LIOB33_X0Y105_IOB_X0Y105_I),
.I1(CLBLM_L_X10Y107_SLICE_X13Y107_CO6),
.I2(RIOB33_X105Y109_IOB_X1Y110_I),
.I3(CLBLM_L_X10Y107_SLICE_X13Y107_DO6),
.I4(LIOB33_X0Y101_IOB_X0Y102_I),
.I5(1'b1),
.O5(CLBLM_R_X11Y107_SLICE_X14Y107_BO5),
.O6(CLBLM_R_X11Y107_SLICE_X14Y107_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h33ff33ff55ff55ff)
  ) CLBLM_R_X11Y107_SLICE_X14Y107_ALUT (
.I0(LIOB33_X0Y105_IOB_X0Y105_I),
.I1(LIOB33_X0Y103_IOB_X0Y104_I),
.I2(1'b1),
.I3(RIOB33_X105Y105_IOB_X1Y105_I),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X11Y107_SLICE_X14Y107_AO5),
.O6(CLBLM_R_X11Y107_SLICE_X14Y107_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h963cf0f0c3960ff0)
  ) CLBLM_R_X11Y107_SLICE_X15Y107_DLUT (
.I0(LIOB33_X0Y103_IOB_X0Y104_I),
.I1(LIOB33_X0Y105_IOB_X0Y105_I),
.I2(CLBLM_R_X11Y107_SLICE_X14Y107_DO6),
.I3(CLBLM_R_X11Y107_SLICE_X14Y107_BO5),
.I4(RIOB33_X105Y109_IOB_X1Y109_I),
.I5(CLBLM_L_X12Y105_SLICE_X17Y105_AO6),
.O5(CLBLM_R_X11Y107_SLICE_X15Y107_DO5),
.O6(CLBLM_R_X11Y107_SLICE_X15Y107_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hf8fe8fef80e0080e)
  ) CLBLM_R_X11Y107_SLICE_X15Y107_CLUT (
.I0(CLBLM_L_X12Y107_SLICE_X16Y107_BO6),
.I1(CLBLM_R_X11Y107_SLICE_X14Y107_AO5),
.I2(CLBLM_L_X12Y108_SLICE_X16Y108_AO6),
.I3(CLBLM_R_X13Y107_SLICE_X18Y107_AO6),
.I4(CLBLM_L_X12Y107_SLICE_X16Y107_AO6),
.I5(CLBLM_R_X11Y111_SLICE_X15Y111_BO6),
.O5(CLBLM_R_X11Y107_SLICE_X15Y107_CO5),
.O6(CLBLM_R_X11Y107_SLICE_X15Y107_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h6996c33c3cc36996)
  ) CLBLM_R_X11Y107_SLICE_X15Y107_BLUT (
.I0(CLBLM_R_X11Y107_SLICE_X14Y107_AO5),
.I1(CLBLM_R_X11Y111_SLICE_X15Y111_BO6),
.I2(CLBLM_L_X12Y107_SLICE_X16Y107_AO6),
.I3(CLBLM_L_X12Y108_SLICE_X16Y108_AO6),
.I4(CLBLM_L_X12Y107_SLICE_X16Y107_BO6),
.I5(CLBLM_R_X13Y107_SLICE_X18Y107_AO6),
.O5(CLBLM_R_X11Y107_SLICE_X15Y107_BO5),
.O6(CLBLM_R_X11Y107_SLICE_X15Y107_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h55ff55ff7f7f1313)
  ) CLBLM_R_X11Y107_SLICE_X15Y107_ALUT (
.I0(RIOB33_X105Y109_IOB_X1Y109_I),
.I1(CLBLM_R_X11Y107_SLICE_X14Y107_DO6),
.I2(LIOB33_X0Y105_IOB_X0Y105_I),
.I3(LIOB33_X0Y103_IOB_X0Y104_I),
.I4(CLBLM_R_X11Y106_SLICE_X15Y106_CO6),
.I5(1'b1),
.O5(CLBLM_R_X11Y107_SLICE_X15Y107_AO5),
.O6(CLBLM_R_X11Y107_SLICE_X15Y107_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h6ac0953f953f6ac0)
  ) CLBLM_R_X11Y108_SLICE_X14Y108_DLUT (
.I0(RIOB33_X105Y103_IOB_X1Y103_I),
.I1(LIOB33_X0Y103_IOB_X0Y104_I),
.I2(RIOB33_X105Y103_IOB_X1Y104_I),
.I3(LIOB33_X0Y105_IOB_X0Y105_I),
.I4(CLBLM_R_X11Y105_SLICE_X15Y105_DO6),
.I5(CLBLM_R_X11Y105_SLICE_X14Y105_DO6),
.O5(CLBLM_R_X11Y108_SLICE_X14Y108_DO5),
.O6(CLBLM_R_X11Y108_SLICE_X14Y108_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h7fff8fff07770888)
  ) CLBLM_R_X11Y108_SLICE_X14Y108_CLUT (
.I0(LIOB33_X0Y103_IOB_X0Y104_I),
.I1(RIOB33_X105Y103_IOB_X1Y104_I),
.I2(RIOB33_X105Y103_IOB_X1Y103_I),
.I3(LIOB33_X0Y105_IOB_X0Y105_I),
.I4(CLBLM_R_X11Y105_SLICE_X15Y105_DO6),
.I5(CLBLM_R_X11Y105_SLICE_X14Y105_DO6),
.O5(CLBLM_R_X11Y108_SLICE_X14Y108_CO5),
.O6(CLBLM_R_X11Y108_SLICE_X14Y108_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h6996996696966666)
  ) CLBLM_R_X11Y108_SLICE_X14Y108_BLUT (
.I0(CLBLM_L_X12Y106_SLICE_X16Y106_CO6),
.I1(CLBLM_R_X11Y105_SLICE_X15Y105_CO6),
.I2(RIOB33_X105Y105_IOB_X1Y105_I),
.I3(RIOB33_X105Y103_IOB_X1Y104_I),
.I4(LIOB33_X0Y103_IOB_X0Y104_I),
.I5(LIOB33_X0Y105_IOB_X0Y105_I),
.O5(CLBLM_R_X11Y108_SLICE_X14Y108_BO5),
.O6(CLBLM_R_X11Y108_SLICE_X14Y108_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hb478787887b48778)
  ) CLBLM_R_X11Y108_SLICE_X14Y108_ALUT (
.I0(RIOB33_X105Y103_IOB_X1Y104_I),
.I1(LIOB33_X0Y105_IOB_X0Y106_I),
.I2(CLBLM_R_X11Y108_SLICE_X15Y108_CO6),
.I3(CLBLM_R_X11Y108_SLICE_X14Y108_BO6),
.I4(RIOB33_X105Y103_IOB_X1Y103_I),
.I5(CLBLM_R_X11Y108_SLICE_X14Y108_CO6),
.O5(CLBLM_R_X11Y108_SLICE_X14Y108_AO5),
.O6(CLBLM_R_X11Y108_SLICE_X14Y108_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h7887877887877878)
  ) CLBLM_R_X11Y108_SLICE_X15Y108_DLUT (
.I0(RIOB33_X105Y107_IOB_X1Y107_I),
.I1(LIOB33_X0Y105_IOB_X0Y105_I),
.I2(CLBLM_L_X12Y107_SLICE_X17Y107_AO5),
.I3(LIOB33_X0Y103_IOB_X0Y104_I),
.I4(CLBLM_L_X12Y107_SLICE_X17Y107_DO6),
.I5(RIOB33_X105Y107_IOB_X1Y108_I),
.O5(CLBLM_R_X11Y108_SLICE_X15Y108_DO5),
.O6(CLBLM_R_X11Y108_SLICE_X15Y108_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h93c96c36cc66cc66)
  ) CLBLM_R_X11Y108_SLICE_X15Y108_CLUT (
.I0(CLBLM_R_X11Y107_SLICE_X14Y107_CO6),
.I1(CLBLM_L_X12Y107_SLICE_X16Y107_CO6),
.I2(RIOB33_X105Y103_IOB_X1Y104_I),
.I3(CLBLM_R_X11Y105_SLICE_X15Y105_CO6),
.I4(RIOB33_X105Y105_IOB_X1Y105_I),
.I5(LIOB33_X0Y105_IOB_X0Y105_I),
.O5(CLBLM_R_X11Y108_SLICE_X15Y108_CO5),
.O6(CLBLM_R_X11Y108_SLICE_X15Y108_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h6996696996966996)
  ) CLBLM_R_X11Y108_SLICE_X15Y108_BLUT (
.I0(CLBLM_R_X11Y111_SLICE_X15Y111_AO5),
.I1(CLBLM_L_X12Y107_SLICE_X16Y107_CO6),
.I2(CLBLM_R_X11Y107_SLICE_X14Y107_AO5),
.I3(CLBLM_R_X11Y105_SLICE_X15Y105_AO5),
.I4(CLBLM_R_X11Y107_SLICE_X14Y107_CO6),
.I5(CLBLM_R_X11Y105_SLICE_X15Y105_CO6),
.O5(CLBLM_R_X11Y108_SLICE_X15Y108_BO5),
.O6(CLBLM_R_X11Y108_SLICE_X15Y108_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'heb82ebeb8282eb82)
  ) CLBLM_R_X11Y108_SLICE_X15Y108_ALUT (
.I0(CLBLM_R_X11Y111_SLICE_X15Y111_AO5),
.I1(CLBLM_L_X12Y107_SLICE_X16Y107_CO6),
.I2(CLBLM_R_X11Y107_SLICE_X14Y107_AO5),
.I3(CLBLM_R_X11Y105_SLICE_X15Y105_AO5),
.I4(CLBLM_R_X11Y107_SLICE_X14Y107_CO6),
.I5(CLBLM_R_X11Y105_SLICE_X15Y105_CO6),
.O5(CLBLM_R_X11Y108_SLICE_X15Y108_AO5),
.O6(CLBLM_R_X11Y108_SLICE_X15Y108_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hedffa5ed84a50084)
  ) CLBLM_R_X11Y109_SLICE_X14Y109_DLUT (
.I0(CLBLM_R_X11Y109_SLICE_X14Y109_AO5),
.I1(CLBLM_L_X10Y109_SLICE_X13Y109_BO6),
.I2(CLBLM_R_X11Y109_SLICE_X15Y109_AO6),
.I3(CLBLM_R_X11Y109_SLICE_X14Y109_CO6),
.I4(CLBLM_R_X11Y110_SLICE_X15Y110_AO6),
.I5(CLBLM_L_X10Y109_SLICE_X13Y109_AO6),
.O5(CLBLM_R_X11Y109_SLICE_X14Y109_DO5),
.O6(CLBLM_R_X11Y109_SLICE_X14Y109_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h69c3963c963c963c)
  ) CLBLM_R_X11Y109_SLICE_X14Y109_CLUT (
.I0(RIOB33_X105Y103_IOB_X1Y103_I),
.I1(CLBLM_R_X11Y108_SLICE_X15Y108_CO6),
.I2(CLBLM_R_X11Y106_SLICE_X14Y106_CO6),
.I3(LIOB33_X0Y107_IOB_X0Y107_I),
.I4(LIOB33_X0Y105_IOB_X0Y106_I),
.I5(RIOB33_X105Y103_IOB_X1Y104_I),
.O5(CLBLM_R_X11Y109_SLICE_X14Y109_CO5),
.O6(CLBLM_R_X11Y109_SLICE_X14Y109_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h788787781ee1e11e)
  ) CLBLM_R_X11Y109_SLICE_X14Y109_BLUT (
.I0(CLBLM_R_X11Y110_SLICE_X15Y110_AO6),
.I1(CLBLM_L_X10Y109_SLICE_X13Y109_BO6),
.I2(CLBLM_R_X11Y109_SLICE_X15Y109_AO6),
.I3(CLBLM_L_X10Y109_SLICE_X13Y109_AO6),
.I4(CLBLM_R_X11Y109_SLICE_X14Y109_AO5),
.I5(CLBLM_R_X11Y109_SLICE_X14Y109_CO6),
.O5(CLBLM_R_X11Y109_SLICE_X14Y109_BO5),
.O6(CLBLM_R_X11Y109_SLICE_X14Y109_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h33ff33ff0fff0fff)
  ) CLBLM_R_X11Y109_SLICE_X14Y109_ALUT (
.I0(1'b1),
.I1(LIOB33_X0Y105_IOB_X0Y106_I),
.I2(LIOB33_X0Y107_IOB_X0Y108_I),
.I3(RIOB33_X105Y103_IOB_X1Y103_I),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X11Y109_SLICE_X14Y109_AO5),
.O6(CLBLM_R_X11Y109_SLICE_X14Y109_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h371177377f55ff7f)
  ) CLBLM_R_X11Y109_SLICE_X15Y109_DLUT (
.I0(CLBLM_L_X12Y109_SLICE_X16Y109_BO6),
.I1(RIOB33_X105Y105_IOB_X1Y105_I),
.I2(LIOB33_X0Y105_IOB_X0Y106_I),
.I3(CLBLM_L_X12Y108_SLICE_X17Y108_DO6),
.I4(CLBLM_R_X11Y108_SLICE_X15Y108_DO6),
.I5(LIOB33_X0Y107_IOB_X0Y107_I),
.O5(CLBLM_R_X11Y109_SLICE_X15Y109_DO5),
.O6(CLBLM_R_X11Y109_SLICE_X15Y109_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h99a569aa69a566aa)
  ) CLBLM_R_X11Y109_SLICE_X15Y109_CLUT (
.I0(CLBLM_L_X12Y109_SLICE_X16Y109_BO6),
.I1(LIOB33_X0Y107_IOB_X0Y107_I),
.I2(CLBLM_L_X12Y108_SLICE_X17Y108_DO6),
.I3(RIOB33_X105Y105_IOB_X1Y105_I),
.I4(CLBLM_R_X11Y108_SLICE_X15Y108_DO6),
.I5(LIOB33_X0Y105_IOB_X0Y106_I),
.O5(CLBLM_R_X11Y109_SLICE_X15Y109_CO5),
.O6(CLBLM_R_X11Y109_SLICE_X15Y109_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h2bbbafff8eee0aaa)
  ) CLBLM_R_X11Y109_SLICE_X15Y109_BLUT (
.I0(CLBLM_R_X11Y106_SLICE_X14Y106_CO6),
.I1(RIOB33_X105Y103_IOB_X1Y104_I),
.I2(LIOB33_X0Y107_IOB_X0Y107_I),
.I3(RIOB33_X105Y103_IOB_X1Y103_I),
.I4(LIOB33_X0Y105_IOB_X0Y106_I),
.I5(CLBLM_R_X11Y108_SLICE_X15Y108_CO6),
.O5(CLBLM_R_X11Y109_SLICE_X15Y109_BO5),
.O6(CLBLM_R_X11Y109_SLICE_X15Y109_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h4bb4d22db44b2dd2)
  ) CLBLM_R_X11Y109_SLICE_X15Y109_ALUT (
.I0(CLBLM_R_X11Y106_SLICE_X14Y106_CO6),
.I1(CLBLM_R_X11Y108_SLICE_X15Y108_BO6),
.I2(CLBLM_R_X11Y108_SLICE_X15Y108_AO6),
.I3(CLBLM_R_X11Y107_SLICE_X15Y107_BO6),
.I4(CLBLM_L_X10Y108_SLICE_X13Y108_BO5),
.I5(CLBLM_R_X11Y111_SLICE_X15Y111_AO6),
.O5(CLBLM_R_X11Y109_SLICE_X15Y109_AO5),
.O6(CLBLM_R_X11Y109_SLICE_X15Y109_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hebeb82eb82eb8282)
  ) CLBLM_R_X11Y110_SLICE_X14Y110_DLUT (
.I0(CLBLM_R_X11Y110_SLICE_X14Y110_AO6),
.I1(CLBLM_R_X11Y110_SLICE_X15Y110_AO5),
.I2(CLBLM_R_X11Y110_SLICE_X15Y110_BO6),
.I3(CLBLM_R_X11Y111_SLICE_X15Y111_CO6),
.I4(CLBLM_R_X11Y109_SLICE_X14Y109_AO5),
.I5(CLBLM_R_X11Y109_SLICE_X15Y109_BO6),
.O5(CLBLM_R_X11Y110_SLICE_X14Y110_DO5),
.O6(CLBLM_R_X11Y110_SLICE_X14Y110_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hd22db4b44bb4b4b4)
  ) CLBLM_R_X11Y110_SLICE_X14Y110_CLUT (
.I0(CLBLM_R_X11Y109_SLICE_X15Y109_BO6),
.I1(CLBLM_R_X11Y111_SLICE_X15Y111_CO6),
.I2(CLBLM_R_X11Y110_SLICE_X15Y110_BO6),
.I3(RIOB33_X105Y103_IOB_X1Y104_I),
.I4(LIOB33_X0Y107_IOB_X0Y108_I),
.I5(RIOB33_X105Y103_IOB_X1Y103_I),
.O5(CLBLM_R_X11Y110_SLICE_X14Y110_CO5),
.O6(CLBLM_R_X11Y110_SLICE_X14Y110_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h69c3963c3c69c396)
  ) CLBLM_R_X11Y110_SLICE_X14Y110_BLUT (
.I0(CLBLM_R_X11Y109_SLICE_X14Y109_AO5),
.I1(CLBLM_R_X11Y110_SLICE_X15Y110_BO6),
.I2(CLBLM_R_X11Y110_SLICE_X15Y110_AO5),
.I3(CLBLM_R_X11Y109_SLICE_X15Y109_BO6),
.I4(CLBLM_R_X11Y110_SLICE_X14Y110_AO6),
.I5(CLBLM_R_X11Y111_SLICE_X15Y111_CO6),
.O5(CLBLM_R_X11Y110_SLICE_X14Y110_BO5),
.O6(CLBLM_R_X11Y110_SLICE_X14Y110_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0fff0fff00ffffff)
  ) CLBLM_R_X11Y110_SLICE_X14Y110_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(LIOB33_X0Y109_IOB_X0Y109_I),
.I3(RIOB33_X105Y103_IOB_X1Y103_I),
.I4(LIOB33_X0Y109_IOB_X0Y110_I),
.I5(1'b1),
.O5(CLBLM_R_X11Y110_SLICE_X14Y110_AO5),
.O6(CLBLM_R_X11Y110_SLICE_X14Y110_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h956aa956ff0033cc)
  ) CLBLM_R_X11Y110_SLICE_X15Y110_DLUT (
.I0(LIOB33_X0Y107_IOB_X0Y107_I),
.I1(CLBLM_L_X12Y109_SLICE_X16Y109_AO5),
.I2(LIOB33_X0Y105_IOB_X0Y106_I),
.I3(CLBLM_L_X12Y108_SLICE_X16Y108_CO6),
.I4(CLBLM_L_X12Y108_SLICE_X16Y108_DO6),
.I5(RIOB33_X105Y107_IOB_X1Y107_I),
.O5(CLBLM_R_X11Y110_SLICE_X15Y110_DO5),
.O6(CLBLM_R_X11Y110_SLICE_X15Y110_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h17ff053f5fff173f)
  ) CLBLM_R_X11Y110_SLICE_X15Y110_CLUT (
.I0(LIOB33_X0Y107_IOB_X0Y107_I),
.I1(CLBLM_L_X12Y109_SLICE_X16Y109_AO5),
.I2(CLBLM_L_X12Y108_SLICE_X16Y108_CO6),
.I3(RIOB33_X105Y107_IOB_X1Y107_I),
.I4(CLBLM_L_X12Y108_SLICE_X16Y108_DO6),
.I5(LIOB33_X0Y105_IOB_X0Y106_I),
.O5(CLBLM_R_X11Y110_SLICE_X15Y110_CO5),
.O6(CLBLM_R_X11Y110_SLICE_X15Y110_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h6a5695a995a96a56)
  ) CLBLM_R_X11Y110_SLICE_X15Y110_BLUT (
.I0(CLBLM_R_X11Y111_SLICE_X15Y111_BO5),
.I1(CLBLM_R_X11Y111_SLICE_X15Y111_AO6),
.I2(CLBLM_R_X11Y108_SLICE_X15Y108_AO6),
.I3(CLBLM_R_X11Y107_SLICE_X15Y107_BO6),
.I4(CLBLM_R_X11Y107_SLICE_X15Y107_CO6),
.I5(CLBLM_L_X12Y109_SLICE_X16Y109_BO6),
.O5(CLBLM_R_X11Y110_SLICE_X15Y110_BO5),
.O6(CLBLM_R_X11Y110_SLICE_X15Y110_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0fff0fff00ffffff)
  ) CLBLM_R_X11Y110_SLICE_X15Y110_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(RIOB33_X105Y101_IOB_X1Y102_I),
.I3(LIOB33_X0Y107_IOB_X0Y108_I),
.I4(RIOB33_X105Y103_IOB_X1Y104_I),
.I5(1'b1),
.O5(CLBLM_R_X11Y110_SLICE_X15Y110_AO5),
.O6(CLBLM_R_X11Y110_SLICE_X15Y110_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h71f3d4fcd4fcd4fc)
  ) CLBLM_R_X11Y111_SLICE_X14Y111_DLUT (
.I0(LIOB33_X0Y107_IOB_X0Y108_I),
.I1(CLBLM_L_X12Y109_SLICE_X16Y109_CO6),
.I2(CLBLM_R_X11Y111_SLICE_X15Y111_DO6),
.I3(RIOB33_X105Y103_IOB_X1Y104_I),
.I4(LIOB33_X0Y107_IOB_X0Y107_I),
.I5(RIOB33_X105Y105_IOB_X1Y105_I),
.O5(CLBLM_R_X11Y111_SLICE_X14Y111_DO5),
.O6(CLBLM_R_X11Y111_SLICE_X14Y111_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h69c3963c963c963c)
  ) CLBLM_R_X11Y111_SLICE_X14Y111_CLUT (
.I0(LIOB33_X0Y107_IOB_X0Y108_I),
.I1(CLBLM_L_X12Y109_SLICE_X16Y109_CO6),
.I2(CLBLM_R_X11Y111_SLICE_X15Y111_DO6),
.I3(RIOB33_X105Y103_IOB_X1Y104_I),
.I4(LIOB33_X0Y107_IOB_X0Y107_I),
.I5(RIOB33_X105Y105_IOB_X1Y105_I),
.O5(CLBLM_R_X11Y111_SLICE_X14Y111_CO5),
.O6(CLBLM_R_X11Y111_SLICE_X14Y111_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h22bbaaff6699aa55)
  ) CLBLM_R_X11Y111_SLICE_X14Y111_BLUT (
.I0(CLBLM_R_X11Y109_SLICE_X15Y109_DO6),
.I1(LIOB33_X0Y107_IOB_X0Y108_I),
.I2(1'b1),
.I3(CLBLM_R_X11Y110_SLICE_X15Y110_DO6),
.I4(RIOB33_X105Y105_IOB_X1Y105_I),
.I5(1'b1),
.O5(CLBLM_R_X11Y111_SLICE_X14Y111_BO5),
.O6(CLBLM_R_X11Y111_SLICE_X14Y111_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0fff0fff2bbb2bbb)
  ) CLBLM_R_X11Y111_SLICE_X14Y111_ALUT (
.I0(CLBLM_R_X11Y111_SLICE_X14Y111_DO6),
.I1(CLBLM_R_X11Y111_SLICE_X14Y111_BO5),
.I2(LIOB33_X0Y109_IOB_X0Y109_I),
.I3(RIOB33_X105Y103_IOB_X1Y104_I),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X11Y111_SLICE_X14Y111_AO5),
.O6(CLBLM_R_X11Y111_SLICE_X14Y111_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h28bebebe88eeeeee)
  ) CLBLM_R_X11Y111_SLICE_X15Y111_DLUT (
.I0(CLBLM_R_X11Y108_SLICE_X15Y108_AO6),
.I1(CLBLM_L_X12Y108_SLICE_X17Y108_AO6),
.I2(LIOB33_X0Y105_IOB_X0Y106_I),
.I3(RIOB33_X105Y103_IOB_X1Y104_I),
.I4(LIOB33_X0Y107_IOB_X0Y107_I),
.I5(RIOB33_X105Y105_IOB_X1Y105_I),
.O5(CLBLM_R_X11Y111_SLICE_X15Y111_DO5),
.O6(CLBLM_R_X11Y111_SLICE_X15Y111_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h6996a55a996655aa)
  ) CLBLM_R_X11Y111_SLICE_X15Y111_CLUT (
.I0(CLBLM_R_X11Y108_SLICE_X15Y108_AO6),
.I1(RIOB33_X105Y103_IOB_X1Y104_I),
.I2(LIOB33_X0Y105_IOB_X0Y106_I),
.I3(CLBLM_L_X12Y108_SLICE_X17Y108_AO6),
.I4(LIOB33_X0Y107_IOB_X0Y107_I),
.I5(RIOB33_X105Y105_IOB_X1Y105_I),
.O5(CLBLM_R_X11Y111_SLICE_X15Y111_CO5),
.O6(CLBLM_R_X11Y111_SLICE_X15Y111_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h55ff55ff0fff0fff)
  ) CLBLM_R_X11Y111_SLICE_X15Y111_BLUT (
.I0(LIOB33_X0Y105_IOB_X0Y106_I),
.I1(1'b1),
.I2(LIOB33_X0Y107_IOB_X0Y107_I),
.I3(RIOB33_X105Y105_IOB_X1Y105_I),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X11Y111_SLICE_X15Y111_BO5),
.O6(CLBLM_R_X11Y111_SLICE_X15Y111_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h3333ffff77777777)
  ) CLBLM_R_X11Y111_SLICE_X15Y111_ALUT (
.I0(LIOB33_X0Y105_IOB_X0Y106_I),
.I1(RIOB33_X105Y103_IOB_X1Y104_I),
.I2(1'b1),
.I3(1'b1),
.I4(LIOB33_X0Y107_IOB_X0Y107_I),
.I5(1'b1),
.O5(CLBLM_R_X11Y111_SLICE_X15Y111_AO5),
.O6(CLBLM_R_X11Y111_SLICE_X15Y111_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X13Y105_SLICE_X18Y105_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X13Y105_SLICE_X18Y105_DO5),
.O6(CLBLM_R_X13Y105_SLICE_X18Y105_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X13Y105_SLICE_X18Y105_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X13Y105_SLICE_X18Y105_CO5),
.O6(CLBLM_R_X13Y105_SLICE_X18Y105_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X13Y105_SLICE_X18Y105_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X13Y105_SLICE_X18Y105_BO5),
.O6(CLBLM_R_X13Y105_SLICE_X18Y105_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hccf3a6f3a53fa53f)
  ) CLBLM_R_X13Y105_SLICE_X18Y105_ALUT (
.I0(RIOB33_X105Y111_IOB_X1Y111_I),
.I1(LIOB33_SING_X0Y100_IOB_X0Y100_I),
.I2(RIOB33_X105Y109_IOB_X1Y109_I),
.I3(RIOB33_X105Y113_IOB_X1Y113_I),
.I4(RIOB33_X105Y111_IOB_X1Y112_I),
.I5(RIOB33_X105Y109_IOB_X1Y110_I),
.O5(CLBLM_R_X13Y105_SLICE_X18Y105_AO5),
.O6(CLBLM_R_X13Y105_SLICE_X18Y105_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X13Y105_SLICE_X19Y105_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X13Y105_SLICE_X19Y105_DO5),
.O6(CLBLM_R_X13Y105_SLICE_X19Y105_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X13Y105_SLICE_X19Y105_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X13Y105_SLICE_X19Y105_CO5),
.O6(CLBLM_R_X13Y105_SLICE_X19Y105_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X13Y105_SLICE_X19Y105_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X13Y105_SLICE_X19Y105_BO5),
.O6(CLBLM_R_X13Y105_SLICE_X19Y105_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X13Y105_SLICE_X19Y105_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X13Y105_SLICE_X19Y105_AO5),
.O6(CLBLM_R_X13Y105_SLICE_X19Y105_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h5aa6a5a659a6a6a6)
  ) CLBLM_R_X13Y106_SLICE_X18Y106_DLUT (
.I0(CLBLM_R_X13Y105_SLICE_X18Y105_AO6),
.I1(CLBLM_R_X13Y106_SLICE_X19Y106_CO6),
.I2(CLBLM_R_X13Y106_SLICE_X19Y106_BO6),
.I3(LIOB33_X0Y101_IOB_X0Y101_I),
.I4(RIOB33_X105Y109_IOB_X1Y109_I),
.I5(RIOB33_X105Y107_IOB_X1Y108_I),
.O5(CLBLM_R_X13Y106_SLICE_X18Y106_DO5),
.O6(CLBLM_R_X13Y106_SLICE_X18Y106_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h59a6a6595aa5a55a)
  ) CLBLM_R_X13Y106_SLICE_X18Y106_CLUT (
.I0(CLBLM_R_X13Y105_SLICE_X18Y105_AO6),
.I1(CLBLM_R_X13Y106_SLICE_X19Y106_CO6),
.I2(CLBLM_R_X13Y106_SLICE_X19Y106_BO6),
.I3(CLBLM_R_X11Y106_SLICE_X15Y106_AO6),
.I4(CLBLM_L_X12Y107_SLICE_X17Y107_AO6),
.I5(CLBLM_L_X12Y106_SLICE_X16Y106_AO6),
.O5(CLBLM_R_X13Y106_SLICE_X18Y106_CO5),
.O6(CLBLM_R_X13Y106_SLICE_X18Y106_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hef8a8aefee8888ee)
  ) CLBLM_R_X13Y106_SLICE_X18Y106_BLUT (
.I0(CLBLM_L_X12Y107_SLICE_X17Y107_AO6),
.I1(CLBLM_R_X13Y106_SLICE_X19Y106_BO6),
.I2(CLBLM_R_X13Y106_SLICE_X19Y106_CO6),
.I3(CLBLM_R_X11Y106_SLICE_X15Y106_AO6),
.I4(CLBLM_R_X13Y105_SLICE_X18Y105_AO6),
.I5(CLBLM_L_X12Y106_SLICE_X16Y106_AO6),
.O5(CLBLM_R_X13Y106_SLICE_X18Y106_BO5),
.O6(CLBLM_R_X13Y106_SLICE_X18Y106_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hc30fc30f3333ffff)
  ) CLBLM_R_X13Y106_SLICE_X18Y106_ALUT (
.I0(1'b1),
.I1(LIOB33_X0Y101_IOB_X0Y101_I),
.I2(CLBLM_R_X13Y105_SLICE_X18Y105_AO6),
.I3(RIOB33_X105Y109_IOB_X1Y109_I),
.I4(RIOB33_X105Y105_IOB_X1Y106_I),
.I5(1'b1),
.O5(CLBLM_R_X13Y106_SLICE_X18Y106_AO5),
.O6(CLBLM_R_X13Y106_SLICE_X18Y106_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X13Y106_SLICE_X19Y106_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X13Y106_SLICE_X19Y106_DO5),
.O6(CLBLM_R_X13Y106_SLICE_X19Y106_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h13a33c004cfc3c00)
  ) CLBLM_R_X13Y106_SLICE_X19Y106_CLUT (
.I0(RIOB33_X105Y111_IOB_X1Y112_I),
.I1(RIOB33_X105Y107_IOB_X1Y108_I),
.I2(RIOB33_X105Y109_IOB_X1Y109_I),
.I3(LIOB33_SING_X0Y100_IOB_X0Y100_I),
.I4(RIOB33_X105Y113_IOB_X1Y113_I),
.I5(RIOB33_X105Y109_IOB_X1Y110_I),
.O5(CLBLM_R_X13Y106_SLICE_X19Y106_CO5),
.O6(CLBLM_R_X13Y106_SLICE_X19Y106_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h13220022b100aa00)
  ) CLBLM_R_X13Y106_SLICE_X19Y106_BLUT (
.I0(RIOB33_X105Y109_IOB_X1Y109_I),
.I1(RIOB33_X105Y107_IOB_X1Y108_I),
.I2(RIOB33_X105Y111_IOB_X1Y112_I),
.I3(RIOB33_X105Y113_IOB_X1Y113_I),
.I4(RIOB33_X105Y109_IOB_X1Y110_I),
.I5(LIOB33_SING_X0Y100_IOB_X0Y100_I),
.O5(CLBLM_R_X13Y106_SLICE_X19Y106_BO5),
.O6(CLBLM_R_X13Y106_SLICE_X19Y106_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hcc0033ffaaaabbff)
  ) CLBLM_R_X13Y106_SLICE_X19Y106_ALUT (
.I0(CLBLM_R_X13Y106_SLICE_X19Y106_BO6),
.I1(RIOB33_X105Y107_IOB_X1Y108_I),
.I2(1'b1),
.I3(LIOB33_X0Y101_IOB_X0Y101_I),
.I4(CLBLM_R_X13Y106_SLICE_X19Y106_CO6),
.I5(1'b1),
.O5(CLBLM_R_X13Y106_SLICE_X19Y106_AO5),
.O6(CLBLM_R_X13Y106_SLICE_X19Y106_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X13Y107_SLICE_X18Y107_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X13Y107_SLICE_X18Y107_DO5),
.O6(CLBLM_R_X13Y107_SLICE_X18Y107_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X13Y107_SLICE_X18Y107_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X13Y107_SLICE_X18Y107_CO5),
.O6(CLBLM_R_X13Y107_SLICE_X18Y107_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X13Y107_SLICE_X18Y107_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X13Y107_SLICE_X18Y107_BO5),
.O6(CLBLM_R_X13Y107_SLICE_X18Y107_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h6999966696669666)
  ) CLBLM_R_X13Y107_SLICE_X18Y107_ALUT (
.I0(CLBLM_R_X13Y106_SLICE_X18Y106_DO6),
.I1(CLBLM_L_X12Y106_SLICE_X17Y106_DO6),
.I2(LIOB33_X0Y101_IOB_X0Y102_I),
.I3(RIOB33_X105Y107_IOB_X1Y108_I),
.I4(RIOB33_X105Y107_IOB_X1Y107_I),
.I5(LIOB33_X0Y103_IOB_X0Y104_I),
.O5(CLBLM_R_X13Y107_SLICE_X18Y107_AO5),
.O6(CLBLM_R_X13Y107_SLICE_X18Y107_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X13Y107_SLICE_X19Y107_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X13Y107_SLICE_X19Y107_DO5),
.O6(CLBLM_R_X13Y107_SLICE_X19Y107_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X13Y107_SLICE_X19Y107_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X13Y107_SLICE_X19Y107_CO5),
.O6(CLBLM_R_X13Y107_SLICE_X19Y107_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X13Y107_SLICE_X19Y107_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X13Y107_SLICE_X19Y107_BO5),
.O6(CLBLM_R_X13Y107_SLICE_X19Y107_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X13Y107_SLICE_X19Y107_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X13Y107_SLICE_X19Y107_AO5),
.O6(CLBLM_R_X13Y107_SLICE_X19Y107_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y101_IOB_X0Y101_IBUF (
.I(LIOB33_X0Y101_IOB_X0Y101_IPAD),
.O(LIOB33_X0Y101_IOB_X0Y101_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y101_IOB_X0Y102_IBUF (
.I(LIOB33_X0Y101_IOB_X0Y102_IPAD),
.O(LIOB33_X0Y101_IOB_X0Y102_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y103_IOB_X0Y103_IBUF (
.I(LIOB33_X0Y103_IOB_X0Y103_IPAD),
.O(LIOB33_X0Y103_IOB_X0Y103_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y103_IOB_X0Y104_IBUF (
.I(LIOB33_X0Y103_IOB_X0Y104_IPAD),
.O(LIOB33_X0Y103_IOB_X0Y104_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y105_IOB_X0Y105_IBUF (
.I(LIOB33_X0Y105_IOB_X0Y105_IPAD),
.O(LIOB33_X0Y105_IOB_X0Y105_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y105_IOB_X0Y106_IBUF (
.I(LIOB33_X0Y105_IOB_X0Y106_IPAD),
.O(LIOB33_X0Y105_IOB_X0Y106_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y107_IOB_X0Y107_IBUF (
.I(LIOB33_X0Y107_IOB_X0Y107_IPAD),
.O(LIOB33_X0Y107_IOB_X0Y107_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y107_IOB_X0Y108_IBUF (
.I(LIOB33_X0Y107_IOB_X0Y108_IPAD),
.O(LIOB33_X0Y107_IOB_X0Y108_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y109_IOB_X0Y109_IBUF (
.I(LIOB33_X0Y109_IOB_X0Y109_IPAD),
.O(LIOB33_X0Y109_IOB_X0Y109_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y109_IOB_X0Y110_IBUF (
.I(LIOB33_X0Y109_IOB_X0Y110_IPAD),
.O(LIOB33_X0Y109_IOB_X0Y110_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y111_IOB_X0Y111_IBUF (
.I(LIOB33_X0Y111_IOB_X0Y111_IPAD),
.O(LIOB33_X0Y111_IOB_X0Y111_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y111_IOB_X0Y112_IBUF (
.I(LIOB33_X0Y111_IOB_X0Y112_IPAD),
.O(LIOB33_X0Y111_IOB_X0Y112_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y113_IOB_X0Y113_IBUF (
.I(LIOB33_X0Y113_IOB_X0Y113_IPAD),
.O(LIOB33_X0Y113_IOB_X0Y113_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y113_IOB_X0Y114_IBUF (
.I(LIOB33_X0Y113_IOB_X0Y114_IPAD),
.O(LIOB33_X0Y113_IOB_X0Y114_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y115_IOB_X0Y115_IBUF (
.I(LIOB33_X0Y115_IOB_X0Y115_IPAD),
.O(LIOB33_X0Y115_IOB_X0Y115_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y115_IOB_X0Y116_IBUF (
.I(LIOB33_X0Y115_IOB_X0Y116_IPAD),
.O(LIOB33_X0Y115_IOB_X0Y116_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y117_IOB_X0Y117_IBUF (
.I(LIOB33_X0Y117_IOB_X0Y117_IPAD),
.O(LIOB33_X0Y117_IOB_X0Y117_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y117_IOB_X0Y118_OBUF (
.I(CLBLL_L_X2Y109_SLICE_X0Y109_AO5),
.O(LIOB33_X0Y117_IOB_X0Y118_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y119_IOB_X0Y119_OBUF (
.I(CLBLL_L_X2Y109_SLICE_X0Y109_AO6),
.O(LIOB33_X0Y119_IOB_X0Y119_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y119_IOB_X0Y120_OBUF (
.I(CLBLM_R_X3Y106_SLICE_X2Y106_AO5),
.O(LIOB33_X0Y119_IOB_X0Y120_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y121_IOB_X0Y121_OBUF (
.I(CLBLL_L_X2Y106_SLICE_X0Y106_AO5),
.O(LIOB33_X0Y121_IOB_X0Y121_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y121_IOB_X0Y122_OBUF (
.I(CLBLL_L_X2Y104_SLICE_X0Y104_AO6),
.O(LIOB33_X0Y121_IOB_X0Y122_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y123_IOB_X0Y123_OBUF (
.I(CLBLL_L_X2Y107_SLICE_X0Y107_AO6),
.O(LIOB33_X0Y123_IOB_X0Y123_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y123_IOB_X0Y124_OBUF (
.I(CLBLM_R_X3Y107_SLICE_X2Y107_AO6),
.O(LIOB33_X0Y123_IOB_X0Y124_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y125_IOB_X0Y125_OBUF (
.I(CLBLM_R_X7Y109_SLICE_X9Y109_AO5),
.O(LIOB33_X0Y125_IOB_X0Y125_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y125_IOB_X0Y126_OBUF (
.I(CLBLM_R_X3Y107_SLICE_X2Y107_CO6),
.O(LIOB33_X0Y125_IOB_X0Y126_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y127_IOB_X0Y127_OBUF (
.I(CLBLM_R_X3Y107_SLICE_X3Y107_AO6),
.O(LIOB33_X0Y127_IOB_X0Y127_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y127_IOB_X0Y128_OBUF (
.I(CLBLM_R_X3Y107_SLICE_X3Y107_BO6),
.O(LIOB33_X0Y127_IOB_X0Y128_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y129_IOB_X0Y129_OBUF (
.I(CLBLM_R_X3Y108_SLICE_X3Y108_AO6),
.O(LIOB33_X0Y129_IOB_X0Y129_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y129_IOB_X0Y130_OBUF (
.I(CLBLL_L_X2Y110_SLICE_X0Y110_AO6),
.O(LIOB33_X0Y129_IOB_X0Y130_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y131_IOB_X0Y131_OBUF (
.I(CLBLL_L_X4Y108_SLICE_X4Y108_AO6),
.O(LIOB33_X0Y131_IOB_X0Y131_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y131_IOB_X0Y132_OBUF (
.I(CLBLL_L_X2Y110_SLICE_X0Y110_AO5),
.O(LIOB33_X0Y131_IOB_X0Y132_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y133_IOB_X0Y133_OBUF (
.I(CLBLM_R_X3Y109_SLICE_X3Y109_AO6),
.O(LIOB33_X0Y133_IOB_X0Y133_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y133_IOB_X0Y134_OBUF (
.I(1'b0),
.O(LIOB33_X0Y133_IOB_X0Y134_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y135_IOB_X0Y135_OBUF (
.I(CLBLL_L_X4Y110_SLICE_X5Y110_AO6),
.O(LIOB33_X0Y135_IOB_X0Y135_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y135_IOB_X0Y136_OBUF (
.I(CLBLL_L_X4Y110_SLICE_X5Y110_AO5),
.O(LIOB33_X0Y135_IOB_X0Y136_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y137_IOB_X0Y137_OBUF (
.I(CLBLL_L_X4Y111_SLICE_X4Y111_AO6),
.O(LIOB33_X0Y137_IOB_X0Y137_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y137_IOB_X0Y138_OBUF (
.I(CLBLL_L_X4Y111_SLICE_X4Y111_AO5),
.O(LIOB33_X0Y137_IOB_X0Y138_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y139_IOB_X0Y139_OBUF (
.I(CLBLL_L_X4Y112_SLICE_X4Y112_AO6),
.O(LIOB33_X0Y139_IOB_X0Y139_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y139_IOB_X0Y140_OBUF (
.I(CLBLL_L_X4Y112_SLICE_X4Y112_AO5),
.O(LIOB33_X0Y139_IOB_X0Y140_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y141_IOB_X0Y141_OBUF (
.I(CLBLL_L_X4Y112_SLICE_X5Y112_DO6),
.O(LIOB33_X0Y141_IOB_X0Y141_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y141_IOB_X0Y142_OBUF (
.I(CLBLL_L_X4Y114_SLICE_X4Y114_DO6),
.O(LIOB33_X0Y141_IOB_X0Y142_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y143_IOB_X0Y143_OBUF (
.I(CLBLL_L_X4Y115_SLICE_X4Y115_DO6),
.O(LIOB33_X0Y143_IOB_X0Y143_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y145_IOB_X0Y145_OBUF (
.I(CLBLL_L_X4Y115_SLICE_X4Y115_AO5),
.O(LIOB33_X0Y145_IOB_X0Y145_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y145_IOB_X0Y146_OBUF (
.I(CLBLL_L_X4Y115_SLICE_X4Y115_CO6),
.O(LIOB33_X0Y145_IOB_X0Y146_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y147_IOB_X0Y147_OBUF (
.I(CLBLM_R_X3Y112_SLICE_X2Y112_AO5),
.O(LIOB33_X0Y147_IOB_X0Y147_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y147_IOB_X0Y148_OBUF (
.I(CLBLM_R_X3Y112_SLICE_X2Y112_CO6),
.O(LIOB33_X0Y147_IOB_X0Y148_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_SING_X0Y100_IOB_X0Y100_IBUF (
.I(LIOB33_SING_X0Y100_IOB_X0Y100_IPAD),
.O(LIOB33_SING_X0Y100_IOB_X0Y100_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_SING_X0Y149_IOB_X0Y149_OBUF (
.I(CLBLM_R_X3Y112_SLICE_X2Y112_DO6),
.O(LIOB33_SING_X0Y149_IOB_X0Y149_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y101_IOB_X1Y101_IBUF (
.I(RIOB33_X105Y101_IOB_X1Y101_IPAD),
.O(RIOB33_X105Y101_IOB_X1Y101_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y101_IOB_X1Y102_IBUF (
.I(RIOB33_X105Y101_IOB_X1Y102_IPAD),
.O(RIOB33_X105Y101_IOB_X1Y102_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y103_IOB_X1Y103_IBUF (
.I(RIOB33_X105Y103_IOB_X1Y103_IPAD),
.O(RIOB33_X105Y103_IOB_X1Y103_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y103_IOB_X1Y104_IBUF (
.I(RIOB33_X105Y103_IOB_X1Y104_IPAD),
.O(RIOB33_X105Y103_IOB_X1Y104_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y105_IOB_X1Y105_IBUF (
.I(RIOB33_X105Y105_IOB_X1Y105_IPAD),
.O(RIOB33_X105Y105_IOB_X1Y105_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y105_IOB_X1Y106_IBUF (
.I(RIOB33_X105Y105_IOB_X1Y106_IPAD),
.O(RIOB33_X105Y105_IOB_X1Y106_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y107_IOB_X1Y107_IBUF (
.I(RIOB33_X105Y107_IOB_X1Y107_IPAD),
.O(RIOB33_X105Y107_IOB_X1Y107_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y107_IOB_X1Y108_IBUF (
.I(RIOB33_X105Y107_IOB_X1Y108_IPAD),
.O(RIOB33_X105Y107_IOB_X1Y108_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y109_IOB_X1Y109_IBUF (
.I(RIOB33_X105Y109_IOB_X1Y109_IPAD),
.O(RIOB33_X105Y109_IOB_X1Y109_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y109_IOB_X1Y110_IBUF (
.I(RIOB33_X105Y109_IOB_X1Y110_IPAD),
.O(RIOB33_X105Y109_IOB_X1Y110_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y111_IOB_X1Y111_IBUF (
.I(RIOB33_X105Y111_IOB_X1Y111_IPAD),
.O(RIOB33_X105Y111_IOB_X1Y111_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y111_IOB_X1Y112_IBUF (
.I(RIOB33_X105Y111_IOB_X1Y112_IPAD),
.O(RIOB33_X105Y111_IOB_X1Y112_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y113_IOB_X1Y113_IBUF (
.I(RIOB33_X105Y113_IOB_X1Y113_IPAD),
.O(RIOB33_X105Y113_IOB_X1Y113_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_SING_X105Y100_IOB_X1Y100_IBUF (
.I(RIOB33_SING_X105Y100_IOB_X1Y100_IPAD),
.O(RIOB33_SING_X105Y100_IOB_X1Y100_I)
  );
  assign CLBLL_L_X2Y104_SLICE_X0Y104_A = CLBLL_L_X2Y104_SLICE_X0Y104_AO6;
  assign CLBLL_L_X2Y104_SLICE_X0Y104_B = CLBLL_L_X2Y104_SLICE_X0Y104_BO6;
  assign CLBLL_L_X2Y104_SLICE_X0Y104_C = CLBLL_L_X2Y104_SLICE_X0Y104_CO6;
  assign CLBLL_L_X2Y104_SLICE_X0Y104_D = CLBLL_L_X2Y104_SLICE_X0Y104_DO6;
  assign CLBLL_L_X2Y104_SLICE_X0Y104_AMUX = CLBLL_L_X2Y104_SLICE_X0Y104_AO5;
  assign CLBLL_L_X2Y104_SLICE_X0Y104_BMUX = CLBLL_L_X2Y104_SLICE_X0Y104_BO6;
  assign CLBLL_L_X2Y104_SLICE_X0Y104_CMUX = CLBLL_L_X2Y104_SLICE_X0Y104_CO6;
  assign CLBLL_L_X2Y104_SLICE_X1Y104_A = CLBLL_L_X2Y104_SLICE_X1Y104_AO6;
  assign CLBLL_L_X2Y104_SLICE_X1Y104_B = CLBLL_L_X2Y104_SLICE_X1Y104_BO6;
  assign CLBLL_L_X2Y104_SLICE_X1Y104_C = CLBLL_L_X2Y104_SLICE_X1Y104_CO6;
  assign CLBLL_L_X2Y104_SLICE_X1Y104_D = CLBLL_L_X2Y104_SLICE_X1Y104_DO6;
  assign CLBLL_L_X2Y104_SLICE_X1Y104_AMUX = CLBLL_L_X2Y104_SLICE_X1Y104_AO5;
  assign CLBLL_L_X2Y106_SLICE_X0Y106_A = CLBLL_L_X2Y106_SLICE_X0Y106_AO6;
  assign CLBLL_L_X2Y106_SLICE_X0Y106_B = CLBLL_L_X2Y106_SLICE_X0Y106_BO6;
  assign CLBLL_L_X2Y106_SLICE_X0Y106_C = CLBLL_L_X2Y106_SLICE_X0Y106_CO6;
  assign CLBLL_L_X2Y106_SLICE_X0Y106_D = CLBLL_L_X2Y106_SLICE_X0Y106_DO6;
  assign CLBLL_L_X2Y106_SLICE_X0Y106_AMUX = CLBLL_L_X2Y106_SLICE_X0Y106_AO5;
  assign CLBLL_L_X2Y106_SLICE_X1Y106_A = CLBLL_L_X2Y106_SLICE_X1Y106_AO6;
  assign CLBLL_L_X2Y106_SLICE_X1Y106_B = CLBLL_L_X2Y106_SLICE_X1Y106_BO6;
  assign CLBLL_L_X2Y106_SLICE_X1Y106_C = CLBLL_L_X2Y106_SLICE_X1Y106_CO6;
  assign CLBLL_L_X2Y106_SLICE_X1Y106_D = CLBLL_L_X2Y106_SLICE_X1Y106_DO6;
  assign CLBLL_L_X2Y106_SLICE_X1Y106_AMUX = CLBLL_L_X2Y106_SLICE_X1Y106_AO5;
  assign CLBLL_L_X2Y106_SLICE_X1Y106_CMUX = CLBLL_L_X2Y106_SLICE_X1Y106_CO6;
  assign CLBLL_L_X2Y107_SLICE_X0Y107_A = CLBLL_L_X2Y107_SLICE_X0Y107_AO6;
  assign CLBLL_L_X2Y107_SLICE_X0Y107_B = CLBLL_L_X2Y107_SLICE_X0Y107_BO6;
  assign CLBLL_L_X2Y107_SLICE_X0Y107_C = CLBLL_L_X2Y107_SLICE_X0Y107_CO6;
  assign CLBLL_L_X2Y107_SLICE_X0Y107_D = CLBLL_L_X2Y107_SLICE_X0Y107_DO6;
  assign CLBLL_L_X2Y107_SLICE_X1Y107_A = CLBLL_L_X2Y107_SLICE_X1Y107_AO6;
  assign CLBLL_L_X2Y107_SLICE_X1Y107_B = CLBLL_L_X2Y107_SLICE_X1Y107_BO6;
  assign CLBLL_L_X2Y107_SLICE_X1Y107_C = CLBLL_L_X2Y107_SLICE_X1Y107_CO6;
  assign CLBLL_L_X2Y107_SLICE_X1Y107_D = CLBLL_L_X2Y107_SLICE_X1Y107_DO6;
  assign CLBLL_L_X2Y109_SLICE_X0Y109_A = CLBLL_L_X2Y109_SLICE_X0Y109_AO6;
  assign CLBLL_L_X2Y109_SLICE_X0Y109_B = CLBLL_L_X2Y109_SLICE_X0Y109_BO6;
  assign CLBLL_L_X2Y109_SLICE_X0Y109_C = CLBLL_L_X2Y109_SLICE_X0Y109_CO6;
  assign CLBLL_L_X2Y109_SLICE_X0Y109_D = CLBLL_L_X2Y109_SLICE_X0Y109_DO6;
  assign CLBLL_L_X2Y109_SLICE_X0Y109_AMUX = CLBLL_L_X2Y109_SLICE_X0Y109_AO5;
  assign CLBLL_L_X2Y109_SLICE_X1Y109_A = CLBLL_L_X2Y109_SLICE_X1Y109_AO6;
  assign CLBLL_L_X2Y109_SLICE_X1Y109_B = CLBLL_L_X2Y109_SLICE_X1Y109_BO6;
  assign CLBLL_L_X2Y109_SLICE_X1Y109_C = CLBLL_L_X2Y109_SLICE_X1Y109_CO6;
  assign CLBLL_L_X2Y109_SLICE_X1Y109_D = CLBLL_L_X2Y109_SLICE_X1Y109_DO6;
  assign CLBLL_L_X2Y110_SLICE_X0Y110_A = CLBLL_L_X2Y110_SLICE_X0Y110_AO6;
  assign CLBLL_L_X2Y110_SLICE_X0Y110_B = CLBLL_L_X2Y110_SLICE_X0Y110_BO6;
  assign CLBLL_L_X2Y110_SLICE_X0Y110_C = CLBLL_L_X2Y110_SLICE_X0Y110_CO6;
  assign CLBLL_L_X2Y110_SLICE_X0Y110_D = CLBLL_L_X2Y110_SLICE_X0Y110_DO6;
  assign CLBLL_L_X2Y110_SLICE_X0Y110_AMUX = CLBLL_L_X2Y110_SLICE_X0Y110_AO5;
  assign CLBLL_L_X2Y110_SLICE_X1Y110_A = CLBLL_L_X2Y110_SLICE_X1Y110_AO6;
  assign CLBLL_L_X2Y110_SLICE_X1Y110_B = CLBLL_L_X2Y110_SLICE_X1Y110_BO6;
  assign CLBLL_L_X2Y110_SLICE_X1Y110_C = CLBLL_L_X2Y110_SLICE_X1Y110_CO6;
  assign CLBLL_L_X2Y110_SLICE_X1Y110_D = CLBLL_L_X2Y110_SLICE_X1Y110_DO6;
  assign CLBLL_L_X4Y103_SLICE_X4Y103_A = CLBLL_L_X4Y103_SLICE_X4Y103_AO6;
  assign CLBLL_L_X4Y103_SLICE_X4Y103_B = CLBLL_L_X4Y103_SLICE_X4Y103_BO6;
  assign CLBLL_L_X4Y103_SLICE_X4Y103_C = CLBLL_L_X4Y103_SLICE_X4Y103_CO6;
  assign CLBLL_L_X4Y103_SLICE_X4Y103_D = CLBLL_L_X4Y103_SLICE_X4Y103_DO6;
  assign CLBLL_L_X4Y103_SLICE_X4Y103_AMUX = CLBLL_L_X4Y103_SLICE_X4Y103_AO5;
  assign CLBLL_L_X4Y103_SLICE_X5Y103_A = CLBLL_L_X4Y103_SLICE_X5Y103_AO6;
  assign CLBLL_L_X4Y103_SLICE_X5Y103_B = CLBLL_L_X4Y103_SLICE_X5Y103_BO6;
  assign CLBLL_L_X4Y103_SLICE_X5Y103_C = CLBLL_L_X4Y103_SLICE_X5Y103_CO6;
  assign CLBLL_L_X4Y103_SLICE_X5Y103_D = CLBLL_L_X4Y103_SLICE_X5Y103_DO6;
  assign CLBLL_L_X4Y103_SLICE_X5Y103_AMUX = CLBLL_L_X4Y103_SLICE_X5Y103_AO5;
  assign CLBLL_L_X4Y104_SLICE_X4Y104_A = CLBLL_L_X4Y104_SLICE_X4Y104_AO6;
  assign CLBLL_L_X4Y104_SLICE_X4Y104_B = CLBLL_L_X4Y104_SLICE_X4Y104_BO6;
  assign CLBLL_L_X4Y104_SLICE_X4Y104_C = CLBLL_L_X4Y104_SLICE_X4Y104_CO6;
  assign CLBLL_L_X4Y104_SLICE_X4Y104_D = CLBLL_L_X4Y104_SLICE_X4Y104_DO6;
  assign CLBLL_L_X4Y104_SLICE_X5Y104_A = CLBLL_L_X4Y104_SLICE_X5Y104_AO6;
  assign CLBLL_L_X4Y104_SLICE_X5Y104_B = CLBLL_L_X4Y104_SLICE_X5Y104_BO6;
  assign CLBLL_L_X4Y104_SLICE_X5Y104_C = CLBLL_L_X4Y104_SLICE_X5Y104_CO6;
  assign CLBLL_L_X4Y104_SLICE_X5Y104_D = CLBLL_L_X4Y104_SLICE_X5Y104_DO6;
  assign CLBLL_L_X4Y104_SLICE_X5Y104_AMUX = CLBLL_L_X4Y104_SLICE_X5Y104_AO5;
  assign CLBLL_L_X4Y105_SLICE_X4Y105_A = CLBLL_L_X4Y105_SLICE_X4Y105_AO6;
  assign CLBLL_L_X4Y105_SLICE_X4Y105_B = CLBLL_L_X4Y105_SLICE_X4Y105_BO6;
  assign CLBLL_L_X4Y105_SLICE_X4Y105_C = CLBLL_L_X4Y105_SLICE_X4Y105_CO6;
  assign CLBLL_L_X4Y105_SLICE_X4Y105_D = CLBLL_L_X4Y105_SLICE_X4Y105_DO6;
  assign CLBLL_L_X4Y105_SLICE_X4Y105_AMUX = CLBLL_L_X4Y105_SLICE_X4Y105_AO6;
  assign CLBLL_L_X4Y105_SLICE_X5Y105_A = CLBLL_L_X4Y105_SLICE_X5Y105_AO6;
  assign CLBLL_L_X4Y105_SLICE_X5Y105_B = CLBLL_L_X4Y105_SLICE_X5Y105_BO6;
  assign CLBLL_L_X4Y105_SLICE_X5Y105_C = CLBLL_L_X4Y105_SLICE_X5Y105_CO6;
  assign CLBLL_L_X4Y105_SLICE_X5Y105_D = CLBLL_L_X4Y105_SLICE_X5Y105_DO6;
  assign CLBLL_L_X4Y106_SLICE_X4Y106_A = CLBLL_L_X4Y106_SLICE_X4Y106_AO6;
  assign CLBLL_L_X4Y106_SLICE_X4Y106_B = CLBLL_L_X4Y106_SLICE_X4Y106_BO6;
  assign CLBLL_L_X4Y106_SLICE_X4Y106_C = CLBLL_L_X4Y106_SLICE_X4Y106_CO6;
  assign CLBLL_L_X4Y106_SLICE_X4Y106_D = CLBLL_L_X4Y106_SLICE_X4Y106_DO6;
  assign CLBLL_L_X4Y106_SLICE_X5Y106_A = CLBLL_L_X4Y106_SLICE_X5Y106_AO6;
  assign CLBLL_L_X4Y106_SLICE_X5Y106_B = CLBLL_L_X4Y106_SLICE_X5Y106_BO6;
  assign CLBLL_L_X4Y106_SLICE_X5Y106_C = CLBLL_L_X4Y106_SLICE_X5Y106_CO6;
  assign CLBLL_L_X4Y106_SLICE_X5Y106_D = CLBLL_L_X4Y106_SLICE_X5Y106_DO6;
  assign CLBLL_L_X4Y107_SLICE_X4Y107_A = CLBLL_L_X4Y107_SLICE_X4Y107_AO6;
  assign CLBLL_L_X4Y107_SLICE_X4Y107_B = CLBLL_L_X4Y107_SLICE_X4Y107_BO6;
  assign CLBLL_L_X4Y107_SLICE_X4Y107_C = CLBLL_L_X4Y107_SLICE_X4Y107_CO6;
  assign CLBLL_L_X4Y107_SLICE_X4Y107_D = CLBLL_L_X4Y107_SLICE_X4Y107_DO6;
  assign CLBLL_L_X4Y107_SLICE_X5Y107_A = CLBLL_L_X4Y107_SLICE_X5Y107_AO6;
  assign CLBLL_L_X4Y107_SLICE_X5Y107_B = CLBLL_L_X4Y107_SLICE_X5Y107_BO6;
  assign CLBLL_L_X4Y107_SLICE_X5Y107_C = CLBLL_L_X4Y107_SLICE_X5Y107_CO6;
  assign CLBLL_L_X4Y107_SLICE_X5Y107_D = CLBLL_L_X4Y107_SLICE_X5Y107_DO6;
  assign CLBLL_L_X4Y107_SLICE_X5Y107_AMUX = CLBLL_L_X4Y107_SLICE_X5Y107_AO5;
  assign CLBLL_L_X4Y107_SLICE_X5Y107_CMUX = CLBLL_L_X4Y107_SLICE_X5Y107_CO6;
  assign CLBLL_L_X4Y108_SLICE_X4Y108_A = CLBLL_L_X4Y108_SLICE_X4Y108_AO6;
  assign CLBLL_L_X4Y108_SLICE_X4Y108_B = CLBLL_L_X4Y108_SLICE_X4Y108_BO6;
  assign CLBLL_L_X4Y108_SLICE_X4Y108_C = CLBLL_L_X4Y108_SLICE_X4Y108_CO6;
  assign CLBLL_L_X4Y108_SLICE_X4Y108_D = CLBLL_L_X4Y108_SLICE_X4Y108_DO6;
  assign CLBLL_L_X4Y108_SLICE_X4Y108_AMUX = CLBLL_L_X4Y108_SLICE_X4Y108_AO5;
  assign CLBLL_L_X4Y108_SLICE_X5Y108_A = CLBLL_L_X4Y108_SLICE_X5Y108_AO6;
  assign CLBLL_L_X4Y108_SLICE_X5Y108_B = CLBLL_L_X4Y108_SLICE_X5Y108_BO6;
  assign CLBLL_L_X4Y108_SLICE_X5Y108_C = CLBLL_L_X4Y108_SLICE_X5Y108_CO6;
  assign CLBLL_L_X4Y108_SLICE_X5Y108_D = CLBLL_L_X4Y108_SLICE_X5Y108_DO6;
  assign CLBLL_L_X4Y109_SLICE_X4Y109_A = CLBLL_L_X4Y109_SLICE_X4Y109_AO6;
  assign CLBLL_L_X4Y109_SLICE_X4Y109_B = CLBLL_L_X4Y109_SLICE_X4Y109_BO6;
  assign CLBLL_L_X4Y109_SLICE_X4Y109_C = CLBLL_L_X4Y109_SLICE_X4Y109_CO6;
  assign CLBLL_L_X4Y109_SLICE_X4Y109_D = CLBLL_L_X4Y109_SLICE_X4Y109_DO6;
  assign CLBLL_L_X4Y109_SLICE_X4Y109_AMUX = CLBLL_L_X4Y109_SLICE_X4Y109_AO5;
  assign CLBLL_L_X4Y109_SLICE_X5Y109_A = CLBLL_L_X4Y109_SLICE_X5Y109_AO6;
  assign CLBLL_L_X4Y109_SLICE_X5Y109_B = CLBLL_L_X4Y109_SLICE_X5Y109_BO6;
  assign CLBLL_L_X4Y109_SLICE_X5Y109_C = CLBLL_L_X4Y109_SLICE_X5Y109_CO6;
  assign CLBLL_L_X4Y109_SLICE_X5Y109_D = CLBLL_L_X4Y109_SLICE_X5Y109_DO6;
  assign CLBLL_L_X4Y109_SLICE_X5Y109_AMUX = CLBLL_L_X4Y109_SLICE_X5Y109_AO5;
  assign CLBLL_L_X4Y110_SLICE_X4Y110_A = CLBLL_L_X4Y110_SLICE_X4Y110_AO6;
  assign CLBLL_L_X4Y110_SLICE_X4Y110_B = CLBLL_L_X4Y110_SLICE_X4Y110_BO6;
  assign CLBLL_L_X4Y110_SLICE_X4Y110_C = CLBLL_L_X4Y110_SLICE_X4Y110_CO6;
  assign CLBLL_L_X4Y110_SLICE_X4Y110_D = CLBLL_L_X4Y110_SLICE_X4Y110_DO6;
  assign CLBLL_L_X4Y110_SLICE_X5Y110_A = CLBLL_L_X4Y110_SLICE_X5Y110_AO6;
  assign CLBLL_L_X4Y110_SLICE_X5Y110_B = CLBLL_L_X4Y110_SLICE_X5Y110_BO6;
  assign CLBLL_L_X4Y110_SLICE_X5Y110_C = CLBLL_L_X4Y110_SLICE_X5Y110_CO6;
  assign CLBLL_L_X4Y110_SLICE_X5Y110_D = CLBLL_L_X4Y110_SLICE_X5Y110_DO6;
  assign CLBLL_L_X4Y110_SLICE_X5Y110_AMUX = CLBLL_L_X4Y110_SLICE_X5Y110_AO5;
  assign CLBLL_L_X4Y110_SLICE_X5Y110_BMUX = CLBLL_L_X4Y110_SLICE_X5Y110_BO5;
  assign CLBLL_L_X4Y111_SLICE_X4Y111_A = CLBLL_L_X4Y111_SLICE_X4Y111_AO6;
  assign CLBLL_L_X4Y111_SLICE_X4Y111_B = CLBLL_L_X4Y111_SLICE_X4Y111_BO6;
  assign CLBLL_L_X4Y111_SLICE_X4Y111_C = CLBLL_L_X4Y111_SLICE_X4Y111_CO6;
  assign CLBLL_L_X4Y111_SLICE_X4Y111_D = CLBLL_L_X4Y111_SLICE_X4Y111_DO6;
  assign CLBLL_L_X4Y111_SLICE_X4Y111_AMUX = CLBLL_L_X4Y111_SLICE_X4Y111_AO5;
  assign CLBLL_L_X4Y111_SLICE_X4Y111_BMUX = CLBLL_L_X4Y111_SLICE_X4Y111_BO6;
  assign CLBLL_L_X4Y111_SLICE_X4Y111_CMUX = CLBLL_L_X4Y111_SLICE_X4Y111_CO6;
  assign CLBLL_L_X4Y111_SLICE_X4Y111_DMUX = CLBLL_L_X4Y111_SLICE_X4Y111_DO6;
  assign CLBLL_L_X4Y111_SLICE_X5Y111_A = CLBLL_L_X4Y111_SLICE_X5Y111_AO6;
  assign CLBLL_L_X4Y111_SLICE_X5Y111_B = CLBLL_L_X4Y111_SLICE_X5Y111_BO6;
  assign CLBLL_L_X4Y111_SLICE_X5Y111_C = CLBLL_L_X4Y111_SLICE_X5Y111_CO6;
  assign CLBLL_L_X4Y111_SLICE_X5Y111_D = CLBLL_L_X4Y111_SLICE_X5Y111_DO6;
  assign CLBLL_L_X4Y111_SLICE_X5Y111_AMUX = CLBLL_L_X4Y111_SLICE_X5Y111_AO5;
  assign CLBLL_L_X4Y112_SLICE_X4Y112_A = CLBLL_L_X4Y112_SLICE_X4Y112_AO6;
  assign CLBLL_L_X4Y112_SLICE_X4Y112_B = CLBLL_L_X4Y112_SLICE_X4Y112_BO6;
  assign CLBLL_L_X4Y112_SLICE_X4Y112_C = CLBLL_L_X4Y112_SLICE_X4Y112_CO6;
  assign CLBLL_L_X4Y112_SLICE_X4Y112_D = CLBLL_L_X4Y112_SLICE_X4Y112_DO6;
  assign CLBLL_L_X4Y112_SLICE_X4Y112_AMUX = CLBLL_L_X4Y112_SLICE_X4Y112_AO5;
  assign CLBLL_L_X4Y112_SLICE_X5Y112_A = CLBLL_L_X4Y112_SLICE_X5Y112_AO6;
  assign CLBLL_L_X4Y112_SLICE_X5Y112_B = CLBLL_L_X4Y112_SLICE_X5Y112_BO6;
  assign CLBLL_L_X4Y112_SLICE_X5Y112_C = CLBLL_L_X4Y112_SLICE_X5Y112_CO6;
  assign CLBLL_L_X4Y112_SLICE_X5Y112_D = CLBLL_L_X4Y112_SLICE_X5Y112_DO6;
  assign CLBLL_L_X4Y112_SLICE_X5Y112_CMUX = CLBLL_L_X4Y112_SLICE_X5Y112_CO6;
  assign CLBLL_L_X4Y113_SLICE_X4Y113_A = CLBLL_L_X4Y113_SLICE_X4Y113_AO6;
  assign CLBLL_L_X4Y113_SLICE_X4Y113_B = CLBLL_L_X4Y113_SLICE_X4Y113_BO6;
  assign CLBLL_L_X4Y113_SLICE_X4Y113_C = CLBLL_L_X4Y113_SLICE_X4Y113_CO6;
  assign CLBLL_L_X4Y113_SLICE_X4Y113_D = CLBLL_L_X4Y113_SLICE_X4Y113_DO6;
  assign CLBLL_L_X4Y113_SLICE_X4Y113_AMUX = CLBLL_L_X4Y113_SLICE_X4Y113_AO5;
  assign CLBLL_L_X4Y113_SLICE_X5Y113_A = CLBLL_L_X4Y113_SLICE_X5Y113_AO6;
  assign CLBLL_L_X4Y113_SLICE_X5Y113_B = CLBLL_L_X4Y113_SLICE_X5Y113_BO6;
  assign CLBLL_L_X4Y113_SLICE_X5Y113_C = CLBLL_L_X4Y113_SLICE_X5Y113_CO6;
  assign CLBLL_L_X4Y113_SLICE_X5Y113_D = CLBLL_L_X4Y113_SLICE_X5Y113_DO6;
  assign CLBLL_L_X4Y113_SLICE_X5Y113_AMUX = CLBLL_L_X4Y113_SLICE_X5Y113_AO5;
  assign CLBLL_L_X4Y114_SLICE_X4Y114_A = CLBLL_L_X4Y114_SLICE_X4Y114_AO6;
  assign CLBLL_L_X4Y114_SLICE_X4Y114_B = CLBLL_L_X4Y114_SLICE_X4Y114_BO6;
  assign CLBLL_L_X4Y114_SLICE_X4Y114_C = CLBLL_L_X4Y114_SLICE_X4Y114_CO6;
  assign CLBLL_L_X4Y114_SLICE_X4Y114_D = CLBLL_L_X4Y114_SLICE_X4Y114_DO6;
  assign CLBLL_L_X4Y114_SLICE_X4Y114_AMUX = CLBLL_L_X4Y114_SLICE_X4Y114_AO5;
  assign CLBLL_L_X4Y114_SLICE_X4Y114_BMUX = CLBLL_L_X4Y114_SLICE_X4Y114_BO5;
  assign CLBLL_L_X4Y114_SLICE_X5Y114_A = CLBLL_L_X4Y114_SLICE_X5Y114_AO6;
  assign CLBLL_L_X4Y114_SLICE_X5Y114_B = CLBLL_L_X4Y114_SLICE_X5Y114_BO6;
  assign CLBLL_L_X4Y114_SLICE_X5Y114_C = CLBLL_L_X4Y114_SLICE_X5Y114_CO6;
  assign CLBLL_L_X4Y114_SLICE_X5Y114_D = CLBLL_L_X4Y114_SLICE_X5Y114_DO6;
  assign CLBLL_L_X4Y115_SLICE_X4Y115_A = CLBLL_L_X4Y115_SLICE_X4Y115_AO6;
  assign CLBLL_L_X4Y115_SLICE_X4Y115_B = CLBLL_L_X4Y115_SLICE_X4Y115_BO6;
  assign CLBLL_L_X4Y115_SLICE_X4Y115_C = CLBLL_L_X4Y115_SLICE_X4Y115_CO6;
  assign CLBLL_L_X4Y115_SLICE_X4Y115_D = CLBLL_L_X4Y115_SLICE_X4Y115_DO6;
  assign CLBLL_L_X4Y115_SLICE_X4Y115_AMUX = CLBLL_L_X4Y115_SLICE_X4Y115_AO5;
  assign CLBLL_L_X4Y115_SLICE_X5Y115_A = CLBLL_L_X4Y115_SLICE_X5Y115_AO6;
  assign CLBLL_L_X4Y115_SLICE_X5Y115_B = CLBLL_L_X4Y115_SLICE_X5Y115_BO6;
  assign CLBLL_L_X4Y115_SLICE_X5Y115_C = CLBLL_L_X4Y115_SLICE_X5Y115_CO6;
  assign CLBLL_L_X4Y115_SLICE_X5Y115_D = CLBLL_L_X4Y115_SLICE_X5Y115_DO6;
  assign CLBLL_L_X4Y116_SLICE_X4Y116_A = CLBLL_L_X4Y116_SLICE_X4Y116_AO6;
  assign CLBLL_L_X4Y116_SLICE_X4Y116_B = CLBLL_L_X4Y116_SLICE_X4Y116_BO6;
  assign CLBLL_L_X4Y116_SLICE_X4Y116_C = CLBLL_L_X4Y116_SLICE_X4Y116_CO6;
  assign CLBLL_L_X4Y116_SLICE_X4Y116_D = CLBLL_L_X4Y116_SLICE_X4Y116_DO6;
  assign CLBLL_L_X4Y116_SLICE_X5Y116_A = CLBLL_L_X4Y116_SLICE_X5Y116_AO6;
  assign CLBLL_L_X4Y116_SLICE_X5Y116_B = CLBLL_L_X4Y116_SLICE_X5Y116_BO6;
  assign CLBLL_L_X4Y116_SLICE_X5Y116_C = CLBLL_L_X4Y116_SLICE_X5Y116_CO6;
  assign CLBLL_L_X4Y116_SLICE_X5Y116_D = CLBLL_L_X4Y116_SLICE_X5Y116_DO6;
  assign CLBLM_L_X8Y103_SLICE_X10Y103_A = CLBLM_L_X8Y103_SLICE_X10Y103_AO6;
  assign CLBLM_L_X8Y103_SLICE_X10Y103_B = CLBLM_L_X8Y103_SLICE_X10Y103_BO6;
  assign CLBLM_L_X8Y103_SLICE_X10Y103_C = CLBLM_L_X8Y103_SLICE_X10Y103_CO6;
  assign CLBLM_L_X8Y103_SLICE_X10Y103_D = CLBLM_L_X8Y103_SLICE_X10Y103_DO6;
  assign CLBLM_L_X8Y103_SLICE_X10Y103_AMUX = CLBLM_L_X8Y103_SLICE_X10Y103_AO5;
  assign CLBLM_L_X8Y103_SLICE_X11Y103_A = CLBLM_L_X8Y103_SLICE_X11Y103_AO6;
  assign CLBLM_L_X8Y103_SLICE_X11Y103_B = CLBLM_L_X8Y103_SLICE_X11Y103_BO6;
  assign CLBLM_L_X8Y103_SLICE_X11Y103_C = CLBLM_L_X8Y103_SLICE_X11Y103_CO6;
  assign CLBLM_L_X8Y103_SLICE_X11Y103_D = CLBLM_L_X8Y103_SLICE_X11Y103_DO6;
  assign CLBLM_L_X8Y103_SLICE_X11Y103_AMUX = CLBLM_L_X8Y103_SLICE_X11Y103_AO6;
  assign CLBLM_L_X8Y104_SLICE_X10Y104_A = CLBLM_L_X8Y104_SLICE_X10Y104_AO6;
  assign CLBLM_L_X8Y104_SLICE_X10Y104_B = CLBLM_L_X8Y104_SLICE_X10Y104_BO6;
  assign CLBLM_L_X8Y104_SLICE_X10Y104_C = CLBLM_L_X8Y104_SLICE_X10Y104_CO6;
  assign CLBLM_L_X8Y104_SLICE_X10Y104_D = CLBLM_L_X8Y104_SLICE_X10Y104_DO6;
  assign CLBLM_L_X8Y104_SLICE_X10Y104_AMUX = CLBLM_L_X8Y104_SLICE_X10Y104_AO5;
  assign CLBLM_L_X8Y104_SLICE_X10Y104_CMUX = CLBLM_L_X8Y104_SLICE_X10Y104_CO6;
  assign CLBLM_L_X8Y104_SLICE_X11Y104_A = CLBLM_L_X8Y104_SLICE_X11Y104_AO6;
  assign CLBLM_L_X8Y104_SLICE_X11Y104_B = CLBLM_L_X8Y104_SLICE_X11Y104_BO6;
  assign CLBLM_L_X8Y104_SLICE_X11Y104_C = CLBLM_L_X8Y104_SLICE_X11Y104_CO6;
  assign CLBLM_L_X8Y104_SLICE_X11Y104_D = CLBLM_L_X8Y104_SLICE_X11Y104_DO6;
  assign CLBLM_L_X8Y105_SLICE_X10Y105_A = CLBLM_L_X8Y105_SLICE_X10Y105_AO6;
  assign CLBLM_L_X8Y105_SLICE_X10Y105_B = CLBLM_L_X8Y105_SLICE_X10Y105_BO6;
  assign CLBLM_L_X8Y105_SLICE_X10Y105_C = CLBLM_L_X8Y105_SLICE_X10Y105_CO6;
  assign CLBLM_L_X8Y105_SLICE_X10Y105_D = CLBLM_L_X8Y105_SLICE_X10Y105_DO6;
  assign CLBLM_L_X8Y105_SLICE_X10Y105_AMUX = CLBLM_L_X8Y105_SLICE_X10Y105_AO5;
  assign CLBLM_L_X8Y105_SLICE_X11Y105_A = CLBLM_L_X8Y105_SLICE_X11Y105_AO6;
  assign CLBLM_L_X8Y105_SLICE_X11Y105_B = CLBLM_L_X8Y105_SLICE_X11Y105_BO6;
  assign CLBLM_L_X8Y105_SLICE_X11Y105_C = CLBLM_L_X8Y105_SLICE_X11Y105_CO6;
  assign CLBLM_L_X8Y105_SLICE_X11Y105_D = CLBLM_L_X8Y105_SLICE_X11Y105_DO6;
  assign CLBLM_L_X8Y105_SLICE_X11Y105_AMUX = CLBLM_L_X8Y105_SLICE_X11Y105_AO5;
  assign CLBLM_L_X8Y105_SLICE_X11Y105_BMUX = CLBLM_L_X8Y105_SLICE_X11Y105_BO6;
  assign CLBLM_L_X8Y106_SLICE_X10Y106_A = CLBLM_L_X8Y106_SLICE_X10Y106_AO6;
  assign CLBLM_L_X8Y106_SLICE_X10Y106_B = CLBLM_L_X8Y106_SLICE_X10Y106_BO6;
  assign CLBLM_L_X8Y106_SLICE_X10Y106_C = CLBLM_L_X8Y106_SLICE_X10Y106_CO6;
  assign CLBLM_L_X8Y106_SLICE_X10Y106_D = CLBLM_L_X8Y106_SLICE_X10Y106_DO6;
  assign CLBLM_L_X8Y106_SLICE_X10Y106_AMUX = CLBLM_L_X8Y106_SLICE_X10Y106_AO5;
  assign CLBLM_L_X8Y106_SLICE_X10Y106_BMUX = CLBLM_L_X8Y106_SLICE_X10Y106_BO6;
  assign CLBLM_L_X8Y106_SLICE_X11Y106_A = CLBLM_L_X8Y106_SLICE_X11Y106_AO6;
  assign CLBLM_L_X8Y106_SLICE_X11Y106_B = CLBLM_L_X8Y106_SLICE_X11Y106_BO6;
  assign CLBLM_L_X8Y106_SLICE_X11Y106_C = CLBLM_L_X8Y106_SLICE_X11Y106_CO6;
  assign CLBLM_L_X8Y106_SLICE_X11Y106_D = CLBLM_L_X8Y106_SLICE_X11Y106_DO6;
  assign CLBLM_L_X8Y107_SLICE_X10Y107_A = CLBLM_L_X8Y107_SLICE_X10Y107_AO6;
  assign CLBLM_L_X8Y107_SLICE_X10Y107_B = CLBLM_L_X8Y107_SLICE_X10Y107_BO6;
  assign CLBLM_L_X8Y107_SLICE_X10Y107_C = CLBLM_L_X8Y107_SLICE_X10Y107_CO6;
  assign CLBLM_L_X8Y107_SLICE_X10Y107_D = CLBLM_L_X8Y107_SLICE_X10Y107_DO6;
  assign CLBLM_L_X8Y107_SLICE_X11Y107_A = CLBLM_L_X8Y107_SLICE_X11Y107_AO6;
  assign CLBLM_L_X8Y107_SLICE_X11Y107_B = CLBLM_L_X8Y107_SLICE_X11Y107_BO6;
  assign CLBLM_L_X8Y107_SLICE_X11Y107_C = CLBLM_L_X8Y107_SLICE_X11Y107_CO6;
  assign CLBLM_L_X8Y107_SLICE_X11Y107_D = CLBLM_L_X8Y107_SLICE_X11Y107_DO6;
  assign CLBLM_L_X8Y107_SLICE_X11Y107_AMUX = CLBLM_L_X8Y107_SLICE_X11Y107_AO5;
  assign CLBLM_L_X8Y107_SLICE_X11Y107_BMUX = CLBLM_L_X8Y107_SLICE_X11Y107_BO5;
  assign CLBLM_L_X8Y107_SLICE_X11Y107_CMUX = CLBLM_L_X8Y107_SLICE_X11Y107_CO6;
  assign CLBLM_L_X8Y108_SLICE_X10Y108_A = CLBLM_L_X8Y108_SLICE_X10Y108_AO6;
  assign CLBLM_L_X8Y108_SLICE_X10Y108_B = CLBLM_L_X8Y108_SLICE_X10Y108_BO6;
  assign CLBLM_L_X8Y108_SLICE_X10Y108_C = CLBLM_L_X8Y108_SLICE_X10Y108_CO6;
  assign CLBLM_L_X8Y108_SLICE_X10Y108_D = CLBLM_L_X8Y108_SLICE_X10Y108_DO6;
  assign CLBLM_L_X8Y108_SLICE_X10Y108_AMUX = CLBLM_L_X8Y108_SLICE_X10Y108_AO5;
  assign CLBLM_L_X8Y108_SLICE_X11Y108_A = CLBLM_L_X8Y108_SLICE_X11Y108_AO6;
  assign CLBLM_L_X8Y108_SLICE_X11Y108_B = CLBLM_L_X8Y108_SLICE_X11Y108_BO6;
  assign CLBLM_L_X8Y108_SLICE_X11Y108_C = CLBLM_L_X8Y108_SLICE_X11Y108_CO6;
  assign CLBLM_L_X8Y108_SLICE_X11Y108_D = CLBLM_L_X8Y108_SLICE_X11Y108_DO6;
  assign CLBLM_L_X8Y109_SLICE_X10Y109_A = CLBLM_L_X8Y109_SLICE_X10Y109_AO6;
  assign CLBLM_L_X8Y109_SLICE_X10Y109_B = CLBLM_L_X8Y109_SLICE_X10Y109_BO6;
  assign CLBLM_L_X8Y109_SLICE_X10Y109_C = CLBLM_L_X8Y109_SLICE_X10Y109_CO6;
  assign CLBLM_L_X8Y109_SLICE_X10Y109_D = CLBLM_L_X8Y109_SLICE_X10Y109_DO6;
  assign CLBLM_L_X8Y109_SLICE_X11Y109_A = CLBLM_L_X8Y109_SLICE_X11Y109_AO6;
  assign CLBLM_L_X8Y109_SLICE_X11Y109_B = CLBLM_L_X8Y109_SLICE_X11Y109_BO6;
  assign CLBLM_L_X8Y109_SLICE_X11Y109_C = CLBLM_L_X8Y109_SLICE_X11Y109_CO6;
  assign CLBLM_L_X8Y109_SLICE_X11Y109_D = CLBLM_L_X8Y109_SLICE_X11Y109_DO6;
  assign CLBLM_L_X8Y110_SLICE_X10Y110_A = CLBLM_L_X8Y110_SLICE_X10Y110_AO6;
  assign CLBLM_L_X8Y110_SLICE_X10Y110_B = CLBLM_L_X8Y110_SLICE_X10Y110_BO6;
  assign CLBLM_L_X8Y110_SLICE_X10Y110_C = CLBLM_L_X8Y110_SLICE_X10Y110_CO6;
  assign CLBLM_L_X8Y110_SLICE_X10Y110_D = CLBLM_L_X8Y110_SLICE_X10Y110_DO6;
  assign CLBLM_L_X8Y110_SLICE_X10Y110_CMUX = CLBLM_L_X8Y110_SLICE_X10Y110_CO6;
  assign CLBLM_L_X8Y110_SLICE_X11Y110_A = CLBLM_L_X8Y110_SLICE_X11Y110_AO6;
  assign CLBLM_L_X8Y110_SLICE_X11Y110_B = CLBLM_L_X8Y110_SLICE_X11Y110_BO6;
  assign CLBLM_L_X8Y110_SLICE_X11Y110_C = CLBLM_L_X8Y110_SLICE_X11Y110_CO6;
  assign CLBLM_L_X8Y110_SLICE_X11Y110_D = CLBLM_L_X8Y110_SLICE_X11Y110_DO6;
  assign CLBLM_L_X8Y110_SLICE_X11Y110_AMUX = CLBLM_L_X8Y110_SLICE_X11Y110_AO5;
  assign CLBLM_L_X8Y110_SLICE_X11Y110_BMUX = CLBLM_L_X8Y110_SLICE_X11Y110_BO6;
  assign CLBLM_L_X8Y111_SLICE_X10Y111_A = CLBLM_L_X8Y111_SLICE_X10Y111_AO6;
  assign CLBLM_L_X8Y111_SLICE_X10Y111_B = CLBLM_L_X8Y111_SLICE_X10Y111_BO6;
  assign CLBLM_L_X8Y111_SLICE_X10Y111_C = CLBLM_L_X8Y111_SLICE_X10Y111_CO6;
  assign CLBLM_L_X8Y111_SLICE_X10Y111_D = CLBLM_L_X8Y111_SLICE_X10Y111_DO6;
  assign CLBLM_L_X8Y111_SLICE_X10Y111_AMUX = CLBLM_L_X8Y111_SLICE_X10Y111_AO5;
  assign CLBLM_L_X8Y111_SLICE_X11Y111_A = CLBLM_L_X8Y111_SLICE_X11Y111_AO6;
  assign CLBLM_L_X8Y111_SLICE_X11Y111_B = CLBLM_L_X8Y111_SLICE_X11Y111_BO6;
  assign CLBLM_L_X8Y111_SLICE_X11Y111_C = CLBLM_L_X8Y111_SLICE_X11Y111_CO6;
  assign CLBLM_L_X8Y111_SLICE_X11Y111_D = CLBLM_L_X8Y111_SLICE_X11Y111_DO6;
  assign CLBLM_L_X8Y111_SLICE_X11Y111_AMUX = CLBLM_L_X8Y111_SLICE_X11Y111_AO5;
  assign CLBLM_L_X8Y112_SLICE_X10Y112_A = CLBLM_L_X8Y112_SLICE_X10Y112_AO6;
  assign CLBLM_L_X8Y112_SLICE_X10Y112_B = CLBLM_L_X8Y112_SLICE_X10Y112_BO6;
  assign CLBLM_L_X8Y112_SLICE_X10Y112_C = CLBLM_L_X8Y112_SLICE_X10Y112_CO6;
  assign CLBLM_L_X8Y112_SLICE_X10Y112_D = CLBLM_L_X8Y112_SLICE_X10Y112_DO6;
  assign CLBLM_L_X8Y112_SLICE_X10Y112_AMUX = CLBLM_L_X8Y112_SLICE_X10Y112_AO5;
  assign CLBLM_L_X8Y112_SLICE_X11Y112_A = CLBLM_L_X8Y112_SLICE_X11Y112_AO6;
  assign CLBLM_L_X8Y112_SLICE_X11Y112_B = CLBLM_L_X8Y112_SLICE_X11Y112_BO6;
  assign CLBLM_L_X8Y112_SLICE_X11Y112_C = CLBLM_L_X8Y112_SLICE_X11Y112_CO6;
  assign CLBLM_L_X8Y112_SLICE_X11Y112_D = CLBLM_L_X8Y112_SLICE_X11Y112_DO6;
  assign CLBLM_L_X8Y113_SLICE_X10Y113_A = CLBLM_L_X8Y113_SLICE_X10Y113_AO6;
  assign CLBLM_L_X8Y113_SLICE_X10Y113_B = CLBLM_L_X8Y113_SLICE_X10Y113_BO6;
  assign CLBLM_L_X8Y113_SLICE_X10Y113_C = CLBLM_L_X8Y113_SLICE_X10Y113_CO6;
  assign CLBLM_L_X8Y113_SLICE_X10Y113_D = CLBLM_L_X8Y113_SLICE_X10Y113_DO6;
  assign CLBLM_L_X8Y113_SLICE_X10Y113_AMUX = CLBLM_L_X8Y113_SLICE_X10Y113_AO5;
  assign CLBLM_L_X8Y113_SLICE_X11Y113_A = CLBLM_L_X8Y113_SLICE_X11Y113_AO6;
  assign CLBLM_L_X8Y113_SLICE_X11Y113_B = CLBLM_L_X8Y113_SLICE_X11Y113_BO6;
  assign CLBLM_L_X8Y113_SLICE_X11Y113_C = CLBLM_L_X8Y113_SLICE_X11Y113_CO6;
  assign CLBLM_L_X8Y113_SLICE_X11Y113_D = CLBLM_L_X8Y113_SLICE_X11Y113_DO6;
  assign CLBLM_L_X10Y102_SLICE_X12Y102_A = CLBLM_L_X10Y102_SLICE_X12Y102_AO6;
  assign CLBLM_L_X10Y102_SLICE_X12Y102_B = CLBLM_L_X10Y102_SLICE_X12Y102_BO6;
  assign CLBLM_L_X10Y102_SLICE_X12Y102_C = CLBLM_L_X10Y102_SLICE_X12Y102_CO6;
  assign CLBLM_L_X10Y102_SLICE_X12Y102_D = CLBLM_L_X10Y102_SLICE_X12Y102_DO6;
  assign CLBLM_L_X10Y102_SLICE_X12Y102_AMUX = CLBLM_L_X10Y102_SLICE_X12Y102_AO5;
  assign CLBLM_L_X10Y102_SLICE_X12Y102_BMUX = CLBLM_L_X10Y102_SLICE_X12Y102_BO6;
  assign CLBLM_L_X10Y102_SLICE_X13Y102_A = CLBLM_L_X10Y102_SLICE_X13Y102_AO6;
  assign CLBLM_L_X10Y102_SLICE_X13Y102_B = CLBLM_L_X10Y102_SLICE_X13Y102_BO6;
  assign CLBLM_L_X10Y102_SLICE_X13Y102_C = CLBLM_L_X10Y102_SLICE_X13Y102_CO6;
  assign CLBLM_L_X10Y102_SLICE_X13Y102_D = CLBLM_L_X10Y102_SLICE_X13Y102_DO6;
  assign CLBLM_L_X10Y103_SLICE_X12Y103_A = CLBLM_L_X10Y103_SLICE_X12Y103_AO6;
  assign CLBLM_L_X10Y103_SLICE_X12Y103_B = CLBLM_L_X10Y103_SLICE_X12Y103_BO6;
  assign CLBLM_L_X10Y103_SLICE_X12Y103_C = CLBLM_L_X10Y103_SLICE_X12Y103_CO6;
  assign CLBLM_L_X10Y103_SLICE_X12Y103_D = CLBLM_L_X10Y103_SLICE_X12Y103_DO6;
  assign CLBLM_L_X10Y103_SLICE_X12Y103_AMUX = CLBLM_L_X10Y103_SLICE_X12Y103_AO5;
  assign CLBLM_L_X10Y103_SLICE_X13Y103_A = CLBLM_L_X10Y103_SLICE_X13Y103_AO6;
  assign CLBLM_L_X10Y103_SLICE_X13Y103_B = CLBLM_L_X10Y103_SLICE_X13Y103_BO6;
  assign CLBLM_L_X10Y103_SLICE_X13Y103_C = CLBLM_L_X10Y103_SLICE_X13Y103_CO6;
  assign CLBLM_L_X10Y103_SLICE_X13Y103_D = CLBLM_L_X10Y103_SLICE_X13Y103_DO6;
  assign CLBLM_L_X10Y104_SLICE_X12Y104_A = CLBLM_L_X10Y104_SLICE_X12Y104_AO6;
  assign CLBLM_L_X10Y104_SLICE_X12Y104_B = CLBLM_L_X10Y104_SLICE_X12Y104_BO6;
  assign CLBLM_L_X10Y104_SLICE_X12Y104_C = CLBLM_L_X10Y104_SLICE_X12Y104_CO6;
  assign CLBLM_L_X10Y104_SLICE_X12Y104_D = CLBLM_L_X10Y104_SLICE_X12Y104_DO6;
  assign CLBLM_L_X10Y104_SLICE_X12Y104_BMUX = CLBLM_L_X10Y104_SLICE_X12Y104_BO6;
  assign CLBLM_L_X10Y104_SLICE_X13Y104_A = CLBLM_L_X10Y104_SLICE_X13Y104_AO6;
  assign CLBLM_L_X10Y104_SLICE_X13Y104_B = CLBLM_L_X10Y104_SLICE_X13Y104_BO6;
  assign CLBLM_L_X10Y104_SLICE_X13Y104_C = CLBLM_L_X10Y104_SLICE_X13Y104_CO6;
  assign CLBLM_L_X10Y104_SLICE_X13Y104_D = CLBLM_L_X10Y104_SLICE_X13Y104_DO6;
  assign CLBLM_L_X10Y104_SLICE_X13Y104_AMUX = CLBLM_L_X10Y104_SLICE_X13Y104_AO5;
  assign CLBLM_L_X10Y105_SLICE_X12Y105_A = CLBLM_L_X10Y105_SLICE_X12Y105_AO6;
  assign CLBLM_L_X10Y105_SLICE_X12Y105_B = CLBLM_L_X10Y105_SLICE_X12Y105_BO6;
  assign CLBLM_L_X10Y105_SLICE_X12Y105_C = CLBLM_L_X10Y105_SLICE_X12Y105_CO6;
  assign CLBLM_L_X10Y105_SLICE_X12Y105_D = CLBLM_L_X10Y105_SLICE_X12Y105_DO6;
  assign CLBLM_L_X10Y105_SLICE_X12Y105_AMUX = CLBLM_L_X10Y105_SLICE_X12Y105_AO5;
  assign CLBLM_L_X10Y105_SLICE_X13Y105_A = CLBLM_L_X10Y105_SLICE_X13Y105_AO6;
  assign CLBLM_L_X10Y105_SLICE_X13Y105_B = CLBLM_L_X10Y105_SLICE_X13Y105_BO6;
  assign CLBLM_L_X10Y105_SLICE_X13Y105_C = CLBLM_L_X10Y105_SLICE_X13Y105_CO6;
  assign CLBLM_L_X10Y105_SLICE_X13Y105_D = CLBLM_L_X10Y105_SLICE_X13Y105_DO6;
  assign CLBLM_L_X10Y105_SLICE_X13Y105_AMUX = CLBLM_L_X10Y105_SLICE_X13Y105_AO5;
  assign CLBLM_L_X10Y106_SLICE_X12Y106_A = CLBLM_L_X10Y106_SLICE_X12Y106_AO6;
  assign CLBLM_L_X10Y106_SLICE_X12Y106_B = CLBLM_L_X10Y106_SLICE_X12Y106_BO6;
  assign CLBLM_L_X10Y106_SLICE_X12Y106_C = CLBLM_L_X10Y106_SLICE_X12Y106_CO6;
  assign CLBLM_L_X10Y106_SLICE_X12Y106_D = CLBLM_L_X10Y106_SLICE_X12Y106_DO6;
  assign CLBLM_L_X10Y106_SLICE_X13Y106_A = CLBLM_L_X10Y106_SLICE_X13Y106_AO6;
  assign CLBLM_L_X10Y106_SLICE_X13Y106_B = CLBLM_L_X10Y106_SLICE_X13Y106_BO6;
  assign CLBLM_L_X10Y106_SLICE_X13Y106_C = CLBLM_L_X10Y106_SLICE_X13Y106_CO6;
  assign CLBLM_L_X10Y106_SLICE_X13Y106_D = CLBLM_L_X10Y106_SLICE_X13Y106_DO6;
  assign CLBLM_L_X10Y107_SLICE_X12Y107_A = CLBLM_L_X10Y107_SLICE_X12Y107_AO6;
  assign CLBLM_L_X10Y107_SLICE_X12Y107_B = CLBLM_L_X10Y107_SLICE_X12Y107_BO6;
  assign CLBLM_L_X10Y107_SLICE_X12Y107_C = CLBLM_L_X10Y107_SLICE_X12Y107_CO6;
  assign CLBLM_L_X10Y107_SLICE_X12Y107_D = CLBLM_L_X10Y107_SLICE_X12Y107_DO6;
  assign CLBLM_L_X10Y107_SLICE_X13Y107_A = CLBLM_L_X10Y107_SLICE_X13Y107_AO6;
  assign CLBLM_L_X10Y107_SLICE_X13Y107_B = CLBLM_L_X10Y107_SLICE_X13Y107_BO6;
  assign CLBLM_L_X10Y107_SLICE_X13Y107_C = CLBLM_L_X10Y107_SLICE_X13Y107_CO6;
  assign CLBLM_L_X10Y107_SLICE_X13Y107_D = CLBLM_L_X10Y107_SLICE_X13Y107_DO6;
  assign CLBLM_L_X10Y107_SLICE_X13Y107_AMUX = CLBLM_L_X10Y107_SLICE_X13Y107_AO6;
  assign CLBLM_L_X10Y108_SLICE_X12Y108_A = CLBLM_L_X10Y108_SLICE_X12Y108_AO6;
  assign CLBLM_L_X10Y108_SLICE_X12Y108_B = CLBLM_L_X10Y108_SLICE_X12Y108_BO6;
  assign CLBLM_L_X10Y108_SLICE_X12Y108_C = CLBLM_L_X10Y108_SLICE_X12Y108_CO6;
  assign CLBLM_L_X10Y108_SLICE_X12Y108_D = CLBLM_L_X10Y108_SLICE_X12Y108_DO6;
  assign CLBLM_L_X10Y108_SLICE_X13Y108_A = CLBLM_L_X10Y108_SLICE_X13Y108_AO6;
  assign CLBLM_L_X10Y108_SLICE_X13Y108_B = CLBLM_L_X10Y108_SLICE_X13Y108_BO6;
  assign CLBLM_L_X10Y108_SLICE_X13Y108_C = CLBLM_L_X10Y108_SLICE_X13Y108_CO6;
  assign CLBLM_L_X10Y108_SLICE_X13Y108_D = CLBLM_L_X10Y108_SLICE_X13Y108_DO6;
  assign CLBLM_L_X10Y108_SLICE_X13Y108_AMUX = CLBLM_L_X10Y108_SLICE_X13Y108_AO5;
  assign CLBLM_L_X10Y108_SLICE_X13Y108_BMUX = CLBLM_L_X10Y108_SLICE_X13Y108_BO5;
  assign CLBLM_L_X10Y108_SLICE_X13Y108_CMUX = CLBLM_L_X10Y108_SLICE_X13Y108_CO6;
  assign CLBLM_L_X10Y109_SLICE_X12Y109_A = CLBLM_L_X10Y109_SLICE_X12Y109_AO6;
  assign CLBLM_L_X10Y109_SLICE_X12Y109_B = CLBLM_L_X10Y109_SLICE_X12Y109_BO6;
  assign CLBLM_L_X10Y109_SLICE_X12Y109_C = CLBLM_L_X10Y109_SLICE_X12Y109_CO6;
  assign CLBLM_L_X10Y109_SLICE_X12Y109_D = CLBLM_L_X10Y109_SLICE_X12Y109_DO6;
  assign CLBLM_L_X10Y109_SLICE_X12Y109_AMUX = CLBLM_L_X10Y109_SLICE_X12Y109_AO6;
  assign CLBLM_L_X10Y109_SLICE_X13Y109_A = CLBLM_L_X10Y109_SLICE_X13Y109_AO6;
  assign CLBLM_L_X10Y109_SLICE_X13Y109_B = CLBLM_L_X10Y109_SLICE_X13Y109_BO6;
  assign CLBLM_L_X10Y109_SLICE_X13Y109_C = CLBLM_L_X10Y109_SLICE_X13Y109_CO6;
  assign CLBLM_L_X10Y109_SLICE_X13Y109_D = CLBLM_L_X10Y109_SLICE_X13Y109_DO6;
  assign CLBLM_L_X10Y109_SLICE_X13Y109_AMUX = CLBLM_L_X10Y109_SLICE_X13Y109_AO5;
  assign CLBLM_L_X10Y110_SLICE_X12Y110_A = CLBLM_L_X10Y110_SLICE_X12Y110_AO6;
  assign CLBLM_L_X10Y110_SLICE_X12Y110_B = CLBLM_L_X10Y110_SLICE_X12Y110_BO6;
  assign CLBLM_L_X10Y110_SLICE_X12Y110_C = CLBLM_L_X10Y110_SLICE_X12Y110_CO6;
  assign CLBLM_L_X10Y110_SLICE_X12Y110_D = CLBLM_L_X10Y110_SLICE_X12Y110_DO6;
  assign CLBLM_L_X10Y110_SLICE_X13Y110_A = CLBLM_L_X10Y110_SLICE_X13Y110_AO6;
  assign CLBLM_L_X10Y110_SLICE_X13Y110_B = CLBLM_L_X10Y110_SLICE_X13Y110_BO6;
  assign CLBLM_L_X10Y110_SLICE_X13Y110_C = CLBLM_L_X10Y110_SLICE_X13Y110_CO6;
  assign CLBLM_L_X10Y110_SLICE_X13Y110_D = CLBLM_L_X10Y110_SLICE_X13Y110_DO6;
  assign CLBLM_L_X10Y110_SLICE_X13Y110_AMUX = CLBLM_L_X10Y110_SLICE_X13Y110_AO5;
  assign CLBLM_L_X10Y111_SLICE_X12Y111_A = CLBLM_L_X10Y111_SLICE_X12Y111_AO6;
  assign CLBLM_L_X10Y111_SLICE_X12Y111_B = CLBLM_L_X10Y111_SLICE_X12Y111_BO6;
  assign CLBLM_L_X10Y111_SLICE_X12Y111_C = CLBLM_L_X10Y111_SLICE_X12Y111_CO6;
  assign CLBLM_L_X10Y111_SLICE_X12Y111_D = CLBLM_L_X10Y111_SLICE_X12Y111_DO6;
  assign CLBLM_L_X10Y111_SLICE_X13Y111_A = CLBLM_L_X10Y111_SLICE_X13Y111_AO6;
  assign CLBLM_L_X10Y111_SLICE_X13Y111_B = CLBLM_L_X10Y111_SLICE_X13Y111_BO6;
  assign CLBLM_L_X10Y111_SLICE_X13Y111_C = CLBLM_L_X10Y111_SLICE_X13Y111_CO6;
  assign CLBLM_L_X10Y111_SLICE_X13Y111_D = CLBLM_L_X10Y111_SLICE_X13Y111_DO6;
  assign CLBLM_L_X10Y111_SLICE_X13Y111_AMUX = CLBLM_L_X10Y111_SLICE_X13Y111_AO5;
  assign CLBLM_L_X10Y111_SLICE_X13Y111_BMUX = CLBLM_L_X10Y111_SLICE_X13Y111_BO6;
  assign CLBLM_L_X10Y112_SLICE_X12Y112_A = CLBLM_L_X10Y112_SLICE_X12Y112_AO6;
  assign CLBLM_L_X10Y112_SLICE_X12Y112_B = CLBLM_L_X10Y112_SLICE_X12Y112_BO6;
  assign CLBLM_L_X10Y112_SLICE_X12Y112_C = CLBLM_L_X10Y112_SLICE_X12Y112_CO6;
  assign CLBLM_L_X10Y112_SLICE_X12Y112_D = CLBLM_L_X10Y112_SLICE_X12Y112_DO6;
  assign CLBLM_L_X10Y112_SLICE_X13Y112_A = CLBLM_L_X10Y112_SLICE_X13Y112_AO6;
  assign CLBLM_L_X10Y112_SLICE_X13Y112_B = CLBLM_L_X10Y112_SLICE_X13Y112_BO6;
  assign CLBLM_L_X10Y112_SLICE_X13Y112_C = CLBLM_L_X10Y112_SLICE_X13Y112_CO6;
  assign CLBLM_L_X10Y112_SLICE_X13Y112_D = CLBLM_L_X10Y112_SLICE_X13Y112_DO6;
  assign CLBLM_L_X10Y112_SLICE_X13Y112_AMUX = CLBLM_L_X10Y112_SLICE_X13Y112_AO5;
  assign CLBLM_L_X12Y104_SLICE_X16Y104_A = CLBLM_L_X12Y104_SLICE_X16Y104_AO6;
  assign CLBLM_L_X12Y104_SLICE_X16Y104_B = CLBLM_L_X12Y104_SLICE_X16Y104_BO6;
  assign CLBLM_L_X12Y104_SLICE_X16Y104_C = CLBLM_L_X12Y104_SLICE_X16Y104_CO6;
  assign CLBLM_L_X12Y104_SLICE_X16Y104_D = CLBLM_L_X12Y104_SLICE_X16Y104_DO6;
  assign CLBLM_L_X12Y104_SLICE_X16Y104_AMUX = CLBLM_L_X12Y104_SLICE_X16Y104_AO5;
  assign CLBLM_L_X12Y104_SLICE_X17Y104_A = CLBLM_L_X12Y104_SLICE_X17Y104_AO6;
  assign CLBLM_L_X12Y104_SLICE_X17Y104_B = CLBLM_L_X12Y104_SLICE_X17Y104_BO6;
  assign CLBLM_L_X12Y104_SLICE_X17Y104_C = CLBLM_L_X12Y104_SLICE_X17Y104_CO6;
  assign CLBLM_L_X12Y104_SLICE_X17Y104_D = CLBLM_L_X12Y104_SLICE_X17Y104_DO6;
  assign CLBLM_L_X12Y105_SLICE_X16Y105_A = CLBLM_L_X12Y105_SLICE_X16Y105_AO6;
  assign CLBLM_L_X12Y105_SLICE_X16Y105_B = CLBLM_L_X12Y105_SLICE_X16Y105_BO6;
  assign CLBLM_L_X12Y105_SLICE_X16Y105_C = CLBLM_L_X12Y105_SLICE_X16Y105_CO6;
  assign CLBLM_L_X12Y105_SLICE_X16Y105_D = CLBLM_L_X12Y105_SLICE_X16Y105_DO6;
  assign CLBLM_L_X12Y105_SLICE_X16Y105_AMUX = CLBLM_L_X12Y105_SLICE_X16Y105_AO5;
  assign CLBLM_L_X12Y105_SLICE_X17Y105_A = CLBLM_L_X12Y105_SLICE_X17Y105_AO6;
  assign CLBLM_L_X12Y105_SLICE_X17Y105_B = CLBLM_L_X12Y105_SLICE_X17Y105_BO6;
  assign CLBLM_L_X12Y105_SLICE_X17Y105_C = CLBLM_L_X12Y105_SLICE_X17Y105_CO6;
  assign CLBLM_L_X12Y105_SLICE_X17Y105_D = CLBLM_L_X12Y105_SLICE_X17Y105_DO6;
  assign CLBLM_L_X12Y106_SLICE_X16Y106_A = CLBLM_L_X12Y106_SLICE_X16Y106_AO6;
  assign CLBLM_L_X12Y106_SLICE_X16Y106_B = CLBLM_L_X12Y106_SLICE_X16Y106_BO6;
  assign CLBLM_L_X12Y106_SLICE_X16Y106_C = CLBLM_L_X12Y106_SLICE_X16Y106_CO6;
  assign CLBLM_L_X12Y106_SLICE_X16Y106_D = CLBLM_L_X12Y106_SLICE_X16Y106_DO6;
  assign CLBLM_L_X12Y106_SLICE_X16Y106_AMUX = CLBLM_L_X12Y106_SLICE_X16Y106_AO5;
  assign CLBLM_L_X12Y106_SLICE_X16Y106_BMUX = CLBLM_L_X12Y106_SLICE_X16Y106_BO5;
  assign CLBLM_L_X12Y106_SLICE_X17Y106_A = CLBLM_L_X12Y106_SLICE_X17Y106_AO6;
  assign CLBLM_L_X12Y106_SLICE_X17Y106_B = CLBLM_L_X12Y106_SLICE_X17Y106_BO6;
  assign CLBLM_L_X12Y106_SLICE_X17Y106_C = CLBLM_L_X12Y106_SLICE_X17Y106_CO6;
  assign CLBLM_L_X12Y106_SLICE_X17Y106_D = CLBLM_L_X12Y106_SLICE_X17Y106_DO6;
  assign CLBLM_L_X12Y106_SLICE_X17Y106_AMUX = CLBLM_L_X12Y106_SLICE_X17Y106_AO5;
  assign CLBLM_L_X12Y107_SLICE_X16Y107_A = CLBLM_L_X12Y107_SLICE_X16Y107_AO6;
  assign CLBLM_L_X12Y107_SLICE_X16Y107_B = CLBLM_L_X12Y107_SLICE_X16Y107_BO6;
  assign CLBLM_L_X12Y107_SLICE_X16Y107_C = CLBLM_L_X12Y107_SLICE_X16Y107_CO6;
  assign CLBLM_L_X12Y107_SLICE_X16Y107_D = CLBLM_L_X12Y107_SLICE_X16Y107_DO6;
  assign CLBLM_L_X12Y107_SLICE_X17Y107_A = CLBLM_L_X12Y107_SLICE_X17Y107_AO6;
  assign CLBLM_L_X12Y107_SLICE_X17Y107_B = CLBLM_L_X12Y107_SLICE_X17Y107_BO6;
  assign CLBLM_L_X12Y107_SLICE_X17Y107_C = CLBLM_L_X12Y107_SLICE_X17Y107_CO6;
  assign CLBLM_L_X12Y107_SLICE_X17Y107_D = CLBLM_L_X12Y107_SLICE_X17Y107_DO6;
  assign CLBLM_L_X12Y107_SLICE_X17Y107_AMUX = CLBLM_L_X12Y107_SLICE_X17Y107_AO5;
  assign CLBLM_L_X12Y108_SLICE_X16Y108_A = CLBLM_L_X12Y108_SLICE_X16Y108_AO6;
  assign CLBLM_L_X12Y108_SLICE_X16Y108_B = CLBLM_L_X12Y108_SLICE_X16Y108_BO6;
  assign CLBLM_L_X12Y108_SLICE_X16Y108_C = CLBLM_L_X12Y108_SLICE_X16Y108_CO6;
  assign CLBLM_L_X12Y108_SLICE_X16Y108_D = CLBLM_L_X12Y108_SLICE_X16Y108_DO6;
  assign CLBLM_L_X12Y108_SLICE_X16Y108_AMUX = CLBLM_L_X12Y108_SLICE_X16Y108_AO5;
  assign CLBLM_L_X12Y108_SLICE_X17Y108_A = CLBLM_L_X12Y108_SLICE_X17Y108_AO6;
  assign CLBLM_L_X12Y108_SLICE_X17Y108_B = CLBLM_L_X12Y108_SLICE_X17Y108_BO6;
  assign CLBLM_L_X12Y108_SLICE_X17Y108_C = CLBLM_L_X12Y108_SLICE_X17Y108_CO6;
  assign CLBLM_L_X12Y108_SLICE_X17Y108_D = CLBLM_L_X12Y108_SLICE_X17Y108_DO6;
  assign CLBLM_L_X12Y109_SLICE_X16Y109_A = CLBLM_L_X12Y109_SLICE_X16Y109_AO6;
  assign CLBLM_L_X12Y109_SLICE_X16Y109_B = CLBLM_L_X12Y109_SLICE_X16Y109_BO6;
  assign CLBLM_L_X12Y109_SLICE_X16Y109_C = CLBLM_L_X12Y109_SLICE_X16Y109_CO6;
  assign CLBLM_L_X12Y109_SLICE_X16Y109_D = CLBLM_L_X12Y109_SLICE_X16Y109_DO6;
  assign CLBLM_L_X12Y109_SLICE_X16Y109_AMUX = CLBLM_L_X12Y109_SLICE_X16Y109_AO5;
  assign CLBLM_L_X12Y109_SLICE_X17Y109_A = CLBLM_L_X12Y109_SLICE_X17Y109_AO6;
  assign CLBLM_L_X12Y109_SLICE_X17Y109_B = CLBLM_L_X12Y109_SLICE_X17Y109_BO6;
  assign CLBLM_L_X12Y109_SLICE_X17Y109_C = CLBLM_L_X12Y109_SLICE_X17Y109_CO6;
  assign CLBLM_L_X12Y109_SLICE_X17Y109_D = CLBLM_L_X12Y109_SLICE_X17Y109_DO6;
  assign CLBLM_L_X12Y109_SLICE_X17Y109_BMUX = CLBLM_L_X12Y109_SLICE_X17Y109_BO6;
  assign CLBLM_L_X12Y110_SLICE_X16Y110_A = CLBLM_L_X12Y110_SLICE_X16Y110_AO6;
  assign CLBLM_L_X12Y110_SLICE_X16Y110_B = CLBLM_L_X12Y110_SLICE_X16Y110_BO6;
  assign CLBLM_L_X12Y110_SLICE_X16Y110_C = CLBLM_L_X12Y110_SLICE_X16Y110_CO6;
  assign CLBLM_L_X12Y110_SLICE_X16Y110_D = CLBLM_L_X12Y110_SLICE_X16Y110_DO6;
  assign CLBLM_L_X12Y110_SLICE_X16Y110_AMUX = CLBLM_L_X12Y110_SLICE_X16Y110_AO5;
  assign CLBLM_L_X12Y110_SLICE_X17Y110_A = CLBLM_L_X12Y110_SLICE_X17Y110_AO6;
  assign CLBLM_L_X12Y110_SLICE_X17Y110_B = CLBLM_L_X12Y110_SLICE_X17Y110_BO6;
  assign CLBLM_L_X12Y110_SLICE_X17Y110_C = CLBLM_L_X12Y110_SLICE_X17Y110_CO6;
  assign CLBLM_L_X12Y110_SLICE_X17Y110_D = CLBLM_L_X12Y110_SLICE_X17Y110_DO6;
  assign CLBLM_R_X3Y103_SLICE_X2Y103_A = CLBLM_R_X3Y103_SLICE_X2Y103_AO6;
  assign CLBLM_R_X3Y103_SLICE_X2Y103_B = CLBLM_R_X3Y103_SLICE_X2Y103_BO6;
  assign CLBLM_R_X3Y103_SLICE_X2Y103_C = CLBLM_R_X3Y103_SLICE_X2Y103_CO6;
  assign CLBLM_R_X3Y103_SLICE_X2Y103_D = CLBLM_R_X3Y103_SLICE_X2Y103_DO6;
  assign CLBLM_R_X3Y103_SLICE_X3Y103_A = CLBLM_R_X3Y103_SLICE_X3Y103_AO6;
  assign CLBLM_R_X3Y103_SLICE_X3Y103_B = CLBLM_R_X3Y103_SLICE_X3Y103_BO6;
  assign CLBLM_R_X3Y103_SLICE_X3Y103_C = CLBLM_R_X3Y103_SLICE_X3Y103_CO6;
  assign CLBLM_R_X3Y103_SLICE_X3Y103_D = CLBLM_R_X3Y103_SLICE_X3Y103_DO6;
  assign CLBLM_R_X3Y103_SLICE_X3Y103_AMUX = CLBLM_R_X3Y103_SLICE_X3Y103_AO5;
  assign CLBLM_R_X3Y104_SLICE_X2Y104_A = CLBLM_R_X3Y104_SLICE_X2Y104_AO6;
  assign CLBLM_R_X3Y104_SLICE_X2Y104_B = CLBLM_R_X3Y104_SLICE_X2Y104_BO6;
  assign CLBLM_R_X3Y104_SLICE_X2Y104_C = CLBLM_R_X3Y104_SLICE_X2Y104_CO6;
  assign CLBLM_R_X3Y104_SLICE_X2Y104_D = CLBLM_R_X3Y104_SLICE_X2Y104_DO6;
  assign CLBLM_R_X3Y104_SLICE_X2Y104_AMUX = CLBLM_R_X3Y104_SLICE_X2Y104_AO5;
  assign CLBLM_R_X3Y104_SLICE_X3Y104_A = CLBLM_R_X3Y104_SLICE_X3Y104_AO6;
  assign CLBLM_R_X3Y104_SLICE_X3Y104_B = CLBLM_R_X3Y104_SLICE_X3Y104_BO6;
  assign CLBLM_R_X3Y104_SLICE_X3Y104_C = CLBLM_R_X3Y104_SLICE_X3Y104_CO6;
  assign CLBLM_R_X3Y104_SLICE_X3Y104_D = CLBLM_R_X3Y104_SLICE_X3Y104_DO6;
  assign CLBLM_R_X3Y104_SLICE_X3Y104_AMUX = CLBLM_R_X3Y104_SLICE_X3Y104_AO5;
  assign CLBLM_R_X3Y105_SLICE_X2Y105_A = CLBLM_R_X3Y105_SLICE_X2Y105_AO6;
  assign CLBLM_R_X3Y105_SLICE_X2Y105_B = CLBLM_R_X3Y105_SLICE_X2Y105_BO6;
  assign CLBLM_R_X3Y105_SLICE_X2Y105_C = CLBLM_R_X3Y105_SLICE_X2Y105_CO6;
  assign CLBLM_R_X3Y105_SLICE_X2Y105_D = CLBLM_R_X3Y105_SLICE_X2Y105_DO6;
  assign CLBLM_R_X3Y105_SLICE_X3Y105_A = CLBLM_R_X3Y105_SLICE_X3Y105_AO6;
  assign CLBLM_R_X3Y105_SLICE_X3Y105_B = CLBLM_R_X3Y105_SLICE_X3Y105_BO6;
  assign CLBLM_R_X3Y105_SLICE_X3Y105_C = CLBLM_R_X3Y105_SLICE_X3Y105_CO6;
  assign CLBLM_R_X3Y105_SLICE_X3Y105_D = CLBLM_R_X3Y105_SLICE_X3Y105_DO6;
  assign CLBLM_R_X3Y106_SLICE_X2Y106_A = CLBLM_R_X3Y106_SLICE_X2Y106_AO6;
  assign CLBLM_R_X3Y106_SLICE_X2Y106_B = CLBLM_R_X3Y106_SLICE_X2Y106_BO6;
  assign CLBLM_R_X3Y106_SLICE_X2Y106_C = CLBLM_R_X3Y106_SLICE_X2Y106_CO6;
  assign CLBLM_R_X3Y106_SLICE_X2Y106_D = CLBLM_R_X3Y106_SLICE_X2Y106_DO6;
  assign CLBLM_R_X3Y106_SLICE_X2Y106_AMUX = CLBLM_R_X3Y106_SLICE_X2Y106_AO5;
  assign CLBLM_R_X3Y106_SLICE_X2Y106_BMUX = CLBLM_R_X3Y106_SLICE_X2Y106_BO5;
  assign CLBLM_R_X3Y106_SLICE_X3Y106_A = CLBLM_R_X3Y106_SLICE_X3Y106_AO6;
  assign CLBLM_R_X3Y106_SLICE_X3Y106_B = CLBLM_R_X3Y106_SLICE_X3Y106_BO6;
  assign CLBLM_R_X3Y106_SLICE_X3Y106_C = CLBLM_R_X3Y106_SLICE_X3Y106_CO6;
  assign CLBLM_R_X3Y106_SLICE_X3Y106_D = CLBLM_R_X3Y106_SLICE_X3Y106_DO6;
  assign CLBLM_R_X3Y106_SLICE_X3Y106_AMUX = CLBLM_R_X3Y106_SLICE_X3Y106_AO5;
  assign CLBLM_R_X3Y107_SLICE_X2Y107_A = CLBLM_R_X3Y107_SLICE_X2Y107_AO6;
  assign CLBLM_R_X3Y107_SLICE_X2Y107_B = CLBLM_R_X3Y107_SLICE_X2Y107_BO6;
  assign CLBLM_R_X3Y107_SLICE_X2Y107_C = CLBLM_R_X3Y107_SLICE_X2Y107_CO6;
  assign CLBLM_R_X3Y107_SLICE_X2Y107_D = CLBLM_R_X3Y107_SLICE_X2Y107_DO6;
  assign CLBLM_R_X3Y107_SLICE_X2Y107_AMUX = CLBLM_R_X3Y107_SLICE_X2Y107_AO5;
  assign CLBLM_R_X3Y107_SLICE_X3Y107_A = CLBLM_R_X3Y107_SLICE_X3Y107_AO6;
  assign CLBLM_R_X3Y107_SLICE_X3Y107_B = CLBLM_R_X3Y107_SLICE_X3Y107_BO6;
  assign CLBLM_R_X3Y107_SLICE_X3Y107_C = CLBLM_R_X3Y107_SLICE_X3Y107_CO6;
  assign CLBLM_R_X3Y107_SLICE_X3Y107_D = CLBLM_R_X3Y107_SLICE_X3Y107_DO6;
  assign CLBLM_R_X3Y107_SLICE_X3Y107_AMUX = CLBLM_R_X3Y107_SLICE_X3Y107_AO5;
  assign CLBLM_R_X3Y107_SLICE_X3Y107_BMUX = CLBLM_R_X3Y107_SLICE_X3Y107_BO5;
  assign CLBLM_R_X3Y107_SLICE_X3Y107_CMUX = CLBLM_R_X3Y107_SLICE_X3Y107_CO6;
  assign CLBLM_R_X3Y108_SLICE_X2Y108_A = CLBLM_R_X3Y108_SLICE_X2Y108_AO6;
  assign CLBLM_R_X3Y108_SLICE_X2Y108_B = CLBLM_R_X3Y108_SLICE_X2Y108_BO6;
  assign CLBLM_R_X3Y108_SLICE_X2Y108_C = CLBLM_R_X3Y108_SLICE_X2Y108_CO6;
  assign CLBLM_R_X3Y108_SLICE_X2Y108_D = CLBLM_R_X3Y108_SLICE_X2Y108_DO6;
  assign CLBLM_R_X3Y108_SLICE_X3Y108_A = CLBLM_R_X3Y108_SLICE_X3Y108_AO6;
  assign CLBLM_R_X3Y108_SLICE_X3Y108_B = CLBLM_R_X3Y108_SLICE_X3Y108_BO6;
  assign CLBLM_R_X3Y108_SLICE_X3Y108_C = CLBLM_R_X3Y108_SLICE_X3Y108_CO6;
  assign CLBLM_R_X3Y108_SLICE_X3Y108_D = CLBLM_R_X3Y108_SLICE_X3Y108_DO6;
  assign CLBLM_R_X3Y109_SLICE_X2Y109_A = CLBLM_R_X3Y109_SLICE_X2Y109_AO6;
  assign CLBLM_R_X3Y109_SLICE_X2Y109_B = CLBLM_R_X3Y109_SLICE_X2Y109_BO6;
  assign CLBLM_R_X3Y109_SLICE_X2Y109_C = CLBLM_R_X3Y109_SLICE_X2Y109_CO6;
  assign CLBLM_R_X3Y109_SLICE_X2Y109_D = CLBLM_R_X3Y109_SLICE_X2Y109_DO6;
  assign CLBLM_R_X3Y109_SLICE_X3Y109_A = CLBLM_R_X3Y109_SLICE_X3Y109_AO6;
  assign CLBLM_R_X3Y109_SLICE_X3Y109_B = CLBLM_R_X3Y109_SLICE_X3Y109_BO6;
  assign CLBLM_R_X3Y109_SLICE_X3Y109_C = CLBLM_R_X3Y109_SLICE_X3Y109_CO6;
  assign CLBLM_R_X3Y109_SLICE_X3Y109_D = CLBLM_R_X3Y109_SLICE_X3Y109_DO6;
  assign CLBLM_R_X3Y112_SLICE_X2Y112_A = CLBLM_R_X3Y112_SLICE_X2Y112_AO6;
  assign CLBLM_R_X3Y112_SLICE_X2Y112_B = CLBLM_R_X3Y112_SLICE_X2Y112_BO6;
  assign CLBLM_R_X3Y112_SLICE_X2Y112_C = CLBLM_R_X3Y112_SLICE_X2Y112_CO6;
  assign CLBLM_R_X3Y112_SLICE_X2Y112_D = CLBLM_R_X3Y112_SLICE_X2Y112_DO6;
  assign CLBLM_R_X3Y112_SLICE_X2Y112_AMUX = CLBLM_R_X3Y112_SLICE_X2Y112_AO5;
  assign CLBLM_R_X3Y112_SLICE_X2Y112_BMUX = CLBLM_R_X3Y112_SLICE_X2Y112_BO6;
  assign CLBLM_R_X3Y112_SLICE_X3Y112_A = CLBLM_R_X3Y112_SLICE_X3Y112_AO6;
  assign CLBLM_R_X3Y112_SLICE_X3Y112_B = CLBLM_R_X3Y112_SLICE_X3Y112_BO6;
  assign CLBLM_R_X3Y112_SLICE_X3Y112_C = CLBLM_R_X3Y112_SLICE_X3Y112_CO6;
  assign CLBLM_R_X3Y112_SLICE_X3Y112_D = CLBLM_R_X3Y112_SLICE_X3Y112_DO6;
  assign CLBLM_R_X3Y112_SLICE_X3Y112_AMUX = CLBLM_R_X3Y112_SLICE_X3Y112_AO5;
  assign CLBLM_R_X5Y104_SLICE_X6Y104_A = CLBLM_R_X5Y104_SLICE_X6Y104_AO6;
  assign CLBLM_R_X5Y104_SLICE_X6Y104_B = CLBLM_R_X5Y104_SLICE_X6Y104_BO6;
  assign CLBLM_R_X5Y104_SLICE_X6Y104_C = CLBLM_R_X5Y104_SLICE_X6Y104_CO6;
  assign CLBLM_R_X5Y104_SLICE_X6Y104_D = CLBLM_R_X5Y104_SLICE_X6Y104_DO6;
  assign CLBLM_R_X5Y104_SLICE_X6Y104_AMUX = CLBLM_R_X5Y104_SLICE_X6Y104_AO5;
  assign CLBLM_R_X5Y104_SLICE_X7Y104_A = CLBLM_R_X5Y104_SLICE_X7Y104_AO6;
  assign CLBLM_R_X5Y104_SLICE_X7Y104_B = CLBLM_R_X5Y104_SLICE_X7Y104_BO6;
  assign CLBLM_R_X5Y104_SLICE_X7Y104_C = CLBLM_R_X5Y104_SLICE_X7Y104_CO6;
  assign CLBLM_R_X5Y104_SLICE_X7Y104_D = CLBLM_R_X5Y104_SLICE_X7Y104_DO6;
  assign CLBLM_R_X5Y105_SLICE_X6Y105_A = CLBLM_R_X5Y105_SLICE_X6Y105_AO6;
  assign CLBLM_R_X5Y105_SLICE_X6Y105_B = CLBLM_R_X5Y105_SLICE_X6Y105_BO6;
  assign CLBLM_R_X5Y105_SLICE_X6Y105_C = CLBLM_R_X5Y105_SLICE_X6Y105_CO6;
  assign CLBLM_R_X5Y105_SLICE_X6Y105_D = CLBLM_R_X5Y105_SLICE_X6Y105_DO6;
  assign CLBLM_R_X5Y105_SLICE_X7Y105_A = CLBLM_R_X5Y105_SLICE_X7Y105_AO6;
  assign CLBLM_R_X5Y105_SLICE_X7Y105_B = CLBLM_R_X5Y105_SLICE_X7Y105_BO6;
  assign CLBLM_R_X5Y105_SLICE_X7Y105_C = CLBLM_R_X5Y105_SLICE_X7Y105_CO6;
  assign CLBLM_R_X5Y105_SLICE_X7Y105_D = CLBLM_R_X5Y105_SLICE_X7Y105_DO6;
  assign CLBLM_R_X5Y105_SLICE_X7Y105_AMUX = CLBLM_R_X5Y105_SLICE_X7Y105_AO5;
  assign CLBLM_R_X5Y106_SLICE_X6Y106_A = CLBLM_R_X5Y106_SLICE_X6Y106_AO6;
  assign CLBLM_R_X5Y106_SLICE_X6Y106_B = CLBLM_R_X5Y106_SLICE_X6Y106_BO6;
  assign CLBLM_R_X5Y106_SLICE_X6Y106_C = CLBLM_R_X5Y106_SLICE_X6Y106_CO6;
  assign CLBLM_R_X5Y106_SLICE_X6Y106_D = CLBLM_R_X5Y106_SLICE_X6Y106_DO6;
  assign CLBLM_R_X5Y106_SLICE_X6Y106_AMUX = CLBLM_R_X5Y106_SLICE_X6Y106_AO5;
  assign CLBLM_R_X5Y106_SLICE_X7Y106_A = CLBLM_R_X5Y106_SLICE_X7Y106_AO6;
  assign CLBLM_R_X5Y106_SLICE_X7Y106_B = CLBLM_R_X5Y106_SLICE_X7Y106_BO6;
  assign CLBLM_R_X5Y106_SLICE_X7Y106_C = CLBLM_R_X5Y106_SLICE_X7Y106_CO6;
  assign CLBLM_R_X5Y106_SLICE_X7Y106_D = CLBLM_R_X5Y106_SLICE_X7Y106_DO6;
  assign CLBLM_R_X5Y106_SLICE_X7Y106_AMUX = CLBLM_R_X5Y106_SLICE_X7Y106_AO5;
  assign CLBLM_R_X5Y106_SLICE_X7Y106_BMUX = CLBLM_R_X5Y106_SLICE_X7Y106_BO5;
  assign CLBLM_R_X5Y107_SLICE_X6Y107_A = CLBLM_R_X5Y107_SLICE_X6Y107_AO6;
  assign CLBLM_R_X5Y107_SLICE_X6Y107_B = CLBLM_R_X5Y107_SLICE_X6Y107_BO6;
  assign CLBLM_R_X5Y107_SLICE_X6Y107_C = CLBLM_R_X5Y107_SLICE_X6Y107_CO6;
  assign CLBLM_R_X5Y107_SLICE_X6Y107_D = CLBLM_R_X5Y107_SLICE_X6Y107_DO6;
  assign CLBLM_R_X5Y107_SLICE_X7Y107_A = CLBLM_R_X5Y107_SLICE_X7Y107_AO6;
  assign CLBLM_R_X5Y107_SLICE_X7Y107_B = CLBLM_R_X5Y107_SLICE_X7Y107_BO6;
  assign CLBLM_R_X5Y107_SLICE_X7Y107_C = CLBLM_R_X5Y107_SLICE_X7Y107_CO6;
  assign CLBLM_R_X5Y107_SLICE_X7Y107_D = CLBLM_R_X5Y107_SLICE_X7Y107_DO6;
  assign CLBLM_R_X5Y107_SLICE_X7Y107_AMUX = CLBLM_R_X5Y107_SLICE_X7Y107_AO5;
  assign CLBLM_R_X5Y108_SLICE_X6Y108_A = CLBLM_R_X5Y108_SLICE_X6Y108_AO6;
  assign CLBLM_R_X5Y108_SLICE_X6Y108_B = CLBLM_R_X5Y108_SLICE_X6Y108_BO6;
  assign CLBLM_R_X5Y108_SLICE_X6Y108_C = CLBLM_R_X5Y108_SLICE_X6Y108_CO6;
  assign CLBLM_R_X5Y108_SLICE_X6Y108_D = CLBLM_R_X5Y108_SLICE_X6Y108_DO6;
  assign CLBLM_R_X5Y108_SLICE_X6Y108_BMUX = CLBLM_R_X5Y108_SLICE_X6Y108_BO6;
  assign CLBLM_R_X5Y108_SLICE_X7Y108_A = CLBLM_R_X5Y108_SLICE_X7Y108_AO6;
  assign CLBLM_R_X5Y108_SLICE_X7Y108_B = CLBLM_R_X5Y108_SLICE_X7Y108_BO6;
  assign CLBLM_R_X5Y108_SLICE_X7Y108_C = CLBLM_R_X5Y108_SLICE_X7Y108_CO6;
  assign CLBLM_R_X5Y108_SLICE_X7Y108_D = CLBLM_R_X5Y108_SLICE_X7Y108_DO6;
  assign CLBLM_R_X5Y108_SLICE_X7Y108_AMUX = CLBLM_R_X5Y108_SLICE_X7Y108_AO5;
  assign CLBLM_R_X5Y109_SLICE_X6Y109_A = CLBLM_R_X5Y109_SLICE_X6Y109_AO6;
  assign CLBLM_R_X5Y109_SLICE_X6Y109_B = CLBLM_R_X5Y109_SLICE_X6Y109_BO6;
  assign CLBLM_R_X5Y109_SLICE_X6Y109_C = CLBLM_R_X5Y109_SLICE_X6Y109_CO6;
  assign CLBLM_R_X5Y109_SLICE_X6Y109_D = CLBLM_R_X5Y109_SLICE_X6Y109_DO6;
  assign CLBLM_R_X5Y109_SLICE_X7Y109_A = CLBLM_R_X5Y109_SLICE_X7Y109_AO6;
  assign CLBLM_R_X5Y109_SLICE_X7Y109_B = CLBLM_R_X5Y109_SLICE_X7Y109_BO6;
  assign CLBLM_R_X5Y109_SLICE_X7Y109_C = CLBLM_R_X5Y109_SLICE_X7Y109_CO6;
  assign CLBLM_R_X5Y109_SLICE_X7Y109_D = CLBLM_R_X5Y109_SLICE_X7Y109_DO6;
  assign CLBLM_R_X5Y110_SLICE_X6Y110_A = CLBLM_R_X5Y110_SLICE_X6Y110_AO6;
  assign CLBLM_R_X5Y110_SLICE_X6Y110_B = CLBLM_R_X5Y110_SLICE_X6Y110_BO6;
  assign CLBLM_R_X5Y110_SLICE_X6Y110_C = CLBLM_R_X5Y110_SLICE_X6Y110_CO6;
  assign CLBLM_R_X5Y110_SLICE_X6Y110_D = CLBLM_R_X5Y110_SLICE_X6Y110_DO6;
  assign CLBLM_R_X5Y110_SLICE_X6Y110_AMUX = CLBLM_R_X5Y110_SLICE_X6Y110_AO5;
  assign CLBLM_R_X5Y110_SLICE_X6Y110_BMUX = CLBLM_R_X5Y110_SLICE_X6Y110_BO5;
  assign CLBLM_R_X5Y110_SLICE_X7Y110_A = CLBLM_R_X5Y110_SLICE_X7Y110_AO6;
  assign CLBLM_R_X5Y110_SLICE_X7Y110_B = CLBLM_R_X5Y110_SLICE_X7Y110_BO6;
  assign CLBLM_R_X5Y110_SLICE_X7Y110_C = CLBLM_R_X5Y110_SLICE_X7Y110_CO6;
  assign CLBLM_R_X5Y110_SLICE_X7Y110_D = CLBLM_R_X5Y110_SLICE_X7Y110_DO6;
  assign CLBLM_R_X5Y110_SLICE_X7Y110_AMUX = CLBLM_R_X5Y110_SLICE_X7Y110_AO5;
  assign CLBLM_R_X5Y110_SLICE_X7Y110_BMUX = CLBLM_R_X5Y110_SLICE_X7Y110_BO5;
  assign CLBLM_R_X5Y110_SLICE_X7Y110_CMUX = CLBLM_R_X5Y110_SLICE_X7Y110_CO6;
  assign CLBLM_R_X5Y111_SLICE_X6Y111_A = CLBLM_R_X5Y111_SLICE_X6Y111_AO6;
  assign CLBLM_R_X5Y111_SLICE_X6Y111_B = CLBLM_R_X5Y111_SLICE_X6Y111_BO6;
  assign CLBLM_R_X5Y111_SLICE_X6Y111_C = CLBLM_R_X5Y111_SLICE_X6Y111_CO6;
  assign CLBLM_R_X5Y111_SLICE_X6Y111_D = CLBLM_R_X5Y111_SLICE_X6Y111_DO6;
  assign CLBLM_R_X5Y111_SLICE_X7Y111_A = CLBLM_R_X5Y111_SLICE_X7Y111_AO6;
  assign CLBLM_R_X5Y111_SLICE_X7Y111_B = CLBLM_R_X5Y111_SLICE_X7Y111_BO6;
  assign CLBLM_R_X5Y111_SLICE_X7Y111_C = CLBLM_R_X5Y111_SLICE_X7Y111_CO6;
  assign CLBLM_R_X5Y111_SLICE_X7Y111_D = CLBLM_R_X5Y111_SLICE_X7Y111_DO6;
  assign CLBLM_R_X5Y112_SLICE_X6Y112_A = CLBLM_R_X5Y112_SLICE_X6Y112_AO6;
  assign CLBLM_R_X5Y112_SLICE_X6Y112_B = CLBLM_R_X5Y112_SLICE_X6Y112_BO6;
  assign CLBLM_R_X5Y112_SLICE_X6Y112_C = CLBLM_R_X5Y112_SLICE_X6Y112_CO6;
  assign CLBLM_R_X5Y112_SLICE_X6Y112_D = CLBLM_R_X5Y112_SLICE_X6Y112_DO6;
  assign CLBLM_R_X5Y112_SLICE_X6Y112_AMUX = CLBLM_R_X5Y112_SLICE_X6Y112_AO5;
  assign CLBLM_R_X5Y112_SLICE_X6Y112_CMUX = CLBLM_R_X5Y112_SLICE_X6Y112_CO6;
  assign CLBLM_R_X5Y112_SLICE_X7Y112_A = CLBLM_R_X5Y112_SLICE_X7Y112_AO6;
  assign CLBLM_R_X5Y112_SLICE_X7Y112_B = CLBLM_R_X5Y112_SLICE_X7Y112_BO6;
  assign CLBLM_R_X5Y112_SLICE_X7Y112_C = CLBLM_R_X5Y112_SLICE_X7Y112_CO6;
  assign CLBLM_R_X5Y112_SLICE_X7Y112_D = CLBLM_R_X5Y112_SLICE_X7Y112_DO6;
  assign CLBLM_R_X5Y112_SLICE_X7Y112_AMUX = CLBLM_R_X5Y112_SLICE_X7Y112_AO5;
  assign CLBLM_R_X5Y113_SLICE_X6Y113_A = CLBLM_R_X5Y113_SLICE_X6Y113_AO6;
  assign CLBLM_R_X5Y113_SLICE_X6Y113_B = CLBLM_R_X5Y113_SLICE_X6Y113_BO6;
  assign CLBLM_R_X5Y113_SLICE_X6Y113_C = CLBLM_R_X5Y113_SLICE_X6Y113_CO6;
  assign CLBLM_R_X5Y113_SLICE_X6Y113_D = CLBLM_R_X5Y113_SLICE_X6Y113_DO6;
  assign CLBLM_R_X5Y113_SLICE_X7Y113_A = CLBLM_R_X5Y113_SLICE_X7Y113_AO6;
  assign CLBLM_R_X5Y113_SLICE_X7Y113_B = CLBLM_R_X5Y113_SLICE_X7Y113_BO6;
  assign CLBLM_R_X5Y113_SLICE_X7Y113_C = CLBLM_R_X5Y113_SLICE_X7Y113_CO6;
  assign CLBLM_R_X5Y113_SLICE_X7Y113_D = CLBLM_R_X5Y113_SLICE_X7Y113_DO6;
  assign CLBLM_R_X5Y113_SLICE_X7Y113_AMUX = CLBLM_R_X5Y113_SLICE_X7Y113_AO5;
  assign CLBLM_R_X7Y103_SLICE_X8Y103_A = CLBLM_R_X7Y103_SLICE_X8Y103_AO6;
  assign CLBLM_R_X7Y103_SLICE_X8Y103_B = CLBLM_R_X7Y103_SLICE_X8Y103_BO6;
  assign CLBLM_R_X7Y103_SLICE_X8Y103_C = CLBLM_R_X7Y103_SLICE_X8Y103_CO6;
  assign CLBLM_R_X7Y103_SLICE_X8Y103_D = CLBLM_R_X7Y103_SLICE_X8Y103_DO6;
  assign CLBLM_R_X7Y103_SLICE_X9Y103_A = CLBLM_R_X7Y103_SLICE_X9Y103_AO6;
  assign CLBLM_R_X7Y103_SLICE_X9Y103_B = CLBLM_R_X7Y103_SLICE_X9Y103_BO6;
  assign CLBLM_R_X7Y103_SLICE_X9Y103_C = CLBLM_R_X7Y103_SLICE_X9Y103_CO6;
  assign CLBLM_R_X7Y103_SLICE_X9Y103_D = CLBLM_R_X7Y103_SLICE_X9Y103_DO6;
  assign CLBLM_R_X7Y104_SLICE_X8Y104_A = CLBLM_R_X7Y104_SLICE_X8Y104_AO6;
  assign CLBLM_R_X7Y104_SLICE_X8Y104_B = CLBLM_R_X7Y104_SLICE_X8Y104_BO6;
  assign CLBLM_R_X7Y104_SLICE_X8Y104_C = CLBLM_R_X7Y104_SLICE_X8Y104_CO6;
  assign CLBLM_R_X7Y104_SLICE_X8Y104_D = CLBLM_R_X7Y104_SLICE_X8Y104_DO6;
  assign CLBLM_R_X7Y104_SLICE_X8Y104_AMUX = CLBLM_R_X7Y104_SLICE_X8Y104_AO5;
  assign CLBLM_R_X7Y104_SLICE_X8Y104_BMUX = CLBLM_R_X7Y104_SLICE_X8Y104_BO5;
  assign CLBLM_R_X7Y104_SLICE_X9Y104_A = CLBLM_R_X7Y104_SLICE_X9Y104_AO6;
  assign CLBLM_R_X7Y104_SLICE_X9Y104_B = CLBLM_R_X7Y104_SLICE_X9Y104_BO6;
  assign CLBLM_R_X7Y104_SLICE_X9Y104_C = CLBLM_R_X7Y104_SLICE_X9Y104_CO6;
  assign CLBLM_R_X7Y104_SLICE_X9Y104_D = CLBLM_R_X7Y104_SLICE_X9Y104_DO6;
  assign CLBLM_R_X7Y104_SLICE_X9Y104_AMUX = CLBLM_R_X7Y104_SLICE_X9Y104_AO5;
  assign CLBLM_R_X7Y105_SLICE_X8Y105_A = CLBLM_R_X7Y105_SLICE_X8Y105_AO6;
  assign CLBLM_R_X7Y105_SLICE_X8Y105_B = CLBLM_R_X7Y105_SLICE_X8Y105_BO6;
  assign CLBLM_R_X7Y105_SLICE_X8Y105_C = CLBLM_R_X7Y105_SLICE_X8Y105_CO6;
  assign CLBLM_R_X7Y105_SLICE_X8Y105_D = CLBLM_R_X7Y105_SLICE_X8Y105_DO6;
  assign CLBLM_R_X7Y105_SLICE_X8Y105_AMUX = CLBLM_R_X7Y105_SLICE_X8Y105_AO5;
  assign CLBLM_R_X7Y105_SLICE_X9Y105_A = CLBLM_R_X7Y105_SLICE_X9Y105_AO6;
  assign CLBLM_R_X7Y105_SLICE_X9Y105_B = CLBLM_R_X7Y105_SLICE_X9Y105_BO6;
  assign CLBLM_R_X7Y105_SLICE_X9Y105_C = CLBLM_R_X7Y105_SLICE_X9Y105_CO6;
  assign CLBLM_R_X7Y105_SLICE_X9Y105_D = CLBLM_R_X7Y105_SLICE_X9Y105_DO6;
  assign CLBLM_R_X7Y106_SLICE_X8Y106_A = CLBLM_R_X7Y106_SLICE_X8Y106_AO6;
  assign CLBLM_R_X7Y106_SLICE_X8Y106_B = CLBLM_R_X7Y106_SLICE_X8Y106_BO6;
  assign CLBLM_R_X7Y106_SLICE_X8Y106_C = CLBLM_R_X7Y106_SLICE_X8Y106_CO6;
  assign CLBLM_R_X7Y106_SLICE_X8Y106_D = CLBLM_R_X7Y106_SLICE_X8Y106_DO6;
  assign CLBLM_R_X7Y106_SLICE_X8Y106_AMUX = CLBLM_R_X7Y106_SLICE_X8Y106_AO5;
  assign CLBLM_R_X7Y106_SLICE_X8Y106_CMUX = CLBLM_R_X7Y106_SLICE_X8Y106_CO6;
  assign CLBLM_R_X7Y106_SLICE_X9Y106_A = CLBLM_R_X7Y106_SLICE_X9Y106_AO6;
  assign CLBLM_R_X7Y106_SLICE_X9Y106_B = CLBLM_R_X7Y106_SLICE_X9Y106_BO6;
  assign CLBLM_R_X7Y106_SLICE_X9Y106_C = CLBLM_R_X7Y106_SLICE_X9Y106_CO6;
  assign CLBLM_R_X7Y106_SLICE_X9Y106_D = CLBLM_R_X7Y106_SLICE_X9Y106_DO6;
  assign CLBLM_R_X7Y107_SLICE_X8Y107_A = CLBLM_R_X7Y107_SLICE_X8Y107_AO6;
  assign CLBLM_R_X7Y107_SLICE_X8Y107_B = CLBLM_R_X7Y107_SLICE_X8Y107_BO6;
  assign CLBLM_R_X7Y107_SLICE_X8Y107_C = CLBLM_R_X7Y107_SLICE_X8Y107_CO6;
  assign CLBLM_R_X7Y107_SLICE_X8Y107_D = CLBLM_R_X7Y107_SLICE_X8Y107_DO6;
  assign CLBLM_R_X7Y107_SLICE_X8Y107_AMUX = CLBLM_R_X7Y107_SLICE_X8Y107_AO6;
  assign CLBLM_R_X7Y107_SLICE_X9Y107_A = CLBLM_R_X7Y107_SLICE_X9Y107_AO6;
  assign CLBLM_R_X7Y107_SLICE_X9Y107_B = CLBLM_R_X7Y107_SLICE_X9Y107_BO6;
  assign CLBLM_R_X7Y107_SLICE_X9Y107_C = CLBLM_R_X7Y107_SLICE_X9Y107_CO6;
  assign CLBLM_R_X7Y107_SLICE_X9Y107_D = CLBLM_R_X7Y107_SLICE_X9Y107_DO6;
  assign CLBLM_R_X7Y107_SLICE_X9Y107_BMUX = CLBLM_R_X7Y107_SLICE_X9Y107_BO6;
  assign CLBLM_R_X7Y107_SLICE_X9Y107_CMUX = CLBLM_R_X7Y107_SLICE_X9Y107_CO6;
  assign CLBLM_R_X7Y108_SLICE_X8Y108_A = CLBLM_R_X7Y108_SLICE_X8Y108_AO6;
  assign CLBLM_R_X7Y108_SLICE_X8Y108_B = CLBLM_R_X7Y108_SLICE_X8Y108_BO6;
  assign CLBLM_R_X7Y108_SLICE_X8Y108_C = CLBLM_R_X7Y108_SLICE_X8Y108_CO6;
  assign CLBLM_R_X7Y108_SLICE_X8Y108_D = CLBLM_R_X7Y108_SLICE_X8Y108_DO6;
  assign CLBLM_R_X7Y108_SLICE_X8Y108_AMUX = CLBLM_R_X7Y108_SLICE_X8Y108_AO5;
  assign CLBLM_R_X7Y108_SLICE_X9Y108_A = CLBLM_R_X7Y108_SLICE_X9Y108_AO6;
  assign CLBLM_R_X7Y108_SLICE_X9Y108_B = CLBLM_R_X7Y108_SLICE_X9Y108_BO6;
  assign CLBLM_R_X7Y108_SLICE_X9Y108_C = CLBLM_R_X7Y108_SLICE_X9Y108_CO6;
  assign CLBLM_R_X7Y108_SLICE_X9Y108_D = CLBLM_R_X7Y108_SLICE_X9Y108_DO6;
  assign CLBLM_R_X7Y108_SLICE_X9Y108_BMUX = CLBLM_R_X7Y108_SLICE_X9Y108_BO6;
  assign CLBLM_R_X7Y109_SLICE_X8Y109_A = CLBLM_R_X7Y109_SLICE_X8Y109_AO6;
  assign CLBLM_R_X7Y109_SLICE_X8Y109_B = CLBLM_R_X7Y109_SLICE_X8Y109_BO6;
  assign CLBLM_R_X7Y109_SLICE_X8Y109_C = CLBLM_R_X7Y109_SLICE_X8Y109_CO6;
  assign CLBLM_R_X7Y109_SLICE_X8Y109_D = CLBLM_R_X7Y109_SLICE_X8Y109_DO6;
  assign CLBLM_R_X7Y109_SLICE_X8Y109_AMUX = CLBLM_R_X7Y109_SLICE_X8Y109_AO5;
  assign CLBLM_R_X7Y109_SLICE_X9Y109_A = CLBLM_R_X7Y109_SLICE_X9Y109_AO6;
  assign CLBLM_R_X7Y109_SLICE_X9Y109_B = CLBLM_R_X7Y109_SLICE_X9Y109_BO6;
  assign CLBLM_R_X7Y109_SLICE_X9Y109_C = CLBLM_R_X7Y109_SLICE_X9Y109_CO6;
  assign CLBLM_R_X7Y109_SLICE_X9Y109_D = CLBLM_R_X7Y109_SLICE_X9Y109_DO6;
  assign CLBLM_R_X7Y109_SLICE_X9Y109_AMUX = CLBLM_R_X7Y109_SLICE_X9Y109_AO5;
  assign CLBLM_R_X7Y110_SLICE_X8Y110_A = CLBLM_R_X7Y110_SLICE_X8Y110_AO6;
  assign CLBLM_R_X7Y110_SLICE_X8Y110_B = CLBLM_R_X7Y110_SLICE_X8Y110_BO6;
  assign CLBLM_R_X7Y110_SLICE_X8Y110_C = CLBLM_R_X7Y110_SLICE_X8Y110_CO6;
  assign CLBLM_R_X7Y110_SLICE_X8Y110_D = CLBLM_R_X7Y110_SLICE_X8Y110_DO6;
  assign CLBLM_R_X7Y110_SLICE_X8Y110_BMUX = CLBLM_R_X7Y110_SLICE_X8Y110_BO6;
  assign CLBLM_R_X7Y110_SLICE_X9Y110_A = CLBLM_R_X7Y110_SLICE_X9Y110_AO6;
  assign CLBLM_R_X7Y110_SLICE_X9Y110_B = CLBLM_R_X7Y110_SLICE_X9Y110_BO6;
  assign CLBLM_R_X7Y110_SLICE_X9Y110_C = CLBLM_R_X7Y110_SLICE_X9Y110_CO6;
  assign CLBLM_R_X7Y110_SLICE_X9Y110_D = CLBLM_R_X7Y110_SLICE_X9Y110_DO6;
  assign CLBLM_R_X7Y110_SLICE_X9Y110_AMUX = CLBLM_R_X7Y110_SLICE_X9Y110_AO5;
  assign CLBLM_R_X7Y110_SLICE_X9Y110_BMUX = CLBLM_R_X7Y110_SLICE_X9Y110_BO5;
  assign CLBLM_R_X7Y110_SLICE_X9Y110_CMUX = CLBLM_R_X7Y110_SLICE_X9Y110_CO6;
  assign CLBLM_R_X7Y111_SLICE_X8Y111_A = CLBLM_R_X7Y111_SLICE_X8Y111_AO6;
  assign CLBLM_R_X7Y111_SLICE_X8Y111_B = CLBLM_R_X7Y111_SLICE_X8Y111_BO6;
  assign CLBLM_R_X7Y111_SLICE_X8Y111_C = CLBLM_R_X7Y111_SLICE_X8Y111_CO6;
  assign CLBLM_R_X7Y111_SLICE_X8Y111_D = CLBLM_R_X7Y111_SLICE_X8Y111_DO6;
  assign CLBLM_R_X7Y111_SLICE_X8Y111_AMUX = CLBLM_R_X7Y111_SLICE_X8Y111_AO5;
  assign CLBLM_R_X7Y111_SLICE_X9Y111_A = CLBLM_R_X7Y111_SLICE_X9Y111_AO6;
  assign CLBLM_R_X7Y111_SLICE_X9Y111_B = CLBLM_R_X7Y111_SLICE_X9Y111_BO6;
  assign CLBLM_R_X7Y111_SLICE_X9Y111_C = CLBLM_R_X7Y111_SLICE_X9Y111_CO6;
  assign CLBLM_R_X7Y111_SLICE_X9Y111_D = CLBLM_R_X7Y111_SLICE_X9Y111_DO6;
  assign CLBLM_R_X7Y111_SLICE_X9Y111_AMUX = CLBLM_R_X7Y111_SLICE_X9Y111_AO5;
  assign CLBLM_R_X7Y112_SLICE_X8Y112_A = CLBLM_R_X7Y112_SLICE_X8Y112_AO6;
  assign CLBLM_R_X7Y112_SLICE_X8Y112_B = CLBLM_R_X7Y112_SLICE_X8Y112_BO6;
  assign CLBLM_R_X7Y112_SLICE_X8Y112_C = CLBLM_R_X7Y112_SLICE_X8Y112_CO6;
  assign CLBLM_R_X7Y112_SLICE_X8Y112_D = CLBLM_R_X7Y112_SLICE_X8Y112_DO6;
  assign CLBLM_R_X7Y112_SLICE_X8Y112_AMUX = CLBLM_R_X7Y112_SLICE_X8Y112_AO5;
  assign CLBLM_R_X7Y112_SLICE_X9Y112_A = CLBLM_R_X7Y112_SLICE_X9Y112_AO6;
  assign CLBLM_R_X7Y112_SLICE_X9Y112_B = CLBLM_R_X7Y112_SLICE_X9Y112_BO6;
  assign CLBLM_R_X7Y112_SLICE_X9Y112_C = CLBLM_R_X7Y112_SLICE_X9Y112_CO6;
  assign CLBLM_R_X7Y112_SLICE_X9Y112_D = CLBLM_R_X7Y112_SLICE_X9Y112_DO6;
  assign CLBLM_R_X7Y113_SLICE_X8Y113_A = CLBLM_R_X7Y113_SLICE_X8Y113_AO6;
  assign CLBLM_R_X7Y113_SLICE_X8Y113_B = CLBLM_R_X7Y113_SLICE_X8Y113_BO6;
  assign CLBLM_R_X7Y113_SLICE_X8Y113_C = CLBLM_R_X7Y113_SLICE_X8Y113_CO6;
  assign CLBLM_R_X7Y113_SLICE_X8Y113_D = CLBLM_R_X7Y113_SLICE_X8Y113_DO6;
  assign CLBLM_R_X7Y113_SLICE_X8Y113_AMUX = CLBLM_R_X7Y113_SLICE_X8Y113_AO5;
  assign CLBLM_R_X7Y113_SLICE_X8Y113_BMUX = CLBLM_R_X7Y113_SLICE_X8Y113_BO5;
  assign CLBLM_R_X7Y113_SLICE_X9Y113_A = CLBLM_R_X7Y113_SLICE_X9Y113_AO6;
  assign CLBLM_R_X7Y113_SLICE_X9Y113_B = CLBLM_R_X7Y113_SLICE_X9Y113_BO6;
  assign CLBLM_R_X7Y113_SLICE_X9Y113_C = CLBLM_R_X7Y113_SLICE_X9Y113_CO6;
  assign CLBLM_R_X7Y113_SLICE_X9Y113_D = CLBLM_R_X7Y113_SLICE_X9Y113_DO6;
  assign CLBLM_R_X7Y114_SLICE_X8Y114_A = CLBLM_R_X7Y114_SLICE_X8Y114_AO6;
  assign CLBLM_R_X7Y114_SLICE_X8Y114_B = CLBLM_R_X7Y114_SLICE_X8Y114_BO6;
  assign CLBLM_R_X7Y114_SLICE_X8Y114_C = CLBLM_R_X7Y114_SLICE_X8Y114_CO6;
  assign CLBLM_R_X7Y114_SLICE_X8Y114_D = CLBLM_R_X7Y114_SLICE_X8Y114_DO6;
  assign CLBLM_R_X7Y114_SLICE_X8Y114_AMUX = CLBLM_R_X7Y114_SLICE_X8Y114_AO5;
  assign CLBLM_R_X7Y114_SLICE_X9Y114_A = CLBLM_R_X7Y114_SLICE_X9Y114_AO6;
  assign CLBLM_R_X7Y114_SLICE_X9Y114_B = CLBLM_R_X7Y114_SLICE_X9Y114_BO6;
  assign CLBLM_R_X7Y114_SLICE_X9Y114_C = CLBLM_R_X7Y114_SLICE_X9Y114_CO6;
  assign CLBLM_R_X7Y114_SLICE_X9Y114_D = CLBLM_R_X7Y114_SLICE_X9Y114_DO6;
  assign CLBLM_R_X11Y104_SLICE_X14Y104_A = CLBLM_R_X11Y104_SLICE_X14Y104_AO6;
  assign CLBLM_R_X11Y104_SLICE_X14Y104_B = CLBLM_R_X11Y104_SLICE_X14Y104_BO6;
  assign CLBLM_R_X11Y104_SLICE_X14Y104_C = CLBLM_R_X11Y104_SLICE_X14Y104_CO6;
  assign CLBLM_R_X11Y104_SLICE_X14Y104_D = CLBLM_R_X11Y104_SLICE_X14Y104_DO6;
  assign CLBLM_R_X11Y104_SLICE_X14Y104_AMUX = CLBLM_R_X11Y104_SLICE_X14Y104_AO5;
  assign CLBLM_R_X11Y104_SLICE_X15Y104_A = CLBLM_R_X11Y104_SLICE_X15Y104_AO6;
  assign CLBLM_R_X11Y104_SLICE_X15Y104_B = CLBLM_R_X11Y104_SLICE_X15Y104_BO6;
  assign CLBLM_R_X11Y104_SLICE_X15Y104_C = CLBLM_R_X11Y104_SLICE_X15Y104_CO6;
  assign CLBLM_R_X11Y104_SLICE_X15Y104_D = CLBLM_R_X11Y104_SLICE_X15Y104_DO6;
  assign CLBLM_R_X11Y104_SLICE_X15Y104_AMUX = CLBLM_R_X11Y104_SLICE_X15Y104_AO5;
  assign CLBLM_R_X11Y104_SLICE_X15Y104_BMUX = CLBLM_R_X11Y104_SLICE_X15Y104_BO6;
  assign CLBLM_R_X11Y105_SLICE_X14Y105_A = CLBLM_R_X11Y105_SLICE_X14Y105_AO6;
  assign CLBLM_R_X11Y105_SLICE_X14Y105_B = CLBLM_R_X11Y105_SLICE_X14Y105_BO6;
  assign CLBLM_R_X11Y105_SLICE_X14Y105_C = CLBLM_R_X11Y105_SLICE_X14Y105_CO6;
  assign CLBLM_R_X11Y105_SLICE_X14Y105_D = CLBLM_R_X11Y105_SLICE_X14Y105_DO6;
  assign CLBLM_R_X11Y105_SLICE_X14Y105_AMUX = CLBLM_R_X11Y105_SLICE_X14Y105_AO5;
  assign CLBLM_R_X11Y105_SLICE_X15Y105_A = CLBLM_R_X11Y105_SLICE_X15Y105_AO6;
  assign CLBLM_R_X11Y105_SLICE_X15Y105_B = CLBLM_R_X11Y105_SLICE_X15Y105_BO6;
  assign CLBLM_R_X11Y105_SLICE_X15Y105_C = CLBLM_R_X11Y105_SLICE_X15Y105_CO6;
  assign CLBLM_R_X11Y105_SLICE_X15Y105_D = CLBLM_R_X11Y105_SLICE_X15Y105_DO6;
  assign CLBLM_R_X11Y105_SLICE_X15Y105_AMUX = CLBLM_R_X11Y105_SLICE_X15Y105_AO5;
  assign CLBLM_R_X11Y106_SLICE_X14Y106_A = CLBLM_R_X11Y106_SLICE_X14Y106_AO6;
  assign CLBLM_R_X11Y106_SLICE_X14Y106_B = CLBLM_R_X11Y106_SLICE_X14Y106_BO6;
  assign CLBLM_R_X11Y106_SLICE_X14Y106_C = CLBLM_R_X11Y106_SLICE_X14Y106_CO6;
  assign CLBLM_R_X11Y106_SLICE_X14Y106_D = CLBLM_R_X11Y106_SLICE_X14Y106_DO6;
  assign CLBLM_R_X11Y106_SLICE_X14Y106_BMUX = CLBLM_R_X11Y106_SLICE_X14Y106_BO6;
  assign CLBLM_R_X11Y106_SLICE_X15Y106_A = CLBLM_R_X11Y106_SLICE_X15Y106_AO6;
  assign CLBLM_R_X11Y106_SLICE_X15Y106_B = CLBLM_R_X11Y106_SLICE_X15Y106_BO6;
  assign CLBLM_R_X11Y106_SLICE_X15Y106_C = CLBLM_R_X11Y106_SLICE_X15Y106_CO6;
  assign CLBLM_R_X11Y106_SLICE_X15Y106_D = CLBLM_R_X11Y106_SLICE_X15Y106_DO6;
  assign CLBLM_R_X11Y106_SLICE_X15Y106_AMUX = CLBLM_R_X11Y106_SLICE_X15Y106_AO5;
  assign CLBLM_R_X11Y107_SLICE_X14Y107_A = CLBLM_R_X11Y107_SLICE_X14Y107_AO6;
  assign CLBLM_R_X11Y107_SLICE_X14Y107_B = CLBLM_R_X11Y107_SLICE_X14Y107_BO6;
  assign CLBLM_R_X11Y107_SLICE_X14Y107_C = CLBLM_R_X11Y107_SLICE_X14Y107_CO6;
  assign CLBLM_R_X11Y107_SLICE_X14Y107_D = CLBLM_R_X11Y107_SLICE_X14Y107_DO6;
  assign CLBLM_R_X11Y107_SLICE_X14Y107_AMUX = CLBLM_R_X11Y107_SLICE_X14Y107_AO5;
  assign CLBLM_R_X11Y107_SLICE_X14Y107_BMUX = CLBLM_R_X11Y107_SLICE_X14Y107_BO5;
  assign CLBLM_R_X11Y107_SLICE_X14Y107_CMUX = CLBLM_R_X11Y107_SLICE_X14Y107_CO6;
  assign CLBLM_R_X11Y107_SLICE_X14Y107_DMUX = CLBLM_R_X11Y107_SLICE_X14Y107_DO6;
  assign CLBLM_R_X11Y107_SLICE_X15Y107_A = CLBLM_R_X11Y107_SLICE_X15Y107_AO6;
  assign CLBLM_R_X11Y107_SLICE_X15Y107_B = CLBLM_R_X11Y107_SLICE_X15Y107_BO6;
  assign CLBLM_R_X11Y107_SLICE_X15Y107_C = CLBLM_R_X11Y107_SLICE_X15Y107_CO6;
  assign CLBLM_R_X11Y107_SLICE_X15Y107_D = CLBLM_R_X11Y107_SLICE_X15Y107_DO6;
  assign CLBLM_R_X11Y107_SLICE_X15Y107_AMUX = CLBLM_R_X11Y107_SLICE_X15Y107_AO5;
  assign CLBLM_R_X11Y108_SLICE_X14Y108_A = CLBLM_R_X11Y108_SLICE_X14Y108_AO6;
  assign CLBLM_R_X11Y108_SLICE_X14Y108_B = CLBLM_R_X11Y108_SLICE_X14Y108_BO6;
  assign CLBLM_R_X11Y108_SLICE_X14Y108_C = CLBLM_R_X11Y108_SLICE_X14Y108_CO6;
  assign CLBLM_R_X11Y108_SLICE_X14Y108_D = CLBLM_R_X11Y108_SLICE_X14Y108_DO6;
  assign CLBLM_R_X11Y108_SLICE_X15Y108_A = CLBLM_R_X11Y108_SLICE_X15Y108_AO6;
  assign CLBLM_R_X11Y108_SLICE_X15Y108_B = CLBLM_R_X11Y108_SLICE_X15Y108_BO6;
  assign CLBLM_R_X11Y108_SLICE_X15Y108_C = CLBLM_R_X11Y108_SLICE_X15Y108_CO6;
  assign CLBLM_R_X11Y108_SLICE_X15Y108_D = CLBLM_R_X11Y108_SLICE_X15Y108_DO6;
  assign CLBLM_R_X11Y108_SLICE_X15Y108_CMUX = CLBLM_R_X11Y108_SLICE_X15Y108_CO6;
  assign CLBLM_R_X11Y109_SLICE_X14Y109_A = CLBLM_R_X11Y109_SLICE_X14Y109_AO6;
  assign CLBLM_R_X11Y109_SLICE_X14Y109_B = CLBLM_R_X11Y109_SLICE_X14Y109_BO6;
  assign CLBLM_R_X11Y109_SLICE_X14Y109_C = CLBLM_R_X11Y109_SLICE_X14Y109_CO6;
  assign CLBLM_R_X11Y109_SLICE_X14Y109_D = CLBLM_R_X11Y109_SLICE_X14Y109_DO6;
  assign CLBLM_R_X11Y109_SLICE_X14Y109_AMUX = CLBLM_R_X11Y109_SLICE_X14Y109_AO5;
  assign CLBLM_R_X11Y109_SLICE_X15Y109_A = CLBLM_R_X11Y109_SLICE_X15Y109_AO6;
  assign CLBLM_R_X11Y109_SLICE_X15Y109_B = CLBLM_R_X11Y109_SLICE_X15Y109_BO6;
  assign CLBLM_R_X11Y109_SLICE_X15Y109_C = CLBLM_R_X11Y109_SLICE_X15Y109_CO6;
  assign CLBLM_R_X11Y109_SLICE_X15Y109_D = CLBLM_R_X11Y109_SLICE_X15Y109_DO6;
  assign CLBLM_R_X11Y109_SLICE_X15Y109_BMUX = CLBLM_R_X11Y109_SLICE_X15Y109_BO6;
  assign CLBLM_R_X11Y110_SLICE_X14Y110_A = CLBLM_R_X11Y110_SLICE_X14Y110_AO6;
  assign CLBLM_R_X11Y110_SLICE_X14Y110_B = CLBLM_R_X11Y110_SLICE_X14Y110_BO6;
  assign CLBLM_R_X11Y110_SLICE_X14Y110_C = CLBLM_R_X11Y110_SLICE_X14Y110_CO6;
  assign CLBLM_R_X11Y110_SLICE_X14Y110_D = CLBLM_R_X11Y110_SLICE_X14Y110_DO6;
  assign CLBLM_R_X11Y110_SLICE_X14Y110_AMUX = CLBLM_R_X11Y110_SLICE_X14Y110_AO5;
  assign CLBLM_R_X11Y110_SLICE_X15Y110_A = CLBLM_R_X11Y110_SLICE_X15Y110_AO6;
  assign CLBLM_R_X11Y110_SLICE_X15Y110_B = CLBLM_R_X11Y110_SLICE_X15Y110_BO6;
  assign CLBLM_R_X11Y110_SLICE_X15Y110_C = CLBLM_R_X11Y110_SLICE_X15Y110_CO6;
  assign CLBLM_R_X11Y110_SLICE_X15Y110_D = CLBLM_R_X11Y110_SLICE_X15Y110_DO6;
  assign CLBLM_R_X11Y110_SLICE_X15Y110_AMUX = CLBLM_R_X11Y110_SLICE_X15Y110_AO5;
  assign CLBLM_R_X11Y110_SLICE_X15Y110_BMUX = CLBLM_R_X11Y110_SLICE_X15Y110_BO6;
  assign CLBLM_R_X11Y111_SLICE_X14Y111_A = CLBLM_R_X11Y111_SLICE_X14Y111_AO6;
  assign CLBLM_R_X11Y111_SLICE_X14Y111_B = CLBLM_R_X11Y111_SLICE_X14Y111_BO6;
  assign CLBLM_R_X11Y111_SLICE_X14Y111_C = CLBLM_R_X11Y111_SLICE_X14Y111_CO6;
  assign CLBLM_R_X11Y111_SLICE_X14Y111_D = CLBLM_R_X11Y111_SLICE_X14Y111_DO6;
  assign CLBLM_R_X11Y111_SLICE_X14Y111_AMUX = CLBLM_R_X11Y111_SLICE_X14Y111_AO5;
  assign CLBLM_R_X11Y111_SLICE_X14Y111_BMUX = CLBLM_R_X11Y111_SLICE_X14Y111_BO5;
  assign CLBLM_R_X11Y111_SLICE_X15Y111_A = CLBLM_R_X11Y111_SLICE_X15Y111_AO6;
  assign CLBLM_R_X11Y111_SLICE_X15Y111_B = CLBLM_R_X11Y111_SLICE_X15Y111_BO6;
  assign CLBLM_R_X11Y111_SLICE_X15Y111_C = CLBLM_R_X11Y111_SLICE_X15Y111_CO6;
  assign CLBLM_R_X11Y111_SLICE_X15Y111_D = CLBLM_R_X11Y111_SLICE_X15Y111_DO6;
  assign CLBLM_R_X11Y111_SLICE_X15Y111_AMUX = CLBLM_R_X11Y111_SLICE_X15Y111_AO5;
  assign CLBLM_R_X11Y111_SLICE_X15Y111_BMUX = CLBLM_R_X11Y111_SLICE_X15Y111_BO5;
  assign CLBLM_R_X13Y105_SLICE_X18Y105_A = CLBLM_R_X13Y105_SLICE_X18Y105_AO6;
  assign CLBLM_R_X13Y105_SLICE_X18Y105_B = CLBLM_R_X13Y105_SLICE_X18Y105_BO6;
  assign CLBLM_R_X13Y105_SLICE_X18Y105_C = CLBLM_R_X13Y105_SLICE_X18Y105_CO6;
  assign CLBLM_R_X13Y105_SLICE_X18Y105_D = CLBLM_R_X13Y105_SLICE_X18Y105_DO6;
  assign CLBLM_R_X13Y105_SLICE_X19Y105_A = CLBLM_R_X13Y105_SLICE_X19Y105_AO6;
  assign CLBLM_R_X13Y105_SLICE_X19Y105_B = CLBLM_R_X13Y105_SLICE_X19Y105_BO6;
  assign CLBLM_R_X13Y105_SLICE_X19Y105_C = CLBLM_R_X13Y105_SLICE_X19Y105_CO6;
  assign CLBLM_R_X13Y105_SLICE_X19Y105_D = CLBLM_R_X13Y105_SLICE_X19Y105_DO6;
  assign CLBLM_R_X13Y106_SLICE_X18Y106_A = CLBLM_R_X13Y106_SLICE_X18Y106_AO6;
  assign CLBLM_R_X13Y106_SLICE_X18Y106_B = CLBLM_R_X13Y106_SLICE_X18Y106_BO6;
  assign CLBLM_R_X13Y106_SLICE_X18Y106_C = CLBLM_R_X13Y106_SLICE_X18Y106_CO6;
  assign CLBLM_R_X13Y106_SLICE_X18Y106_D = CLBLM_R_X13Y106_SLICE_X18Y106_DO6;
  assign CLBLM_R_X13Y106_SLICE_X18Y106_AMUX = CLBLM_R_X13Y106_SLICE_X18Y106_AO5;
  assign CLBLM_R_X13Y106_SLICE_X19Y106_A = CLBLM_R_X13Y106_SLICE_X19Y106_AO6;
  assign CLBLM_R_X13Y106_SLICE_X19Y106_B = CLBLM_R_X13Y106_SLICE_X19Y106_BO6;
  assign CLBLM_R_X13Y106_SLICE_X19Y106_C = CLBLM_R_X13Y106_SLICE_X19Y106_CO6;
  assign CLBLM_R_X13Y106_SLICE_X19Y106_D = CLBLM_R_X13Y106_SLICE_X19Y106_DO6;
  assign CLBLM_R_X13Y106_SLICE_X19Y106_AMUX = CLBLM_R_X13Y106_SLICE_X19Y106_AO5;
  assign CLBLM_R_X13Y106_SLICE_X19Y106_BMUX = CLBLM_R_X13Y106_SLICE_X19Y106_BO6;
  assign CLBLM_R_X13Y106_SLICE_X19Y106_CMUX = CLBLM_R_X13Y106_SLICE_X19Y106_CO6;
  assign CLBLM_R_X13Y107_SLICE_X18Y107_A = CLBLM_R_X13Y107_SLICE_X18Y107_AO6;
  assign CLBLM_R_X13Y107_SLICE_X18Y107_B = CLBLM_R_X13Y107_SLICE_X18Y107_BO6;
  assign CLBLM_R_X13Y107_SLICE_X18Y107_C = CLBLM_R_X13Y107_SLICE_X18Y107_CO6;
  assign CLBLM_R_X13Y107_SLICE_X18Y107_D = CLBLM_R_X13Y107_SLICE_X18Y107_DO6;
  assign CLBLM_R_X13Y107_SLICE_X19Y107_A = CLBLM_R_X13Y107_SLICE_X19Y107_AO6;
  assign CLBLM_R_X13Y107_SLICE_X19Y107_B = CLBLM_R_X13Y107_SLICE_X19Y107_BO6;
  assign CLBLM_R_X13Y107_SLICE_X19Y107_C = CLBLM_R_X13Y107_SLICE_X19Y107_CO6;
  assign CLBLM_R_X13Y107_SLICE_X19Y107_D = CLBLM_R_X13Y107_SLICE_X19Y107_DO6;
  assign LIOI3_X0Y101_ILOGIC_X0Y102_O = LIOB33_X0Y101_IOB_X0Y102_I;
  assign LIOI3_X0Y101_ILOGIC_X0Y101_O = LIOB33_X0Y101_IOB_X0Y101_I;
  assign LIOI3_X0Y103_ILOGIC_X0Y104_O = LIOB33_X0Y103_IOB_X0Y104_I;
  assign LIOI3_X0Y103_ILOGIC_X0Y103_O = LIOB33_X0Y103_IOB_X0Y103_I;
  assign LIOI3_X0Y105_ILOGIC_X0Y106_O = LIOB33_X0Y105_IOB_X0Y106_I;
  assign LIOI3_X0Y105_ILOGIC_X0Y105_O = LIOB33_X0Y105_IOB_X0Y105_I;
  assign LIOI3_X0Y109_ILOGIC_X0Y110_O = LIOB33_X0Y109_IOB_X0Y110_I;
  assign LIOI3_X0Y109_ILOGIC_X0Y109_O = LIOB33_X0Y109_IOB_X0Y109_I;
  assign LIOI3_X0Y111_ILOGIC_X0Y112_O = LIOB33_X0Y111_IOB_X0Y112_I;
  assign LIOI3_X0Y111_ILOGIC_X0Y111_O = LIOB33_X0Y111_IOB_X0Y111_I;
  assign LIOI3_X0Y115_ILOGIC_X0Y116_O = LIOB33_X0Y115_IOB_X0Y116_I;
  assign LIOI3_X0Y115_ILOGIC_X0Y115_O = LIOB33_X0Y115_IOB_X0Y115_I;
  assign LIOI3_X0Y117_ILOGIC_X0Y117_O = LIOB33_X0Y117_IOB_X0Y117_I;
  assign LIOI3_X0Y117_OLOGIC_X0Y118_OQ = CLBLL_L_X2Y109_SLICE_X0Y109_AO5;
  assign LIOI3_X0Y117_OLOGIC_X0Y118_TQ = 1'b1;
  assign LIOI3_X0Y121_OLOGIC_X0Y122_OQ = CLBLL_L_X2Y104_SLICE_X0Y104_AO6;
  assign LIOI3_X0Y121_OLOGIC_X0Y122_TQ = 1'b1;
  assign LIOI3_X0Y121_OLOGIC_X0Y121_OQ = CLBLL_L_X2Y106_SLICE_X0Y106_AO5;
  assign LIOI3_X0Y121_OLOGIC_X0Y121_TQ = 1'b1;
  assign LIOI3_X0Y123_OLOGIC_X0Y124_OQ = CLBLM_R_X3Y107_SLICE_X2Y107_AO6;
  assign LIOI3_X0Y123_OLOGIC_X0Y124_TQ = 1'b1;
  assign LIOI3_X0Y123_OLOGIC_X0Y123_OQ = CLBLL_L_X2Y107_SLICE_X0Y107_AO6;
  assign LIOI3_X0Y123_OLOGIC_X0Y123_TQ = 1'b1;
  assign LIOI3_X0Y125_OLOGIC_X0Y126_OQ = CLBLM_R_X3Y107_SLICE_X2Y107_CO6;
  assign LIOI3_X0Y125_OLOGIC_X0Y126_TQ = 1'b1;
  assign LIOI3_X0Y125_OLOGIC_X0Y125_OQ = CLBLM_R_X7Y109_SLICE_X9Y109_AO5;
  assign LIOI3_X0Y125_OLOGIC_X0Y125_TQ = 1'b1;
  assign LIOI3_X0Y127_OLOGIC_X0Y128_OQ = CLBLM_R_X3Y107_SLICE_X3Y107_BO6;
  assign LIOI3_X0Y127_OLOGIC_X0Y128_TQ = 1'b1;
  assign LIOI3_X0Y127_OLOGIC_X0Y127_OQ = CLBLM_R_X3Y107_SLICE_X3Y107_AO6;
  assign LIOI3_X0Y127_OLOGIC_X0Y127_TQ = 1'b1;
  assign LIOI3_X0Y129_OLOGIC_X0Y130_OQ = CLBLL_L_X2Y110_SLICE_X0Y110_AO6;
  assign LIOI3_X0Y129_OLOGIC_X0Y130_TQ = 1'b1;
  assign LIOI3_X0Y129_OLOGIC_X0Y129_OQ = CLBLM_R_X3Y108_SLICE_X3Y108_AO6;
  assign LIOI3_X0Y129_OLOGIC_X0Y129_TQ = 1'b1;
  assign LIOI3_X0Y133_OLOGIC_X0Y134_OQ = 1'b0;
  assign LIOI3_X0Y133_OLOGIC_X0Y134_TQ = 1'b1;
  assign LIOI3_X0Y133_OLOGIC_X0Y133_OQ = CLBLM_R_X3Y109_SLICE_X3Y109_AO6;
  assign LIOI3_X0Y133_OLOGIC_X0Y133_TQ = 1'b1;
  assign LIOI3_X0Y135_OLOGIC_X0Y136_OQ = CLBLL_L_X4Y110_SLICE_X5Y110_AO5;
  assign LIOI3_X0Y135_OLOGIC_X0Y136_TQ = 1'b1;
  assign LIOI3_X0Y135_OLOGIC_X0Y135_OQ = CLBLL_L_X4Y110_SLICE_X5Y110_AO6;
  assign LIOI3_X0Y135_OLOGIC_X0Y135_TQ = 1'b1;
  assign LIOI3_X0Y139_OLOGIC_X0Y140_OQ = CLBLL_L_X4Y112_SLICE_X4Y112_AO5;
  assign LIOI3_X0Y139_OLOGIC_X0Y140_TQ = 1'b1;
  assign LIOI3_X0Y139_OLOGIC_X0Y139_OQ = CLBLL_L_X4Y112_SLICE_X4Y112_AO6;
  assign LIOI3_X0Y139_OLOGIC_X0Y139_TQ = 1'b1;
  assign LIOI3_X0Y141_OLOGIC_X0Y142_OQ = CLBLL_L_X4Y114_SLICE_X4Y114_DO6;
  assign LIOI3_X0Y141_OLOGIC_X0Y142_TQ = 1'b1;
  assign LIOI3_X0Y141_OLOGIC_X0Y141_OQ = CLBLL_L_X4Y112_SLICE_X5Y112_DO6;
  assign LIOI3_X0Y141_OLOGIC_X0Y141_TQ = 1'b1;
  assign LIOI3_X0Y145_OLOGIC_X0Y146_OQ = CLBLL_L_X4Y115_SLICE_X4Y115_CO6;
  assign LIOI3_X0Y145_OLOGIC_X0Y146_TQ = 1'b1;
  assign LIOI3_X0Y145_OLOGIC_X0Y145_OQ = CLBLL_L_X4Y115_SLICE_X4Y115_AO5;
  assign LIOI3_X0Y145_OLOGIC_X0Y145_TQ = 1'b1;
  assign LIOI3_X0Y147_OLOGIC_X0Y148_OQ = CLBLM_R_X3Y112_SLICE_X2Y112_CO6;
  assign LIOI3_X0Y147_OLOGIC_X0Y148_TQ = 1'b1;
  assign LIOI3_X0Y147_OLOGIC_X0Y147_OQ = CLBLM_R_X3Y112_SLICE_X2Y112_AO5;
  assign LIOI3_X0Y147_OLOGIC_X0Y147_TQ = 1'b1;
  assign LIOI3_SING_X0Y100_ILOGIC_X0Y100_O = LIOB33_SING_X0Y100_IOB_X0Y100_I;
  assign LIOI3_SING_X0Y149_OLOGIC_X0Y149_OQ = CLBLM_R_X3Y112_SLICE_X2Y112_DO6;
  assign LIOI3_SING_X0Y149_OLOGIC_X0Y149_TQ = 1'b1;
  assign LIOI3_TBYTESRC_X0Y107_ILOGIC_X0Y108_O = LIOB33_X0Y107_IOB_X0Y108_I;
  assign LIOI3_TBYTESRC_X0Y107_ILOGIC_X0Y107_O = LIOB33_X0Y107_IOB_X0Y107_I;
  assign LIOI3_TBYTESRC_X0Y119_OLOGIC_X0Y120_OQ = CLBLM_R_X3Y106_SLICE_X2Y106_AO5;
  assign LIOI3_TBYTESRC_X0Y119_OLOGIC_X0Y120_TQ = 1'b1;
  assign LIOI3_TBYTESRC_X0Y119_OLOGIC_X0Y119_OQ = CLBLL_L_X2Y109_SLICE_X0Y109_AO6;
  assign LIOI3_TBYTESRC_X0Y119_OLOGIC_X0Y119_TQ = 1'b1;
  assign LIOI3_TBYTESRC_X0Y131_OLOGIC_X0Y132_OQ = CLBLL_L_X2Y110_SLICE_X0Y110_AO5;
  assign LIOI3_TBYTESRC_X0Y131_OLOGIC_X0Y132_TQ = 1'b1;
  assign LIOI3_TBYTESRC_X0Y131_OLOGIC_X0Y131_OQ = CLBLL_L_X4Y108_SLICE_X4Y108_AO6;
  assign LIOI3_TBYTESRC_X0Y131_OLOGIC_X0Y131_TQ = 1'b1;
  assign LIOI3_TBYTESRC_X0Y143_OLOGIC_X0Y144_OQ = CLBLL_L_X4Y116_SLICE_X4Y116_AO6;
  assign LIOI3_TBYTESRC_X0Y143_OLOGIC_X0Y144_TQ = 1'b1;
  assign LIOI3_TBYTESRC_X0Y143_OLOGIC_X0Y143_OQ = CLBLL_L_X4Y115_SLICE_X4Y115_DO6;
  assign LIOI3_TBYTESRC_X0Y143_OLOGIC_X0Y143_TQ = 1'b1;
  assign LIOI3_TBYTETERM_X0Y113_ILOGIC_X0Y114_O = LIOB33_X0Y113_IOB_X0Y114_I;
  assign LIOI3_TBYTETERM_X0Y113_ILOGIC_X0Y113_O = LIOB33_X0Y113_IOB_X0Y113_I;
  assign LIOI3_TBYTETERM_X0Y137_OLOGIC_X0Y138_OQ = CLBLL_L_X4Y111_SLICE_X4Y111_AO5;
  assign LIOI3_TBYTETERM_X0Y137_OLOGIC_X0Y138_TQ = 1'b1;
  assign LIOI3_TBYTETERM_X0Y137_OLOGIC_X0Y137_OQ = CLBLL_L_X4Y111_SLICE_X4Y111_AO6;
  assign LIOI3_TBYTETERM_X0Y137_OLOGIC_X0Y137_TQ = 1'b1;
  assign RIOI3_X105Y101_ILOGIC_X1Y102_O = RIOB33_X105Y101_IOB_X1Y102_I;
  assign RIOI3_X105Y101_ILOGIC_X1Y101_O = RIOB33_X105Y101_IOB_X1Y101_I;
  assign RIOI3_X105Y103_ILOGIC_X1Y104_O = RIOB33_X105Y103_IOB_X1Y104_I;
  assign RIOI3_X105Y103_ILOGIC_X1Y103_O = RIOB33_X105Y103_IOB_X1Y103_I;
  assign RIOI3_X105Y105_ILOGIC_X1Y106_O = RIOB33_X105Y105_IOB_X1Y106_I;
  assign RIOI3_X105Y105_ILOGIC_X1Y105_O = RIOB33_X105Y105_IOB_X1Y105_I;
  assign RIOI3_X105Y109_ILOGIC_X1Y110_O = RIOB33_X105Y109_IOB_X1Y110_I;
  assign RIOI3_X105Y109_ILOGIC_X1Y109_O = RIOB33_X105Y109_IOB_X1Y109_I;
  assign RIOI3_X105Y111_ILOGIC_X1Y112_O = RIOB33_X105Y111_IOB_X1Y112_I;
  assign RIOI3_X105Y111_ILOGIC_X1Y111_O = RIOB33_X105Y111_IOB_X1Y111_I;
  assign RIOI3_SING_X105Y100_ILOGIC_X1Y100_O = RIOB33_SING_X105Y100_IOB_X1Y100_I;
  assign RIOI3_TBYTESRC_X105Y107_ILOGIC_X1Y108_O = RIOB33_X105Y107_IOB_X1Y108_I;
  assign RIOI3_TBYTESRC_X105Y107_ILOGIC_X1Y107_O = RIOB33_X105Y107_IOB_X1Y107_I;
  assign RIOI3_TBYTETERM_X105Y113_ILOGIC_X1Y113_O = RIOB33_X105Y113_IOB_X1Y113_I;
  assign CLBLM_L_X10Y103_SLICE_X12Y103_C6 = CLBLM_L_X10Y103_SLICE_X12Y103_BO6;
  assign CLBLM_L_X10Y103_SLICE_X12Y103_D1 = RIOB33_X105Y101_IOB_X1Y101_I;
  assign CLBLM_L_X10Y103_SLICE_X12Y103_D2 = CLBLM_L_X8Y104_SLICE_X10Y104_CO6;
  assign CLBLM_L_X10Y103_SLICE_X12Y103_D3 = RIOB33_X105Y101_IOB_X1Y102_I;
  assign CLBLM_L_X10Y103_SLICE_X12Y103_D4 = CLBLM_L_X10Y103_SLICE_X12Y103_CO6;
  assign CLBLM_L_X10Y103_SLICE_X12Y103_D5 = LIOB33_X0Y101_IOB_X0Y102_I;
  assign CLBLM_L_X10Y103_SLICE_X12Y103_D6 = LIOB33_X0Y103_IOB_X0Y104_I;
  assign CLBLM_R_X7Y109_SLICE_X9Y109_A4 = CLBLM_R_X3Y107_SLICE_X2Y107_BO6;
  assign CLBLM_R_X7Y109_SLICE_X9Y109_A5 = RIOB33_X105Y109_IOB_X1Y110_I;
  assign LIOB33_X0Y147_IOB_X0Y147_O = CLBLM_R_X3Y112_SLICE_X2Y112_AO5;
  assign LIOB33_X0Y147_IOB_X0Y148_O = CLBLM_R_X3Y112_SLICE_X2Y112_CO6;
  assign CLBLM_R_X7Y109_SLICE_X9Y109_A6 = 1'b1;
  assign CLBLL_L_X2Y106_SLICE_X1Y106_B6 = RIOB33_SING_X105Y100_IOB_X1Y100_I;
  assign CLBLM_R_X13Y107_SLICE_X19Y107_A1 = 1'b1;
  assign CLBLM_R_X13Y107_SLICE_X19Y107_A2 = 1'b1;
  assign CLBLM_R_X13Y107_SLICE_X19Y107_A3 = 1'b1;
  assign CLBLM_R_X13Y107_SLICE_X19Y107_A4 = 1'b1;
  assign CLBLM_R_X13Y107_SLICE_X19Y107_A5 = 1'b1;
  assign CLBLM_R_X13Y107_SLICE_X19Y107_A6 = 1'b1;
  assign CLBLM_R_X13Y107_SLICE_X19Y107_B1 = 1'b1;
  assign CLBLM_R_X13Y107_SLICE_X19Y107_B2 = 1'b1;
  assign CLBLM_R_X13Y107_SLICE_X19Y107_B3 = 1'b1;
  assign CLBLM_R_X13Y107_SLICE_X19Y107_B4 = 1'b1;
  assign CLBLM_R_X13Y107_SLICE_X19Y107_B5 = 1'b1;
  assign CLBLM_R_X13Y107_SLICE_X19Y107_B6 = 1'b1;
  assign CLBLM_R_X13Y107_SLICE_X19Y107_C1 = 1'b1;
  assign CLBLM_R_X13Y107_SLICE_X19Y107_C2 = 1'b1;
  assign CLBLM_R_X13Y107_SLICE_X19Y107_C3 = 1'b1;
  assign CLBLM_R_X13Y107_SLICE_X19Y107_C4 = 1'b1;
  assign CLBLM_R_X13Y107_SLICE_X19Y107_C5 = 1'b1;
  assign CLBLM_R_X13Y107_SLICE_X19Y107_C6 = 1'b1;
  assign CLBLM_R_X13Y107_SLICE_X19Y107_D1 = 1'b1;
  assign CLBLM_R_X13Y107_SLICE_X19Y107_D2 = 1'b1;
  assign CLBLM_R_X13Y107_SLICE_X19Y107_D3 = 1'b1;
  assign CLBLM_R_X13Y107_SLICE_X19Y107_D4 = 1'b1;
  assign CLBLM_R_X13Y107_SLICE_X19Y107_D5 = 1'b1;
  assign CLBLM_R_X13Y107_SLICE_X19Y107_D6 = 1'b1;
  assign CLBLM_R_X13Y107_SLICE_X18Y107_A1 = CLBLM_R_X13Y106_SLICE_X18Y106_DO6;
  assign CLBLM_R_X13Y107_SLICE_X18Y107_A2 = CLBLM_L_X12Y106_SLICE_X17Y106_DO6;
  assign CLBLM_R_X13Y107_SLICE_X18Y107_A3 = LIOB33_X0Y101_IOB_X0Y102_I;
  assign CLBLM_R_X13Y107_SLICE_X18Y107_A4 = RIOB33_X105Y107_IOB_X1Y108_I;
  assign CLBLM_R_X13Y107_SLICE_X18Y107_A5 = RIOB33_X105Y107_IOB_X1Y107_I;
  assign CLBLM_R_X13Y107_SLICE_X18Y107_A6 = LIOB33_X0Y103_IOB_X0Y104_I;
  assign CLBLM_R_X13Y107_SLICE_X18Y107_B1 = 1'b1;
  assign CLBLM_R_X13Y107_SLICE_X18Y107_B2 = 1'b1;
  assign CLBLM_R_X13Y107_SLICE_X18Y107_B3 = 1'b1;
  assign CLBLM_R_X13Y107_SLICE_X18Y107_B4 = 1'b1;
  assign CLBLM_R_X13Y107_SLICE_X18Y107_B5 = 1'b1;
  assign CLBLM_R_X13Y107_SLICE_X18Y107_B6 = 1'b1;
  assign CLBLM_R_X13Y107_SLICE_X18Y107_C1 = 1'b1;
  assign CLBLM_R_X13Y107_SLICE_X18Y107_C2 = 1'b1;
  assign CLBLM_R_X13Y107_SLICE_X18Y107_C3 = 1'b1;
  assign CLBLM_R_X13Y107_SLICE_X18Y107_C4 = 1'b1;
  assign CLBLM_R_X13Y107_SLICE_X18Y107_C5 = 1'b1;
  assign CLBLM_R_X13Y107_SLICE_X18Y107_C6 = 1'b1;
  assign CLBLM_R_X13Y107_SLICE_X18Y107_D1 = 1'b1;
  assign CLBLM_R_X13Y107_SLICE_X18Y107_D2 = 1'b1;
  assign CLBLM_R_X13Y107_SLICE_X18Y107_D3 = 1'b1;
  assign CLBLM_R_X13Y107_SLICE_X18Y107_D4 = 1'b1;
  assign CLBLM_R_X13Y107_SLICE_X18Y107_D5 = 1'b1;
  assign CLBLM_R_X13Y107_SLICE_X18Y107_D6 = 1'b1;
  assign CLBLM_L_X10Y104_SLICE_X13Y104_A1 = LIOB33_X0Y101_IOB_X0Y101_I;
  assign CLBLM_L_X10Y104_SLICE_X13Y104_A2 = 1'b1;
  assign CLBLM_L_X10Y104_SLICE_X13Y104_A3 = LIOB33_X0Y101_IOB_X0Y102_I;
  assign CLBLM_L_X10Y104_SLICE_X13Y104_A4 = RIOB33_X105Y103_IOB_X1Y103_I;
  assign CLBLM_L_X10Y104_SLICE_X13Y104_A5 = 1'b1;
  assign CLBLM_L_X10Y104_SLICE_X13Y104_A6 = 1'b1;
  assign CLBLM_L_X10Y104_SLICE_X13Y104_B1 = CLBLM_R_X11Y104_SLICE_X15Y104_BO6;
  assign CLBLM_L_X10Y104_SLICE_X13Y104_B2 = CLBLM_L_X10Y104_SLICE_X12Y104_BO6;
  assign CLBLM_L_X10Y104_SLICE_X13Y104_B3 = CLBLM_L_X10Y104_SLICE_X13Y104_AO6;
  assign CLBLM_L_X10Y104_SLICE_X13Y104_B4 = CLBLM_L_X10Y104_SLICE_X12Y104_DO6;
  assign CLBLM_L_X10Y104_SLICE_X13Y104_B5 = CLBLM_R_X11Y104_SLICE_X14Y104_AO6;
  assign CLBLM_L_X10Y104_SLICE_X13Y104_B6 = CLBLM_L_X10Y104_SLICE_X13Y104_AO5;
  assign CLBLM_L_X10Y104_SLICE_X13Y104_C1 = RIOB33_X105Y103_IOB_X1Y104_I;
  assign CLBLM_L_X10Y104_SLICE_X13Y104_C2 = RIOB33_X105Y103_IOB_X1Y103_I;
  assign CLBLM_L_X10Y104_SLICE_X13Y104_C3 = CLBLM_L_X10Y104_SLICE_X12Y104_BO6;
  assign CLBLM_L_X10Y104_SLICE_X13Y104_C4 = CLBLM_R_X11Y104_SLICE_X15Y104_BO6;
  assign CLBLM_L_X10Y104_SLICE_X13Y104_C5 = LIOB33_X0Y101_IOB_X0Y101_I;
  assign CLBLM_L_X10Y104_SLICE_X13Y104_C6 = CLBLM_L_X10Y104_SLICE_X12Y104_DO6;
  assign CLBLM_L_X10Y104_SLICE_X13Y104_D1 = CLBLM_R_X11Y104_SLICE_X14Y104_AO6;
  assign CLBLM_L_X10Y104_SLICE_X13Y104_D2 = CLBLM_R_X11Y104_SLICE_X15Y104_BO6;
  assign CLBLM_L_X10Y104_SLICE_X13Y104_D3 = CLBLM_L_X10Y104_SLICE_X12Y104_BO6;
  assign CLBLM_L_X10Y104_SLICE_X13Y104_D4 = CLBLM_L_X10Y104_SLICE_X13Y104_AO5;
  assign CLBLM_L_X10Y104_SLICE_X13Y104_D5 = CLBLM_L_X10Y104_SLICE_X13Y104_AO6;
  assign CLBLM_L_X10Y104_SLICE_X13Y104_D6 = CLBLM_L_X10Y104_SLICE_X12Y104_DO6;
  assign CLBLM_L_X10Y104_SLICE_X12Y104_A1 = RIOB33_X105Y101_IOB_X1Y102_I;
  assign CLBLM_L_X10Y104_SLICE_X12Y104_A2 = RIOB33_X105Y111_IOB_X1Y112_I;
  assign CLBLM_L_X10Y104_SLICE_X12Y104_A3 = RIOB33_X105Y113_IOB_X1Y113_I;
  assign CLBLM_L_X10Y104_SLICE_X12Y104_A4 = RIOB33_X105Y103_IOB_X1Y104_I;
  assign CLBLM_L_X10Y104_SLICE_X12Y104_A5 = RIOB33_X105Y103_IOB_X1Y103_I;
  assign CLBLM_L_X10Y104_SLICE_X12Y104_A6 = LIOB33_SING_X0Y100_IOB_X0Y100_I;
  assign CLBLM_L_X10Y104_SLICE_X12Y104_B1 = RIOB33_X105Y103_IOB_X1Y104_I;
  assign CLBLM_L_X10Y104_SLICE_X12Y104_B2 = RIOB33_X105Y103_IOB_X1Y103_I;
  assign CLBLM_L_X10Y104_SLICE_X12Y104_B3 = RIOB33_X105Y111_IOB_X1Y112_I;
  assign CLBLM_L_X10Y104_SLICE_X12Y104_B4 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X10Y104_SLICE_X12Y104_B5 = RIOB33_X105Y113_IOB_X1Y113_I;
  assign CLBLM_L_X10Y104_SLICE_X12Y104_B6 = LIOB33_SING_X0Y100_IOB_X0Y100_I;
  assign CLBLM_L_X10Y104_SLICE_X12Y104_C1 = CLBLM_L_X10Y105_SLICE_X13Y105_AO6;
  assign CLBLM_L_X10Y104_SLICE_X12Y104_C2 = CLBLM_L_X8Y104_SLICE_X10Y104_CO6;
  assign CLBLM_L_X10Y104_SLICE_X12Y104_C3 = CLBLM_L_X10Y102_SLICE_X12Y102_BO6;
  assign CLBLM_L_X10Y104_SLICE_X12Y104_C4 = CLBLM_L_X10Y102_SLICE_X12Y102_CO6;
  assign CLBLM_L_X10Y104_SLICE_X12Y104_C5 = CLBLM_L_X10Y104_SLICE_X13Y104_BO6;
  assign CLBLM_L_X10Y104_SLICE_X12Y104_C6 = CLBLM_L_X8Y105_SLICE_X11Y105_AO6;
  assign CLBLM_L_X10Y104_SLICE_X12Y104_D1 = RIOB33_X105Y113_IOB_X1Y113_I;
  assign CLBLM_L_X10Y104_SLICE_X12Y104_D2 = LIOB33_SING_X0Y100_IOB_X0Y100_I;
  assign CLBLM_L_X10Y104_SLICE_X12Y104_D3 = RIOB33_X105Y103_IOB_X1Y103_I;
  assign CLBLM_L_X10Y104_SLICE_X12Y104_D4 = RIOB33_X105Y111_IOB_X1Y112_I;
  assign CLBLM_L_X10Y104_SLICE_X12Y104_D5 = RIOB33_X105Y103_IOB_X1Y104_I;
  assign CLBLM_L_X10Y104_SLICE_X12Y104_D6 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X10Y105_SLICE_X13Y105_A1 = RIOB33_X105Y101_IOB_X1Y102_I;
  assign CLBLM_L_X10Y105_SLICE_X13Y105_A2 = LIOB33_X0Y105_IOB_X0Y105_I;
  assign CLBLM_L_X10Y105_SLICE_X13Y105_A3 = 1'b1;
  assign CLBLM_L_X10Y105_SLICE_X13Y105_A4 = LIOB33_X0Y103_IOB_X0Y104_I;
  assign CLBLM_L_X10Y105_SLICE_X13Y105_A5 = 1'b1;
  assign CLBLM_L_X10Y105_SLICE_X13Y105_A6 = 1'b1;
  assign CLBLM_L_X10Y105_SLICE_X13Y105_B1 = CLBLM_L_X10Y104_SLICE_X13Y104_DO6;
  assign CLBLM_L_X10Y105_SLICE_X13Y105_B2 = CLBLM_R_X11Y105_SLICE_X14Y105_AO6;
  assign CLBLM_L_X10Y105_SLICE_X13Y105_B3 = CLBLM_L_X10Y104_SLICE_X13Y104_BO6;
  assign CLBLM_L_X10Y105_SLICE_X13Y105_B4 = CLBLM_R_X11Y104_SLICE_X14Y104_BO6;
  assign CLBLM_L_X10Y105_SLICE_X13Y105_B5 = CLBLM_L_X10Y105_SLICE_X13Y105_AO6;
  assign CLBLM_L_X10Y105_SLICE_X13Y105_B6 = CLBLM_L_X10Y102_SLICE_X12Y102_CO6;
  assign CLBLM_L_X8Y103_SLICE_X10Y103_C2 = 1'b1;
  assign CLBLM_L_X8Y103_SLICE_X10Y103_C3 = 1'b1;
  assign CLBLM_L_X10Y105_SLICE_X13Y105_C1 = LIOB33_X0Y103_IOB_X0Y104_I;
  assign CLBLM_L_X10Y105_SLICE_X13Y105_C2 = CLBLM_L_X10Y102_SLICE_X12Y102_CO6;
  assign CLBLM_L_X10Y105_SLICE_X13Y105_C3 = RIOB33_X105Y103_IOB_X1Y103_I;
  assign CLBLM_L_X10Y105_SLICE_X13Y105_C4 = CLBLM_L_X10Y104_SLICE_X13Y104_CO6;
  assign CLBLM_L_X10Y105_SLICE_X13Y105_C5 = RIOB33_X105Y101_IOB_X1Y102_I;
  assign CLBLM_L_X10Y105_SLICE_X13Y105_C6 = LIOB33_X0Y101_IOB_X0Y102_I;
  assign CLBLM_L_X8Y103_SLICE_X10Y103_C4 = 1'b1;
  assign CLBLM_L_X10Y105_SLICE_X13Y105_D1 = LIOB33_X0Y103_IOB_X0Y104_I;
  assign CLBLM_L_X10Y105_SLICE_X13Y105_D2 = LIOB33_X0Y105_IOB_X0Y105_I;
  assign CLBLM_L_X10Y105_SLICE_X13Y105_D3 = CLBLM_L_X10Y105_SLICE_X12Y105_DO6;
  assign CLBLM_L_X10Y105_SLICE_X13Y105_D4 = CLBLM_L_X10Y105_SLICE_X13Y105_CO6;
  assign CLBLM_L_X10Y105_SLICE_X13Y105_D5 = RIOB33_X105Y101_IOB_X1Y102_I;
  assign CLBLM_L_X10Y105_SLICE_X13Y105_D6 = RIOB33_X105Y103_IOB_X1Y103_I;
  assign CLBLM_L_X10Y105_SLICE_X12Y105_A1 = RIOB33_X105Y103_IOB_X1Y103_I;
  assign CLBLM_L_X10Y105_SLICE_X12Y105_A2 = CLBLM_L_X10Y104_SLICE_X12Y104_BO6;
  assign CLBLM_L_X10Y105_SLICE_X12Y105_A3 = LIOB33_X0Y101_IOB_X0Y101_I;
  assign CLBLM_L_X10Y105_SLICE_X12Y105_A4 = CLBLM_L_X10Y104_SLICE_X12Y104_DO6;
  assign CLBLM_L_X10Y105_SLICE_X12Y105_A5 = 1'b1;
  assign CLBLM_L_X10Y105_SLICE_X12Y105_A6 = 1'b1;
  assign CLBLM_L_X10Y105_SLICE_X12Y105_B1 = RIOB33_X105Y101_IOB_X1Y102_I;
  assign CLBLM_L_X10Y105_SLICE_X12Y105_B2 = LIOB33_X0Y101_IOB_X0Y102_I;
  assign CLBLM_L_X10Y105_SLICE_X12Y105_B3 = CLBLM_L_X10Y104_SLICE_X13Y104_CO6;
  assign CLBLM_L_X10Y105_SLICE_X12Y105_B4 = RIOB33_X105Y103_IOB_X1Y103_I;
  assign CLBLM_L_X10Y105_SLICE_X12Y105_B5 = CLBLM_L_X10Y105_SLICE_X12Y105_AO6;
  assign CLBLM_L_X10Y105_SLICE_X12Y105_B6 = CLBLM_L_X10Y103_SLICE_X12Y103_AO5;
  assign CLBLM_L_X10Y105_SLICE_X12Y105_C1 = LIOB33_X0Y103_IOB_X0Y104_I;
  assign CLBLM_L_X10Y105_SLICE_X12Y105_C2 = RIOB33_X105Y103_IOB_X1Y103_I;
  assign CLBLM_L_X10Y105_SLICE_X12Y105_C3 = RIOB33_X105Y101_IOB_X1Y102_I;
  assign CLBLM_L_X10Y105_SLICE_X12Y105_C4 = CLBLM_L_X10Y102_SLICE_X12Y102_CO6;
  assign CLBLM_L_X10Y105_SLICE_X12Y105_C5 = LIOB33_X0Y101_IOB_X0Y102_I;
  assign CLBLM_L_X10Y105_SLICE_X12Y105_C6 = CLBLM_L_X10Y104_SLICE_X13Y104_CO6;
  assign CLBLM_L_X10Y105_SLICE_X12Y105_D1 = CLBLM_R_X11Y104_SLICE_X15Y104_AO6;
  assign CLBLM_L_X10Y105_SLICE_X12Y105_D2 = RIOB33_X105Y103_IOB_X1Y104_I;
  assign CLBLM_L_X10Y105_SLICE_X12Y105_D3 = CLBLM_R_X11Y104_SLICE_X14Y104_DO6;
  assign CLBLM_L_X10Y105_SLICE_X12Y105_D4 = CLBLM_L_X10Y105_SLICE_X12Y105_AO5;
  assign CLBLM_L_X10Y105_SLICE_X12Y105_D5 = LIOB33_X0Y101_IOB_X0Y102_I;
  assign CLBLM_L_X10Y105_SLICE_X12Y105_D6 = RIOB33_X105Y103_IOB_X1Y103_I;
  assign CLBLM_L_X10Y106_SLICE_X13Y106_A1 = LIOB33_X0Y105_IOB_X0Y105_I;
  assign CLBLM_L_X10Y106_SLICE_X13Y106_A2 = CLBLM_R_X11Y105_SLICE_X14Y105_CO6;
  assign CLBLM_L_X10Y106_SLICE_X13Y106_A3 = RIOB33_X105Y101_IOB_X1Y102_I;
  assign CLBLM_L_X10Y106_SLICE_X13Y106_A4 = CLBLM_R_X11Y105_SLICE_X14Y105_BO6;
  assign CLBLM_L_X10Y106_SLICE_X13Y106_A5 = CLBLM_L_X10Y105_SLICE_X13Y105_CO6;
  assign CLBLM_L_X10Y106_SLICE_X13Y106_A6 = RIOB33_X105Y103_IOB_X1Y103_I;
  assign CLBLM_L_X10Y106_SLICE_X13Y106_B1 = RIOB33_X105Y103_IOB_X1Y103_I;
  assign CLBLM_L_X10Y106_SLICE_X13Y106_B2 = CLBLM_L_X10Y105_SLICE_X12Y105_DO6;
  assign CLBLM_L_X10Y106_SLICE_X13Y106_B3 = RIOB33_X105Y101_IOB_X1Y102_I;
  assign CLBLM_L_X10Y106_SLICE_X13Y106_B4 = CLBLM_L_X10Y105_SLICE_X13Y105_CO6;
  assign CLBLM_L_X10Y106_SLICE_X13Y106_B5 = LIOB33_X0Y105_IOB_X0Y105_I;
  assign CLBLM_L_X10Y106_SLICE_X13Y106_B6 = LIOB33_X0Y103_IOB_X0Y104_I;
  assign CLBLM_L_X10Y106_SLICE_X13Y106_C1 = CLBLM_R_X11Y105_SLICE_X14Y105_BO6;
  assign CLBLM_L_X10Y106_SLICE_X13Y106_C2 = CLBLM_R_X11Y105_SLICE_X14Y105_CO6;
  assign CLBLM_L_X10Y106_SLICE_X13Y106_C3 = CLBLM_R_X11Y105_SLICE_X14Y105_AO5;
  assign CLBLM_L_X10Y106_SLICE_X13Y106_C4 = CLBLM_L_X10Y108_SLICE_X13Y108_AO5;
  assign CLBLM_L_X10Y106_SLICE_X13Y106_C5 = CLBLM_L_X10Y105_SLICE_X13Y105_AO5;
  assign CLBLM_L_X10Y106_SLICE_X13Y106_C6 = CLBLM_L_X10Y105_SLICE_X13Y105_CO6;
  assign CLBLM_L_X10Y106_SLICE_X13Y106_D1 = CLBLM_R_X11Y105_SLICE_X14Y105_BO6;
  assign CLBLM_L_X10Y106_SLICE_X13Y106_D2 = CLBLM_R_X11Y105_SLICE_X14Y105_CO6;
  assign CLBLM_L_X10Y106_SLICE_X13Y106_D3 = CLBLM_L_X10Y105_SLICE_X13Y105_AO5;
  assign CLBLM_L_X10Y106_SLICE_X13Y106_D4 = CLBLM_L_X10Y108_SLICE_X13Y108_AO5;
  assign CLBLM_L_X10Y106_SLICE_X13Y106_D5 = CLBLM_R_X11Y105_SLICE_X14Y105_AO5;
  assign CLBLM_L_X10Y106_SLICE_X13Y106_D6 = CLBLM_L_X10Y105_SLICE_X13Y105_CO6;
  assign CLBLM_L_X10Y106_SLICE_X12Y106_A1 = RIOB33_X105Y101_IOB_X1Y101_I;
  assign CLBLM_L_X10Y106_SLICE_X12Y106_A2 = LIOB33_X0Y107_IOB_X0Y107_I;
  assign CLBLM_L_X10Y106_SLICE_X12Y106_A3 = CLBLM_L_X10Y106_SLICE_X13Y106_AO6;
  assign CLBLM_L_X10Y106_SLICE_X12Y106_A4 = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLM_L_X10Y106_SLICE_X12Y106_A5 = RIOB33_X105Y101_IOB_X1Y102_I;
  assign CLBLM_L_X10Y106_SLICE_X12Y106_A6 = CLBLM_L_X8Y105_SLICE_X11Y105_CO6;
  assign CLBLM_L_X10Y106_SLICE_X12Y106_B1 = RIOB33_X105Y101_IOB_X1Y101_I;
  assign CLBLM_L_X10Y106_SLICE_X12Y106_B2 = CLBLM_L_X10Y106_SLICE_X13Y106_BO6;
  assign CLBLM_L_X10Y106_SLICE_X12Y106_B3 = CLBLM_L_X10Y106_SLICE_X13Y106_AO6;
  assign CLBLM_L_X10Y106_SLICE_X12Y106_B4 = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLM_L_X10Y106_SLICE_X12Y106_B5 = RIOB33_X105Y101_IOB_X1Y102_I;
  assign CLBLM_L_X10Y106_SLICE_X12Y106_B6 = CLBLM_L_X10Y106_SLICE_X12Y106_CO6;
  assign CLBLM_L_X10Y106_SLICE_X12Y106_C1 = RIOB33_X105Y101_IOB_X1Y102_I;
  assign CLBLM_L_X10Y106_SLICE_X12Y106_C2 = LIOB33_X0Y103_IOB_X0Y104_I;
  assign CLBLM_L_X10Y106_SLICE_X12Y106_C3 = LIOB33_X0Y105_IOB_X0Y105_I;
  assign CLBLM_L_X10Y106_SLICE_X12Y106_C4 = CLBLM_L_X10Y103_SLICE_X12Y103_DO6;
  assign CLBLM_L_X10Y106_SLICE_X12Y106_C5 = RIOB33_X105Y101_IOB_X1Y101_I;
  assign CLBLM_L_X10Y106_SLICE_X12Y106_C6 = CLBLM_L_X10Y105_SLICE_X12Y105_BO6;
  assign CLBLM_L_X10Y106_SLICE_X12Y106_D1 = RIOB33_X105Y101_IOB_X1Y102_I;
  assign CLBLM_L_X10Y106_SLICE_X12Y106_D2 = CLBLM_L_X10Y106_SLICE_X13Y106_AO6;
  assign CLBLM_L_X10Y106_SLICE_X12Y106_D3 = LIOB33_X0Y107_IOB_X0Y107_I;
  assign CLBLM_L_X10Y106_SLICE_X12Y106_D4 = CLBLM_L_X8Y105_SLICE_X11Y105_CO6;
  assign CLBLM_L_X10Y106_SLICE_X12Y106_D5 = RIOB33_X105Y101_IOB_X1Y101_I;
  assign CLBLM_L_X10Y106_SLICE_X12Y106_D6 = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLM_L_X10Y107_SLICE_X13Y107_A1 = LIOB33_X0Y105_IOB_X0Y105_I;
  assign CLBLM_L_X10Y107_SLICE_X13Y107_A2 = CLBLM_R_X11Y107_SLICE_X15Y107_AO5;
  assign CLBLM_L_X10Y107_SLICE_X13Y107_A3 = RIOB33_X105Y109_IOB_X1Y109_I;
  assign CLBLM_L_X10Y107_SLICE_X13Y107_A4 = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLM_L_X10Y107_SLICE_X13Y107_A5 = RIOB33_X105Y109_IOB_X1Y110_I;
  assign CLBLM_L_X10Y107_SLICE_X13Y107_A6 = CLBLM_L_X10Y107_SLICE_X13Y107_CO6;
  assign CLBLM_L_X10Y107_SLICE_X13Y107_B1 = CLBLM_L_X10Y108_SLICE_X13Y108_DO6;
  assign CLBLM_L_X10Y107_SLICE_X13Y107_B2 = CLBLM_R_X11Y107_SLICE_X15Y107_AO5;
  assign CLBLM_L_X10Y107_SLICE_X13Y107_B3 = LIOB33_X0Y107_IOB_X0Y107_I;
  assign CLBLM_L_X10Y107_SLICE_X13Y107_B4 = RIOB33_X105Y109_IOB_X1Y109_I;
  assign CLBLM_L_X10Y107_SLICE_X13Y107_B5 = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLM_L_X10Y107_SLICE_X13Y107_B6 = CLBLM_R_X11Y107_SLICE_X14Y107_BO6;
  assign CLBLM_L_X10Y107_SLICE_X13Y107_C1 = LIOB33_X0Y101_IOB_X0Y102_I;
  assign CLBLM_L_X10Y107_SLICE_X13Y107_C2 = CLBLM_L_X10Y107_SLICE_X12Y107_CO6;
  assign CLBLM_L_X10Y107_SLICE_X13Y107_C3 = RIOB33_X105Y109_IOB_X1Y110_I;
  assign CLBLM_L_X10Y107_SLICE_X13Y107_C4 = RIOB33_X105Y111_IOB_X1Y111_I;
  assign CLBLM_L_X10Y107_SLICE_X13Y107_C5 = LIOB33_X0Y103_IOB_X0Y104_I;
  assign CLBLM_L_X10Y107_SLICE_X13Y107_C6 = LIOB33_X0Y101_IOB_X0Y101_I;
  assign CLBLM_L_X10Y107_SLICE_X13Y107_D1 = LIOB33_X0Y101_IOB_X0Y101_I;
  assign CLBLM_L_X10Y107_SLICE_X13Y107_D2 = RIOB33_X105Y113_IOB_X1Y113_I;
  assign CLBLM_L_X10Y107_SLICE_X13Y107_D3 = RIOB33_X105Y111_IOB_X1Y111_I;
  assign CLBLM_L_X10Y107_SLICE_X13Y107_D4 = RIOB33_X105Y109_IOB_X1Y110_I;
  assign CLBLM_L_X10Y107_SLICE_X13Y107_D5 = LIOB33_SING_X0Y100_IOB_X0Y100_I;
  assign CLBLM_L_X10Y107_SLICE_X13Y107_D6 = RIOB33_X105Y111_IOB_X1Y112_I;
  assign CLBLM_L_X10Y107_SLICE_X12Y107_A1 = CLBLM_L_X10Y106_SLICE_X13Y106_DO6;
  assign CLBLM_L_X10Y107_SLICE_X12Y107_A2 = CLBLM_L_X10Y108_SLICE_X13Y108_BO6;
  assign CLBLM_L_X10Y107_SLICE_X12Y107_A3 = CLBLM_L_X10Y106_SLICE_X13Y106_CO6;
  assign CLBLM_L_X10Y107_SLICE_X12Y107_A4 = CLBLM_L_X10Y108_SLICE_X13Y108_AO6;
  assign CLBLM_L_X10Y107_SLICE_X12Y107_A5 = CLBLM_R_X11Y106_SLICE_X14Y106_AO6;
  assign CLBLM_L_X10Y107_SLICE_X12Y107_A6 = CLBLM_L_X8Y105_SLICE_X11Y105_CO6;
  assign CLBLM_L_X10Y107_SLICE_X12Y107_B1 = RIOB33_X105Y109_IOB_X1Y110_I;
  assign CLBLM_L_X10Y107_SLICE_X12Y107_B2 = LIOB33_X0Y101_IOB_X0Y101_I;
  assign CLBLM_L_X10Y107_SLICE_X12Y107_B3 = LIOB33_X0Y101_IOB_X0Y102_I;
  assign CLBLM_L_X10Y107_SLICE_X12Y107_B4 = RIOB33_X105Y111_IOB_X1Y111_I;
  assign CLBLM_L_X10Y107_SLICE_X12Y107_B5 = LIOB33_X0Y103_IOB_X0Y104_I;
  assign CLBLM_L_X10Y107_SLICE_X12Y107_B6 = CLBLM_L_X10Y107_SLICE_X12Y107_CO6;
  assign CLBLM_L_X10Y107_SLICE_X12Y107_C1 = LIOB33_SING_X0Y100_IOB_X0Y100_I;
  assign CLBLM_L_X10Y107_SLICE_X12Y107_C2 = RIOB33_X105Y109_IOB_X1Y110_I;
  assign CLBLM_L_X10Y107_SLICE_X12Y107_C3 = RIOB33_X105Y111_IOB_X1Y111_I;
  assign CLBLM_L_X10Y107_SLICE_X12Y107_C4 = RIOB33_X105Y113_IOB_X1Y113_I;
  assign CLBLM_L_X10Y107_SLICE_X12Y107_C5 = LIOB33_X0Y101_IOB_X0Y101_I;
  assign CLBLM_L_X10Y107_SLICE_X12Y107_C6 = RIOB33_X105Y111_IOB_X1Y112_I;
  assign CLBLM_L_X10Y107_SLICE_X12Y107_D1 = 1'b1;
  assign CLBLM_L_X10Y107_SLICE_X12Y107_D2 = 1'b1;
  assign CLBLM_L_X10Y107_SLICE_X12Y107_D3 = 1'b1;
  assign CLBLM_L_X10Y107_SLICE_X12Y107_D4 = 1'b1;
  assign CLBLM_L_X10Y107_SLICE_X12Y107_D5 = 1'b1;
  assign CLBLM_L_X10Y107_SLICE_X12Y107_D6 = 1'b1;
  assign CLBLL_L_X4Y103_SLICE_X4Y103_A1 = LIOB33_X0Y101_IOB_X0Y101_I;
  assign CLBLL_L_X4Y103_SLICE_X4Y103_A2 = 1'b1;
  assign CLBLL_L_X4Y103_SLICE_X4Y103_A3 = 1'b1;
  assign CLBLL_L_X4Y103_SLICE_X4Y103_A4 = LIOB33_X0Y115_IOB_X0Y116_I;
  assign CLBLL_L_X4Y103_SLICE_X4Y103_A5 = LIOB33_X0Y103_IOB_X0Y103_I;
  assign CLBLL_L_X4Y103_SLICE_X4Y103_A6 = 1'b1;
  assign CLBLL_L_X4Y103_SLICE_X4Y103_B1 = LIOB33_X0Y101_IOB_X0Y101_I;
  assign CLBLL_L_X4Y103_SLICE_X4Y103_B2 = CLBLL_L_X4Y104_SLICE_X5Y104_BO6;
  assign CLBLL_L_X4Y103_SLICE_X4Y103_B3 = CLBLM_R_X3Y103_SLICE_X3Y103_BO6;
  assign CLBLL_L_X4Y103_SLICE_X4Y103_B4 = CLBLM_R_X3Y103_SLICE_X2Y103_BO6;
  assign CLBLL_L_X4Y103_SLICE_X4Y103_B5 = LIOB33_X0Y113_IOB_X0Y114_I;
  assign CLBLL_L_X4Y103_SLICE_X4Y103_B6 = LIOB33_X0Y115_IOB_X0Y116_I;
  assign CLBLL_L_X4Y103_SLICE_X4Y103_C1 = CLBLM_R_X3Y103_SLICE_X3Y103_BO6;
  assign CLBLL_L_X4Y103_SLICE_X4Y103_C2 = CLBLL_L_X4Y103_SLICE_X5Y103_AO5;
  assign CLBLL_L_X4Y103_SLICE_X4Y103_C3 = CLBLL_L_X4Y104_SLICE_X5Y104_BO6;
  assign CLBLL_L_X4Y103_SLICE_X4Y103_C4 = CLBLL_L_X4Y103_SLICE_X4Y103_AO5;
  assign CLBLL_L_X4Y103_SLICE_X4Y103_C5 = CLBLM_R_X3Y106_SLICE_X2Y106_BO5;
  assign CLBLL_L_X4Y103_SLICE_X4Y103_C6 = CLBLM_R_X3Y103_SLICE_X2Y103_BO6;
  assign CLBLL_L_X4Y103_SLICE_X4Y103_D1 = CLBLM_R_X3Y103_SLICE_X3Y103_BO6;
  assign CLBLL_L_X4Y103_SLICE_X4Y103_D2 = CLBLL_L_X4Y103_SLICE_X5Y103_AO5;
  assign CLBLL_L_X4Y103_SLICE_X4Y103_D3 = CLBLL_L_X4Y104_SLICE_X5Y104_BO6;
  assign CLBLL_L_X4Y103_SLICE_X4Y103_D4 = CLBLL_L_X4Y103_SLICE_X4Y103_AO5;
  assign CLBLL_L_X4Y103_SLICE_X4Y103_D5 = CLBLM_R_X3Y106_SLICE_X2Y106_BO5;
  assign CLBLL_L_X4Y103_SLICE_X4Y103_D6 = CLBLM_R_X3Y103_SLICE_X2Y103_BO6;
  assign CLBLL_L_X4Y103_SLICE_X5Y103_A1 = LIOB33_X0Y113_IOB_X0Y114_I;
  assign CLBLL_L_X4Y103_SLICE_X5Y103_A2 = LIOB33_X0Y115_IOB_X0Y116_I;
  assign CLBLL_L_X4Y103_SLICE_X5Y103_A3 = LIOB33_X0Y101_IOB_X0Y102_I;
  assign CLBLL_L_X4Y103_SLICE_X5Y103_A4 = 1'b1;
  assign CLBLL_L_X4Y103_SLICE_X5Y103_A5 = 1'b1;
  assign CLBLL_L_X4Y103_SLICE_X5Y103_A6 = 1'b1;
  assign CLBLL_L_X4Y103_SLICE_X5Y103_B1 = CLBLM_R_X7Y103_SLICE_X8Y103_AO6;
  assign CLBLL_L_X4Y103_SLICE_X5Y103_B2 = CLBLM_R_X7Y104_SLICE_X8Y104_AO6;
  assign CLBLL_L_X4Y103_SLICE_X5Y103_B3 = CLBLL_L_X4Y103_SLICE_X4Y103_AO5;
  assign CLBLL_L_X4Y103_SLICE_X5Y103_B4 = CLBLM_R_X5Y104_SLICE_X6Y104_BO6;
  assign CLBLL_L_X4Y103_SLICE_X5Y103_B5 = CLBLL_L_X4Y103_SLICE_X5Y103_AO6;
  assign CLBLL_L_X4Y103_SLICE_X5Y103_B6 = CLBLL_L_X4Y104_SLICE_X5Y104_BO6;
  assign CLBLL_L_X4Y103_SLICE_X5Y103_C1 = CLBLL_L_X4Y103_SLICE_X5Y103_AO6;
  assign CLBLL_L_X4Y103_SLICE_X5Y103_C2 = CLBLM_R_X5Y104_SLICE_X6Y104_BO6;
  assign CLBLL_L_X4Y103_SLICE_X5Y103_C3 = CLBLM_R_X7Y104_SLICE_X8Y104_AO6;
  assign CLBLL_L_X4Y103_SLICE_X5Y103_C4 = CLBLL_L_X4Y104_SLICE_X5Y104_BO6;
  assign CLBLL_L_X4Y103_SLICE_X5Y103_C5 = CLBLM_R_X7Y103_SLICE_X8Y103_AO6;
  assign CLBLL_L_X4Y103_SLICE_X5Y103_C6 = CLBLL_L_X4Y103_SLICE_X4Y103_AO5;
  assign CLBLL_L_X4Y103_SLICE_X5Y103_D1 = 1'b1;
  assign CLBLL_L_X4Y103_SLICE_X5Y103_D2 = 1'b1;
  assign CLBLL_L_X4Y103_SLICE_X5Y103_D3 = 1'b1;
  assign CLBLL_L_X4Y103_SLICE_X5Y103_D4 = 1'b1;
  assign CLBLL_L_X4Y103_SLICE_X5Y103_D5 = 1'b1;
  assign CLBLL_L_X4Y103_SLICE_X5Y103_D6 = 1'b1;
  assign CLBLM_R_X11Y108_SLICE_X15Y108_B1 = CLBLM_R_X11Y111_SLICE_X15Y111_AO5;
  assign CLBLM_R_X11Y108_SLICE_X15Y108_B2 = CLBLM_L_X12Y107_SLICE_X16Y107_CO6;
  assign CLBLM_R_X11Y108_SLICE_X15Y108_B3 = CLBLM_R_X11Y107_SLICE_X14Y107_AO5;
  assign CLBLM_L_X10Y108_SLICE_X13Y108_A1 = 1'b1;
  assign CLBLM_L_X10Y108_SLICE_X13Y108_A2 = 1'b1;
  assign CLBLM_L_X10Y108_SLICE_X13Y108_A3 = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLM_L_X10Y108_SLICE_X13Y108_A4 = LIOB33_X0Y107_IOB_X0Y107_I;
  assign CLBLM_L_X10Y108_SLICE_X13Y108_A5 = RIOB33_X105Y101_IOB_X1Y102_I;
  assign CLBLM_L_X10Y108_SLICE_X13Y108_A6 = 1'b1;
  assign CLBLM_L_X10Y108_SLICE_X13Y108_B1 = 1'b1;
  assign CLBLM_L_X10Y108_SLICE_X13Y108_B2 = LIOB33_X0Y107_IOB_X0Y107_I;
  assign CLBLM_L_X10Y108_SLICE_X13Y108_B3 = 1'b1;
  assign CLBLM_L_X10Y108_SLICE_X13Y108_B4 = RIOB33_X105Y103_IOB_X1Y103_I;
  assign CLBLM_L_X10Y108_SLICE_X13Y108_B5 = RIOB33_X105Y101_IOB_X1Y101_I;
  assign CLBLM_L_X10Y108_SLICE_X13Y108_B6 = 1'b1;
  assign CLBLM_R_X11Y108_SLICE_X15Y108_C3 = RIOB33_X105Y103_IOB_X1Y104_I;
  assign CLBLM_L_X10Y108_SLICE_X13Y108_C1 = CLBLM_L_X10Y108_SLICE_X13Y108_AO6;
  assign CLBLM_L_X10Y108_SLICE_X13Y108_C2 = CLBLM_R_X11Y108_SLICE_X15Y108_BO6;
  assign CLBLM_L_X10Y108_SLICE_X13Y108_C3 = CLBLM_R_X11Y106_SLICE_X14Y106_AO6;
  assign CLBLM_L_X10Y108_SLICE_X13Y108_C4 = CLBLM_L_X10Y106_SLICE_X13Y106_CO6;
  assign CLBLM_L_X10Y108_SLICE_X13Y108_C5 = CLBLM_L_X10Y108_SLICE_X13Y108_BO5;
  assign CLBLM_L_X10Y108_SLICE_X13Y108_C6 = CLBLM_R_X11Y106_SLICE_X14Y106_CO6;
  assign CLBLM_R_X11Y108_SLICE_X15Y108_C4 = CLBLM_R_X11Y105_SLICE_X15Y105_CO6;
  assign CLBLM_L_X10Y108_SLICE_X13Y108_D1 = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLM_L_X10Y108_SLICE_X13Y108_D2 = RIOB33_X105Y109_IOB_X1Y110_I;
  assign CLBLM_L_X10Y108_SLICE_X13Y108_D3 = RIOB33_X105Y111_IOB_X1Y111_I;
  assign CLBLM_L_X10Y108_SLICE_X13Y108_D4 = LIOB33_X0Y103_IOB_X0Y104_I;
  assign CLBLM_L_X10Y108_SLICE_X13Y108_D5 = LIOB33_X0Y105_IOB_X0Y105_I;
  assign CLBLM_L_X10Y108_SLICE_X13Y108_D6 = CLBLM_L_X10Y107_SLICE_X12Y107_BO6;
  assign CLBLM_L_X10Y108_SLICE_X12Y108_A1 = CLBLM_L_X10Y109_SLICE_X13Y109_AO5;
  assign CLBLM_L_X10Y108_SLICE_X12Y108_A2 = CLBLM_L_X8Y107_SLICE_X11Y107_AO5;
  assign CLBLM_L_X10Y108_SLICE_X12Y108_A3 = CLBLM_L_X10Y108_SLICE_X13Y108_CO6;
  assign CLBLM_L_X10Y108_SLICE_X12Y108_A4 = CLBLM_R_X11Y110_SLICE_X15Y110_AO6;
  assign CLBLM_L_X10Y108_SLICE_X12Y108_A5 = CLBLM_L_X10Y106_SLICE_X12Y106_DO6;
  assign CLBLM_L_X10Y108_SLICE_X12Y108_A6 = CLBLM_L_X10Y108_SLICE_X12Y108_CO6;
  assign CLBLM_L_X10Y108_SLICE_X12Y108_B1 = LIOB33_X0Y107_IOB_X0Y108_I;
  assign CLBLM_L_X10Y108_SLICE_X12Y108_B2 = RIOB33_X105Y101_IOB_X1Y101_I;
  assign CLBLM_L_X10Y108_SLICE_X12Y108_B3 = CLBLM_L_X10Y108_SLICE_X13Y108_CO6;
  assign CLBLM_L_X10Y108_SLICE_X12Y108_B4 = RIOB33_X105Y101_IOB_X1Y102_I;
  assign CLBLM_L_X10Y108_SLICE_X12Y108_B5 = CLBLM_L_X10Y106_SLICE_X12Y106_DO6;
  assign CLBLM_L_X10Y108_SLICE_X12Y108_B6 = CLBLM_L_X10Y108_SLICE_X12Y108_CO6;
  assign CLBLM_L_X10Y108_SLICE_X12Y108_C1 = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLM_L_X10Y108_SLICE_X12Y108_C2 = CLBLM_R_X11Y106_SLICE_X14Y106_DO6;
  assign CLBLM_L_X10Y108_SLICE_X12Y108_C3 = RIOB33_X105Y101_IOB_X1Y102_I;
  assign CLBLM_L_X10Y108_SLICE_X12Y108_C4 = CLBLM_L_X10Y106_SLICE_X13Y106_CO6;
  assign CLBLM_L_X10Y108_SLICE_X12Y108_C5 = RIOB33_X105Y103_IOB_X1Y103_I;
  assign CLBLM_L_X10Y108_SLICE_X12Y108_C6 = LIOB33_X0Y107_IOB_X0Y107_I;
  assign CLBLM_L_X10Y108_SLICE_X12Y108_D1 = CLBLM_L_X10Y106_SLICE_X12Y106_DO6;
  assign CLBLM_L_X10Y108_SLICE_X12Y108_D2 = CLBLM_L_X10Y108_SLICE_X13Y108_CO6;
  assign CLBLM_L_X10Y108_SLICE_X12Y108_D3 = CLBLM_L_X8Y107_SLICE_X11Y107_AO5;
  assign CLBLM_L_X10Y108_SLICE_X12Y108_D4 = CLBLM_L_X10Y108_SLICE_X12Y108_CO6;
  assign CLBLM_L_X10Y108_SLICE_X12Y108_D5 = CLBLM_L_X10Y109_SLICE_X13Y109_AO5;
  assign CLBLM_L_X10Y108_SLICE_X12Y108_D6 = CLBLM_R_X11Y110_SLICE_X15Y110_AO6;
  assign CLBLL_L_X4Y104_SLICE_X4Y104_A1 = CLBLL_L_X2Y104_SLICE_X0Y104_AO5;
  assign CLBLL_L_X4Y104_SLICE_X4Y104_A2 = CLBLM_R_X5Y104_SLICE_X6Y104_AO6;
  assign CLBLL_L_X4Y104_SLICE_X4Y104_A3 = CLBLL_L_X4Y103_SLICE_X4Y103_CO6;
  assign CLBLL_L_X4Y104_SLICE_X4Y104_A4 = CLBLL_L_X4Y103_SLICE_X4Y103_DO6;
  assign CLBLL_L_X4Y104_SLICE_X4Y104_A5 = CLBLL_L_X4Y103_SLICE_X5Y103_BO6;
  assign CLBLL_L_X4Y104_SLICE_X4Y104_A6 = CLBLM_R_X3Y104_SLICE_X3Y104_DO6;
  assign CLBLL_L_X4Y104_SLICE_X4Y104_B1 = CLBLL_L_X4Y103_SLICE_X4Y103_BO6;
  assign CLBLL_L_X4Y104_SLICE_X4Y104_B2 = LIOB33_X0Y103_IOB_X0Y103_I;
  assign CLBLL_L_X4Y104_SLICE_X4Y104_B3 = LIOB33_X0Y103_IOB_X0Y104_I;
  assign CLBLL_L_X4Y104_SLICE_X4Y104_B4 = LIOB33_X0Y113_IOB_X0Y114_I;
  assign CLBLL_L_X4Y104_SLICE_X4Y104_B5 = LIOB33_X0Y101_IOB_X0Y102_I;
  assign CLBLL_L_X4Y104_SLICE_X4Y104_B6 = CLBLM_R_X3Y104_SLICE_X3Y104_DO6;
  assign CLBLL_L_X4Y104_SLICE_X4Y104_C1 = LIOB33_X0Y101_IOB_X0Y102_I;
  assign CLBLL_L_X4Y104_SLICE_X4Y104_C2 = LIOB33_X0Y113_IOB_X0Y114_I;
  assign CLBLL_L_X4Y104_SLICE_X4Y104_C3 = CLBLL_L_X4Y103_SLICE_X4Y103_BO6;
  assign CLBLL_L_X4Y104_SLICE_X4Y104_C4 = LIOB33_X0Y103_IOB_X0Y104_I;
  assign CLBLL_L_X4Y104_SLICE_X4Y104_C5 = LIOB33_X0Y103_IOB_X0Y103_I;
  assign CLBLL_L_X4Y104_SLICE_X4Y104_C6 = CLBLM_R_X3Y104_SLICE_X3Y104_DO6;
  assign CLBLL_L_X4Y104_SLICE_X4Y104_D1 = LIOB33_X0Y115_IOB_X0Y116_I;
  assign CLBLL_L_X4Y104_SLICE_X4Y104_D2 = CLBLL_L_X4Y104_SLICE_X5Y104_CO6;
  assign CLBLL_L_X4Y104_SLICE_X4Y104_D3 = CLBLL_L_X4Y104_SLICE_X5Y104_AO6;
  assign CLBLL_L_X4Y104_SLICE_X4Y104_D4 = LIOB33_X0Y113_IOB_X0Y114_I;
  assign CLBLL_L_X4Y104_SLICE_X4Y104_D5 = LIOB33_X0Y101_IOB_X0Y102_I;
  assign CLBLL_L_X4Y104_SLICE_X4Y104_D6 = CLBLM_R_X3Y103_SLICE_X3Y103_AO5;
  assign CLBLL_L_X4Y104_SLICE_X5Y104_A1 = 1'b1;
  assign CLBLL_L_X4Y104_SLICE_X5Y104_A2 = LIOB33_X0Y101_IOB_X0Y101_I;
  assign CLBLL_L_X4Y104_SLICE_X5Y104_A3 = LIOB33_X0Y115_IOB_X0Y116_I;
  assign CLBLL_L_X4Y104_SLICE_X5Y104_A4 = CLBLL_L_X4Y104_SLICE_X5Y104_BO6;
  assign CLBLL_L_X4Y104_SLICE_X5Y104_A5 = CLBLM_R_X5Y104_SLICE_X6Y104_BO6;
  assign CLBLL_L_X4Y104_SLICE_X5Y104_A6 = 1'b1;
  assign CLBLL_L_X4Y104_SLICE_X5Y104_B1 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLL_L_X4Y104_SLICE_X5Y104_B2 = RIOB33_X105Y111_IOB_X1Y112_I;
  assign CLBLL_L_X4Y104_SLICE_X5Y104_B3 = LIOB33_SING_X0Y100_IOB_X0Y100_I;
  assign CLBLL_L_X4Y104_SLICE_X5Y104_B4 = RIOB33_X105Y113_IOB_X1Y113_I;
  assign CLBLL_L_X4Y104_SLICE_X5Y104_B5 = LIOB33_X0Y115_IOB_X0Y116_I;
  assign CLBLL_L_X4Y104_SLICE_X5Y104_B6 = RIOB33_X105Y101_IOB_X1Y101_I;
  assign CLBLL_L_X4Y104_SLICE_X5Y104_C1 = CLBLM_R_X5Y104_SLICE_X6Y104_BO6;
  assign CLBLL_L_X4Y104_SLICE_X5Y104_C2 = CLBLM_R_X7Y103_SLICE_X8Y103_AO6;
  assign CLBLL_L_X4Y104_SLICE_X5Y104_C3 = LIOB33_X0Y101_IOB_X0Y101_I;
  assign CLBLL_L_X4Y104_SLICE_X5Y104_C4 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLL_L_X4Y104_SLICE_X5Y104_C5 = LIOB33_X0Y115_IOB_X0Y116_I;
  assign CLBLL_L_X4Y104_SLICE_X5Y104_C6 = CLBLL_L_X4Y104_SLICE_X5Y104_BO6;
  assign CLBLL_L_X4Y104_SLICE_X5Y104_D1 = CLBLM_R_X5Y104_SLICE_X6Y104_AO6;
  assign CLBLL_L_X4Y104_SLICE_X5Y104_D2 = CLBLL_L_X4Y103_SLICE_X4Y103_DO6;
  assign CLBLL_L_X4Y104_SLICE_X5Y104_D3 = CLBLL_L_X4Y103_SLICE_X5Y103_BO6;
  assign CLBLL_L_X4Y104_SLICE_X5Y104_D4 = CLBLL_L_X4Y103_SLICE_X5Y103_CO6;
  assign CLBLL_L_X4Y104_SLICE_X5Y104_D5 = CLBLM_R_X5Y104_SLICE_X6Y104_AO5;
  assign CLBLL_L_X4Y104_SLICE_X5Y104_D6 = CLBLM_R_X7Y104_SLICE_X8Y104_CO6;
  assign LIOI3_X0Y101_ILOGIC_X0Y102_D = LIOB33_X0Y101_IOB_X0Y102_I;
  assign LIOI3_X0Y101_ILOGIC_X0Y101_D = LIOB33_X0Y101_IOB_X0Y101_I;
  assign CLBLM_L_X10Y109_SLICE_X13Y109_A1 = 1'b1;
  assign CLBLM_L_X10Y109_SLICE_X13Y109_A2 = 1'b1;
  assign CLBLM_L_X10Y109_SLICE_X13Y109_A3 = RIOB33_X105Y101_IOB_X1Y101_I;
  assign CLBLM_L_X10Y109_SLICE_X13Y109_A4 = LIOB33_X0Y109_IOB_X0Y109_I;
  assign CLBLM_L_X10Y109_SLICE_X13Y109_A5 = RIOB33_X105Y101_IOB_X1Y102_I;
  assign CLBLM_L_X10Y109_SLICE_X13Y109_A6 = 1'b1;
  assign CLBLM_L_X10Y109_SLICE_X13Y109_B1 = RIOB33_X105Y101_IOB_X1Y102_I;
  assign CLBLM_L_X10Y109_SLICE_X13Y109_B2 = CLBLM_R_X11Y106_SLICE_X14Y106_DO6;
  assign CLBLM_L_X10Y109_SLICE_X13Y109_B3 = RIOB33_X105Y103_IOB_X1Y103_I;
  assign CLBLM_L_X10Y109_SLICE_X13Y109_B4 = LIOB33_X0Y107_IOB_X0Y107_I;
  assign CLBLM_L_X10Y109_SLICE_X13Y109_B5 = CLBLM_L_X10Y106_SLICE_X13Y106_CO6;
  assign CLBLM_L_X10Y109_SLICE_X13Y109_B6 = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLM_L_X10Y109_SLICE_X13Y109_C1 = RIOB33_X105Y101_IOB_X1Y102_I;
  assign CLBLM_L_X10Y109_SLICE_X13Y109_C2 = CLBLM_R_X11Y106_SLICE_X14Y106_DO6;
  assign CLBLM_L_X10Y109_SLICE_X13Y109_C3 = CLBLM_L_X10Y105_SLICE_X13Y105_DO6;
  assign CLBLM_L_X10Y109_SLICE_X13Y109_C4 = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLM_L_X10Y109_SLICE_X13Y109_C5 = CLBLM_R_X11Y108_SLICE_X14Y108_DO6;
  assign CLBLM_L_X10Y109_SLICE_X13Y109_C6 = RIOB33_X105Y103_IOB_X1Y103_I;
  assign CLBLM_L_X10Y109_SLICE_X13Y109_D1 = CLBLM_R_X11Y109_SLICE_X15Y109_AO6;
  assign CLBLM_L_X10Y109_SLICE_X13Y109_D2 = RIOB33_X105Y103_IOB_X1Y103_I;
  assign CLBLM_L_X10Y109_SLICE_X13Y109_D3 = LIOB33_X0Y107_IOB_X0Y108_I;
  assign CLBLM_L_X10Y109_SLICE_X13Y109_D4 = CLBLM_R_X11Y109_SLICE_X14Y109_CO6;
  assign CLBLM_L_X10Y109_SLICE_X13Y109_D5 = RIOB33_X105Y101_IOB_X1Y102_I;
  assign CLBLM_L_X10Y109_SLICE_X13Y109_D6 = CLBLM_L_X10Y109_SLICE_X13Y109_BO6;
  assign CLBLM_L_X10Y109_SLICE_X12Y109_A1 = LIOB33_X0Y107_IOB_X0Y108_I;
  assign CLBLM_L_X10Y109_SLICE_X12Y109_A2 = CLBLM_L_X10Y106_SLICE_X12Y106_DO6;
  assign CLBLM_L_X10Y109_SLICE_X12Y109_A3 = RIOB33_X105Y101_IOB_X1Y102_I;
  assign CLBLM_L_X10Y109_SLICE_X12Y109_A4 = CLBLM_L_X10Y109_SLICE_X13Y109_CO6;
  assign CLBLM_L_X10Y109_SLICE_X12Y109_A5 = RIOB33_X105Y101_IOB_X1Y101_I;
  assign CLBLM_L_X10Y109_SLICE_X12Y109_A6 = LIOB33_X0Y107_IOB_X0Y107_I;
  assign CLBLM_L_X10Y109_SLICE_X12Y109_B1 = LIOB33_X0Y107_IOB_X0Y108_I;
  assign CLBLM_L_X10Y109_SLICE_X12Y109_B2 = CLBLM_L_X10Y106_SLICE_X12Y106_DO6;
  assign CLBLM_L_X10Y109_SLICE_X12Y109_B3 = RIOB33_X105Y101_IOB_X1Y102_I;
  assign CLBLM_L_X10Y109_SLICE_X12Y109_B4 = CLBLM_L_X10Y109_SLICE_X13Y109_CO6;
  assign CLBLM_L_X10Y109_SLICE_X12Y109_B5 = RIOB33_X105Y101_IOB_X1Y101_I;
  assign CLBLM_L_X10Y109_SLICE_X12Y109_B6 = LIOB33_X0Y107_IOB_X0Y107_I;
  assign CLBLM_L_X10Y109_SLICE_X12Y109_C1 = CLBLM_L_X10Y107_SLICE_X12Y107_BO6;
  assign CLBLM_L_X10Y109_SLICE_X12Y109_C2 = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLM_L_X10Y109_SLICE_X12Y109_C3 = LIOB33_X0Y105_IOB_X0Y105_I;
  assign CLBLM_L_X10Y109_SLICE_X12Y109_C4 = RIOB33_X105Y111_IOB_X1Y111_I;
  assign CLBLM_L_X10Y109_SLICE_X12Y109_C5 = RIOB33_X105Y109_IOB_X1Y110_I;
  assign CLBLM_L_X10Y109_SLICE_X12Y109_C6 = LIOB33_X0Y103_IOB_X0Y104_I;
  assign CLBLM_L_X10Y109_SLICE_X12Y109_D1 = CLBLM_L_X10Y107_SLICE_X12Y107_BO6;
  assign CLBLM_L_X10Y109_SLICE_X12Y109_D2 = RIOB33_X105Y109_IOB_X1Y110_I;
  assign CLBLM_L_X10Y109_SLICE_X12Y109_D3 = LIOB33_X0Y105_IOB_X0Y105_I;
  assign CLBLM_L_X10Y109_SLICE_X12Y109_D4 = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLM_L_X10Y109_SLICE_X12Y109_D5 = RIOB33_X105Y111_IOB_X1Y111_I;
  assign CLBLL_L_X4Y105_SLICE_X4Y105_A1 = CLBLL_L_X4Y104_SLICE_X5Y104_DO6;
  assign CLBLL_L_X4Y105_SLICE_X4Y105_A2 = LIOB33_X0Y113_IOB_X0Y114_I;
  assign CLBLL_L_X4Y105_SLICE_X4Y105_A3 = LIOB33_X0Y105_IOB_X0Y105_I;
  assign CLBLL_L_X4Y105_SLICE_X4Y105_A4 = CLBLL_L_X4Y105_SLICE_X4Y105_BO6;
  assign CLBLL_L_X4Y105_SLICE_X4Y105_A5 = LIOB33_X0Y103_IOB_X0Y103_I;
  assign CLBLL_L_X4Y105_SLICE_X4Y105_A6 = CLBLL_L_X4Y104_SLICE_X4Y104_CO6;
  assign CLBLM_L_X10Y109_SLICE_X12Y109_D6 = LIOB33_X0Y103_IOB_X0Y104_I;
  assign CLBLL_L_X4Y105_SLICE_X4Y105_B1 = LIOB33_X0Y101_IOB_X0Y102_I;
  assign CLBLL_L_X4Y105_SLICE_X4Y105_B2 = LIOB33_X0Y103_IOB_X0Y104_I;
  assign CLBLL_L_X4Y105_SLICE_X4Y105_B3 = CLBLL_L_X4Y103_SLICE_X4Y103_DO6;
  assign CLBLL_L_X4Y105_SLICE_X4Y105_B4 = LIOB33_X0Y113_IOB_X0Y114_I;
  assign CLBLL_L_X4Y105_SLICE_X4Y105_B5 = LIOB33_X0Y115_IOB_X0Y116_I;
  assign CLBLL_L_X4Y105_SLICE_X4Y105_B6 = CLBLL_L_X4Y104_SLICE_X5Y104_CO6;
  assign CLBLL_L_X4Y105_SLICE_X4Y105_C1 = 1'b1;
  assign CLBLL_L_X4Y105_SLICE_X4Y105_C2 = 1'b1;
  assign CLBLL_L_X4Y105_SLICE_X4Y105_C3 = 1'b1;
  assign CLBLL_L_X4Y105_SLICE_X4Y105_C4 = 1'b1;
  assign CLBLL_L_X4Y105_SLICE_X4Y105_C5 = 1'b1;
  assign CLBLL_L_X4Y105_SLICE_X4Y105_C6 = 1'b1;
  assign CLBLL_L_X4Y105_SLICE_X4Y105_D1 = 1'b1;
  assign CLBLL_L_X4Y105_SLICE_X4Y105_D2 = 1'b1;
  assign CLBLL_L_X4Y105_SLICE_X4Y105_D3 = 1'b1;
  assign CLBLL_L_X4Y105_SLICE_X4Y105_D4 = 1'b1;
  assign CLBLL_L_X4Y105_SLICE_X4Y105_D5 = 1'b1;
  assign CLBLL_L_X4Y105_SLICE_X4Y105_D6 = 1'b1;
  assign LIOI3_TBYTETERM_X0Y137_OLOGIC_X0Y138_D1 = CLBLL_L_X4Y111_SLICE_X4Y111_AO5;
  assign CLBLL_L_X4Y105_SLICE_X5Y105_A1 = LIOB33_X0Y101_IOB_X0Y102_I;
  assign CLBLL_L_X4Y105_SLICE_X5Y105_A2 = LIOB33_X0Y103_IOB_X0Y104_I;
  assign CLBLL_L_X4Y105_SLICE_X5Y105_A3 = LIOB33_X0Y115_IOB_X0Y116_I;
  assign CLBLL_L_X4Y105_SLICE_X5Y105_A4 = LIOB33_X0Y113_IOB_X0Y114_I;
  assign CLBLL_L_X4Y105_SLICE_X5Y105_A5 = CLBLL_L_X4Y103_SLICE_X4Y103_DO6;
  assign CLBLL_L_X4Y105_SLICE_X5Y105_A6 = CLBLL_L_X4Y104_SLICE_X5Y104_CO6;
  assign CLBLL_L_X4Y105_SLICE_X5Y105_B1 = CLBLL_L_X4Y104_SLICE_X5Y104_DO6;
  assign CLBLL_L_X4Y105_SLICE_X5Y105_B2 = CLBLL_L_X4Y105_SLICE_X4Y105_BO6;
  assign CLBLL_L_X4Y105_SLICE_X5Y105_B3 = CLBLM_R_X3Y106_SLICE_X3Y106_AO6;
  assign CLBLL_L_X4Y105_SLICE_X5Y105_B4 = CLBLL_L_X4Y104_SLICE_X4Y104_CO6;
  assign CLBLL_L_X4Y105_SLICE_X5Y105_B5 = CLBLM_R_X5Y106_SLICE_X7Y106_AO5;
  assign CLBLL_L_X4Y105_SLICE_X5Y105_B6 = CLBLM_R_X5Y105_SLICE_X7Y105_AO5;
  assign CLBLL_L_X4Y105_SLICE_X5Y105_C1 = 1'b1;
  assign CLBLL_L_X4Y105_SLICE_X5Y105_C2 = 1'b1;
  assign CLBLL_L_X4Y105_SLICE_X5Y105_C3 = 1'b1;
  assign CLBLL_L_X4Y105_SLICE_X5Y105_C4 = 1'b1;
  assign CLBLL_L_X4Y105_SLICE_X5Y105_C5 = 1'b1;
  assign CLBLL_L_X4Y105_SLICE_X5Y105_C6 = 1'b1;
  assign CLBLL_L_X4Y105_SLICE_X5Y105_D1 = 1'b1;
  assign CLBLL_L_X4Y105_SLICE_X5Y105_D2 = 1'b1;
  assign CLBLL_L_X4Y105_SLICE_X5Y105_D3 = 1'b1;
  assign CLBLL_L_X4Y105_SLICE_X5Y105_D4 = 1'b1;
  assign CLBLL_L_X4Y105_SLICE_X5Y105_D5 = 1'b1;
  assign CLBLL_L_X4Y105_SLICE_X5Y105_D6 = 1'b1;
  assign LIOI3_TBYTETERM_X0Y137_OLOGIC_X0Y138_T1 = 1'b1;
  assign CLBLM_L_X8Y104_SLICE_X10Y104_A2 = 1'b1;
  assign LIOI3_TBYTETERM_X0Y137_OLOGIC_X0Y137_D1 = CLBLL_L_X4Y111_SLICE_X4Y111_AO6;
  assign CLBLM_L_X8Y104_SLICE_X10Y104_B4 = CLBLM_L_X10Y102_SLICE_X12Y102_AO6;
  assign CLBLM_L_X8Y104_SLICE_X10Y104_B6 = CLBLM_L_X8Y104_SLICE_X10Y104_AO5;
  assign CLBLM_L_X10Y110_SLICE_X13Y110_A1 = LIOB33_X0Y109_IOB_X0Y110_I;
  assign CLBLM_L_X10Y110_SLICE_X13Y110_A2 = 1'b1;
  assign CLBLM_L_X10Y110_SLICE_X13Y110_A3 = 1'b1;
  assign CLBLM_L_X10Y110_SLICE_X13Y110_A4 = RIOB33_X105Y101_IOB_X1Y101_I;
  assign CLBLM_L_X10Y110_SLICE_X13Y110_A5 = RIOB33_X105Y101_IOB_X1Y102_I;
  assign CLBLM_L_X10Y110_SLICE_X13Y110_A6 = 1'b1;
  assign CLBLM_L_X10Y110_SLICE_X13Y110_B1 = CLBLM_L_X10Y108_SLICE_X12Y108_DO6;
  assign CLBLM_L_X10Y110_SLICE_X13Y110_B2 = CLBLM_R_X11Y110_SLICE_X14Y110_BO6;
  assign CLBLM_L_X10Y110_SLICE_X13Y110_B3 = CLBLM_R_X11Y109_SLICE_X14Y109_DO6;
  assign CLBLM_L_X10Y110_SLICE_X13Y110_B4 = CLBLM_R_X11Y109_SLICE_X14Y109_BO6;
  assign CLBLM_L_X10Y110_SLICE_X13Y110_B5 = CLBLM_L_X10Y110_SLICE_X13Y110_AO6;
  assign CLBLM_L_X10Y110_SLICE_X13Y110_B6 = CLBLM_L_X10Y110_SLICE_X13Y110_AO5;
  assign CLBLM_L_X10Y110_SLICE_X13Y110_C1 = CLBLM_R_X11Y110_SLICE_X14Y110_BO6;
  assign CLBLM_L_X10Y110_SLICE_X13Y110_C2 = CLBLM_R_X11Y110_SLICE_X14Y110_AO5;
  assign CLBLM_L_X10Y110_SLICE_X13Y110_C3 = CLBLM_L_X10Y111_SLICE_X13Y111_BO6;
  assign CLBLM_L_X10Y110_SLICE_X13Y110_C4 = CLBLM_L_X10Y110_SLICE_X13Y110_AO5;
  assign CLBLM_L_X10Y110_SLICE_X13Y110_C5 = CLBLM_R_X11Y109_SLICE_X14Y109_DO6;
  assign CLBLM_L_X10Y110_SLICE_X13Y110_C6 = CLBLM_R_X11Y110_SLICE_X14Y110_DO6;
  assign CLBLM_L_X10Y110_SLICE_X13Y110_D1 = CLBLM_L_X12Y108_SLICE_X16Y108_BO6;
  assign CLBLM_L_X10Y110_SLICE_X13Y110_D2 = LIOB33_X0Y107_IOB_X0Y107_I;
  assign CLBLM_L_X10Y110_SLICE_X13Y110_D3 = LIOB33_X0Y107_IOB_X0Y108_I;
  assign CLBLM_L_X10Y110_SLICE_X13Y110_D4 = CLBLM_L_X10Y107_SLICE_X13Y107_AO6;
  assign CLBLM_L_X10Y110_SLICE_X13Y110_D5 = RIOB33_X105Y107_IOB_X1Y108_I;
  assign CLBLM_L_X10Y110_SLICE_X13Y110_D6 = CLBLM_L_X10Y107_SLICE_X13Y107_BO6;
  assign CLBLM_L_X10Y110_SLICE_X12Y110_A1 = LIOB33_X0Y107_IOB_X0Y108_I;
  assign CLBLM_L_X10Y110_SLICE_X12Y110_A2 = CLBLM_R_X11Y108_SLICE_X14Y108_AO6;
  assign CLBLM_L_X10Y110_SLICE_X12Y110_A3 = RIOB33_X105Y103_IOB_X1Y103_I;
  assign CLBLM_L_X10Y110_SLICE_X12Y110_A4 = CLBLM_L_X10Y109_SLICE_X13Y109_BO6;
  assign CLBLM_L_X10Y110_SLICE_X12Y110_A5 = RIOB33_X105Y101_IOB_X1Y102_I;
  assign CLBLM_L_X10Y110_SLICE_X12Y110_A6 = LIOB33_X0Y107_IOB_X0Y107_I;
  assign CLBLM_L_X10Y110_SLICE_X12Y110_B1 = RIOB33_X105Y101_IOB_X1Y101_I;
  assign CLBLM_L_X10Y110_SLICE_X12Y110_B2 = CLBLM_L_X10Y109_SLICE_X12Y109_AO6;
  assign CLBLM_L_X10Y110_SLICE_X12Y110_B3 = RIOB33_X105Y101_IOB_X1Y102_I;
  assign CLBLM_L_X10Y110_SLICE_X12Y110_B4 = LIOB33_X0Y109_IOB_X0Y109_I;
  assign CLBLM_L_X10Y110_SLICE_X12Y110_B5 = CLBLM_L_X10Y110_SLICE_X12Y110_AO6;
  assign CLBLM_L_X10Y110_SLICE_X12Y110_B6 = CLBLM_L_X10Y109_SLICE_X13Y109_DO6;
  assign CLBLM_L_X10Y110_SLICE_X12Y110_C1 = RIOB33_X105Y101_IOB_X1Y102_I;
  assign CLBLM_L_X10Y110_SLICE_X12Y110_C2 = LIOB33_X0Y107_IOB_X0Y107_I;
  assign CLBLM_L_X10Y110_SLICE_X12Y110_C3 = LIOB33_X0Y107_IOB_X0Y108_I;
  assign CLBLM_L_X10Y110_SLICE_X12Y110_C4 = CLBLM_R_X11Y108_SLICE_X14Y108_AO6;
  assign CLBLM_L_X10Y110_SLICE_X12Y110_C5 = RIOB33_X105Y103_IOB_X1Y103_I;
  assign CLBLM_L_X10Y110_SLICE_X12Y110_C6 = CLBLM_L_X10Y109_SLICE_X13Y109_BO6;
  assign CLBLL_L_X4Y106_SLICE_X4Y106_A1 = CLBLL_L_X4Y104_SLICE_X4Y104_DO6;
  assign CLBLL_L_X4Y106_SLICE_X4Y106_A2 = LIOB33_X0Y103_IOB_X0Y104_I;
  assign CLBLL_L_X4Y106_SLICE_X4Y106_A3 = LIOB33_X0Y105_IOB_X0Y105_I;
  assign CLBLL_L_X4Y106_SLICE_X4Y106_A4 = LIOB33_X0Y113_IOB_X0Y114_I;
  assign CLBLL_L_X4Y106_SLICE_X4Y106_A5 = LIOB33_X0Y103_IOB_X0Y103_I;
  assign CLBLL_L_X4Y106_SLICE_X4Y106_A6 = CLBLL_L_X4Y104_SLICE_X4Y104_CO6;
  assign CLBLM_L_X10Y110_SLICE_X12Y110_D1 = RIOB33_X105Y101_IOB_X1Y102_I;
  assign CLBLM_L_X10Y110_SLICE_X12Y110_D2 = LIOB33_X0Y109_IOB_X0Y109_I;
  assign CLBLM_L_X10Y110_SLICE_X12Y110_D3 = CLBLM_R_X11Y110_SLICE_X14Y110_CO6;
  assign CLBLL_L_X4Y106_SLICE_X4Y106_B1 = CLBLL_L_X4Y106_SLICE_X4Y106_DO6;
  assign CLBLL_L_X4Y106_SLICE_X4Y106_B2 = CLBLM_R_X5Y105_SLICE_X6Y105_BO6;
  assign CLBLL_L_X4Y106_SLICE_X4Y106_B3 = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLL_L_X4Y106_SLICE_X4Y106_B4 = LIOB33_X0Y103_IOB_X0Y103_I;
  assign CLBLL_L_X4Y106_SLICE_X4Y106_B5 = CLBLM_R_X5Y105_SLICE_X6Y105_AO6;
  assign CLBLL_L_X4Y106_SLICE_X4Y106_B6 = LIOB33_X0Y113_IOB_X0Y114_I;
  assign CLBLL_L_X4Y106_SLICE_X4Y106_C1 = LIOB33_X0Y103_IOB_X0Y103_I;
  assign CLBLL_L_X4Y106_SLICE_X4Y106_C2 = CLBLL_L_X4Y105_SLICE_X4Y105_AO6;
  assign CLBLL_L_X4Y106_SLICE_X4Y106_C3 = RIOB33_X105Y105_IOB_X1Y106_I;
  assign CLBLL_L_X4Y106_SLICE_X4Y106_C4 = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLL_L_X4Y106_SLICE_X4Y106_C5 = LIOB33_X0Y107_IOB_X0Y107_I;
  assign CLBLL_L_X4Y106_SLICE_X4Y106_C6 = CLBLM_R_X3Y106_SLICE_X3Y106_DO6;
  assign CLBLL_L_X4Y106_SLICE_X4Y106_D1 = LIOB33_X0Y105_IOB_X0Y105_I;
  assign CLBLL_L_X4Y106_SLICE_X4Y106_D2 = LIOB33_X0Y103_IOB_X0Y103_I;
  assign CLBLL_L_X4Y106_SLICE_X4Y106_D3 = CLBLL_L_X4Y104_SLICE_X4Y104_DO6;
  assign CLBLL_L_X4Y106_SLICE_X4Y106_D4 = CLBLL_L_X4Y104_SLICE_X4Y104_CO6;
  assign CLBLL_L_X4Y106_SLICE_X4Y106_D5 = LIOB33_X0Y103_IOB_X0Y104_I;
  assign CLBLL_L_X4Y106_SLICE_X4Y106_D6 = LIOB33_X0Y113_IOB_X0Y114_I;
  assign CLBLM_R_X11Y104_SLICE_X15Y104_A1 = RIOB33_X105Y103_IOB_X1Y104_I;
  assign CLBLM_R_X11Y104_SLICE_X15Y104_A2 = 1'b1;
  assign CLBLM_R_X11Y104_SLICE_X15Y104_A3 = LIOB33_X0Y101_IOB_X0Y101_I;
  assign CLBLM_R_X11Y104_SLICE_X15Y104_A4 = CLBLM_R_X11Y104_SLICE_X15Y104_BO6;
  assign CLBLM_R_X11Y104_SLICE_X15Y104_A5 = CLBLM_R_X11Y104_SLICE_X15Y104_DO6;
  assign CLBLM_R_X11Y104_SLICE_X15Y104_A6 = 1'b1;
  assign CLBLL_L_X4Y106_SLICE_X5Y106_A1 = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLL_L_X4Y106_SLICE_X5Y106_A2 = LIOB33_X0Y113_IOB_X0Y114_I;
  assign CLBLL_L_X4Y106_SLICE_X5Y106_A3 = CLBLM_R_X5Y105_SLICE_X6Y105_AO6;
  assign CLBLL_L_X4Y106_SLICE_X5Y106_A4 = CLBLL_L_X4Y105_SLICE_X5Y105_BO6;
  assign CLBLL_L_X4Y106_SLICE_X5Y106_A5 = LIOB33_X0Y107_IOB_X0Y107_I;
  assign CLBLL_L_X4Y106_SLICE_X5Y106_A6 = LIOB33_X0Y103_IOB_X0Y103_I;
  assign CLBLM_R_X11Y104_SLICE_X15Y104_B1 = RIOB33_X105Y107_IOB_X1Y107_I;
  assign CLBLM_R_X11Y104_SLICE_X15Y104_B2 = RIOB33_X105Y111_IOB_X1Y112_I;
  assign CLBLM_R_X11Y104_SLICE_X15Y104_B3 = RIOB33_X105Y103_IOB_X1Y104_I;
  assign CLBLL_L_X4Y106_SLICE_X5Y106_B1 = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLL_L_X4Y106_SLICE_X5Y106_B2 = CLBLL_L_X4Y105_SLICE_X5Y105_BO6;
  assign CLBLL_L_X4Y106_SLICE_X5Y106_B3 = CLBLM_R_X5Y105_SLICE_X6Y105_AO6;
  assign CLBLL_L_X4Y106_SLICE_X5Y106_B4 = LIOB33_X0Y113_IOB_X0Y114_I;
  assign CLBLL_L_X4Y106_SLICE_X5Y106_B5 = LIOB33_X0Y107_IOB_X0Y107_I;
  assign CLBLL_L_X4Y106_SLICE_X5Y106_B6 = LIOB33_X0Y103_IOB_X0Y103_I;
  assign CLBLM_R_X11Y104_SLICE_X15Y104_C1 = LIOB33_SING_X0Y100_IOB_X0Y100_I;
  assign CLBLM_R_X11Y104_SLICE_X15Y104_C2 = RIOB33_X105Y113_IOB_X1Y113_I;
  assign CLBLL_L_X4Y106_SLICE_X5Y106_C1 = LIOB33_X0Y107_IOB_X0Y107_I;
  assign CLBLL_L_X4Y106_SLICE_X5Y106_C2 = CLBLM_R_X5Y105_SLICE_X6Y105_CO6;
  assign CLBLL_L_X4Y106_SLICE_X5Y106_C3 = LIOB33_X0Y113_IOB_X0Y114_I;
  assign CLBLL_L_X4Y106_SLICE_X5Y106_C4 = LIOB33_X0Y107_IOB_X0Y108_I;
  assign CLBLL_L_X4Y106_SLICE_X5Y106_C5 = LIOB33_X0Y103_IOB_X0Y103_I;
  assign CLBLL_L_X4Y106_SLICE_X5Y106_C6 = CLBLL_L_X4Y106_SLICE_X5Y106_BO6;
  assign CLBLM_R_X11Y104_SLICE_X15Y104_D1 = RIOB33_X105Y113_IOB_X1Y113_I;
  assign CLBLM_R_X11Y104_SLICE_X15Y104_D2 = LIOB33_SING_X0Y100_IOB_X0Y100_I;
  assign CLBLM_R_X11Y104_SLICE_X15Y104_D3 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X11Y104_SLICE_X15Y104_D4 = RIOB33_X105Y107_IOB_X1Y107_I;
  assign CLBLM_R_X11Y104_SLICE_X15Y104_D5 = RIOB33_X105Y103_IOB_X1Y104_I;
  assign CLBLM_R_X11Y104_SLICE_X15Y104_D6 = RIOB33_X105Y111_IOB_X1Y112_I;
  assign CLBLL_L_X4Y106_SLICE_X5Y106_D1 = LIOB33_X0Y113_IOB_X0Y114_I;
  assign CLBLL_L_X4Y106_SLICE_X5Y106_D2 = CLBLM_R_X5Y105_SLICE_X6Y105_CO6;
  assign CLBLL_L_X4Y106_SLICE_X5Y106_D3 = LIOB33_X0Y107_IOB_X0Y107_I;
  assign CLBLL_L_X4Y106_SLICE_X5Y106_D4 = LIOB33_X0Y107_IOB_X0Y108_I;
  assign CLBLL_L_X4Y106_SLICE_X5Y106_D5 = LIOB33_X0Y103_IOB_X0Y103_I;
  assign CLBLL_L_X4Y106_SLICE_X5Y106_D6 = CLBLL_L_X4Y106_SLICE_X5Y106_BO6;
  assign CLBLM_R_X11Y104_SLICE_X14Y104_A1 = 1'b1;
  assign CLBLM_R_X11Y104_SLICE_X14Y104_A2 = LIOB33_X0Y101_IOB_X0Y101_I;
  assign CLBLM_R_X11Y104_SLICE_X14Y104_A3 = 1'b1;
  assign CLBLM_R_X11Y104_SLICE_X14Y104_A4 = LIOB33_X0Y101_IOB_X0Y102_I;
  assign CLBLM_R_X11Y104_SLICE_X14Y104_A5 = RIOB33_X105Y103_IOB_X1Y104_I;
  assign CLBLM_R_X11Y104_SLICE_X14Y104_A6 = 1'b1;
  assign CLBLM_R_X11Y104_SLICE_X14Y104_B1 = CLBLM_R_X11Y104_SLICE_X15Y104_CO6;
  assign CLBLM_R_X11Y104_SLICE_X14Y104_B2 = CLBLM_R_X11Y104_SLICE_X15Y104_BO6;
  assign CLBLM_R_X11Y104_SLICE_X14Y104_B3 = CLBLM_R_X11Y104_SLICE_X15Y104_DO6;
  assign CLBLM_R_X11Y104_SLICE_X14Y104_B4 = CLBLM_L_X12Y104_SLICE_X16Y104_AO6;
  assign CLBLM_R_X11Y104_SLICE_X14Y104_B5 = CLBLM_R_X11Y104_SLICE_X14Y104_AO6;
  assign CLBLM_R_X11Y104_SLICE_X14Y104_B6 = CLBLM_R_X11Y104_SLICE_X14Y104_AO5;
  assign CLBLM_R_X11Y104_SLICE_X14Y104_C1 = CLBLM_R_X11Y104_SLICE_X14Y104_AO6;
  assign CLBLM_R_X11Y104_SLICE_X14Y104_C2 = CLBLM_R_X11Y104_SLICE_X15Y104_CO6;
  assign CLBLM_R_X11Y104_SLICE_X14Y104_C3 = CLBLM_R_X11Y104_SLICE_X15Y104_DO6;
  assign CLBLM_R_X11Y104_SLICE_X14Y104_C4 = CLBLM_R_X11Y104_SLICE_X14Y104_AO5;
  assign CLBLM_R_X11Y104_SLICE_X14Y104_C5 = CLBLM_R_X11Y104_SLICE_X15Y104_BO6;
  assign CLBLM_R_X11Y104_SLICE_X14Y104_C6 = CLBLM_L_X12Y104_SLICE_X16Y104_AO6;
  assign CLBLM_R_X11Y104_SLICE_X14Y104_D1 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X11Y104_SLICE_X14Y104_D2 = CLBLM_R_X11Y104_SLICE_X15Y104_CO6;
  assign CLBLM_R_X11Y104_SLICE_X14Y104_D3 = CLBLM_R_X11Y104_SLICE_X15Y104_DO6;
  assign CLBLM_R_X11Y104_SLICE_X14Y104_D4 = CLBLM_R_X11Y104_SLICE_X15Y104_BO6;
  assign CLBLM_R_X11Y104_SLICE_X14Y104_D5 = RIOB33_X105Y103_IOB_X1Y104_I;
  assign CLBLM_R_X11Y104_SLICE_X14Y104_D6 = LIOB33_X0Y101_IOB_X0Y101_I;
  assign CLBLM_L_X10Y111_SLICE_X13Y111_A1 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X10Y111_SLICE_X13Y111_A2 = LIOB33_X0Y107_IOB_X0Y108_I;
  assign CLBLM_L_X10Y111_SLICE_X13Y111_A3 = LIOB33_X0Y109_IOB_X0Y110_I;
  assign CLBLM_L_X10Y111_SLICE_X13Y111_A4 = 1'b1;
  assign CLBLM_L_X10Y111_SLICE_X13Y111_A5 = 1'b1;
  assign CLBLM_L_X10Y111_SLICE_X13Y111_A6 = 1'b1;
  assign CLBLM_L_X10Y111_SLICE_X13Y111_B1 = CLBLM_R_X11Y111_SLICE_X15Y111_DO6;
  assign CLBLM_L_X10Y111_SLICE_X13Y111_B2 = CLBLM_R_X11Y110_SLICE_X15Y110_AO5;
  assign CLBLM_L_X10Y111_SLICE_X13Y111_B3 = CLBLM_R_X11Y109_SLICE_X15Y109_CO6;
  assign CLBLM_L_X10Y111_SLICE_X13Y111_B4 = CLBLM_R_X11Y111_SLICE_X14Y111_AO6;
  assign CLBLM_L_X10Y111_SLICE_X13Y111_B5 = CLBLM_L_X10Y111_SLICE_X13Y111_AO6;
  assign CLBLM_L_X10Y111_SLICE_X13Y111_B6 = CLBLM_L_X12Y110_SLICE_X16Y110_DO6;
  assign CLBLM_L_X10Y111_SLICE_X13Y111_C1 = RIOB33_X105Y103_IOB_X1Y104_I;
  assign CLBLM_L_X10Y111_SLICE_X13Y111_C2 = RIOB33_X105Y103_IOB_X1Y103_I;
  assign CLBLM_L_X10Y111_SLICE_X13Y111_C3 = LIOB33_X0Y109_IOB_X0Y109_I;
  assign CLBLM_L_X10Y111_SLICE_X13Y111_C4 = CLBLM_L_X12Y110_SLICE_X16Y110_CO6;
  assign CLBLM_L_X10Y111_SLICE_X13Y111_C5 = CLBLM_L_X10Y111_SLICE_X13Y111_DO6;
  assign CLBLM_L_X10Y111_SLICE_X13Y111_C6 = CLBLM_R_X11Y111_SLICE_X14Y111_CO6;
  assign CLBLM_L_X10Y111_SLICE_X13Y111_D1 = LIOB33_X0Y107_IOB_X0Y108_I;
  assign CLBLM_L_X10Y111_SLICE_X13Y111_D2 = CLBLM_R_X11Y109_SLICE_X15Y109_CO6;
  assign CLBLM_L_X10Y111_SLICE_X13Y111_D3 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X10Y111_SLICE_X13Y111_D4 = CLBLM_R_X11Y111_SLICE_X15Y111_DO6;
  assign CLBLM_L_X10Y111_SLICE_X13Y111_D5 = CLBLM_L_X12Y110_SLICE_X16Y110_DO6;
  assign CLBLM_L_X10Y111_SLICE_X13Y111_D6 = RIOB33_X105Y103_IOB_X1Y104_I;
  assign CLBLM_L_X10Y111_SLICE_X12Y111_A1 = LIOB33_X0Y109_IOB_X0Y109_I;
  assign CLBLM_L_X10Y111_SLICE_X12Y111_A2 = CLBLM_L_X10Y111_SLICE_X13Y111_BO6;
  assign CLBLM_L_X10Y111_SLICE_X12Y111_A3 = LIOB33_X0Y109_IOB_X0Y110_I;
  assign CLBLM_L_X10Y111_SLICE_X12Y111_A4 = CLBLM_R_X11Y111_SLICE_X14Y111_CO6;
  assign CLBLM_L_X10Y111_SLICE_X12Y111_A5 = RIOB33_X105Y103_IOB_X1Y103_I;
  assign CLBLM_L_X10Y111_SLICE_X12Y111_A6 = CLBLM_L_X12Y110_SLICE_X16Y110_CO6;
  assign CLBLM_L_X10Y111_SLICE_X12Y111_B1 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X10Y111_SLICE_X12Y111_B2 = LIOB33_X0Y109_IOB_X0Y109_I;
  assign CLBLM_L_X10Y111_SLICE_X12Y111_B3 = CLBLM_R_X11Y111_SLICE_X14Y111_BO6;
  assign CLBLM_L_X10Y111_SLICE_X12Y111_B4 = LIOB33_X0Y107_IOB_X0Y108_I;
  assign CLBLM_L_X10Y111_SLICE_X12Y111_B5 = RIOB33_X105Y107_IOB_X1Y107_I;
  assign CLBLM_L_X10Y111_SLICE_X12Y111_B6 = CLBLM_L_X10Y112_SLICE_X13Y112_AO5;
  assign CLBLM_L_X10Y111_SLICE_X12Y111_C1 = LIOB33_X0Y109_IOB_X0Y110_I;
  assign CLBLM_L_X10Y111_SLICE_X12Y111_C2 = RIOB33_X105Y103_IOB_X1Y103_I;
  assign CLBLM_L_X10Y111_SLICE_X12Y111_C3 = CLBLM_L_X10Y111_SLICE_X13Y111_BO6;
  assign CLBLM_L_X10Y111_SLICE_X12Y111_C4 = CLBLM_L_X12Y110_SLICE_X16Y110_CO6;
  assign CLBLM_L_X10Y111_SLICE_X12Y111_C5 = LIOB33_X0Y109_IOB_X0Y109_I;
  assign CLBLM_L_X10Y111_SLICE_X12Y111_C6 = CLBLM_R_X11Y111_SLICE_X14Y111_CO6;
  assign CLBLL_L_X4Y107_SLICE_X4Y107_A1 = LIOB33_X0Y103_IOB_X0Y103_I;
  assign CLBLL_L_X4Y107_SLICE_X4Y107_A2 = CLBLL_L_X4Y106_SLICE_X4Y106_CO6;
  assign CLBLL_L_X4Y107_SLICE_X4Y107_A3 = LIOB33_X0Y107_IOB_X0Y107_I;
  assign CLBLL_L_X4Y107_SLICE_X4Y107_A4 = RIOB33_X105Y105_IOB_X1Y106_I;
  assign CLBLL_L_X4Y107_SLICE_X4Y107_A5 = CLBLL_L_X4Y106_SLICE_X4Y106_BO6;
  assign CLBLM_L_X10Y111_SLICE_X12Y111_D1 = CLBLM_R_X11Y111_SLICE_X14Y111_BO6;
  assign CLBLL_L_X4Y107_SLICE_X4Y107_A6 = LIOB33_X0Y107_IOB_X0Y108_I;
  assign CLBLM_L_X10Y111_SLICE_X12Y111_D4 = CLBLM_L_X10Y112_SLICE_X13Y112_AO5;
  assign CLBLL_L_X4Y107_SLICE_X4Y107_B1 = RIOB33_SING_X105Y100_IOB_X1Y100_I;
  assign CLBLL_L_X4Y107_SLICE_X4Y107_B2 = CLBLM_R_X3Y107_SLICE_X3Y107_CO6;
  assign CLBLL_L_X4Y107_SLICE_X4Y107_B3 = CLBLL_L_X4Y107_SLICE_X5Y107_CO6;
  assign CLBLL_L_X4Y107_SLICE_X4Y107_B4 = LIOB33_X0Y109_IOB_X0Y109_I;
  assign CLBLL_L_X4Y107_SLICE_X4Y107_B5 = CLBLL_L_X4Y107_SLICE_X4Y107_AO6;
  assign CLBLL_L_X4Y107_SLICE_X4Y107_B6 = LIOB33_X0Y109_IOB_X0Y110_I;
  assign CLBLM_L_X10Y111_SLICE_X12Y111_D3 = RIOB33_X105Y107_IOB_X1Y107_I;
  assign CLBLM_L_X10Y111_SLICE_X12Y111_D5 = LIOB33_X0Y107_IOB_X0Y108_I;
  assign CLBLM_L_X10Y111_SLICE_X12Y111_D6 = LIOB33_X0Y109_IOB_X0Y109_I;
  assign CLBLL_L_X4Y107_SLICE_X4Y107_C1 = LIOB33_X0Y107_IOB_X0Y107_I;
  assign CLBLL_L_X4Y107_SLICE_X4Y107_C2 = CLBLL_L_X4Y106_SLICE_X4Y106_CO6;
  assign CLBLL_L_X4Y107_SLICE_X4Y107_C3 = RIOB33_X105Y105_IOB_X1Y106_I;
  assign CLBLL_L_X4Y107_SLICE_X4Y107_C4 = LIOB33_X0Y107_IOB_X0Y108_I;
  assign CLBLL_L_X4Y107_SLICE_X4Y107_C5 = LIOB33_X0Y103_IOB_X0Y103_I;
  assign CLBLL_L_X4Y107_SLICE_X4Y107_C6 = CLBLL_L_X4Y106_SLICE_X4Y106_BO6;
  assign CLBLL_L_X4Y107_SLICE_X4Y107_D1 = 1'b1;
  assign CLBLL_L_X4Y107_SLICE_X4Y107_D2 = 1'b1;
  assign CLBLL_L_X4Y107_SLICE_X4Y107_D3 = 1'b1;
  assign CLBLL_L_X4Y107_SLICE_X4Y107_D4 = 1'b1;
  assign CLBLL_L_X4Y107_SLICE_X4Y107_D5 = 1'b1;
  assign CLBLL_L_X4Y107_SLICE_X4Y107_D6 = 1'b1;
  assign CLBLM_R_X11Y105_SLICE_X15Y105_A1 = 1'b1;
  assign CLBLM_R_X11Y105_SLICE_X15Y105_A2 = RIOB33_X105Y103_IOB_X1Y104_I;
  assign CLBLM_R_X11Y105_SLICE_X15Y105_A3 = LIOB33_X0Y103_IOB_X0Y104_I;
  assign CLBLM_R_X11Y105_SLICE_X15Y105_A4 = LIOB33_X0Y105_IOB_X0Y105_I;
  assign CLBLM_R_X11Y105_SLICE_X15Y105_A5 = 1'b1;
  assign CLBLL_L_X4Y107_SLICE_X5Y107_A1 = LIOB33_X0Y103_IOB_X0Y103_I;
  assign CLBLL_L_X4Y107_SLICE_X5Y107_A2 = RIOB33_X105Y105_IOB_X1Y106_I;
  assign CLBLL_L_X4Y107_SLICE_X5Y107_A3 = 1'b1;
  assign CLBLL_L_X4Y107_SLICE_X5Y107_A4 = LIOB33_X0Y107_IOB_X0Y108_I;
  assign CLBLL_L_X4Y107_SLICE_X5Y107_A5 = 1'b1;
  assign CLBLL_L_X4Y107_SLICE_X5Y107_A6 = 1'b1;
  assign CLBLM_R_X11Y105_SLICE_X15Y105_A6 = 1'b1;
  assign CLBLM_R_X11Y105_SLICE_X15Y105_B3 = LIOB33_X0Y103_IOB_X0Y104_I;
  assign CLBLM_R_X11Y105_SLICE_X15Y105_B4 = RIOB33_X105Y103_IOB_X1Y104_I;
  assign CLBLL_L_X4Y107_SLICE_X5Y107_B1 = LIOB33_X0Y103_IOB_X0Y103_I;
  assign CLBLL_L_X4Y107_SLICE_X5Y107_B2 = CLBLM_R_X5Y106_SLICE_X7Y106_CO6;
  assign CLBLL_L_X4Y107_SLICE_X5Y107_B3 = LIOB33_X0Y107_IOB_X0Y108_I;
  assign CLBLL_L_X4Y107_SLICE_X5Y107_B4 = CLBLL_L_X4Y106_SLICE_X4Y106_CO6;
  assign CLBLL_L_X4Y107_SLICE_X5Y107_B5 = CLBLL_L_X4Y106_SLICE_X5Y106_AO6;
  assign CLBLL_L_X4Y107_SLICE_X5Y107_B6 = RIOB33_X105Y105_IOB_X1Y106_I;
  assign CLBLM_R_X11Y105_SLICE_X15Y105_B6 = LIOB33_X0Y101_IOB_X0Y102_I;
  assign CLBLM_R_X11Y105_SLICE_X15Y105_C3 = RIOB33_X105Y103_IOB_X1Y104_I;
  assign CLBLM_R_X11Y105_SLICE_X15Y105_C4 = LIOB33_X0Y101_IOB_X0Y102_I;
  assign CLBLL_L_X4Y107_SLICE_X5Y107_C1 = CLBLL_L_X4Y107_SLICE_X5Y107_AO6;
  assign CLBLL_L_X4Y107_SLICE_X5Y107_C2 = CLBLM_R_X5Y106_SLICE_X7Y106_CO6;
  assign CLBLL_L_X4Y107_SLICE_X5Y107_C3 = CLBLM_R_X3Y107_SLICE_X3Y107_AO5;
  assign CLBLL_L_X4Y107_SLICE_X5Y107_C4 = CLBLL_L_X4Y107_SLICE_X5Y107_AO5;
  assign CLBLL_L_X4Y107_SLICE_X5Y107_C5 = CLBLL_L_X4Y106_SLICE_X5Y106_AO6;
  assign CLBLL_L_X4Y107_SLICE_X5Y107_C6 = CLBLL_L_X4Y106_SLICE_X4Y106_CO6;
  assign CLBLM_R_X11Y105_SLICE_X15Y105_C5 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X11Y105_SLICE_X15Y105_C6 = CLBLM_L_X12Y105_SLICE_X16Y105_CO6;
  assign CLBLM_R_X11Y105_SLICE_X15Y105_D1 = RIOB33_X105Y103_IOB_X1Y104_I;
  assign CLBLM_R_X11Y105_SLICE_X15Y105_D2 = CLBLM_R_X11Y104_SLICE_X15Y104_AO5;
  assign CLBLM_R_X11Y105_SLICE_X15Y105_D3 = LIOB33_X0Y101_IOB_X0Y102_I;
  assign CLBLM_R_X11Y105_SLICE_X15Y105_D4 = CLBLM_L_X12Y105_SLICE_X16Y105_AO5;
  assign CLBLL_L_X4Y107_SLICE_X5Y107_D1 = CLBLL_L_X4Y107_SLICE_X5Y107_AO6;
  assign CLBLL_L_X4Y107_SLICE_X5Y107_D2 = CLBLM_R_X5Y106_SLICE_X7Y106_CO6;
  assign CLBLL_L_X4Y107_SLICE_X5Y107_D3 = CLBLM_R_X3Y107_SLICE_X3Y107_AO5;
  assign CLBLL_L_X4Y107_SLICE_X5Y107_D4 = CLBLL_L_X4Y107_SLICE_X5Y107_AO5;
  assign CLBLL_L_X4Y107_SLICE_X5Y107_D5 = CLBLL_L_X4Y106_SLICE_X5Y106_AO6;
  assign CLBLL_L_X4Y107_SLICE_X5Y107_D6 = CLBLL_L_X4Y106_SLICE_X4Y106_CO6;
  assign CLBLM_R_X11Y105_SLICE_X15Y105_D5 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X11Y105_SLICE_X14Y105_A1 = 1'b1;
  assign CLBLL_L_X4Y110_SLICE_X4Y110_C1 = 1'b1;
  assign CLBLM_R_X11Y105_SLICE_X14Y105_A2 = RIOB33_X105Y103_IOB_X1Y103_I;
  assign CLBLM_R_X11Y105_SLICE_X14Y105_A3 = LIOB33_X0Y103_IOB_X0Y104_I;
  assign CLBLM_R_X11Y105_SLICE_X14Y105_A4 = LIOB33_X0Y105_IOB_X0Y105_I;
  assign CLBLM_R_X11Y105_SLICE_X14Y105_A5 = 1'b1;
  assign CLBLM_R_X11Y105_SLICE_X14Y105_A6 = 1'b1;
  assign CLBLM_R_X11Y105_SLICE_X14Y105_B1 = CLBLM_L_X12Y104_SLICE_X16Y104_BO6;
  assign CLBLM_R_X11Y105_SLICE_X14Y105_B2 = CLBLM_R_X11Y104_SLICE_X14Y104_CO6;
  assign CLBLM_R_X11Y105_SLICE_X14Y105_B3 = CLBLM_R_X11Y105_SLICE_X15Y105_AO6;
  assign CLBLM_R_X11Y105_SLICE_X14Y105_B4 = CLBLM_R_X11Y104_SLICE_X14Y104_BO6;
  assign CLBLM_R_X11Y105_SLICE_X14Y105_B5 = CLBLM_R_X11Y105_SLICE_X14Y105_AO6;
  assign CLBLM_R_X11Y105_SLICE_X14Y105_B6 = CLBLM_L_X10Y104_SLICE_X13Y104_DO6;
  assign CLBLM_R_X11Y105_SLICE_X14Y105_C1 = RIOB33_X105Y103_IOB_X1Y103_I;
  assign CLBLM_R_X11Y105_SLICE_X14Y105_C2 = LIOB33_X0Y101_IOB_X0Y102_I;
  assign CLBLM_R_X11Y105_SLICE_X14Y105_C3 = CLBLM_R_X11Y104_SLICE_X14Y104_DO6;
  assign CLBLM_R_X11Y105_SLICE_X14Y105_C4 = LIOB33_X0Y103_IOB_X0Y104_I;
  assign CLBLM_R_X11Y105_SLICE_X14Y105_C5 = RIOB33_X105Y103_IOB_X1Y104_I;
  assign CLBLM_R_X11Y105_SLICE_X14Y105_C6 = CLBLM_L_X10Y104_SLICE_X13Y104_DO6;
  assign CLBLM_R_X11Y105_SLICE_X14Y105_D1 = RIOB33_X105Y103_IOB_X1Y103_I;
  assign CLBLM_R_X11Y105_SLICE_X14Y105_D2 = LIOB33_X0Y101_IOB_X0Y102_I;
  assign CLBLM_R_X11Y105_SLICE_X14Y105_D3 = CLBLM_R_X11Y104_SLICE_X14Y104_DO6;
  assign CLBLM_R_X11Y105_SLICE_X14Y105_D4 = LIOB33_X0Y103_IOB_X0Y104_I;
  assign CLBLM_R_X11Y105_SLICE_X14Y105_D5 = RIOB33_X105Y103_IOB_X1Y104_I;
  assign CLBLM_R_X11Y105_SLICE_X14Y105_D6 = CLBLM_L_X10Y104_SLICE_X13Y104_DO6;
  assign CLBLM_L_X10Y112_SLICE_X13Y112_A1 = CLBLM_R_X11Y110_SLICE_X15Y110_CO6;
  assign CLBLM_L_X10Y112_SLICE_X13Y112_A2 = CLBLM_L_X10Y107_SLICE_X13Y107_AO6;
  assign CLBLM_L_X10Y112_SLICE_X13Y112_A3 = RIOB33_X105Y107_IOB_X1Y108_I;
  assign CLBLM_L_X10Y112_SLICE_X13Y112_A4 = CLBLM_L_X12Y108_SLICE_X16Y108_BO6;
  assign CLBLM_L_X10Y112_SLICE_X13Y112_A5 = LIOB33_X0Y107_IOB_X0Y107_I;
  assign CLBLM_L_X10Y112_SLICE_X13Y112_A6 = 1'b1;
  assign CLBLM_L_X10Y112_SLICE_X13Y112_B1 = CLBLM_L_X10Y112_SLICE_X13Y112_DO6;
  assign CLBLM_L_X10Y112_SLICE_X13Y112_B2 = RIOB33_X105Y107_IOB_X1Y107_I;
  assign CLBLM_L_X10Y112_SLICE_X13Y112_B3 = LIOB33_X0Y109_IOB_X0Y109_I;
  assign CLBLM_L_X10Y112_SLICE_X13Y112_B4 = LIOB33_X0Y107_IOB_X0Y108_I;
  assign CLBLM_L_X10Y112_SLICE_X13Y112_B5 = CLBLM_L_X10Y112_SLICE_X13Y112_AO6;
  assign CLBLM_L_X10Y112_SLICE_X13Y112_B6 = CLBLM_R_X11Y110_SLICE_X15Y110_CO6;
  assign CLBLM_L_X10Y112_SLICE_X13Y112_C1 = CLBLM_L_X10Y112_SLICE_X13Y112_AO6;
  assign CLBLM_L_X10Y112_SLICE_X13Y112_C2 = RIOB33_X105Y107_IOB_X1Y107_I;
  assign CLBLM_L_X10Y112_SLICE_X13Y112_C3 = CLBLM_R_X11Y110_SLICE_X15Y110_CO6;
  assign CLBLM_L_X10Y112_SLICE_X13Y112_C4 = LIOB33_X0Y107_IOB_X0Y108_I;
  assign CLBLM_L_X10Y112_SLICE_X13Y112_C5 = CLBLM_L_X10Y112_SLICE_X13Y112_DO6;
  assign CLBLM_L_X10Y112_SLICE_X13Y112_C6 = LIOB33_X0Y109_IOB_X0Y109_I;
  assign CLBLM_L_X10Y112_SLICE_X13Y112_D1 = CLBLM_L_X12Y108_SLICE_X16Y108_BO6;
  assign CLBLM_L_X10Y112_SLICE_X13Y112_D2 = CLBLM_L_X10Y107_SLICE_X13Y107_AO6;
  assign CLBLM_L_X10Y112_SLICE_X13Y112_D3 = LIOB33_X0Y107_IOB_X0Y108_I;
  assign CLBLM_L_X10Y112_SLICE_X13Y112_D4 = LIOB33_X0Y107_IOB_X0Y107_I;
  assign CLBLM_L_X10Y112_SLICE_X13Y112_D5 = RIOB33_X105Y107_IOB_X1Y108_I;
  assign CLBLM_L_X10Y112_SLICE_X13Y112_D6 = CLBLM_L_X10Y107_SLICE_X13Y107_BO6;
  assign CLBLM_L_X10Y112_SLICE_X12Y112_A1 = CLBLM_R_X11Y110_SLICE_X14Y110_BO6;
  assign CLBLM_L_X10Y112_SLICE_X12Y112_A2 = LIOB33_X0Y109_IOB_X0Y109_I;
  assign CLBLM_L_X10Y112_SLICE_X12Y112_A3 = RIOB33_X105Y101_IOB_X1Y102_I;
  assign CLBLM_L_X10Y112_SLICE_X12Y112_A4 = CLBLM_L_X12Y110_SLICE_X16Y110_BO6;
  assign CLBLM_L_X10Y112_SLICE_X12Y112_A5 = LIOB33_X0Y109_IOB_X0Y110_I;
  assign CLBLM_L_X10Y112_SLICE_X12Y112_A6 = CLBLM_L_X10Y110_SLICE_X12Y110_CO6;
  assign CLBLM_L_X10Y112_SLICE_X12Y112_B1 = CLBLM_R_X11Y110_SLICE_X14Y110_BO6;
  assign CLBLM_L_X10Y112_SLICE_X12Y112_B2 = CLBLM_L_X12Y110_SLICE_X16Y110_BO6;
  assign CLBLM_L_X10Y112_SLICE_X12Y112_B3 = RIOB33_X105Y101_IOB_X1Y102_I;
  assign CLBLM_L_X10Y112_SLICE_X12Y112_B4 = CLBLM_L_X10Y110_SLICE_X12Y110_CO6;
  assign CLBLM_L_X10Y112_SLICE_X12Y112_B5 = LIOB33_X0Y109_IOB_X0Y110_I;
  assign CLBLM_L_X10Y112_SLICE_X12Y112_B6 = LIOB33_X0Y109_IOB_X0Y109_I;
  assign CLBLM_L_X10Y112_SLICE_X12Y112_C1 = 1'b1;
  assign CLBLM_L_X10Y112_SLICE_X12Y112_C2 = 1'b1;
  assign CLBLM_L_X10Y112_SLICE_X12Y112_C3 = 1'b1;
  assign CLBLM_L_X10Y112_SLICE_X12Y112_C4 = 1'b1;
  assign CLBLM_L_X10Y112_SLICE_X12Y112_C5 = 1'b1;
  assign CLBLM_L_X10Y112_SLICE_X12Y112_C6 = 1'b1;
  assign CLBLL_L_X4Y108_SLICE_X4Y108_A1 = CLBLM_R_X5Y108_SLICE_X6Y108_AO6;
  assign CLBLL_L_X4Y108_SLICE_X4Y108_A2 = RIOB33_X105Y105_IOB_X1Y106_I;
  assign CLBLL_L_X4Y108_SLICE_X4Y108_A3 = LIOB33_X0Y111_IOB_X0Y112_I;
  assign CLBLL_L_X4Y108_SLICE_X4Y108_A4 = CLBLL_L_X4Y108_SLICE_X4Y108_BO6;
  assign CLBLL_L_X4Y108_SLICE_X4Y108_A5 = RIOB33_SING_X105Y100_IOB_X1Y100_I;
  assign CLBLL_L_X4Y108_SLICE_X4Y108_A6 = 1'b1;
  assign CLBLM_L_X10Y112_SLICE_X12Y112_D1 = 1'b1;
  assign CLBLM_L_X10Y112_SLICE_X12Y112_D2 = 1'b1;
  assign CLBLM_L_X10Y112_SLICE_X12Y112_D3 = 1'b1;
  assign CLBLM_L_X10Y112_SLICE_X12Y112_D4 = 1'b1;
  assign CLBLM_L_X10Y112_SLICE_X12Y112_D5 = 1'b1;
  assign CLBLM_L_X10Y112_SLICE_X12Y112_D6 = 1'b1;
  assign CLBLL_L_X4Y108_SLICE_X4Y108_B1 = LIOB33_X0Y111_IOB_X0Y111_I;
  assign CLBLL_L_X4Y108_SLICE_X4Y108_B2 = LIOB33_X0Y109_IOB_X0Y110_I;
  assign CLBLL_L_X4Y108_SLICE_X4Y108_B3 = RIOB33_X105Y105_IOB_X1Y106_I;
  assign CLBLL_L_X4Y108_SLICE_X4Y108_B4 = CLBLL_L_X4Y107_SLICE_X4Y107_BO6;
  assign CLBLL_L_X4Y108_SLICE_X4Y108_B5 = CLBLM_R_X5Y107_SLICE_X6Y107_AO6;
  assign CLBLL_L_X4Y108_SLICE_X4Y108_B6 = RIOB33_SING_X105Y100_IOB_X1Y100_I;
  assign CLBLL_L_X4Y108_SLICE_X4Y108_C1 = CLBLM_R_X5Y108_SLICE_X6Y108_BO6;
  assign CLBLL_L_X4Y108_SLICE_X4Y108_C2 = CLBLM_R_X5Y110_SLICE_X7Y110_AO6;
  assign CLBLL_L_X4Y108_SLICE_X4Y108_C3 = CLBLM_R_X7Y107_SLICE_X8Y107_AO6;
  assign CLBLL_L_X4Y108_SLICE_X4Y108_C4 = CLBLL_L_X4Y108_SLICE_X4Y108_AO5;
  assign CLBLL_L_X4Y108_SLICE_X4Y108_C5 = CLBLM_R_X5Y108_SLICE_X6Y108_AO6;
  assign CLBLL_L_X4Y108_SLICE_X4Y108_C6 = CLBLL_L_X4Y108_SLICE_X4Y108_BO6;
  assign CLBLL_L_X4Y108_SLICE_X4Y108_D1 = RIOB33_SING_X105Y100_IOB_X1Y100_I;
  assign CLBLL_L_X4Y108_SLICE_X4Y108_D2 = CLBLM_R_X5Y108_SLICE_X6Y108_CO6;
  assign CLBLL_L_X4Y108_SLICE_X4Y108_D3 = CLBLM_R_X7Y107_SLICE_X8Y107_AO6;
  assign CLBLL_L_X4Y108_SLICE_X4Y108_D4 = CLBLL_L_X4Y108_SLICE_X4Y108_AO5;
  assign CLBLL_L_X4Y108_SLICE_X4Y108_D5 = LIOB33_X0Y113_IOB_X0Y113_I;
  assign CLBLL_L_X4Y108_SLICE_X4Y108_D6 = CLBLM_R_X5Y108_SLICE_X6Y108_BO6;
  assign CLBLL_L_X4Y108_SLICE_X5Y108_A1 = CLBLM_R_X7Y107_SLICE_X8Y107_AO6;
  assign CLBLL_L_X4Y108_SLICE_X5Y108_A2 = LIOB33_X0Y111_IOB_X0Y112_I;
  assign CLBLL_L_X4Y108_SLICE_X5Y108_A3 = LIOB33_X0Y103_IOB_X0Y103_I;
  assign CLBLL_L_X4Y108_SLICE_X5Y108_A4 = CLBLM_R_X7Y107_SLICE_X8Y107_BO6;
  assign CLBLL_L_X4Y108_SLICE_X5Y108_A5 = RIOB33_X105Y105_IOB_X1Y106_I;
  assign CLBLL_L_X4Y108_SLICE_X5Y108_A6 = CLBLM_R_X5Y108_SLICE_X6Y108_BO6;
  assign CLBLM_R_X11Y106_SLICE_X15Y106_A1 = CLBLM_R_X11Y106_SLICE_X15Y106_DO6;
  assign CLBLM_R_X11Y106_SLICE_X15Y106_A2 = RIOB33_X105Y109_IOB_X1Y109_I;
  assign CLBLM_R_X11Y106_SLICE_X15Y106_A3 = LIOB33_X0Y107_IOB_X0Y107_I;
  assign CLBLL_L_X4Y108_SLICE_X5Y108_B1 = LIOB33_X0Y113_IOB_X0Y113_I;
  assign CLBLL_L_X4Y108_SLICE_X5Y108_B2 = CLBLM_R_X7Y107_SLICE_X8Y107_CO6;
  assign CLBLL_L_X4Y108_SLICE_X5Y108_B3 = LIOB33_X0Y103_IOB_X0Y103_I;
  assign CLBLL_L_X4Y108_SLICE_X5Y108_B4 = CLBLM_R_X5Y108_SLICE_X7Y108_CO6;
  assign CLBLL_L_X4Y108_SLICE_X5Y108_B5 = CLBLM_R_X7Y108_SLICE_X8Y108_BO6;
  assign CLBLL_L_X4Y108_SLICE_X5Y108_B6 = LIOB33_X0Y111_IOB_X0Y112_I;
  assign CLBLM_R_X11Y106_SLICE_X15Y106_B1 = RIOB33_X105Y109_IOB_X1Y110_I;
  assign CLBLM_R_X11Y106_SLICE_X15Y106_B2 = LIOB33_X0Y103_IOB_X0Y104_I;
  assign CLBLL_L_X4Y108_SLICE_X5Y108_C1 = CLBLM_R_X7Y108_SLICE_X8Y108_BO6;
  assign CLBLL_L_X4Y108_SLICE_X5Y108_C2 = CLBLM_R_X7Y107_SLICE_X8Y107_CO6;
  assign CLBLL_L_X4Y108_SLICE_X5Y108_C3 = LIOB33_X0Y113_IOB_X0Y113_I;
  assign CLBLL_L_X4Y108_SLICE_X5Y108_C4 = LIOB33_X0Y111_IOB_X0Y112_I;
  assign CLBLL_L_X4Y108_SLICE_X5Y108_C5 = LIOB33_X0Y103_IOB_X0Y103_I;
  assign CLBLL_L_X4Y108_SLICE_X5Y108_C6 = CLBLM_R_X5Y108_SLICE_X7Y108_CO6;
  assign CLBLM_R_X11Y106_SLICE_X15Y106_C1 = RIOB33_X105Y109_IOB_X1Y109_I;
  assign CLBLM_R_X11Y106_SLICE_X15Y106_C2 = CLBLM_L_X12Y105_SLICE_X17Y105_AO6;
  assign CLBLM_R_X11Y106_SLICE_X15Y106_C3 = LIOB33_X0Y101_IOB_X0Y102_I;
  assign CLBLM_R_X11Y106_SLICE_X15Y106_C4 = CLBLM_L_X10Y107_SLICE_X13Y107_DO6;
  assign CLBLM_R_X11Y106_SLICE_X15Y106_C5 = RIOB33_X105Y109_IOB_X1Y110_I;
  assign CLBLM_R_X11Y106_SLICE_X15Y106_C6 = LIOB33_X0Y103_IOB_X0Y104_I;
  assign CLBLL_L_X4Y108_SLICE_X5Y108_D1 = LIOB33_X0Y113_IOB_X0Y114_I;
  assign CLBLL_L_X4Y108_SLICE_X5Y108_D2 = CLBLM_R_X7Y107_SLICE_X8Y107_CO6;
  assign CLBLL_L_X4Y108_SLICE_X5Y108_D3 = LIOB33_X0Y111_IOB_X0Y112_I;
  assign CLBLL_L_X4Y108_SLICE_X5Y108_D4 = CLBLM_R_X7Y108_SLICE_X8Y108_CO6;
  assign CLBLL_L_X4Y108_SLICE_X5Y108_D5 = LIOB33_X0Y103_IOB_X0Y103_I;
  assign CLBLL_L_X4Y108_SLICE_X5Y108_D6 = CLBLM_R_X5Y108_SLICE_X7Y108_CO6;
  assign CLBLM_R_X11Y106_SLICE_X15Y106_D1 = RIOB33_X105Y109_IOB_X1Y109_I;
  assign CLBLM_R_X11Y106_SLICE_X15Y106_D2 = LIOB33_X0Y105_IOB_X0Y105_I;
  assign CLBLM_R_X11Y106_SLICE_X15Y106_D3 = CLBLM_R_X11Y107_SLICE_X15Y107_AO5;
  assign CLBLM_R_X11Y106_SLICE_X15Y106_D4 = RIOB33_X105Y109_IOB_X1Y110_I;
  assign CLBLM_R_X11Y106_SLICE_X15Y106_D5 = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLM_R_X11Y106_SLICE_X15Y106_D6 = CLBLM_L_X10Y107_SLICE_X13Y107_CO6;
  assign CLBLM_R_X11Y106_SLICE_X14Y106_A1 = CLBLM_R_X11Y106_SLICE_X14Y106_BO6;
  assign CLBLM_R_X11Y106_SLICE_X14Y106_A2 = CLBLM_R_X11Y105_SLICE_X15Y105_AO5;
  assign CLBLM_R_X11Y106_SLICE_X14Y106_A3 = CLBLM_R_X11Y109_SLICE_X14Y109_AO6;
  assign CLBLM_R_X11Y106_SLICE_X14Y106_A4 = CLBLM_R_X11Y105_SLICE_X14Y105_DO6;
  assign CLBLM_R_X11Y106_SLICE_X14Y106_A5 = CLBLM_R_X11Y105_SLICE_X15Y105_BO6;
  assign CLBLM_R_X11Y106_SLICE_X14Y106_A6 = CLBLM_R_X11Y105_SLICE_X14Y105_AO5;
  assign CLBLM_R_X11Y106_SLICE_X14Y106_B1 = CLBLM_R_X11Y105_SLICE_X15Y105_AO6;
  assign CLBLM_R_X11Y106_SLICE_X14Y106_B2 = CLBLM_L_X12Y106_SLICE_X17Y106_BO6;
  assign CLBLM_R_X11Y106_SLICE_X14Y106_B3 = CLBLM_L_X12Y104_SLICE_X16Y104_BO6;
  assign CLBLM_R_X11Y106_SLICE_X14Y106_B4 = CLBLM_R_X11Y107_SLICE_X14Y107_AO6;
  assign CLBLM_R_X11Y106_SLICE_X14Y106_B5 = CLBLM_R_X11Y104_SLICE_X14Y104_CO6;
  assign CLBLM_R_X11Y106_SLICE_X14Y106_B6 = CLBLM_L_X12Y104_SLICE_X16Y104_DO6;
  assign CLBLM_R_X11Y106_SLICE_X14Y106_C1 = CLBLM_R_X11Y109_SLICE_X14Y109_AO6;
  assign CLBLM_R_X11Y106_SLICE_X14Y106_C2 = CLBLM_R_X11Y105_SLICE_X14Y105_AO5;
  assign CLBLM_R_X11Y106_SLICE_X14Y106_C3 = CLBLM_R_X11Y105_SLICE_X15Y105_AO5;
  assign CLBLM_R_X11Y106_SLICE_X14Y106_C4 = CLBLM_R_X11Y105_SLICE_X14Y105_DO6;
  assign CLBLM_R_X11Y106_SLICE_X14Y106_C5 = CLBLM_R_X11Y105_SLICE_X15Y105_BO6;
  assign CLBLM_R_X11Y106_SLICE_X14Y106_C6 = CLBLM_R_X11Y106_SLICE_X14Y106_BO6;
  assign CLBLM_R_X11Y106_SLICE_X14Y106_D1 = CLBLM_R_X11Y105_SLICE_X15Y105_BO6;
  assign CLBLM_R_X11Y106_SLICE_X14Y106_D2 = RIOB33_X105Y103_IOB_X1Y103_I;
  assign CLBLM_R_X11Y106_SLICE_X14Y106_D3 = RIOB33_X105Y103_IOB_X1Y104_I;
  assign CLBLM_R_X11Y106_SLICE_X14Y106_D4 = CLBLM_R_X11Y105_SLICE_X14Y105_DO6;
  assign CLBLM_R_X11Y106_SLICE_X14Y106_D5 = LIOB33_X0Y105_IOB_X0Y105_I;
  assign CLBLM_R_X11Y106_SLICE_X14Y106_D6 = CLBLM_R_X11Y106_SLICE_X14Y106_BO6;
  assign CLBLL_L_X4Y110_SLICE_X5Y110_C3 = CLBLL_L_X4Y109_SLICE_X4Y109_BO6;
  assign CLBLL_L_X4Y110_SLICE_X5Y110_C6 = CLBLL_L_X4Y110_SLICE_X5Y110_BO6;
  assign CLBLM_L_X8Y103_SLICE_X11Y103_A1 = RIOB33_X105Y101_IOB_X1Y101_I;
  assign CLBLM_L_X8Y103_SLICE_X11Y103_A2 = LIOB33_X0Y103_IOB_X0Y104_I;
  assign CLBLM_L_X8Y103_SLICE_X11Y103_A3 = CLBLM_L_X8Y104_SLICE_X10Y104_CO6;
  assign CLBLM_L_X8Y103_SLICE_X11Y103_A4 = LIOB33_X0Y101_IOB_X0Y102_I;
  assign CLBLM_L_X8Y103_SLICE_X11Y103_A5 = RIOB33_X105Y101_IOB_X1Y102_I;
  assign CLBLM_L_X8Y103_SLICE_X11Y103_A6 = CLBLM_L_X10Y103_SLICE_X12Y103_CO6;
  assign CLBLM_L_X8Y103_SLICE_X11Y103_B1 = RIOB33_X105Y101_IOB_X1Y101_I;
  assign CLBLM_L_X8Y103_SLICE_X11Y103_B2 = LIOB33_X0Y101_IOB_X0Y102_I;
  assign CLBLM_L_X8Y103_SLICE_X11Y103_B3 = CLBLM_L_X8Y103_SLICE_X10Y103_AO5;
  assign CLBLM_L_X8Y103_SLICE_X11Y103_B4 = RIOB33_X105Y101_IOB_X1Y102_I;
  assign CLBLM_L_X8Y103_SLICE_X11Y103_B5 = CLBLM_L_X10Y103_SLICE_X12Y103_AO6;
  assign CLBLM_L_X8Y103_SLICE_X11Y103_B6 = CLBLM_L_X10Y103_SLICE_X12Y103_CO6;
  assign CLBLM_L_X8Y103_SLICE_X11Y103_C1 = 1'b1;
  assign CLBLM_L_X8Y103_SLICE_X11Y103_C2 = 1'b1;
  assign CLBLM_L_X8Y103_SLICE_X11Y103_C3 = 1'b1;
  assign CLBLM_L_X8Y103_SLICE_X11Y103_C4 = 1'b1;
  assign CLBLM_L_X8Y103_SLICE_X11Y103_C5 = 1'b1;
  assign CLBLM_L_X8Y103_SLICE_X11Y103_C6 = 1'b1;
  assign CLBLM_L_X8Y103_SLICE_X11Y103_D1 = 1'b1;
  assign CLBLM_L_X8Y103_SLICE_X11Y103_D2 = 1'b1;
  assign CLBLM_L_X8Y103_SLICE_X11Y103_D3 = 1'b1;
  assign CLBLM_L_X8Y103_SLICE_X11Y103_D4 = 1'b1;
  assign CLBLM_L_X8Y103_SLICE_X11Y103_D5 = 1'b1;
  assign CLBLM_L_X8Y103_SLICE_X11Y103_D6 = 1'b1;
  assign CLBLM_L_X8Y103_SLICE_X10Y103_A1 = LIOB33_X0Y101_IOB_X0Y101_I;
  assign CLBLM_L_X8Y103_SLICE_X10Y103_A2 = 1'b1;
  assign CLBLM_L_X8Y103_SLICE_X10Y103_A3 = RIOB33_X105Y101_IOB_X1Y101_I;
  assign CLBLL_L_X4Y109_SLICE_X4Y109_A1 = 1'b1;
  assign CLBLM_L_X8Y103_SLICE_X10Y103_A5 = CLBLM_R_X7Y103_SLICE_X8Y103_BO6;
  assign CLBLM_L_X8Y103_SLICE_X10Y103_A6 = 1'b1;
  assign CLBLL_L_X4Y109_SLICE_X4Y109_A2 = LIOB33_X0Y115_IOB_X0Y115_I;
  assign CLBLL_L_X4Y109_SLICE_X4Y109_A3 = RIOB33_X105Y105_IOB_X1Y106_I;
  assign CLBLL_L_X4Y109_SLICE_X4Y109_A4 = RIOB33_SING_X105Y100_IOB_X1Y100_I;
  assign CLBLL_L_X4Y109_SLICE_X4Y109_A5 = 1'b1;
  assign CLBLL_L_X4Y109_SLICE_X4Y109_A6 = 1'b1;
  assign CLBLM_L_X8Y103_SLICE_X10Y103_A4 = CLBLM_L_X8Y103_SLICE_X10Y103_BO6;
  assign CLBLM_L_X8Y103_SLICE_X10Y103_B1 = LIOB33_SING_X0Y100_IOB_X0Y100_I;
  assign CLBLM_L_X8Y103_SLICE_X10Y103_B2 = RIOB33_X105Y101_IOB_X1Y102_I;
  assign CLBLM_L_X8Y103_SLICE_X10Y103_B3 = RIOB33_X105Y101_IOB_X1Y101_I;
  assign CLBLM_L_X8Y103_SLICE_X10Y103_B4 = RIOB33_X105Y113_IOB_X1Y113_I;
  assign CLBLM_L_X8Y103_SLICE_X10Y103_B5 = RIOB33_X105Y111_IOB_X1Y112_I;
  assign CLBLM_L_X8Y103_SLICE_X10Y103_B6 = RIOB33_X105Y103_IOB_X1Y103_I;
  assign CLBLL_L_X4Y109_SLICE_X4Y109_B1 = CLBLL_L_X4Y109_SLICE_X4Y109_DO6;
  assign CLBLL_L_X4Y109_SLICE_X4Y109_B2 = CLBLL_L_X4Y109_SLICE_X4Y109_AO5;
  assign CLBLM_L_X8Y103_SLICE_X10Y103_C1 = 1'b1;
  assign CLBLL_L_X4Y109_SLICE_X4Y109_B3 = CLBLL_L_X4Y108_SLICE_X5Y108_BO6;
  assign CLBLL_L_X4Y109_SLICE_X4Y109_B4 = CLBLL_L_X4Y108_SLICE_X4Y108_DO6;
  assign CLBLL_L_X4Y109_SLICE_X4Y109_B5 = CLBLL_L_X4Y109_SLICE_X4Y109_AO6;
  assign CLBLL_L_X4Y109_SLICE_X4Y109_B6 = CLBLL_L_X4Y109_SLICE_X4Y109_CO6;
  assign CLBLL_L_X4Y109_SLICE_X4Y109_C1 = RIOB33_X105Y105_IOB_X1Y106_I;
  assign CLBLL_L_X4Y109_SLICE_X4Y109_C2 = CLBLM_R_X5Y108_SLICE_X6Y108_BO6;
  assign CLBLL_L_X4Y109_SLICE_X4Y109_C3 = LIOB33_X0Y113_IOB_X0Y113_I;
  assign CLBLL_L_X4Y109_SLICE_X4Y109_C4 = CLBLM_R_X7Y107_SLICE_X8Y107_DO6;
  assign CLBLL_L_X4Y109_SLICE_X4Y109_C5 = LIOB33_X0Y111_IOB_X0Y112_I;
  assign CLBLL_L_X4Y109_SLICE_X4Y109_C6 = CLBLM_R_X7Y107_SLICE_X8Y107_AO6;
  assign CLBLM_L_X8Y103_SLICE_X10Y103_C5 = 1'b1;
  assign CLBLM_L_X8Y103_SLICE_X10Y103_C6 = 1'b1;
  assign CLBLL_L_X4Y109_SLICE_X4Y109_D1 = RIOB33_X105Y105_IOB_X1Y106_I;
  assign CLBLL_L_X4Y109_SLICE_X4Y109_D2 = CLBLM_R_X5Y108_SLICE_X6Y108_BO6;
  assign CLBLL_L_X4Y109_SLICE_X4Y109_D3 = LIOB33_X0Y113_IOB_X0Y113_I;
  assign CLBLL_L_X4Y109_SLICE_X4Y109_D4 = CLBLM_R_X7Y107_SLICE_X8Y107_DO6;
  assign CLBLL_L_X4Y109_SLICE_X4Y109_D5 = LIOB33_X0Y111_IOB_X0Y112_I;
  assign CLBLL_L_X4Y109_SLICE_X4Y109_D6 = CLBLM_R_X7Y107_SLICE_X8Y107_AO6;
  assign CLBLM_L_X8Y103_SLICE_X10Y103_D1 = 1'b1;
  assign CLBLM_L_X8Y103_SLICE_X10Y103_D2 = 1'b1;
  assign CLBLM_L_X8Y103_SLICE_X10Y103_D3 = 1'b1;
  assign CLBLM_L_X8Y103_SLICE_X10Y103_D4 = 1'b1;
  assign CLBLM_L_X8Y103_SLICE_X10Y103_D5 = 1'b1;
  assign CLBLM_L_X8Y103_SLICE_X10Y103_D6 = 1'b1;
  assign CLBLL_L_X4Y109_SLICE_X5Y109_A1 = LIOB33_X0Y113_IOB_X0Y113_I;
  assign CLBLL_L_X4Y109_SLICE_X5Y109_A2 = CLBLM_R_X5Y109_SLICE_X7Y109_AO6;
  assign CLBLL_L_X4Y109_SLICE_X5Y109_A3 = LIOB33_X0Y113_IOB_X0Y114_I;
  assign CLBLL_L_X4Y109_SLICE_X5Y109_A4 = CLBLM_R_X5Y110_SLICE_X7Y110_CO6;
  assign CLBLL_L_X4Y109_SLICE_X5Y109_A5 = RIOB33_X105Y101_IOB_X1Y102_I;
  assign CLBLL_L_X4Y109_SLICE_X5Y109_A6 = 1'b1;
  assign CLBLM_R_X11Y107_SLICE_X15Y107_A1 = RIOB33_X105Y109_IOB_X1Y109_I;
  assign CLBLM_R_X11Y107_SLICE_X15Y107_A3 = LIOB33_X0Y105_IOB_X0Y105_I;
  assign CLBLM_R_X11Y107_SLICE_X15Y107_A4 = LIOB33_X0Y103_IOB_X0Y104_I;
  assign CLBLL_L_X4Y109_SLICE_X5Y109_B1 = LIOB33_X0Y113_IOB_X0Y113_I;
  assign CLBLL_L_X4Y109_SLICE_X5Y109_B2 = CLBLM_R_X5Y109_SLICE_X7Y109_AO6;
  assign CLBLL_L_X4Y109_SLICE_X5Y109_B3 = LIOB33_X0Y113_IOB_X0Y114_I;
  assign CLBLL_L_X4Y109_SLICE_X5Y109_B4 = LIOB33_X0Y103_IOB_X0Y103_I;
  assign CLBLL_L_X4Y109_SLICE_X5Y109_B5 = LIOB33_X0Y115_IOB_X0Y115_I;
  assign CLBLL_L_X4Y109_SLICE_X5Y109_B6 = CLBLL_L_X4Y108_SLICE_X5Y108_CO6;
  assign CLBLM_R_X11Y107_SLICE_X15Y107_A6 = 1'b1;
  assign CLBLM_R_X11Y107_SLICE_X15Y107_A5 = CLBLM_R_X11Y106_SLICE_X15Y106_CO6;
  assign CLBLL_L_X4Y109_SLICE_X5Y109_C1 = LIOB33_X0Y115_IOB_X0Y115_I;
  assign CLBLL_L_X4Y109_SLICE_X5Y109_C2 = CLBLL_L_X4Y109_SLICE_X4Y109_CO6;
  assign CLBLL_L_X4Y109_SLICE_X5Y109_C3 = LIOB33_X0Y113_IOB_X0Y113_I;
  assign CLBLL_L_X4Y109_SLICE_X5Y109_C4 = RIOB33_X105Y105_IOB_X1Y106_I;
  assign CLBLL_L_X4Y109_SLICE_X5Y109_C5 = CLBLL_L_X4Y108_SLICE_X5Y108_DO6;
  assign CLBLL_L_X4Y109_SLICE_X5Y109_C6 = LIOB33_X0Y103_IOB_X0Y103_I;
  assign CLBLM_R_X11Y107_SLICE_X15Y107_B6 = CLBLM_R_X13Y107_SLICE_X18Y107_AO6;
  assign CLBLM_R_X11Y107_SLICE_X15Y107_C1 = CLBLM_L_X12Y107_SLICE_X16Y107_BO6;
  assign CLBLM_R_X11Y107_SLICE_X15Y107_C2 = CLBLM_R_X11Y107_SLICE_X14Y107_AO5;
  assign CLBLM_R_X11Y107_SLICE_X15Y107_C3 = CLBLM_L_X12Y108_SLICE_X16Y108_AO6;
  assign CLBLM_R_X11Y107_SLICE_X15Y107_C5 = CLBLM_L_X12Y107_SLICE_X16Y107_AO6;
  assign CLBLM_R_X11Y107_SLICE_X15Y107_C4 = CLBLM_R_X13Y107_SLICE_X18Y107_AO6;
  assign CLBLM_R_X11Y107_SLICE_X15Y107_C6 = CLBLM_R_X11Y111_SLICE_X15Y111_BO6;
  assign CLBLL_L_X4Y109_SLICE_X5Y109_D1 = LIOB33_X0Y115_IOB_X0Y115_I;
  assign CLBLL_L_X4Y109_SLICE_X5Y109_D2 = CLBLL_L_X4Y108_SLICE_X5Y108_CO6;
  assign CLBLL_L_X4Y109_SLICE_X5Y109_D3 = LIOB33_X0Y113_IOB_X0Y113_I;
  assign CLBLL_L_X4Y109_SLICE_X5Y109_D4 = LIOB33_X0Y113_IOB_X0Y114_I;
  assign CLBLL_L_X4Y109_SLICE_X5Y109_D5 = LIOB33_X0Y103_IOB_X0Y103_I;
  assign CLBLL_L_X4Y109_SLICE_X5Y109_D6 = CLBLM_R_X5Y109_SLICE_X7Y109_AO6;
  assign CLBLM_R_X11Y107_SLICE_X15Y107_D3 = CLBLM_R_X11Y107_SLICE_X14Y107_DO6;
  assign CLBLM_R_X11Y107_SLICE_X15Y107_D1 = LIOB33_X0Y103_IOB_X0Y104_I;
  assign CLBLM_R_X11Y107_SLICE_X15Y107_D5 = RIOB33_X105Y109_IOB_X1Y109_I;
  assign CLBLM_R_X11Y107_SLICE_X15Y107_D6 = CLBLM_L_X12Y105_SLICE_X17Y105_AO6;
  assign CLBLM_R_X11Y107_SLICE_X15Y107_D2 = LIOB33_X0Y105_IOB_X0Y105_I;
  assign CLBLM_R_X11Y107_SLICE_X15Y107_D4 = CLBLM_R_X11Y107_SLICE_X14Y107_BO5;
  assign CLBLM_R_X11Y107_SLICE_X14Y107_A1 = LIOB33_X0Y105_IOB_X0Y105_I;
  assign CLBLM_R_X11Y107_SLICE_X14Y107_A2 = LIOB33_X0Y103_IOB_X0Y104_I;
  assign CLBLM_R_X11Y107_SLICE_X14Y107_A3 = 1'b1;
  assign CLBLM_R_X11Y107_SLICE_X14Y107_A4 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X11Y107_SLICE_X14Y107_A5 = 1'b1;
  assign CLBLM_R_X11Y107_SLICE_X14Y107_A6 = 1'b1;
  assign LIOI3_X0Y105_ILOGIC_X0Y106_D = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLM_R_X11Y107_SLICE_X14Y107_B1 = LIOB33_X0Y105_IOB_X0Y105_I;
  assign CLBLM_R_X11Y107_SLICE_X14Y107_B2 = CLBLM_L_X10Y107_SLICE_X13Y107_CO6;
  assign CLBLM_R_X11Y107_SLICE_X14Y107_B3 = RIOB33_X105Y109_IOB_X1Y110_I;
  assign CLBLM_R_X11Y107_SLICE_X14Y107_B4 = CLBLM_L_X10Y107_SLICE_X13Y107_DO6;
  assign CLBLM_R_X11Y107_SLICE_X14Y107_B5 = LIOB33_X0Y101_IOB_X0Y102_I;
  assign CLBLM_R_X11Y107_SLICE_X14Y107_B6 = 1'b1;
  assign LIOI3_X0Y105_ILOGIC_X0Y105_D = LIOB33_X0Y105_IOB_X0Y105_I;
  assign CLBLM_R_X11Y107_SLICE_X14Y107_C1 = LIOB33_X0Y101_IOB_X0Y102_I;
  assign CLBLM_R_X11Y107_SLICE_X14Y107_C2 = CLBLM_L_X12Y104_SLICE_X16Y104_DO6;
  assign CLBLM_R_X11Y107_SLICE_X14Y107_C3 = CLBLM_L_X12Y106_SLICE_X16Y106_DO6;
  assign CLBLM_R_X11Y107_SLICE_X14Y107_C4 = RIOB33_X105Y107_IOB_X1Y107_I;
  assign CLBLM_R_X11Y107_SLICE_X14Y107_C5 = LIOB33_X0Y103_IOB_X0Y104_I;
  assign CLBLM_R_X11Y107_SLICE_X14Y107_C6 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X7Y111_SLICE_X9Y111_C6 = LIOB33_X0Y107_IOB_X0Y107_I;
  assign CLBLM_R_X11Y107_SLICE_X14Y107_D1 = LIOB33_X0Y101_IOB_X0Y101_I;
  assign CLBLM_R_X11Y107_SLICE_X14Y107_D2 = LIOB33_X0Y103_IOB_X0Y104_I;
  assign CLBLM_R_X11Y107_SLICE_X14Y107_D3 = CLBLM_L_X10Y107_SLICE_X12Y107_CO6;
  assign CLBLM_R_X11Y107_SLICE_X14Y107_D4 = LIOB33_X0Y101_IOB_X0Y102_I;
  assign CLBLM_R_X11Y107_SLICE_X14Y107_D5 = RIOB33_X105Y111_IOB_X1Y111_I;
  assign CLBLM_R_X11Y107_SLICE_X14Y107_D6 = RIOB33_X105Y109_IOB_X1Y110_I;
  assign LIOI3_TBYTETERM_X0Y113_ILOGIC_X0Y114_D = LIOB33_X0Y113_IOB_X0Y114_I;
  assign LIOI3_TBYTETERM_X0Y113_ILOGIC_X0Y113_D = LIOB33_X0Y113_IOB_X0Y113_I;
  assign CLBLM_L_X8Y104_SLICE_X11Y104_A1 = CLBLM_R_X7Y105_SLICE_X8Y105_AO6;
  assign CLBLM_L_X8Y104_SLICE_X11Y104_A2 = CLBLM_R_X7Y104_SLICE_X9Y104_AO5;
  assign CLBLM_L_X8Y104_SLICE_X11Y104_A3 = CLBLM_L_X10Y104_SLICE_X12Y104_CO6;
  assign CLBLM_L_X8Y104_SLICE_X11Y104_A4 = CLBLM_L_X8Y104_SLICE_X11Y104_BO6;
  assign CLBLM_L_X8Y104_SLICE_X11Y104_A5 = CLBLM_L_X8Y103_SLICE_X11Y103_AO6;
  assign CLBLM_L_X8Y104_SLICE_X11Y104_A6 = CLBLM_L_X8Y105_SLICE_X11Y105_AO5;
  assign CLBLM_L_X8Y104_SLICE_X11Y104_B1 = RIOB33_X105Y101_IOB_X1Y101_I;
  assign CLBLM_L_X8Y104_SLICE_X11Y104_B2 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLM_L_X8Y104_SLICE_X11Y104_B3 = LIOB33_X0Y101_IOB_X0Y102_I;
  assign CLBLM_L_X8Y104_SLICE_X11Y104_B4 = CLBLM_R_X7Y104_SLICE_X8Y104_DO6;
  assign CLBLM_L_X8Y104_SLICE_X11Y104_B5 = CLBLM_L_X8Y104_SLICE_X10Y104_DO6;
  assign CLBLM_L_X8Y104_SLICE_X11Y104_B6 = LIOB33_X0Y103_IOB_X0Y104_I;
  assign CLBLM_L_X8Y104_SLICE_X11Y104_C1 = RIOB33_X105Y101_IOB_X1Y101_I;
  assign CLBLM_L_X8Y104_SLICE_X11Y104_C2 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLM_L_X8Y104_SLICE_X11Y104_C3 = LIOB33_X0Y105_IOB_X0Y105_I;
  assign CLBLM_L_X8Y104_SLICE_X11Y104_C4 = LIOB33_X0Y103_IOB_X0Y104_I;
  assign CLBLM_L_X8Y104_SLICE_X11Y104_C5 = CLBLM_L_X8Y103_SLICE_X11Y103_BO6;
  assign CLBLM_L_X8Y104_SLICE_X11Y104_C6 = CLBLM_L_X8Y104_SLICE_X11Y104_BO6;
  assign CLBLM_L_X8Y104_SLICE_X11Y104_D1 = CLBLM_L_X8Y103_SLICE_X11Y103_AO6;
  assign CLBLM_L_X8Y104_SLICE_X11Y104_D2 = CLBLM_L_X8Y105_SLICE_X11Y105_AO5;
  assign CLBLM_L_X8Y104_SLICE_X11Y104_D3 = CLBLM_R_X7Y104_SLICE_X9Y104_AO5;
  assign CLBLM_L_X8Y104_SLICE_X11Y104_D4 = CLBLM_R_X7Y105_SLICE_X8Y105_AO6;
  assign CLBLM_L_X8Y104_SLICE_X11Y104_D5 = CLBLM_L_X10Y104_SLICE_X12Y104_CO6;
  assign CLBLM_L_X8Y104_SLICE_X11Y104_D6 = CLBLM_L_X8Y104_SLICE_X11Y104_BO6;
  assign CLBLL_L_X4Y110_SLICE_X4Y110_A1 = LIOB33_X0Y113_IOB_X0Y113_I;
  assign CLBLL_L_X4Y110_SLICE_X4Y110_A2 = CLBLM_R_X7Y110_SLICE_X8Y110_AO6;
  assign CLBLL_L_X4Y110_SLICE_X4Y110_A3 = CLBLM_R_X5Y109_SLICE_X7Y109_BO6;
  assign CLBLL_L_X4Y110_SLICE_X4Y110_A4 = LIOB33_X0Y113_IOB_X0Y114_I;
  assign CLBLM_L_X8Y104_SLICE_X10Y104_A3 = RIOB33_X105Y101_IOB_X1Y101_I;
  assign CLBLL_L_X4Y110_SLICE_X4Y110_A5 = LIOB33_X0Y115_IOB_X0Y116_I;
  assign CLBLM_L_X8Y104_SLICE_X10Y104_A4 = 1'b1;
  assign CLBLM_L_X8Y104_SLICE_X10Y104_A5 = LIOB33_X0Y101_IOB_X0Y102_I;
  assign CLBLM_L_X8Y104_SLICE_X10Y104_A6 = 1'b1;
  assign CLBLL_L_X4Y110_SLICE_X4Y110_A6 = LIOB33_X0Y115_IOB_X0Y115_I;
  assign CLBLL_L_X4Y110_SLICE_X4Y110_B1 = LIOB33_X0Y113_IOB_X0Y113_I;
  assign CLBLM_L_X8Y104_SLICE_X10Y104_A1 = LIOB33_X0Y101_IOB_X0Y101_I;
  assign CLBLL_L_X4Y110_SLICE_X4Y110_B3 = CLBLM_R_X5Y109_SLICE_X7Y109_BO6;
  assign CLBLL_L_X4Y110_SLICE_X4Y110_B2 = LIOB33_X0Y115_IOB_X0Y116_I;
  assign CLBLL_L_X4Y110_SLICE_X4Y110_B4 = LIOB33_X0Y113_IOB_X0Y114_I;
  assign CLBLL_L_X4Y110_SLICE_X4Y110_B5 = CLBLM_R_X7Y110_SLICE_X8Y110_AO6;
  assign CLBLL_L_X4Y110_SLICE_X4Y110_B6 = LIOB33_X0Y115_IOB_X0Y115_I;
  assign CLBLM_L_X8Y104_SLICE_X10Y104_B1 = CLBLM_L_X8Y103_SLICE_X10Y103_BO6;
  assign CLBLM_L_X8Y104_SLICE_X10Y104_B2 = CLBLM_L_X10Y104_SLICE_X12Y104_AO6;
  assign CLBLL_L_X4Y110_SLICE_X4Y110_C2 = 1'b1;
  assign CLBLL_L_X4Y110_SLICE_X4Y110_C3 = 1'b1;
  assign CLBLM_L_X8Y104_SLICE_X10Y104_B3 = CLBLM_R_X7Y103_SLICE_X8Y103_BO6;
  assign CLBLL_L_X4Y110_SLICE_X4Y110_C5 = 1'b1;
  assign CLBLL_L_X4Y110_SLICE_X4Y110_C6 = 1'b1;
  assign CLBLM_L_X8Y104_SLICE_X10Y104_B5 = CLBLM_L_X8Y104_SLICE_X10Y104_AO6;
  assign CLBLM_L_X8Y104_SLICE_X10Y104_C4 = CLBLM_L_X8Y104_SLICE_X10Y104_AO5;
  assign CLBLM_L_X8Y104_SLICE_X10Y104_C5 = CLBLM_L_X8Y104_SLICE_X10Y104_AO6;
  assign CLBLM_L_X8Y104_SLICE_X10Y104_C6 = CLBLM_L_X8Y103_SLICE_X10Y103_BO6;
  assign CLBLL_L_X4Y110_SLICE_X4Y110_C4 = 1'b1;
  assign CLBLM_L_X8Y104_SLICE_X10Y104_C1 = CLBLM_R_X7Y103_SLICE_X8Y103_BO6;
  assign CLBLM_L_X8Y104_SLICE_X10Y104_C2 = CLBLM_L_X10Y102_SLICE_X12Y102_AO6;
  assign CLBLM_L_X8Y104_SLICE_X10Y104_C3 = CLBLM_L_X10Y104_SLICE_X12Y104_AO6;
  assign CLBLL_L_X4Y110_SLICE_X4Y110_D1 = 1'b1;
  assign CLBLL_L_X4Y110_SLICE_X4Y110_D2 = 1'b1;
  assign CLBLL_L_X4Y110_SLICE_X4Y110_D3 = 1'b1;
  assign CLBLL_L_X4Y110_SLICE_X4Y110_D4 = 1'b1;
  assign CLBLL_L_X4Y110_SLICE_X4Y110_D5 = 1'b1;
  assign CLBLM_L_X8Y104_SLICE_X10Y104_D1 = CLBLM_R_X7Y103_SLICE_X8Y103_BO6;
  assign CLBLM_L_X8Y104_SLICE_X10Y104_D2 = RIOB33_X105Y101_IOB_X1Y102_I;
  assign CLBLM_L_X8Y104_SLICE_X10Y104_D3 = LIOB33_X0Y101_IOB_X0Y101_I;
  assign CLBLM_L_X8Y104_SLICE_X10Y104_D4 = CLBLM_L_X10Y104_SLICE_X12Y104_AO6;
  assign CLBLM_L_X8Y104_SLICE_X10Y104_D5 = RIOB33_X105Y101_IOB_X1Y101_I;
  assign CLBLM_L_X8Y104_SLICE_X10Y104_D6 = CLBLM_L_X8Y103_SLICE_X10Y103_BO6;
  assign CLBLL_L_X4Y110_SLICE_X4Y110_D6 = 1'b1;
  assign CLBLL_L_X4Y110_SLICE_X5Y110_A1 = CLBLL_L_X4Y109_SLICE_X5Y109_DO6;
  assign CLBLL_L_X4Y110_SLICE_X5Y110_A2 = CLBLL_L_X4Y109_SLICE_X4Y109_BO6;
  assign CLBLL_L_X4Y110_SLICE_X5Y110_A3 = CLBLL_L_X4Y109_SLICE_X5Y109_BO6;
  assign CLBLL_L_X4Y110_SLICE_X5Y110_A4 = CLBLL_L_X4Y109_SLICE_X5Y109_CO6;
  assign CLBLL_L_X4Y110_SLICE_X5Y110_A5 = CLBLL_L_X4Y110_SLICE_X4Y110_AO6;
  assign CLBLL_L_X4Y110_SLICE_X5Y110_A6 = 1'b1;
  assign CLBLM_R_X11Y108_SLICE_X15Y108_A1 = CLBLM_R_X11Y111_SLICE_X15Y111_AO5;
  assign CLBLM_R_X11Y108_SLICE_X15Y108_A2 = CLBLM_L_X12Y107_SLICE_X16Y107_CO6;
  assign CLBLM_R_X11Y108_SLICE_X15Y108_A3 = CLBLM_R_X11Y107_SLICE_X14Y107_AO5;
  assign CLBLM_R_X11Y108_SLICE_X15Y108_A4 = CLBLM_R_X11Y105_SLICE_X15Y105_AO5;
  assign CLBLM_R_X11Y108_SLICE_X15Y108_A5 = CLBLM_R_X11Y107_SLICE_X14Y107_CO6;
  assign CLBLM_R_X11Y108_SLICE_X15Y108_A6 = CLBLM_R_X11Y105_SLICE_X15Y105_CO6;
  assign CLBLL_L_X4Y110_SLICE_X5Y110_B1 = LIOB33_X0Y115_IOB_X0Y115_I;
  assign CLBLL_L_X4Y110_SLICE_X5Y110_B2 = LIOB33_X0Y113_IOB_X0Y114_I;
  assign CLBLL_L_X4Y110_SLICE_X5Y110_B3 = 1'b1;
  assign CLBLL_L_X4Y110_SLICE_X5Y110_B4 = 1'b1;
  assign CLBLL_L_X4Y110_SLICE_X5Y110_B5 = LIOB33_X0Y103_IOB_X0Y103_I;
  assign CLBLL_L_X4Y110_SLICE_X5Y110_B6 = 1'b1;
  assign CLBLM_R_X5Y113_SLICE_X7Y113_D6 = 1'b1;
  assign CLBLM_R_X11Y108_SLICE_X15Y108_B4 = CLBLM_R_X11Y105_SLICE_X15Y105_AO5;
  assign CLBLM_R_X11Y108_SLICE_X15Y108_B5 = CLBLM_R_X11Y107_SLICE_X14Y107_CO6;
  assign CLBLM_R_X11Y108_SLICE_X15Y108_B6 = CLBLM_R_X11Y105_SLICE_X15Y105_CO6;
  assign CLBLL_L_X4Y110_SLICE_X5Y110_C1 = CLBLL_L_X4Y109_SLICE_X5Y109_AO6;
  assign CLBLL_L_X4Y110_SLICE_X5Y110_C2 = CLBLL_L_X4Y108_SLICE_X5Y108_CO6;
  assign CLBLM_R_X11Y108_SLICE_X15Y108_C1 = CLBLM_R_X11Y107_SLICE_X14Y107_CO6;
  assign CLBLM_R_X11Y108_SLICE_X15Y108_C2 = CLBLM_L_X12Y107_SLICE_X16Y107_CO6;
  assign CLBLL_L_X4Y110_SLICE_X5Y110_C4 = CLBLL_L_X4Y109_SLICE_X5Y109_CO6;
  assign CLBLL_L_X4Y110_SLICE_X5Y110_C5 = CLBLL_L_X4Y110_SLICE_X4Y110_AO6;
  assign CLBLM_R_X11Y108_SLICE_X15Y108_C5 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLL_L_X4Y110_SLICE_X5Y110_D1 = CLBLL_L_X4Y109_SLICE_X5Y109_CO6;
  assign CLBLL_L_X4Y110_SLICE_X5Y110_D2 = CLBLL_L_X4Y109_SLICE_X5Y109_BO6;
  assign CLBLL_L_X4Y110_SLICE_X5Y110_D3 = CLBLL_L_X4Y109_SLICE_X5Y109_DO6;
  assign CLBLL_L_X4Y110_SLICE_X5Y110_D4 = CLBLL_L_X4Y110_SLICE_X4Y110_AO6;
  assign CLBLL_L_X4Y110_SLICE_X5Y110_D5 = CLBLL_L_X4Y112_SLICE_X4Y112_DO6;
  assign CLBLL_L_X4Y110_SLICE_X5Y110_D6 = CLBLL_L_X4Y109_SLICE_X4Y109_BO6;
  assign CLBLM_R_X11Y108_SLICE_X15Y108_C6 = LIOB33_X0Y105_IOB_X0Y105_I;
  assign CLBLM_R_X11Y108_SLICE_X15Y108_D1 = RIOB33_X105Y107_IOB_X1Y107_I;
  assign CLBLM_R_X11Y108_SLICE_X15Y108_D2 = LIOB33_X0Y105_IOB_X0Y105_I;
  assign CLBLM_R_X11Y108_SLICE_X15Y108_D3 = CLBLM_L_X12Y107_SLICE_X17Y107_AO5;
  assign CLBLM_R_X11Y108_SLICE_X15Y108_D4 = LIOB33_X0Y103_IOB_X0Y104_I;
  assign CLBLM_R_X11Y108_SLICE_X15Y108_D5 = CLBLM_L_X12Y107_SLICE_X17Y107_DO6;
  assign CLBLM_R_X11Y108_SLICE_X15Y108_D6 = RIOB33_X105Y107_IOB_X1Y108_I;
  assign CLBLM_R_X11Y108_SLICE_X14Y108_A1 = RIOB33_X105Y103_IOB_X1Y104_I;
  assign CLBLM_R_X11Y108_SLICE_X14Y108_A2 = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLM_R_X11Y108_SLICE_X14Y108_A3 = CLBLM_R_X11Y108_SLICE_X15Y108_CO6;
  assign CLBLM_R_X11Y108_SLICE_X14Y108_A4 = CLBLM_R_X11Y108_SLICE_X14Y108_BO6;
  assign CLBLM_R_X11Y108_SLICE_X14Y108_A5 = RIOB33_X105Y103_IOB_X1Y103_I;
  assign CLBLM_R_X11Y108_SLICE_X14Y108_A6 = CLBLM_R_X11Y108_SLICE_X14Y108_CO6;
  assign CLBLM_R_X11Y108_SLICE_X14Y108_B1 = CLBLM_L_X12Y106_SLICE_X16Y106_CO6;
  assign CLBLM_R_X11Y108_SLICE_X14Y108_B2 = CLBLM_R_X11Y105_SLICE_X15Y105_CO6;
  assign CLBLM_R_X11Y108_SLICE_X14Y108_B3 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X11Y108_SLICE_X14Y108_B4 = RIOB33_X105Y103_IOB_X1Y104_I;
  assign CLBLM_R_X11Y108_SLICE_X14Y108_B5 = LIOB33_X0Y103_IOB_X0Y104_I;
  assign CLBLM_R_X11Y108_SLICE_X14Y108_B6 = LIOB33_X0Y105_IOB_X0Y105_I;
  assign CLBLM_R_X11Y108_SLICE_X14Y108_C1 = LIOB33_X0Y103_IOB_X0Y104_I;
  assign CLBLM_R_X11Y108_SLICE_X14Y108_C2 = RIOB33_X105Y103_IOB_X1Y104_I;
  assign CLBLM_R_X11Y108_SLICE_X14Y108_C3 = RIOB33_X105Y103_IOB_X1Y103_I;
  assign CLBLM_R_X11Y108_SLICE_X14Y108_C4 = LIOB33_X0Y105_IOB_X0Y105_I;
  assign CLBLM_R_X11Y108_SLICE_X14Y108_C5 = CLBLM_R_X11Y105_SLICE_X15Y105_DO6;
  assign CLBLM_R_X11Y108_SLICE_X14Y108_C6 = CLBLM_R_X11Y105_SLICE_X14Y105_DO6;
  assign CLBLM_R_X11Y108_SLICE_X14Y108_D1 = RIOB33_X105Y103_IOB_X1Y103_I;
  assign CLBLM_R_X11Y108_SLICE_X14Y108_D2 = LIOB33_X0Y103_IOB_X0Y104_I;
  assign CLBLM_R_X11Y108_SLICE_X14Y108_D3 = RIOB33_X105Y103_IOB_X1Y104_I;
  assign CLBLM_R_X11Y108_SLICE_X14Y108_D4 = LIOB33_X0Y105_IOB_X0Y105_I;
  assign CLBLM_R_X11Y108_SLICE_X14Y108_D5 = CLBLM_R_X11Y105_SLICE_X15Y105_DO6;
  assign CLBLM_R_X11Y108_SLICE_X14Y108_D6 = CLBLM_R_X11Y105_SLICE_X14Y105_DO6;
  assign CLBLM_R_X5Y113_SLICE_X6Y113_B6 = 1'b1;
  assign CLBLM_R_X5Y113_SLICE_X6Y113_C4 = 1'b1;
  assign CLBLM_R_X5Y113_SLICE_X6Y113_C5 = 1'b1;
  assign CLBLM_R_X5Y113_SLICE_X6Y113_C6 = 1'b1;
  assign CLBLM_L_X8Y105_SLICE_X11Y105_A1 = 1'b1;
  assign CLBLM_L_X8Y105_SLICE_X11Y105_A2 = LIOB33_X0Y103_IOB_X0Y104_I;
  assign CLBLM_L_X8Y105_SLICE_X11Y105_A3 = LIOB33_X0Y105_IOB_X0Y105_I;
  assign CLBLM_L_X8Y105_SLICE_X11Y105_A4 = RIOB33_X105Y101_IOB_X1Y101_I;
  assign CLBLM_L_X8Y105_SLICE_X11Y105_A5 = 1'b1;
  assign CLBLM_L_X8Y105_SLICE_X11Y105_A6 = 1'b1;
  assign CLBLM_L_X8Y105_SLICE_X11Y105_B1 = CLBLM_L_X10Y105_SLICE_X12Y105_CO6;
  assign CLBLM_L_X8Y105_SLICE_X11Y105_B2 = CLBLM_L_X10Y105_SLICE_X13Y105_BO6;
  assign CLBLM_L_X8Y105_SLICE_X11Y105_B3 = CLBLM_L_X8Y105_SLICE_X10Y105_AO5;
  assign CLBLM_L_X8Y105_SLICE_X11Y105_B4 = CLBLM_L_X10Y103_SLICE_X12Y103_DO6;
  assign CLBLM_L_X8Y105_SLICE_X11Y105_B5 = CLBLM_L_X10Y105_SLICE_X13Y105_AO5;
  assign CLBLM_L_X8Y105_SLICE_X11Y105_B6 = CLBLM_L_X8Y105_SLICE_X11Y105_AO5;
  assign CLBLM_L_X8Y105_SLICE_X11Y105_C1 = CLBLM_L_X10Y105_SLICE_X13Y105_AO5;
  assign CLBLM_L_X8Y105_SLICE_X11Y105_C2 = CLBLM_L_X10Y105_SLICE_X13Y105_BO6;
  assign CLBLM_L_X8Y105_SLICE_X11Y105_C3 = CLBLM_L_X8Y105_SLICE_X11Y105_AO5;
  assign CLBLM_L_X8Y105_SLICE_X11Y105_C4 = CLBLM_L_X10Y105_SLICE_X12Y105_CO6;
  assign CLBLM_L_X8Y105_SLICE_X11Y105_C5 = CLBLM_L_X10Y103_SLICE_X12Y103_DO6;
  assign CLBLM_L_X8Y105_SLICE_X11Y105_C6 = CLBLM_L_X8Y105_SLICE_X10Y105_AO5;
  assign CLBLM_L_X8Y105_SLICE_X11Y105_D1 = RIOB33_X105Y101_IOB_X1Y102_I;
  assign CLBLM_L_X8Y105_SLICE_X11Y105_D2 = CLBLM_L_X10Y105_SLICE_X13Y105_BO6;
  assign CLBLM_L_X8Y105_SLICE_X11Y105_D3 = RIOB33_X105Y101_IOB_X1Y101_I;
  assign CLBLM_L_X8Y105_SLICE_X11Y105_D4 = CLBLM_L_X10Y103_SLICE_X12Y103_DO6;
  assign CLBLM_L_X8Y105_SLICE_X11Y105_D5 = CLBLM_L_X10Y105_SLICE_X12Y105_CO6;
  assign CLBLM_L_X8Y105_SLICE_X11Y105_D6 = LIOB33_X0Y105_IOB_X0Y105_I;
  assign CLBLL_L_X4Y111_SLICE_X4Y111_A1 = CLBLL_L_X4Y111_SLICE_X4Y111_BO6;
  assign CLBLL_L_X4Y111_SLICE_X4Y111_A2 = CLBLL_L_X4Y110_SLICE_X4Y110_BO6;
  assign CLBLL_L_X4Y111_SLICE_X4Y111_A3 = CLBLL_L_X4Y110_SLICE_X5Y110_CO6;
  assign CLBLL_L_X4Y111_SLICE_X4Y111_A4 = CLBLL_L_X4Y112_SLICE_X4Y112_BO6;
  assign CLBLL_L_X4Y111_SLICE_X4Y111_A5 = CLBLL_L_X4Y111_SLICE_X4Y111_CO6;
  assign CLBLL_L_X4Y111_SLICE_X4Y111_A6 = 1'b1;
  assign CLBLM_L_X8Y105_SLICE_X10Y105_A1 = RIOB33_X105Y101_IOB_X1Y101_I;
  assign CLBLM_L_X8Y105_SLICE_X10Y105_A3 = LIOB33_X0Y115_IOB_X0Y116_I;
  assign CLBLM_L_X8Y105_SLICE_X10Y105_A4 = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLM_L_X8Y105_SLICE_X10Y105_A5 = 1'b1;
  assign CLBLM_L_X8Y105_SLICE_X10Y105_A6 = 1'b1;
  assign CLBLL_L_X4Y111_SLICE_X4Y111_B4 = CLBLM_R_X7Y112_SLICE_X9Y112_AO6;
  assign CLBLL_L_X4Y111_SLICE_X4Y111_B5 = LIOB33_X0Y115_IOB_X0Y115_I;
  assign CLBLL_L_X4Y111_SLICE_X4Y111_B6 = LIOB33_X0Y113_IOB_X0Y113_I;
  assign CLBLM_L_X8Y105_SLICE_X10Y105_A2 = 1'b1;
  assign CLBLL_L_X4Y111_SLICE_X4Y111_B1 = CLBLM_R_X7Y112_SLICE_X9Y112_BO6;
  assign CLBLL_L_X4Y111_SLICE_X4Y111_B2 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLL_L_X4Y111_SLICE_X4Y111_C2 = CLBLM_R_X7Y112_SLICE_X9Y112_AO6;
  assign CLBLL_L_X4Y111_SLICE_X4Y111_C3 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLM_L_X8Y105_SLICE_X10Y105_B1 = CLBLM_R_X7Y105_SLICE_X8Y105_AO6;
  assign CLBLL_L_X4Y111_SLICE_X4Y111_C5 = CLBLM_R_X7Y112_SLICE_X9Y112_BO6;
  assign CLBLM_L_X8Y105_SLICE_X10Y105_B2 = CLBLM_L_X8Y104_SLICE_X11Y104_CO6;
  assign CLBLL_L_X4Y111_SLICE_X4Y111_C1 = LIOB33_X0Y115_IOB_X0Y115_I;
  assign CLBLM_L_X8Y105_SLICE_X10Y105_B3 = LIOB33_X0Y115_IOB_X0Y116_I;
  assign CLBLM_L_X8Y105_SLICE_X10Y105_B4 = LIOB33_X0Y107_IOB_X0Y107_I;
  assign CLBLL_L_X4Y111_SLICE_X4Y111_C4 = LIOB33_X0Y113_IOB_X0Y113_I;
  assign CLBLM_L_X8Y105_SLICE_X10Y105_B5 = CLBLM_R_X7Y105_SLICE_X9Y105_BO6;
  assign CLBLL_L_X4Y111_SLICE_X4Y111_C6 = LIOB33_X0Y115_IOB_X0Y116_I;
  assign CLBLM_L_X8Y105_SLICE_X10Y105_B6 = CLBLM_L_X8Y106_SLICE_X11Y106_AO6;
  assign CLBLL_L_X4Y111_SLICE_X4Y111_D1 = CLBLM_L_X8Y112_SLICE_X10Y112_DO6;
  assign CLBLL_L_X4Y111_SLICE_X4Y111_D2 = CLBLL_L_X4Y110_SLICE_X5Y110_CO6;
  assign CLBLL_L_X4Y111_SLICE_X4Y111_D3 = CLBLM_R_X7Y112_SLICE_X9Y112_BO6;
  assign CLBLM_L_X8Y105_SLICE_X10Y105_C1 = 1'b1;
  assign CLBLM_L_X8Y105_SLICE_X10Y105_C2 = 1'b1;
  assign CLBLM_L_X8Y105_SLICE_X10Y105_C3 = 1'b1;
  assign CLBLM_L_X8Y105_SLICE_X10Y105_C4 = 1'b1;
  assign CLBLM_L_X8Y105_SLICE_X10Y105_C5 = 1'b1;
  assign CLBLM_L_X8Y105_SLICE_X10Y105_C6 = 1'b1;
  assign CLBLL_L_X4Y111_SLICE_X4Y111_D4 = CLBLL_L_X4Y114_SLICE_X4Y114_AO6;
  assign CLBLL_L_X4Y111_SLICE_X4Y111_D5 = CLBLL_L_X4Y110_SLICE_X4Y110_BO6;
  assign CLBLL_L_X4Y111_SLICE_X4Y111_D6 = CLBLL_L_X4Y112_SLICE_X4Y112_BO6;
  assign CLBLM_L_X8Y105_SLICE_X10Y105_D1 = 1'b1;
  assign CLBLM_L_X8Y105_SLICE_X10Y105_D2 = 1'b1;
  assign CLBLM_L_X8Y105_SLICE_X10Y105_D3 = 1'b1;
  assign CLBLM_L_X8Y105_SLICE_X10Y105_D4 = 1'b1;
  assign CLBLM_L_X8Y105_SLICE_X10Y105_D5 = 1'b1;
  assign CLBLM_L_X8Y105_SLICE_X10Y105_D6 = 1'b1;
  assign CLBLL_L_X4Y111_SLICE_X5Y111_A1 = CLBLM_R_X7Y112_SLICE_X8Y112_CO6;
  assign CLBLL_L_X4Y111_SLICE_X5Y111_A2 = 1'b1;
  assign CLBLL_L_X4Y111_SLICE_X5Y111_A3 = RIOB33_X105Y101_IOB_X1Y101_I;
  assign CLBLL_L_X4Y111_SLICE_X5Y111_A4 = CLBLL_L_X4Y109_SLICE_X5Y109_AO5;
  assign CLBLL_L_X4Y111_SLICE_X5Y111_A5 = LIOB33_X0Y115_IOB_X0Y115_I;
  assign CLBLL_L_X4Y111_SLICE_X5Y111_A6 = 1'b1;
  assign CLBLL_L_X4Y111_SLICE_X5Y111_B1 = CLBLM_R_X7Y112_SLICE_X8Y112_CO6;
  assign CLBLL_L_X4Y111_SLICE_X5Y111_B2 = CLBLL_L_X4Y111_SLICE_X4Y111_DO6;
  assign CLBLL_L_X4Y111_SLICE_X5Y111_B3 = CLBLL_L_X4Y109_SLICE_X5Y109_AO5;
  assign CLBLL_L_X4Y111_SLICE_X5Y111_B4 = CLBLM_R_X5Y112_SLICE_X6Y112_BO6;
  assign CLBLL_L_X4Y111_SLICE_X5Y111_B5 = CLBLL_L_X4Y112_SLICE_X4Y112_CO6;
  assign CLBLL_L_X4Y111_SLICE_X5Y111_B6 = CLBLL_L_X4Y111_SLICE_X5Y111_AO5;
  assign CLBLM_R_X11Y109_SLICE_X15Y109_A1 = CLBLM_R_X11Y106_SLICE_X14Y106_CO6;
  assign CLBLM_R_X11Y109_SLICE_X15Y109_A2 = CLBLM_R_X11Y108_SLICE_X15Y108_BO6;
  assign CLBLM_R_X11Y109_SLICE_X15Y109_A3 = CLBLM_R_X11Y108_SLICE_X15Y108_AO6;
  assign CLBLL_L_X4Y111_SLICE_X5Y111_C1 = CLBLM_L_X8Y112_SLICE_X10Y112_DO6;
  assign CLBLL_L_X4Y111_SLICE_X5Y111_C2 = CLBLL_L_X4Y114_SLICE_X4Y114_AO6;
  assign CLBLL_L_X4Y111_SLICE_X5Y111_C3 = CLBLM_R_X7Y112_SLICE_X9Y112_DO6;
  assign CLBLL_L_X4Y111_SLICE_X5Y111_C4 = CLBLM_R_X7Y112_SLICE_X9Y112_BO6;
  assign CLBLL_L_X4Y111_SLICE_X5Y111_C5 = CLBLL_L_X4Y110_SLICE_X5Y110_BO5;
  assign CLBLL_L_X4Y111_SLICE_X5Y111_C6 = CLBLM_R_X5Y109_SLICE_X7Y109_BO6;
  assign CLBLM_R_X11Y109_SLICE_X15Y109_A4 = CLBLM_R_X11Y107_SLICE_X15Y107_BO6;
  assign CLBLM_R_X11Y109_SLICE_X15Y109_A5 = CLBLM_L_X10Y108_SLICE_X13Y108_BO5;
  assign CLBLM_R_X11Y109_SLICE_X15Y109_A6 = CLBLM_R_X11Y111_SLICE_X15Y111_AO6;
  assign CLBLM_R_X11Y109_SLICE_X15Y109_B5 = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLM_R_X11Y109_SLICE_X15Y109_B6 = CLBLM_R_X11Y108_SLICE_X15Y108_CO6;
  assign CLBLM_R_X11Y109_SLICE_X15Y109_B1 = CLBLM_R_X11Y106_SLICE_X14Y106_CO6;
  assign CLBLM_R_X11Y109_SLICE_X15Y109_B2 = RIOB33_X105Y103_IOB_X1Y104_I;
  assign CLBLM_R_X11Y109_SLICE_X15Y109_B3 = LIOB33_X0Y107_IOB_X0Y107_I;
  assign CLBLM_R_X11Y109_SLICE_X15Y109_B4 = RIOB33_X105Y103_IOB_X1Y103_I;
  assign CLBLL_L_X4Y111_SLICE_X5Y111_D1 = CLBLM_R_X5Y111_SLICE_X6Y111_AO6;
  assign CLBLL_L_X4Y111_SLICE_X5Y111_D2 = CLBLL_L_X4Y111_SLICE_X4Y111_CO6;
  assign CLBLL_L_X4Y111_SLICE_X5Y111_D3 = CLBLL_L_X4Y112_SLICE_X4Y112_CO6;
  assign CLBLL_L_X4Y111_SLICE_X5Y111_D4 = CLBLL_L_X4Y111_SLICE_X5Y111_CO6;
  assign CLBLL_L_X4Y111_SLICE_X5Y111_D5 = CLBLL_L_X4Y110_SLICE_X5Y110_DO6;
  assign CLBLL_L_X4Y111_SLICE_X5Y111_D6 = CLBLL_L_X4Y112_SLICE_X4Y112_BO6;
  assign CLBLM_R_X11Y109_SLICE_X15Y109_C1 = CLBLM_L_X12Y109_SLICE_X16Y109_BO6;
  assign CLBLM_R_X11Y109_SLICE_X15Y109_C2 = LIOB33_X0Y107_IOB_X0Y107_I;
  assign CLBLM_R_X11Y109_SLICE_X15Y109_C3 = CLBLM_L_X12Y108_SLICE_X17Y108_DO6;
  assign CLBLM_R_X11Y109_SLICE_X15Y109_C4 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X11Y109_SLICE_X15Y109_C5 = CLBLM_R_X11Y108_SLICE_X15Y108_DO6;
  assign CLBLM_R_X11Y109_SLICE_X15Y109_C6 = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLM_R_X11Y109_SLICE_X15Y109_D1 = CLBLM_L_X12Y109_SLICE_X16Y109_BO6;
  assign CLBLM_R_X11Y109_SLICE_X15Y109_D2 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X11Y109_SLICE_X15Y109_D3 = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLM_R_X11Y109_SLICE_X15Y109_D4 = CLBLM_L_X12Y108_SLICE_X17Y108_DO6;
  assign CLBLM_R_X11Y109_SLICE_X15Y109_D5 = CLBLM_R_X11Y108_SLICE_X15Y108_DO6;
  assign CLBLM_R_X11Y109_SLICE_X15Y109_D6 = LIOB33_X0Y107_IOB_X0Y107_I;
  assign LIOI3_TBYTETERM_X0Y137_OLOGIC_X0Y137_T1 = 1'b1;
  assign CLBLM_R_X11Y109_SLICE_X14Y109_A1 = 1'b1;
  assign CLBLM_R_X11Y109_SLICE_X14Y109_A2 = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLM_R_X11Y109_SLICE_X14Y109_A3 = LIOB33_X0Y107_IOB_X0Y108_I;
  assign CLBLM_R_X11Y109_SLICE_X14Y109_A4 = RIOB33_X105Y103_IOB_X1Y103_I;
  assign CLBLM_R_X11Y109_SLICE_X14Y109_A5 = 1'b1;
  assign CLBLM_R_X11Y109_SLICE_X14Y109_A6 = 1'b1;
  assign CLBLM_R_X11Y109_SLICE_X14Y109_B1 = CLBLM_R_X11Y110_SLICE_X15Y110_AO6;
  assign CLBLM_R_X11Y109_SLICE_X14Y109_B2 = CLBLM_L_X10Y109_SLICE_X13Y109_BO6;
  assign CLBLM_R_X11Y109_SLICE_X14Y109_B3 = CLBLM_R_X11Y109_SLICE_X15Y109_AO6;
  assign CLBLM_R_X11Y109_SLICE_X14Y109_B4 = CLBLM_L_X10Y109_SLICE_X13Y109_AO6;
  assign CLBLM_R_X11Y109_SLICE_X14Y109_B5 = CLBLM_R_X11Y109_SLICE_X14Y109_AO5;
  assign CLBLM_R_X11Y109_SLICE_X14Y109_B6 = CLBLM_R_X11Y109_SLICE_X14Y109_CO6;
  assign CLBLM_R_X11Y109_SLICE_X14Y109_C1 = RIOB33_X105Y103_IOB_X1Y103_I;
  assign CLBLM_R_X11Y109_SLICE_X14Y109_C2 = CLBLM_R_X11Y108_SLICE_X15Y108_CO6;
  assign CLBLM_R_X11Y109_SLICE_X14Y109_C3 = CLBLM_R_X11Y106_SLICE_X14Y106_CO6;
  assign CLBLM_R_X11Y109_SLICE_X14Y109_C4 = LIOB33_X0Y107_IOB_X0Y107_I;
  assign CLBLM_R_X11Y109_SLICE_X14Y109_C5 = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLM_R_X11Y109_SLICE_X14Y109_C6 = RIOB33_X105Y103_IOB_X1Y104_I;
  assign CLBLM_R_X11Y109_SLICE_X14Y109_D1 = CLBLM_R_X11Y109_SLICE_X14Y109_AO5;
  assign CLBLM_R_X11Y109_SLICE_X14Y109_D2 = CLBLM_L_X10Y109_SLICE_X13Y109_BO6;
  assign CLBLM_R_X11Y109_SLICE_X14Y109_D3 = CLBLM_R_X11Y109_SLICE_X15Y109_AO6;
  assign CLBLM_R_X11Y109_SLICE_X14Y109_D4 = CLBLM_R_X11Y109_SLICE_X14Y109_CO6;
  assign CLBLM_R_X11Y109_SLICE_X14Y109_D5 = CLBLM_R_X11Y110_SLICE_X15Y110_AO6;
  assign CLBLM_R_X11Y109_SLICE_X14Y109_D6 = CLBLM_L_X10Y109_SLICE_X13Y109_AO6;
  assign LIOI3_X0Y109_ILOGIC_X0Y110_D = LIOB33_X0Y109_IOB_X0Y110_I;
  assign LIOI3_X0Y109_ILOGIC_X0Y109_D = LIOB33_X0Y109_IOB_X0Y109_I;
  assign CLBLM_L_X8Y106_SLICE_X11Y106_A1 = LIOB33_X0Y105_IOB_X0Y105_I;
  assign CLBLM_L_X8Y106_SLICE_X11Y106_A2 = CLBLM_L_X10Y103_SLICE_X12Y103_DO6;
  assign CLBLM_L_X8Y106_SLICE_X11Y106_A3 = RIOB33_X105Y101_IOB_X1Y102_I;
  assign CLBLM_L_X8Y106_SLICE_X11Y106_A4 = LIOB33_X0Y103_IOB_X0Y104_I;
  assign CLBLM_L_X8Y106_SLICE_X11Y106_A5 = CLBLM_L_X10Y105_SLICE_X12Y105_BO6;
  assign CLBLM_L_X8Y106_SLICE_X11Y106_A6 = RIOB33_X105Y101_IOB_X1Y101_I;
  assign CLBLM_L_X8Y106_SLICE_X11Y106_B1 = CLBLM_L_X8Y107_SLICE_X11Y107_BO5;
  assign CLBLM_L_X8Y106_SLICE_X11Y106_B2 = CLBLM_L_X8Y107_SLICE_X11Y107_AO6;
  assign CLBLM_L_X8Y106_SLICE_X11Y106_B3 = CLBLM_R_X7Y106_SLICE_X8Y106_AO6;
  assign CLBLM_L_X8Y106_SLICE_X11Y106_B4 = CLBLM_L_X8Y105_SLICE_X10Y105_BO6;
  assign CLBLM_L_X8Y106_SLICE_X11Y106_B5 = CLBLM_L_X8Y106_SLICE_X10Y106_BO6;
  assign CLBLM_L_X8Y106_SLICE_X11Y106_B6 = CLBLM_L_X8Y106_SLICE_X11Y106_CO6;
  assign CLBLM_L_X8Y106_SLICE_X11Y106_C1 = CLBLM_L_X10Y108_SLICE_X13Y108_BO6;
  assign CLBLM_L_X8Y106_SLICE_X11Y106_C2 = CLBLM_L_X8Y106_SLICE_X10Y106_AO5;
  assign CLBLM_L_X8Y106_SLICE_X11Y106_C3 = CLBLM_L_X10Y106_SLICE_X13Y106_DO6;
  assign CLBLM_L_X8Y106_SLICE_X11Y106_C4 = CLBLM_L_X8Y105_SLICE_X11Y105_CO6;
  assign CLBLM_L_X8Y106_SLICE_X11Y106_C5 = CLBLM_L_X8Y104_SLICE_X11Y104_DO6;
  assign CLBLM_L_X8Y106_SLICE_X11Y106_C6 = CLBLM_L_X8Y105_SLICE_X11Y105_BO6;
  assign CLBLM_L_X8Y106_SLICE_X11Y106_D1 = CLBLM_R_X7Y106_SLICE_X8Y106_AO6;
  assign CLBLL_L_X4Y112_SLICE_X4Y112_A1 = CLBLL_L_X4Y111_SLICE_X4Y111_DO6;
  assign CLBLM_L_X8Y106_SLICE_X11Y106_D3 = CLBLM_L_X8Y106_SLICE_X10Y106_BO6;
  assign CLBLM_L_X8Y106_SLICE_X11Y106_D4 = CLBLM_L_X8Y106_SLICE_X11Y106_CO6;
  assign CLBLM_L_X8Y106_SLICE_X11Y106_D5 = CLBLM_L_X8Y107_SLICE_X11Y107_BO5;
  assign CLBLM_L_X8Y106_SLICE_X11Y106_D6 = CLBLM_L_X8Y105_SLICE_X10Y105_BO6;
  assign CLBLL_L_X4Y112_SLICE_X4Y112_A2 = CLBLL_L_X4Y112_SLICE_X4Y112_CO6;
  assign CLBLL_L_X4Y112_SLICE_X4Y112_A3 = CLBLM_R_X5Y112_SLICE_X6Y112_BO6;
  assign CLBLL_L_X4Y112_SLICE_X4Y112_A4 = CLBLL_L_X4Y111_SLICE_X5Y111_AO6;
  assign CLBLL_L_X4Y112_SLICE_X4Y112_A5 = CLBLM_R_X5Y111_SLICE_X6Y111_AO6;
  assign CLBLL_L_X4Y112_SLICE_X4Y112_A6 = 1'b1;
  assign CLBLM_L_X8Y106_SLICE_X10Y106_A1 = 1'b1;
  assign CLBLM_L_X8Y106_SLICE_X10Y106_A2 = LIOB33_X0Y107_IOB_X0Y107_I;
  assign CLBLM_L_X8Y106_SLICE_X10Y106_A3 = LIOB33_X0Y115_IOB_X0Y116_I;
  assign CLBLM_L_X8Y106_SLICE_X10Y106_A4 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLL_L_X4Y112_SLICE_X4Y112_B1 = CLBLM_R_X7Y112_SLICE_X8Y112_AO5;
  assign CLBLL_L_X4Y112_SLICE_X4Y112_B2 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLM_L_X8Y106_SLICE_X10Y106_A5 = 1'b1;
  assign CLBLM_L_X8Y106_SLICE_X10Y106_A6 = 1'b1;
  assign CLBLL_L_X4Y112_SLICE_X4Y112_C1 = LIOB33_X0Y115_IOB_X0Y115_I;
  assign CLBLL_L_X4Y112_SLICE_X4Y112_C2 = RIOB33_X105Y101_IOB_X1Y101_I;
  assign CLBLL_L_X4Y112_SLICE_X4Y112_C3 = CLBLM_R_X7Y112_SLICE_X9Y112_CO6;
  assign CLBLL_L_X4Y112_SLICE_X4Y112_C4 = LIOB33_X0Y113_IOB_X0Y113_I;
  assign CLBLL_L_X4Y112_SLICE_X4Y112_C5 = CLBLM_R_X7Y112_SLICE_X8Y112_AO5;
  assign CLBLL_L_X4Y112_SLICE_X4Y112_C6 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLM_L_X8Y106_SLICE_X10Y106_B1 = LIOB33_X0Y107_IOB_X0Y107_I;
  assign CLBLM_L_X8Y106_SLICE_X10Y106_B2 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLM_L_X8Y106_SLICE_X10Y106_B3 = CLBLM_L_X8Y106_SLICE_X11Y106_AO6;
  assign CLBLM_L_X8Y106_SLICE_X10Y106_B4 = CLBLM_L_X8Y105_SLICE_X11Y105_BO6;
  assign CLBLM_L_X8Y106_SLICE_X10Y106_B5 = CLBLM_L_X8Y104_SLICE_X11Y104_CO6;
  assign CLBLM_L_X8Y106_SLICE_X10Y106_B6 = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLL_L_X4Y112_SLICE_X4Y112_D1 = CLBLL_L_X4Y114_SLICE_X4Y114_AO6;
  assign CLBLL_L_X4Y112_SLICE_X4Y112_D2 = CLBLM_R_X7Y112_SLICE_X9Y112_DO6;
  assign CLBLL_L_X4Y112_SLICE_X4Y112_D3 = CLBLL_L_X4Y110_SLICE_X5Y110_BO5;
  assign CLBLL_L_X4Y112_SLICE_X4Y112_D4 = CLBLM_R_X5Y109_SLICE_X7Y109_BO6;
  assign CLBLL_L_X4Y112_SLICE_X4Y112_D5 = CLBLM_L_X8Y112_SLICE_X10Y112_DO6;
  assign CLBLL_L_X4Y112_SLICE_X4Y112_D6 = CLBLM_R_X7Y112_SLICE_X9Y112_BO6;
  assign CLBLM_L_X8Y106_SLICE_X10Y106_C1 = CLBLM_L_X8Y104_SLICE_X11Y104_CO6;
  assign CLBLM_L_X8Y106_SLICE_X10Y106_C2 = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLM_L_X8Y106_SLICE_X10Y106_C3 = CLBLM_L_X8Y106_SLICE_X11Y106_AO6;
  assign CLBLM_L_X8Y106_SLICE_X10Y106_C4 = CLBLM_L_X8Y105_SLICE_X11Y105_BO6;
  assign CLBLM_L_X8Y106_SLICE_X10Y106_C5 = LIOB33_X0Y107_IOB_X0Y107_I;
  assign CLBLM_L_X8Y106_SLICE_X10Y106_C6 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLM_L_X8Y106_SLICE_X10Y106_D1 = CLBLM_L_X8Y104_SLICE_X11Y104_AO6;
  assign CLBLM_L_X8Y106_SLICE_X10Y106_D2 = CLBLM_L_X8Y106_SLICE_X10Y106_AO6;
  assign CLBLM_L_X8Y106_SLICE_X10Y106_D3 = CLBLM_L_X8Y104_SLICE_X11Y104_DO6;
  assign CLBLM_L_X8Y106_SLICE_X10Y106_D4 = CLBLM_L_X8Y106_SLICE_X10Y106_AO5;
  assign CLBLM_L_X8Y106_SLICE_X10Y106_D5 = CLBLM_R_X7Y105_SLICE_X9Y105_BO6;
  assign CLBLM_L_X8Y106_SLICE_X10Y106_D6 = CLBLM_L_X8Y105_SLICE_X11Y105_BO6;
  assign CLBLL_L_X4Y112_SLICE_X5Y112_A1 = CLBLM_R_X5Y110_SLICE_X7Y110_DO6;
  assign CLBLL_L_X4Y112_SLICE_X5Y112_A2 = LIOB33_X0Y115_IOB_X0Y115_I;
  assign CLBLL_L_X4Y112_SLICE_X5Y112_A3 = RIOB33_X105Y101_IOB_X1Y102_I;
  assign CLBLL_L_X4Y112_SLICE_X5Y112_A4 = RIOB33_X105Y103_IOB_X1Y103_I;
  assign CLBLL_L_X4Y112_SLICE_X5Y112_A5 = CLBLM_R_X5Y111_SLICE_X6Y111_DO6;
  assign CLBLL_L_X4Y112_SLICE_X5Y112_A6 = LIOB33_X0Y113_IOB_X0Y113_I;
  assign CLBLL_L_X4Y112_SLICE_X5Y112_B1 = CLBLM_R_X5Y110_SLICE_X7Y110_DO6;
  assign CLBLL_L_X4Y112_SLICE_X5Y112_B2 = CLBLL_L_X4Y113_SLICE_X5Y113_AO6;
  assign CLBLL_L_X4Y112_SLICE_X5Y112_B3 = CLBLM_R_X5Y112_SLICE_X6Y112_AO6;
  assign CLBLL_L_X4Y112_SLICE_X5Y112_B4 = CLBLM_R_X5Y112_SLICE_X7Y112_AO5;
  assign CLBLL_L_X4Y112_SLICE_X5Y112_B5 = CLBLL_L_X4Y111_SLICE_X5Y111_AO6;
  assign CLBLL_L_X4Y112_SLICE_X5Y112_B6 = CLBLL_L_X4Y111_SLICE_X5Y111_DO6;
  assign CLBLL_L_X4Y111_SLICE_X4Y111_B3 = LIOB33_X0Y115_IOB_X0Y116_I;
  assign CLBLL_L_X4Y112_SLICE_X5Y112_C1 = CLBLL_L_X4Y112_SLICE_X5Y112_AO6;
  assign CLBLL_L_X4Y112_SLICE_X5Y112_C2 = CLBLL_L_X4Y113_SLICE_X5Y113_AO6;
  assign CLBLL_L_X4Y112_SLICE_X5Y112_C3 = CLBLL_L_X4Y111_SLICE_X5Y111_DO6;
  assign CLBLL_L_X4Y112_SLICE_X5Y112_C4 = CLBLM_R_X5Y112_SLICE_X6Y112_BO6;
  assign CLBLL_L_X4Y112_SLICE_X5Y112_C5 = CLBLL_L_X4Y113_SLICE_X5Y113_BO6;
  assign CLBLL_L_X4Y112_SLICE_X5Y112_C6 = CLBLL_L_X4Y111_SLICE_X5Y111_AO6;
  assign CLBLM_R_X11Y110_SLICE_X15Y110_A1 = 1'b1;
  assign CLBLM_R_X11Y110_SLICE_X15Y110_A2 = 1'b1;
  assign CLBLM_R_X11Y110_SLICE_X15Y110_A3 = RIOB33_X105Y101_IOB_X1Y102_I;
  assign CLBLM_R_X11Y110_SLICE_X15Y110_A4 = LIOB33_X0Y107_IOB_X0Y108_I;
  assign CLBLM_R_X11Y110_SLICE_X15Y110_A5 = RIOB33_X105Y103_IOB_X1Y104_I;
  assign CLBLM_R_X11Y110_SLICE_X15Y110_A6 = 1'b1;
  assign CLBLM_R_X11Y110_SLICE_X15Y110_B1 = CLBLM_R_X11Y111_SLICE_X15Y111_BO5;
  assign CLBLL_L_X4Y112_SLICE_X5Y112_D1 = CLBLL_L_X4Y112_SLICE_X5Y112_AO6;
  assign CLBLL_L_X4Y112_SLICE_X5Y112_D2 = CLBLL_L_X4Y113_SLICE_X5Y113_AO6;
  assign CLBLL_L_X4Y112_SLICE_X5Y112_D3 = 1'b1;
  assign CLBLL_L_X4Y112_SLICE_X5Y112_D4 = 1'b1;
  assign CLBLL_L_X4Y112_SLICE_X5Y112_D5 = 1'b1;
  assign CLBLL_L_X4Y112_SLICE_X5Y112_D6 = CLBLL_L_X4Y111_SLICE_X5Y111_BO6;
  assign CLBLM_R_X11Y110_SLICE_X15Y110_B3 = CLBLM_R_X11Y108_SLICE_X15Y108_AO6;
  assign CLBLM_R_X11Y110_SLICE_X15Y110_B4 = CLBLM_R_X11Y107_SLICE_X15Y107_BO6;
  assign CLBLM_R_X11Y110_SLICE_X15Y110_B6 = CLBLM_L_X12Y109_SLICE_X16Y109_BO6;
  assign CLBLM_R_X11Y110_SLICE_X15Y110_C1 = LIOB33_X0Y107_IOB_X0Y107_I;
  assign CLBLM_R_X11Y110_SLICE_X15Y110_C2 = CLBLM_L_X12Y109_SLICE_X16Y109_AO5;
  assign CLBLM_R_X11Y110_SLICE_X15Y110_C3 = CLBLM_L_X12Y108_SLICE_X16Y108_CO6;
  assign CLBLM_R_X11Y110_SLICE_X15Y110_C4 = RIOB33_X105Y107_IOB_X1Y107_I;
  assign CLBLM_R_X11Y110_SLICE_X15Y110_C5 = CLBLM_L_X12Y108_SLICE_X16Y108_DO6;
  assign CLBLM_R_X11Y110_SLICE_X15Y110_C6 = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLM_R_X11Y110_SLICE_X15Y110_D1 = LIOB33_X0Y107_IOB_X0Y107_I;
  assign CLBLM_R_X11Y110_SLICE_X15Y110_D2 = CLBLM_L_X12Y109_SLICE_X16Y109_AO5;
  assign CLBLM_R_X11Y110_SLICE_X15Y110_D3 = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLM_R_X11Y110_SLICE_X15Y110_D4 = CLBLM_L_X12Y108_SLICE_X16Y108_CO6;
  assign CLBLM_R_X11Y110_SLICE_X15Y110_D5 = CLBLM_L_X12Y108_SLICE_X16Y108_DO6;
  assign CLBLM_R_X11Y110_SLICE_X15Y110_D6 = RIOB33_X105Y107_IOB_X1Y107_I;
  assign CLBLM_R_X11Y110_SLICE_X14Y110_A1 = 1'b1;
  assign CLBLM_R_X11Y110_SLICE_X14Y110_A2 = 1'b1;
  assign CLBLM_R_X11Y110_SLICE_X14Y110_A3 = LIOB33_X0Y109_IOB_X0Y109_I;
  assign CLBLM_R_X11Y110_SLICE_X14Y110_A4 = RIOB33_X105Y103_IOB_X1Y103_I;
  assign CLBLM_R_X11Y110_SLICE_X14Y110_A5 = LIOB33_X0Y109_IOB_X0Y110_I;
  assign CLBLM_R_X11Y110_SLICE_X14Y110_A6 = 1'b1;
  assign CLBLM_R_X11Y110_SLICE_X14Y110_B1 = CLBLM_R_X11Y109_SLICE_X14Y109_AO5;
  assign CLBLM_R_X11Y110_SLICE_X14Y110_B2 = CLBLM_R_X11Y110_SLICE_X15Y110_BO6;
  assign CLBLM_R_X11Y110_SLICE_X14Y110_B3 = CLBLM_R_X11Y110_SLICE_X15Y110_AO5;
  assign CLBLM_R_X11Y110_SLICE_X14Y110_B4 = CLBLM_R_X11Y109_SLICE_X15Y109_BO6;
  assign CLBLM_R_X11Y110_SLICE_X14Y110_B5 = CLBLM_R_X11Y110_SLICE_X14Y110_AO6;
  assign CLBLM_R_X11Y110_SLICE_X14Y110_B6 = CLBLM_R_X11Y111_SLICE_X15Y111_CO6;
  assign CLBLM_R_X11Y110_SLICE_X14Y110_C1 = CLBLM_R_X11Y109_SLICE_X15Y109_BO6;
  assign CLBLM_R_X11Y110_SLICE_X14Y110_C2 = CLBLM_R_X11Y111_SLICE_X15Y111_CO6;
  assign CLBLM_R_X11Y110_SLICE_X14Y110_C3 = CLBLM_R_X11Y110_SLICE_X15Y110_BO6;
  assign CLBLM_R_X11Y110_SLICE_X14Y110_C4 = RIOB33_X105Y103_IOB_X1Y104_I;
  assign CLBLM_R_X11Y110_SLICE_X14Y110_C5 = LIOB33_X0Y107_IOB_X0Y108_I;
  assign CLBLM_R_X11Y110_SLICE_X14Y110_C6 = RIOB33_X105Y103_IOB_X1Y103_I;
  assign CLBLM_R_X11Y110_SLICE_X14Y110_D1 = CLBLM_R_X11Y110_SLICE_X14Y110_AO6;
  assign CLBLM_R_X11Y110_SLICE_X14Y110_D2 = CLBLM_R_X11Y110_SLICE_X15Y110_AO5;
  assign CLBLM_R_X11Y110_SLICE_X14Y110_D3 = CLBLM_R_X11Y110_SLICE_X15Y110_BO6;
  assign CLBLM_R_X11Y110_SLICE_X14Y110_D4 = CLBLM_R_X11Y111_SLICE_X15Y111_CO6;
  assign CLBLM_R_X11Y110_SLICE_X14Y110_D5 = CLBLM_R_X11Y109_SLICE_X14Y109_AO5;
  assign CLBLM_R_X11Y110_SLICE_X14Y110_D6 = CLBLM_R_X11Y109_SLICE_X15Y109_BO6;
  assign CLBLM_L_X8Y107_SLICE_X11Y107_A1 = RIOB33_X105Y101_IOB_X1Y101_I;
  assign CLBLM_L_X8Y107_SLICE_X11Y107_A2 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLM_L_X8Y107_SLICE_X11Y107_A3 = 1'b1;
  assign CLBLM_L_X8Y107_SLICE_X11Y107_A4 = LIOB33_X0Y107_IOB_X0Y108_I;
  assign CLBLM_L_X8Y107_SLICE_X11Y107_A5 = 1'b1;
  assign CLBLM_L_X8Y107_SLICE_X11Y107_A6 = 1'b1;
  assign CLBLM_L_X8Y107_SLICE_X11Y107_B1 = LIOB33_X0Y115_IOB_X0Y116_I;
  assign CLBLM_L_X8Y107_SLICE_X11Y107_B2 = LIOB33_X0Y109_IOB_X0Y109_I;
  assign CLBLM_L_X8Y107_SLICE_X11Y107_B3 = 1'b1;
  assign CLBLM_L_X8Y107_SLICE_X11Y107_B4 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLM_L_X8Y107_SLICE_X11Y107_B5 = 1'b1;
  assign CLBLM_L_X8Y107_SLICE_X11Y107_B6 = 1'b1;
  assign CLBLM_L_X8Y107_SLICE_X11Y107_C1 = CLBLM_L_X10Y106_SLICE_X12Y106_AO6;
  assign CLBLM_L_X8Y107_SLICE_X11Y107_C2 = CLBLM_L_X10Y107_SLICE_X12Y107_AO6;
  assign CLBLM_L_X8Y107_SLICE_X11Y107_C3 = CLBLM_L_X8Y106_SLICE_X10Y106_CO6;
  assign CLBLM_L_X8Y107_SLICE_X11Y107_C4 = CLBLM_L_X8Y107_SLICE_X11Y107_AO5;
  assign CLBLM_L_X8Y107_SLICE_X11Y107_C5 = CLBLM_L_X8Y107_SLICE_X11Y107_AO6;
  assign CLBLM_L_X8Y107_SLICE_X11Y107_C6 = CLBLM_L_X8Y107_SLICE_X11Y107_BO6;
  assign CLBLL_L_X4Y113_SLICE_X4Y113_A1 = RIOB33_X105Y107_IOB_X1Y108_I;
  assign CLBLL_L_X4Y113_SLICE_X4Y113_A2 = CLBLM_R_X5Y113_SLICE_X7Y113_BO6;
  assign CLBLL_L_X4Y113_SLICE_X4Y113_A3 = LIOB33_X0Y115_IOB_X0Y115_I;
  assign CLBLL_L_X4Y113_SLICE_X4Y113_A4 = CLBLM_R_X5Y110_SLICE_X6Y110_CO6;
  assign CLBLL_L_X4Y113_SLICE_X4Y113_A5 = CLBLM_R_X5Y112_SLICE_X6Y112_DO6;
  assign CLBLL_L_X4Y113_SLICE_X4Y113_A6 = 1'b1;
  assign CLBLM_L_X8Y107_SLICE_X11Y107_D1 = CLBLM_L_X8Y106_SLICE_X10Y106_CO6;
  assign CLBLM_L_X8Y107_SLICE_X11Y107_D4 = CLBLM_L_X8Y107_SLICE_X11Y107_AO5;
  assign CLBLL_L_X4Y113_SLICE_X4Y113_B1 = CLBLM_R_X7Y113_SLICE_X8Y113_DO6;
  assign CLBLL_L_X4Y113_SLICE_X4Y113_B2 = CLBLM_R_X5Y113_SLICE_X7Y113_BO6;
  assign CLBLL_L_X4Y113_SLICE_X4Y113_B3 = CLBLL_L_X4Y113_SLICE_X4Y113_DO6;
  assign CLBLL_L_X4Y113_SLICE_X4Y113_B4 = CLBLM_R_X5Y110_SLICE_X6Y110_CO6;
  assign CLBLL_L_X4Y113_SLICE_X4Y113_B5 = CLBLM_R_X5Y112_SLICE_X6Y112_DO6;
  assign CLBLL_L_X4Y113_SLICE_X4Y113_B6 = CLBLL_L_X4Y113_SLICE_X4Y113_CO6;
  assign CLBLM_L_X8Y107_SLICE_X11Y107_D5 = CLBLM_L_X8Y107_SLICE_X11Y107_AO6;
  assign CLBLM_L_X8Y107_SLICE_X10Y107_A1 = CLBLM_L_X8Y106_SLICE_X10Y106_CO6;
  assign CLBLM_L_X8Y107_SLICE_X10Y107_A2 = CLBLM_L_X10Y106_SLICE_X12Y106_AO6;
  assign CLBLL_L_X4Y113_SLICE_X4Y113_C1 = CLBLL_L_X4Y112_SLICE_X5Y112_CO6;
  assign CLBLL_L_X4Y113_SLICE_X4Y113_C2 = CLBLL_L_X4Y113_SLICE_X5Y113_CO6;
  assign CLBLL_L_X4Y113_SLICE_X4Y113_C3 = CLBLM_R_X7Y114_SLICE_X8Y114_CO6;
  assign CLBLL_L_X4Y113_SLICE_X4Y113_C4 = CLBLM_R_X7Y114_SLICE_X8Y114_DO6;
  assign CLBLL_L_X4Y113_SLICE_X4Y113_C5 = CLBLL_L_X4Y114_SLICE_X4Y114_BO6;
  assign CLBLL_L_X4Y113_SLICE_X4Y113_C6 = CLBLM_R_X7Y113_SLICE_X8Y113_CO6;
  assign CLBLM_L_X8Y107_SLICE_X10Y107_A3 = CLBLM_L_X8Y107_SLICE_X11Y107_AO6;
  assign CLBLM_L_X8Y107_SLICE_X10Y107_A4 = CLBLM_R_X7Y106_SLICE_X8Y106_AO6;
  assign CLBLM_L_X8Y107_SLICE_X10Y107_A5 = CLBLM_L_X8Y105_SLICE_X10Y105_BO6;
  assign CLBLM_L_X8Y107_SLICE_X10Y107_A6 = CLBLM_L_X8Y106_SLICE_X10Y106_BO6;
  assign CLBLM_L_X8Y107_SLICE_X10Y107_B1 = CLBLM_R_X7Y106_SLICE_X9Y106_DO6;
  assign CLBLM_L_X8Y107_SLICE_X10Y107_B2 = CLBLM_L_X8Y106_SLICE_X11Y106_DO6;
  assign CLBLM_L_X8Y107_SLICE_X10Y107_B3 = CLBLM_L_X8Y107_SLICE_X11Y107_CO6;
  assign CLBLL_L_X4Y113_SLICE_X4Y113_D1 = LIOB33_X0Y115_IOB_X0Y115_I;
  assign CLBLL_L_X4Y113_SLICE_X4Y113_D2 = 1'b1;
  assign CLBLL_L_X4Y113_SLICE_X4Y113_D3 = 1'b1;
  assign CLBLL_L_X4Y113_SLICE_X4Y113_D4 = 1'b1;
  assign CLBLL_L_X4Y113_SLICE_X4Y113_D5 = 1'b1;
  assign CLBLL_L_X4Y113_SLICE_X4Y113_D6 = RIOB33_X105Y107_IOB_X1Y108_I;
  assign CLBLM_L_X8Y107_SLICE_X10Y107_B5 = CLBLM_L_X8Y106_SLICE_X11Y106_BO6;
  assign CLBLM_L_X8Y107_SLICE_X10Y107_B6 = CLBLM_L_X8Y108_SLICE_X10Y108_AO5;
  assign CLBLM_L_X8Y107_SLICE_X10Y107_C1 = CLBLM_L_X8Y106_SLICE_X10Y106_CO6;
  assign CLBLM_L_X8Y107_SLICE_X10Y107_C2 = RIOB33_X105Y101_IOB_X1Y101_I;
  assign CLBLM_L_X8Y107_SLICE_X10Y107_C3 = CLBLM_L_X10Y106_SLICE_X12Y106_AO6;
  assign CLBLM_L_X8Y107_SLICE_X10Y107_C4 = CLBLM_L_X10Y107_SLICE_X12Y107_AO6;
  assign CLBLM_L_X8Y107_SLICE_X10Y107_C5 = LIOB33_X0Y107_IOB_X0Y108_I;
  assign CLBLM_L_X8Y107_SLICE_X10Y107_C6 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLM_L_X8Y107_SLICE_X10Y107_D1 = CLBLM_L_X8Y105_SLICE_X10Y105_BO6;
  assign CLBLM_L_X8Y107_SLICE_X10Y107_D2 = CLBLM_L_X8Y107_SLICE_X11Y107_AO6;
  assign CLBLM_L_X8Y107_SLICE_X10Y107_D3 = CLBLM_L_X10Y106_SLICE_X12Y106_AO6;
  assign CLBLM_L_X8Y107_SLICE_X10Y107_D4 = CLBLM_L_X8Y106_SLICE_X10Y106_BO6;
  assign CLBLM_L_X8Y107_SLICE_X10Y107_D5 = CLBLM_L_X8Y106_SLICE_X10Y106_CO6;
  assign CLBLM_L_X8Y107_SLICE_X10Y107_D6 = CLBLM_R_X7Y106_SLICE_X8Y106_AO6;
  assign CLBLL_L_X4Y113_SLICE_X5Y113_A1 = 1'b1;
  assign CLBLL_L_X4Y113_SLICE_X5Y113_A2 = CLBLM_R_X5Y111_SLICE_X6Y111_BO6;
  assign CLBLL_L_X4Y113_SLICE_X5Y113_A3 = RIOB33_X105Y103_IOB_X1Y103_I;
  assign CLBLL_L_X4Y113_SLICE_X5Y113_A4 = CLBLM_R_X5Y113_SLICE_X7Y113_AO6;
  assign CLBLL_L_X4Y113_SLICE_X5Y113_A5 = LIOB33_X0Y115_IOB_X0Y115_I;
  assign CLBLL_L_X4Y113_SLICE_X5Y113_A6 = 1'b1;
  assign CLBLL_L_X4Y113_SLICE_X5Y113_B1 = RIOB33_X105Y103_IOB_X1Y104_I;
  assign CLBLL_L_X4Y113_SLICE_X5Y113_B2 = CLBLM_R_X7Y114_SLICE_X8Y114_BO6;
  assign CLBLL_L_X4Y113_SLICE_X5Y113_B3 = RIOB33_X105Y103_IOB_X1Y103_I;
  assign CLBLL_L_X4Y113_SLICE_X5Y113_B4 = CLBLM_R_X5Y113_SLICE_X7Y113_AO6;
  assign CLBLL_L_X4Y113_SLICE_X5Y113_B5 = LIOB33_X0Y115_IOB_X0Y115_I;
  assign CLBLL_L_X4Y113_SLICE_X5Y113_B6 = CLBLM_R_X5Y111_SLICE_X6Y111_BO6;
  assign CLBLL_L_X4Y113_SLICE_X5Y113_C1 = LIOB33_X0Y115_IOB_X0Y115_I;
  assign CLBLL_L_X4Y113_SLICE_X5Y113_C2 = CLBLM_R_X7Y114_SLICE_X8Y114_BO6;
  assign CLBLL_L_X4Y113_SLICE_X5Y113_C3 = RIOB33_X105Y103_IOB_X1Y104_I;
  assign CLBLL_L_X4Y113_SLICE_X5Y113_C4 = CLBLM_R_X5Y111_SLICE_X6Y111_BO6;
  assign CLBLL_L_X4Y113_SLICE_X5Y113_C5 = RIOB33_X105Y103_IOB_X1Y103_I;
  assign CLBLL_L_X4Y113_SLICE_X5Y113_C6 = CLBLM_R_X5Y113_SLICE_X7Y113_AO6;
  assign CLBLM_R_X11Y111_SLICE_X15Y111_A1 = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLM_R_X11Y111_SLICE_X15Y111_A2 = RIOB33_X105Y103_IOB_X1Y104_I;
  assign CLBLM_R_X11Y111_SLICE_X15Y111_A3 = 1'b1;
  assign CLBLM_R_X11Y111_SLICE_X15Y111_A4 = 1'b1;
  assign CLBLM_R_X11Y111_SLICE_X15Y111_A5 = LIOB33_X0Y107_IOB_X0Y107_I;
  assign CLBLM_R_X11Y111_SLICE_X15Y111_A6 = 1'b1;
  assign CLBLL_L_X4Y113_SLICE_X5Y113_D1 = 1'b1;
  assign CLBLL_L_X4Y113_SLICE_X5Y113_D2 = 1'b1;
  assign CLBLL_L_X4Y113_SLICE_X5Y113_D3 = 1'b1;
  assign CLBLL_L_X4Y113_SLICE_X5Y113_D4 = 1'b1;
  assign CLBLL_L_X4Y113_SLICE_X5Y113_D5 = 1'b1;
  assign CLBLL_L_X4Y113_SLICE_X5Y113_D6 = 1'b1;
  assign CLBLM_R_X11Y111_SLICE_X15Y111_B1 = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLM_R_X11Y111_SLICE_X15Y111_B2 = 1'b1;
  assign CLBLM_R_X11Y111_SLICE_X15Y111_B3 = LIOB33_X0Y107_IOB_X0Y107_I;
  assign CLBLM_R_X11Y111_SLICE_X15Y111_B4 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X11Y111_SLICE_X15Y111_B5 = 1'b1;
  assign CLBLM_R_X11Y111_SLICE_X15Y111_B6 = 1'b1;
  assign CLBLM_R_X11Y111_SLICE_X15Y111_C1 = CLBLM_R_X11Y108_SLICE_X15Y108_AO6;
  assign CLBLM_R_X11Y111_SLICE_X15Y111_C2 = RIOB33_X105Y103_IOB_X1Y104_I;
  assign CLBLM_R_X11Y111_SLICE_X15Y111_C3 = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLM_R_X11Y111_SLICE_X15Y111_C4 = CLBLM_L_X12Y108_SLICE_X17Y108_AO6;
  assign CLBLM_R_X11Y111_SLICE_X15Y111_C5 = LIOB33_X0Y107_IOB_X0Y107_I;
  assign CLBLM_R_X11Y111_SLICE_X15Y111_C6 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X11Y111_SLICE_X15Y111_D1 = CLBLM_R_X11Y108_SLICE_X15Y108_AO6;
  assign CLBLM_R_X11Y111_SLICE_X15Y111_D2 = CLBLM_L_X12Y108_SLICE_X17Y108_AO6;
  assign CLBLM_R_X11Y111_SLICE_X15Y111_D3 = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLM_R_X11Y111_SLICE_X15Y111_D4 = RIOB33_X105Y103_IOB_X1Y104_I;
  assign CLBLM_R_X11Y111_SLICE_X15Y111_D5 = LIOB33_X0Y107_IOB_X0Y107_I;
  assign CLBLM_R_X11Y111_SLICE_X15Y111_D6 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X11Y111_SLICE_X14Y111_A1 = CLBLM_R_X11Y111_SLICE_X14Y111_DO6;
  assign CLBLM_R_X11Y111_SLICE_X14Y111_A2 = CLBLM_R_X11Y111_SLICE_X14Y111_BO5;
  assign CLBLM_R_X11Y111_SLICE_X14Y111_A3 = LIOB33_X0Y109_IOB_X0Y109_I;
  assign CLBLM_R_X11Y111_SLICE_X14Y111_A4 = RIOB33_X105Y103_IOB_X1Y104_I;
  assign CLBLM_R_X11Y111_SLICE_X14Y111_A5 = 1'b1;
  assign CLBLM_R_X11Y111_SLICE_X14Y111_A6 = 1'b1;
  assign CLBLM_R_X11Y111_SLICE_X14Y111_B1 = CLBLM_R_X11Y109_SLICE_X15Y109_DO6;
  assign CLBLM_R_X11Y111_SLICE_X14Y111_B2 = LIOB33_X0Y107_IOB_X0Y108_I;
  assign CLBLM_R_X11Y111_SLICE_X14Y111_B3 = 1'b1;
  assign CLBLM_R_X11Y111_SLICE_X14Y111_B4 = CLBLM_R_X11Y110_SLICE_X15Y110_DO6;
  assign CLBLM_R_X11Y111_SLICE_X14Y111_B5 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X11Y111_SLICE_X14Y111_B6 = 1'b1;
  assign CLBLM_R_X11Y111_SLICE_X14Y111_C1 = LIOB33_X0Y107_IOB_X0Y108_I;
  assign CLBLM_R_X11Y111_SLICE_X14Y111_C2 = CLBLM_L_X12Y109_SLICE_X16Y109_CO6;
  assign CLBLM_R_X11Y111_SLICE_X14Y111_C3 = CLBLM_R_X11Y111_SLICE_X15Y111_DO6;
  assign CLBLM_R_X11Y111_SLICE_X14Y111_C4 = RIOB33_X105Y103_IOB_X1Y104_I;
  assign CLBLM_R_X11Y111_SLICE_X14Y111_C5 = LIOB33_X0Y107_IOB_X0Y107_I;
  assign CLBLM_R_X11Y111_SLICE_X14Y111_C6 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X11Y111_SLICE_X14Y111_D1 = LIOB33_X0Y107_IOB_X0Y108_I;
  assign CLBLM_R_X11Y111_SLICE_X14Y111_D2 = CLBLM_L_X12Y109_SLICE_X16Y109_CO6;
  assign CLBLM_R_X11Y111_SLICE_X14Y111_D3 = CLBLM_R_X11Y111_SLICE_X15Y111_DO6;
  assign CLBLM_R_X11Y111_SLICE_X14Y111_D4 = RIOB33_X105Y103_IOB_X1Y104_I;
  assign CLBLM_R_X11Y111_SLICE_X14Y111_D5 = LIOB33_X0Y107_IOB_X0Y107_I;
  assign CLBLM_R_X11Y111_SLICE_X14Y111_D6 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X11Y110_SLICE_X15Y110_B2 = CLBLM_R_X11Y111_SLICE_X15Y111_AO6;
  assign CLBLM_R_X11Y110_SLICE_X15Y110_B5 = CLBLM_R_X11Y107_SLICE_X15Y107_CO6;
  assign CLBLM_L_X8Y108_SLICE_X11Y108_A1 = CLBLM_L_X8Y108_SLICE_X11Y108_DO6;
  assign CLBLM_L_X8Y108_SLICE_X11Y108_A2 = LIOB33_X0Y109_IOB_X0Y110_I;
  assign CLBLM_L_X8Y108_SLICE_X11Y108_A3 = LIOB33_X0Y109_IOB_X0Y109_I;
  assign CLBLM_L_X8Y108_SLICE_X11Y108_A4 = CLBLM_L_X10Y109_SLICE_X12Y109_BO6;
  assign CLBLM_L_X8Y108_SLICE_X11Y108_A5 = CLBLM_L_X10Y108_SLICE_X12Y108_AO6;
  assign CLBLM_L_X8Y108_SLICE_X11Y108_A6 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLM_L_X8Y108_SLICE_X11Y108_B1 = CLBLM_L_X8Y108_SLICE_X11Y108_DO6;
  assign CLBLM_L_X8Y108_SLICE_X11Y108_B2 = LIOB33_X0Y109_IOB_X0Y110_I;
  assign CLBLM_L_X8Y108_SLICE_X11Y108_B3 = LIOB33_X0Y109_IOB_X0Y109_I;
  assign CLBLM_L_X8Y108_SLICE_X11Y108_B4 = CLBLM_L_X10Y108_SLICE_X12Y108_AO6;
  assign CLBLM_L_X8Y108_SLICE_X11Y108_B5 = CLBLM_L_X10Y109_SLICE_X12Y109_BO6;
  assign CLBLM_L_X8Y108_SLICE_X11Y108_B6 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLM_L_X8Y108_SLICE_X11Y108_C1 = LIOB33_X0Y109_IOB_X0Y109_I;
  assign CLBLM_L_X8Y108_SLICE_X11Y108_C2 = CLBLM_L_X10Y108_SLICE_X12Y108_BO6;
  assign CLBLM_L_X8Y108_SLICE_X11Y108_C3 = CLBLM_L_X10Y109_SLICE_X12Y109_BO6;
  assign CLBLM_L_X8Y108_SLICE_X11Y108_C4 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLM_L_X8Y108_SLICE_X11Y108_C5 = CLBLM_L_X8Y108_SLICE_X11Y108_DO6;
  assign CLBLM_L_X8Y108_SLICE_X11Y108_C6 = RIOB33_X105Y101_IOB_X1Y101_I;
  assign CLBLL_L_X4Y114_SLICE_X4Y114_A1 = 1'b1;
  assign CLBLL_L_X4Y114_SLICE_X4Y114_A2 = LIOB33_X0Y115_IOB_X0Y116_I;
  assign CLBLL_L_X4Y114_SLICE_X4Y114_A3 = LIOB33_X0Y115_IOB_X0Y115_I;
  assign CLBLL_L_X4Y114_SLICE_X4Y114_A4 = 1'b1;
  assign CLBLL_L_X4Y114_SLICE_X4Y114_A5 = RIOB33_X105Y103_IOB_X1Y104_I;
  assign CLBLL_L_X4Y114_SLICE_X4Y114_A6 = 1'b1;
  assign CLBLM_L_X8Y108_SLICE_X11Y108_D1 = CLBLM_L_X10Y106_SLICE_X12Y106_BO6;
  assign CLBLL_L_X4Y114_SLICE_X4Y114_B1 = CLBLM_R_X7Y114_SLICE_X8Y114_AO5;
  assign CLBLL_L_X4Y114_SLICE_X4Y114_B2 = CLBLM_R_X7Y114_SLICE_X8Y114_BO6;
  assign CLBLM_L_X8Y108_SLICE_X11Y108_D4 = LIOB33_X0Y107_IOB_X0Y107_I;
  assign CLBLL_L_X4Y114_SLICE_X4Y114_B3 = LIOB33_X0Y115_IOB_X0Y115_I;
  assign CLBLM_L_X8Y108_SLICE_X11Y108_D5 = CLBLM_L_X8Y106_SLICE_X10Y106_CO6;
  assign CLBLM_L_X8Y108_SLICE_X11Y108_D6 = RIOB33_X105Y101_IOB_X1Y101_I;
  assign CLBLL_L_X4Y114_SLICE_X4Y114_B4 = CLBLM_R_X5Y113_SLICE_X7Y113_AO5;
  assign CLBLL_L_X4Y114_SLICE_X4Y114_B5 = RIOB33_X105Y103_IOB_X1Y104_I;
  assign CLBLL_L_X4Y114_SLICE_X4Y114_B6 = 1'b1;
  assign CLBLM_L_X8Y108_SLICE_X11Y108_D3 = LIOB33_X0Y107_IOB_X0Y108_I;
  assign CLBLL_L_X4Y114_SLICE_X4Y114_C1 = CLBLM_R_X7Y114_SLICE_X8Y114_CO6;
  assign CLBLL_L_X4Y114_SLICE_X4Y114_C2 = CLBLL_L_X4Y113_SLICE_X5Y113_AO5;
  assign CLBLL_L_X4Y114_SLICE_X4Y114_C3 = CLBLM_R_X7Y114_SLICE_X8Y114_AO5;
  assign CLBLL_L_X4Y114_SLICE_X4Y114_C4 = CLBLL_L_X4Y114_SLICE_X4Y114_AO5;
  assign CLBLL_L_X4Y114_SLICE_X4Y114_C5 = CLBLL_L_X4Y112_SLICE_X5Y112_BO6;
  assign CLBLL_L_X4Y114_SLICE_X4Y114_C6 = CLBLM_R_X5Y113_SLICE_X7Y113_AO5;
  assign CLBLM_L_X8Y108_SLICE_X10Y108_A1 = LIOB33_X0Y115_IOB_X0Y116_I;
  assign CLBLM_L_X8Y108_SLICE_X10Y108_A2 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLM_L_X8Y108_SLICE_X10Y108_A3 = 1'b1;
  assign CLBLM_L_X8Y108_SLICE_X10Y108_A4 = LIOB33_X0Y109_IOB_X0Y110_I;
  assign CLBLM_L_X8Y108_SLICE_X10Y108_A5 = 1'b1;
  assign CLBLM_L_X8Y108_SLICE_X10Y108_A6 = 1'b1;
  assign CLBLM_L_X8Y108_SLICE_X10Y108_B2 = LIOB33_X0Y107_IOB_X0Y107_I;
  assign CLBLM_L_X8Y108_SLICE_X10Y108_B3 = CLBLM_L_X10Y106_SLICE_X12Y106_BO6;
  assign CLBLM_L_X8Y108_SLICE_X10Y108_B4 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLM_L_X8Y108_SLICE_X10Y108_B5 = CLBLM_L_X8Y106_SLICE_X10Y106_CO6;
  assign CLBLM_L_X8Y108_SLICE_X10Y108_B6 = RIOB33_X105Y101_IOB_X1Y101_I;
  assign CLBLM_L_X8Y108_SLICE_X10Y108_B1 = LIOB33_X0Y107_IOB_X0Y108_I;
  assign CLBLL_L_X4Y114_SLICE_X4Y114_D1 = CLBLL_L_X4Y113_SLICE_X5Y113_BO6;
  assign CLBLL_L_X4Y114_SLICE_X4Y114_D2 = 1'b1;
  assign CLBLL_L_X4Y114_SLICE_X4Y114_D3 = 1'b1;
  assign CLBLL_L_X4Y114_SLICE_X4Y114_D4 = 1'b1;
  assign CLBLL_L_X4Y114_SLICE_X4Y114_D5 = 1'b1;
  assign CLBLL_L_X4Y114_SLICE_X4Y114_D6 = CLBLL_L_X4Y112_SLICE_X5Y112_BO6;
  assign CLBLM_L_X8Y108_SLICE_X10Y108_C1 = CLBLM_L_X8Y108_SLICE_X10Y108_AO6;
  assign CLBLM_L_X8Y108_SLICE_X10Y108_C2 = CLBLM_L_X8Y107_SLICE_X11Y107_CO6;
  assign CLBLM_L_X8Y108_SLICE_X10Y108_C3 = CLBLM_L_X10Y108_SLICE_X12Y108_AO6;
  assign CLBLM_L_X8Y108_SLICE_X10Y108_C4 = CLBLM_L_X8Y108_SLICE_X10Y108_AO5;
  assign CLBLM_L_X8Y108_SLICE_X10Y108_C5 = CLBLM_L_X8Y106_SLICE_X11Y106_DO6;
  assign CLBLM_L_X8Y108_SLICE_X10Y108_C6 = CLBLM_L_X8Y107_SLICE_X11Y107_DO6;
  assign CLBLM_L_X8Y108_SLICE_X10Y108_D1 = CLBLM_L_X8Y108_SLICE_X10Y108_AO6;
  assign CLBLM_L_X8Y108_SLICE_X10Y108_D2 = CLBLM_R_X11Y109_SLICE_X14Y109_BO6;
  assign CLBLM_L_X8Y108_SLICE_X10Y108_D3 = CLBLM_L_X10Y110_SLICE_X13Y110_AO6;
  assign CLBLM_L_X8Y108_SLICE_X10Y108_D4 = CLBLM_L_X10Y108_SLICE_X12Y108_AO6;
  assign CLBLM_L_X8Y108_SLICE_X10Y108_D5 = CLBLM_L_X10Y108_SLICE_X12Y108_DO6;
  assign CLBLM_L_X8Y108_SLICE_X10Y108_D6 = CLBLM_L_X8Y107_SLICE_X11Y107_DO6;
  assign CLBLL_L_X4Y114_SLICE_X5Y114_A1 = 1'b1;
  assign CLBLL_L_X4Y114_SLICE_X5Y114_A2 = 1'b1;
  assign CLBLL_L_X4Y114_SLICE_X5Y114_A3 = 1'b1;
  assign CLBLL_L_X4Y114_SLICE_X5Y114_A4 = 1'b1;
  assign CLBLL_L_X4Y114_SLICE_X5Y114_A5 = 1'b1;
  assign CLBLL_L_X4Y114_SLICE_X5Y114_A6 = 1'b1;
  assign LIOI3_X0Y111_ILOGIC_X0Y112_D = LIOB33_X0Y111_IOB_X0Y112_I;
  assign LIOI3_X0Y111_ILOGIC_X0Y111_D = LIOB33_X0Y111_IOB_X0Y111_I;
  assign CLBLL_L_X4Y114_SLICE_X5Y114_B1 = 1'b1;
  assign CLBLL_L_X4Y114_SLICE_X5Y114_B2 = 1'b1;
  assign CLBLL_L_X4Y114_SLICE_X5Y114_B3 = 1'b1;
  assign CLBLL_L_X4Y114_SLICE_X5Y114_B4 = 1'b1;
  assign CLBLL_L_X4Y114_SLICE_X5Y114_B5 = 1'b1;
  assign CLBLL_L_X4Y114_SLICE_X5Y114_B6 = 1'b1;
  assign CLBLL_L_X4Y114_SLICE_X5Y114_C1 = 1'b1;
  assign CLBLL_L_X4Y114_SLICE_X5Y114_C2 = 1'b1;
  assign CLBLL_L_X4Y114_SLICE_X5Y114_C3 = 1'b1;
  assign CLBLL_L_X4Y114_SLICE_X5Y114_C4 = 1'b1;
  assign CLBLL_L_X4Y114_SLICE_X5Y114_C5 = 1'b1;
  assign CLBLL_L_X4Y114_SLICE_X5Y114_C6 = 1'b1;
  assign CLBLL_L_X4Y114_SLICE_X5Y114_D1 = 1'b1;
  assign CLBLL_L_X4Y114_SLICE_X5Y114_D2 = 1'b1;
  assign CLBLL_L_X4Y114_SLICE_X5Y114_D3 = 1'b1;
  assign CLBLL_L_X4Y114_SLICE_X5Y114_D4 = 1'b1;
  assign CLBLL_L_X4Y114_SLICE_X5Y114_D5 = 1'b1;
  assign CLBLL_L_X4Y114_SLICE_X5Y114_D6 = 1'b1;
  assign CLBLM_R_X7Y112_SLICE_X9Y112_B3 = CLBLM_L_X8Y110_SLICE_X10Y110_BO6;
  assign CLBLM_R_X7Y112_SLICE_X9Y112_B4 = CLBLM_L_X8Y111_SLICE_X10Y111_BO6;
  assign CLBLM_L_X8Y109_SLICE_X11Y109_A1 = 1'b1;
  assign CLBLM_L_X8Y109_SLICE_X11Y109_A2 = 1'b1;
  assign CLBLM_L_X8Y109_SLICE_X11Y109_A3 = 1'b1;
  assign CLBLM_L_X8Y109_SLICE_X11Y109_A4 = 1'b1;
  assign CLBLM_L_X8Y109_SLICE_X11Y109_A5 = 1'b1;
  assign CLBLM_L_X8Y109_SLICE_X11Y109_A6 = 1'b1;
  assign CLBLM_L_X8Y109_SLICE_X11Y109_B1 = 1'b1;
  assign CLBLM_L_X8Y109_SLICE_X11Y109_B2 = 1'b1;
  assign CLBLM_L_X8Y109_SLICE_X11Y109_B3 = 1'b1;
  assign CLBLM_L_X8Y109_SLICE_X11Y109_B4 = 1'b1;
  assign CLBLM_L_X8Y109_SLICE_X11Y109_B5 = 1'b1;
  assign CLBLM_L_X8Y109_SLICE_X11Y109_B6 = 1'b1;
  assign CLBLM_L_X8Y109_SLICE_X11Y109_C1 = 1'b1;
  assign CLBLL_L_X4Y115_SLICE_X4Y115_A1 = CLBLM_R_X7Y113_SLICE_X8Y113_DO6;
  assign CLBLL_L_X4Y115_SLICE_X4Y115_A2 = CLBLM_R_X7Y114_SLICE_X8Y114_DO6;
  assign CLBLL_L_X4Y115_SLICE_X4Y115_A3 = CLBLL_L_X4Y113_SLICE_X4Y113_AO6;
  assign CLBLM_L_X8Y109_SLICE_X11Y109_C5 = 1'b1;
  assign CLBLM_L_X8Y109_SLICE_X11Y109_C6 = 1'b1;
  assign CLBLL_L_X4Y115_SLICE_X4Y115_A4 = CLBLL_L_X4Y115_SLICE_X4Y115_BO6;
  assign CLBLL_L_X4Y115_SLICE_X4Y115_A5 = CLBLM_R_X7Y113_SLICE_X8Y113_CO6;
  assign CLBLL_L_X4Y115_SLICE_X4Y115_A6 = 1'b1;
  assign CLBLM_L_X8Y109_SLICE_X11Y109_C2 = 1'b1;
  assign CLBLM_L_X8Y109_SLICE_X11Y109_C3 = 1'b1;
  assign CLBLM_L_X8Y109_SLICE_X11Y109_C4 = 1'b1;
  assign CLBLL_L_X4Y115_SLICE_X4Y115_B1 = CLBLL_L_X4Y112_SLICE_X5Y112_BO6;
  assign CLBLL_L_X4Y115_SLICE_X4Y115_B2 = CLBLL_L_X4Y114_SLICE_X4Y114_BO6;
  assign CLBLL_L_X4Y115_SLICE_X4Y115_B3 = CLBLM_R_X7Y114_SLICE_X8Y114_CO6;
  assign CLBLL_L_X4Y115_SLICE_X4Y115_B4 = CLBLL_L_X4Y114_SLICE_X4Y114_BO5;
  assign CLBLM_L_X8Y109_SLICE_X11Y109_D3 = 1'b1;
  assign CLBLL_L_X4Y115_SLICE_X4Y115_B5 = CLBLL_L_X4Y115_SLICE_X4Y115_AO6;
  assign CLBLM_L_X8Y109_SLICE_X11Y109_D5 = 1'b1;
  assign CLBLM_L_X8Y109_SLICE_X11Y109_D6 = 1'b1;
  assign CLBLL_L_X4Y115_SLICE_X4Y115_B6 = CLBLL_L_X4Y113_SLICE_X5Y113_AO5;
  assign CLBLM_L_X8Y109_SLICE_X11Y109_D1 = 1'b1;
  assign CLBLL_L_X4Y115_SLICE_X4Y115_C1 = CLBLL_L_X4Y113_SLICE_X4Y113_AO6;
  assign CLBLL_L_X4Y115_SLICE_X4Y115_C2 = CLBLM_R_X7Y113_SLICE_X8Y113_CO6;
  assign CLBLL_L_X4Y115_SLICE_X4Y115_C3 = CLBLM_R_X7Y114_SLICE_X8Y114_DO6;
  assign CLBLL_L_X4Y115_SLICE_X4Y115_C4 = CLBLL_L_X4Y113_SLICE_X4Y113_AO5;
  assign CLBLL_L_X4Y115_SLICE_X4Y115_C5 = CLBLM_R_X7Y113_SLICE_X8Y113_DO6;
  assign CLBLL_L_X4Y115_SLICE_X4Y115_C6 = CLBLL_L_X4Y115_SLICE_X4Y115_BO6;
  assign CLBLM_L_X8Y109_SLICE_X10Y109_A1 = CLBLM_L_X8Y109_SLICE_X10Y109_DO6;
  assign CLBLM_L_X8Y109_SLICE_X10Y109_A2 = LIOB33_X0Y107_IOB_X0Y108_I;
  assign CLBLM_L_X8Y109_SLICE_X10Y109_A3 = RIOB33_X105Y109_IOB_X1Y109_I;
  assign CLBLM_L_X8Y109_SLICE_X10Y109_A4 = CLBLM_R_X7Y109_SLICE_X9Y109_AO6;
  assign CLBLM_L_X8Y109_SLICE_X10Y109_A5 = LIOB33_X0Y109_IOB_X0Y109_I;
  assign CLBLM_L_X8Y109_SLICE_X10Y109_A6 = CLBLM_R_X11Y106_SLICE_X15Y106_AO5;
  assign CLBLL_L_X4Y115_SLICE_X4Y115_D1 = CLBLL_L_X4Y112_SLICE_X5Y112_BO6;
  assign CLBLL_L_X4Y115_SLICE_X4Y115_D2 = CLBLM_R_X7Y114_SLICE_X8Y114_CO6;
  assign CLBLL_L_X4Y115_SLICE_X4Y115_D3 = CLBLL_L_X4Y114_SLICE_X4Y114_BO6;
  assign CLBLL_L_X4Y115_SLICE_X4Y115_D4 = CLBLL_L_X4Y113_SLICE_X5Y113_AO5;
  assign CLBLL_L_X4Y115_SLICE_X4Y115_D5 = 1'b1;
  assign CLBLL_L_X4Y115_SLICE_X4Y115_D6 = CLBLL_L_X4Y114_SLICE_X4Y114_BO5;
  assign CLBLM_L_X8Y109_SLICE_X10Y109_B1 = RIOB33_X105Y109_IOB_X1Y110_I;
  assign CLBLM_L_X8Y109_SLICE_X10Y109_B2 = LIOB33_X0Y107_IOB_X0Y108_I;
  assign CLBLM_L_X8Y109_SLICE_X10Y109_B3 = CLBLM_L_X10Y109_SLICE_X12Y109_CO6;
  assign CLBLM_L_X8Y109_SLICE_X10Y109_B4 = RIOB33_X105Y109_IOB_X1Y109_I;
  assign CLBLM_L_X8Y109_SLICE_X10Y109_B5 = LIOB33_X0Y107_IOB_X0Y107_I;
  assign CLBLM_L_X8Y109_SLICE_X10Y109_B6 = CLBLM_R_X11Y106_SLICE_X15Y106_AO5;
  assign CLBLM_L_X8Y109_SLICE_X10Y109_C1 = LIOB33_X0Y109_IOB_X0Y109_I;
  assign CLBLM_L_X8Y109_SLICE_X10Y109_C2 = CLBLM_R_X7Y109_SLICE_X9Y109_AO6;
  assign CLBLM_L_X8Y109_SLICE_X10Y109_C3 = LIOB33_X0Y107_IOB_X0Y108_I;
  assign CLBLM_L_X8Y109_SLICE_X10Y109_C4 = RIOB33_X105Y109_IOB_X1Y109_I;
  assign CLBLM_L_X8Y109_SLICE_X10Y109_C5 = CLBLM_L_X8Y109_SLICE_X10Y109_DO6;
  assign CLBLM_L_X8Y109_SLICE_X10Y109_C6 = CLBLM_R_X11Y106_SLICE_X15Y106_AO5;
  assign CLBLM_L_X8Y109_SLICE_X10Y109_D1 = LIOB33_X0Y107_IOB_X0Y108_I;
  assign CLBLM_L_X8Y109_SLICE_X10Y109_D2 = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLM_L_X8Y109_SLICE_X10Y109_D3 = RIOB33_X105Y109_IOB_X1Y110_I;
  assign CLBLM_L_X8Y109_SLICE_X10Y109_D4 = RIOB33_X105Y111_IOB_X1Y111_I;
  assign CLBLM_L_X8Y109_SLICE_X10Y109_D5 = CLBLM_L_X10Y109_SLICE_X12Y109_DO6;
  assign CLBLL_L_X4Y115_SLICE_X5Y115_A1 = 1'b1;
  assign CLBLL_L_X4Y115_SLICE_X5Y115_A2 = 1'b1;
  assign CLBLL_L_X4Y115_SLICE_X5Y115_A3 = 1'b1;
  assign CLBLL_L_X4Y115_SLICE_X5Y115_A4 = 1'b1;
  assign CLBLL_L_X4Y115_SLICE_X5Y115_A5 = 1'b1;
  assign CLBLL_L_X4Y115_SLICE_X5Y115_A6 = 1'b1;
  assign CLBLM_L_X8Y109_SLICE_X10Y109_D6 = LIOB33_X0Y107_IOB_X0Y107_I;
  assign CLBLL_L_X4Y115_SLICE_X5Y115_B1 = 1'b1;
  assign CLBLL_L_X4Y115_SLICE_X5Y115_B2 = 1'b1;
  assign CLBLL_L_X4Y115_SLICE_X5Y115_B3 = 1'b1;
  assign CLBLL_L_X4Y115_SLICE_X5Y115_B4 = 1'b1;
  assign CLBLL_L_X4Y115_SLICE_X5Y115_B5 = 1'b1;
  assign CLBLL_L_X4Y115_SLICE_X5Y115_B6 = 1'b1;
  assign CLBLL_L_X4Y115_SLICE_X5Y115_C1 = 1'b1;
  assign CLBLL_L_X4Y115_SLICE_X5Y115_C2 = 1'b1;
  assign CLBLL_L_X4Y115_SLICE_X5Y115_C3 = 1'b1;
  assign CLBLL_L_X4Y115_SLICE_X5Y115_C4 = 1'b1;
  assign CLBLL_L_X4Y115_SLICE_X5Y115_C5 = 1'b1;
  assign CLBLL_L_X4Y115_SLICE_X5Y115_C6 = 1'b1;
  assign CLBLL_L_X4Y115_SLICE_X5Y115_D1 = 1'b1;
  assign CLBLL_L_X4Y115_SLICE_X5Y115_D2 = 1'b1;
  assign CLBLL_L_X4Y115_SLICE_X5Y115_D3 = 1'b1;
  assign CLBLL_L_X4Y115_SLICE_X5Y115_D4 = 1'b1;
  assign CLBLL_L_X4Y115_SLICE_X5Y115_D5 = 1'b1;
  assign CLBLL_L_X4Y115_SLICE_X5Y115_D6 = 1'b1;
  assign CLBLM_R_X7Y103_SLICE_X9Y103_A1 = 1'b1;
  assign CLBLM_R_X7Y103_SLICE_X9Y103_A2 = 1'b1;
  assign CLBLM_R_X7Y103_SLICE_X9Y103_A3 = 1'b1;
  assign CLBLM_R_X7Y103_SLICE_X9Y103_A4 = 1'b1;
  assign CLBLM_R_X7Y103_SLICE_X9Y103_A5 = 1'b1;
  assign CLBLM_R_X7Y103_SLICE_X9Y103_A6 = 1'b1;
  assign CLBLM_R_X7Y103_SLICE_X9Y103_B1 = 1'b1;
  assign CLBLM_R_X7Y103_SLICE_X9Y103_B2 = 1'b1;
  assign CLBLM_R_X7Y103_SLICE_X9Y103_B3 = 1'b1;
  assign CLBLM_R_X7Y103_SLICE_X9Y103_B4 = 1'b1;
  assign CLBLM_R_X7Y103_SLICE_X9Y103_B5 = 1'b1;
  assign CLBLM_R_X7Y103_SLICE_X9Y103_B6 = 1'b1;
  assign CLBLM_L_X8Y106_SLICE_X11Y106_D2 = CLBLM_L_X8Y107_SLICE_X11Y107_AO6;
  assign CLBLM_R_X7Y103_SLICE_X9Y103_C1 = 1'b1;
  assign CLBLM_R_X7Y103_SLICE_X9Y103_C2 = 1'b1;
  assign CLBLM_R_X7Y103_SLICE_X9Y103_C3 = 1'b1;
  assign CLBLM_R_X7Y103_SLICE_X9Y103_C4 = 1'b1;
  assign CLBLM_R_X7Y103_SLICE_X9Y103_C5 = 1'b1;
  assign CLBLM_R_X7Y103_SLICE_X9Y103_C6 = 1'b1;
  assign CLBLM_R_X7Y103_SLICE_X9Y103_D1 = 1'b1;
  assign CLBLM_R_X7Y103_SLICE_X9Y103_D2 = 1'b1;
  assign CLBLM_R_X7Y103_SLICE_X9Y103_D3 = 1'b1;
  assign CLBLM_R_X7Y103_SLICE_X9Y103_D4 = 1'b1;
  assign CLBLM_R_X7Y103_SLICE_X9Y103_D5 = 1'b1;
  assign CLBLM_R_X7Y103_SLICE_X9Y103_D6 = 1'b1;
  assign CLBLM_R_X7Y103_SLICE_X8Y103_A1 = RIOB33_X105Y101_IOB_X1Y101_I;
  assign CLBLM_R_X7Y103_SLICE_X8Y103_A2 = RIOB33_X105Y101_IOB_X1Y102_I;
  assign CLBLM_R_X7Y103_SLICE_X8Y103_A3 = RIOB33_X105Y113_IOB_X1Y113_I;
  assign CLBLM_R_X7Y103_SLICE_X8Y103_A4 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLM_R_X7Y103_SLICE_X8Y103_A5 = RIOB33_X105Y111_IOB_X1Y112_I;
  assign CLBLM_R_X7Y103_SLICE_X8Y103_A6 = LIOB33_SING_X0Y100_IOB_X0Y100_I;
  assign CLBLM_R_X7Y103_SLICE_X8Y103_B1 = RIOB33_X105Y101_IOB_X1Y101_I;
  assign CLBLM_R_X7Y103_SLICE_X8Y103_B2 = RIOB33_X105Y101_IOB_X1Y102_I;
  assign CLBLM_R_X7Y103_SLICE_X8Y103_B3 = RIOB33_X105Y113_IOB_X1Y113_I;
  assign CLBLM_R_X7Y103_SLICE_X8Y103_B4 = RIOB33_X105Y111_IOB_X1Y112_I;
  assign CLBLM_R_X7Y103_SLICE_X8Y103_B5 = RIOB33_X105Y103_IOB_X1Y103_I;
  assign CLBLM_R_X7Y103_SLICE_X8Y103_B6 = LIOB33_SING_X0Y100_IOB_X0Y100_I;
  assign CLBLM_R_X7Y103_SLICE_X8Y103_C1 = RIOB33_X105Y113_IOB_X1Y113_I;
  assign CLBLM_R_X7Y103_SLICE_X8Y103_C2 = LIOB33_SING_X0Y100_IOB_X0Y100_I;
  assign CLBLM_R_X7Y103_SLICE_X8Y103_C3 = RIOB33_X105Y101_IOB_X1Y102_I;
  assign CLBLM_R_X7Y103_SLICE_X8Y103_C4 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLM_R_X7Y103_SLICE_X8Y103_C5 = RIOB33_X105Y101_IOB_X1Y101_I;
  assign CLBLM_R_X7Y103_SLICE_X8Y103_C6 = RIOB33_X105Y111_IOB_X1Y112_I;
  assign CLBLM_R_X7Y103_SLICE_X8Y103_D1 = CLBLM_R_X7Y103_SLICE_X8Y103_AO6;
  assign CLBLM_R_X7Y103_SLICE_X8Y103_D2 = LIOB33_X0Y101_IOB_X0Y101_I;
  assign CLBLM_R_X7Y103_SLICE_X8Y103_D3 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLM_R_X7Y103_SLICE_X8Y103_D4 = CLBLM_R_X7Y103_SLICE_X8Y103_CO6;
  assign CLBLM_R_X7Y103_SLICE_X8Y103_D5 = RIOB33_X105Y101_IOB_X1Y101_I;
  assign CLBLM_R_X7Y103_SLICE_X8Y103_D6 = CLBLM_R_X7Y103_SLICE_X8Y103_BO6;
  assign CLBLM_L_X8Y110_SLICE_X11Y110_A1 = 1'b1;
  assign CLBLM_L_X8Y110_SLICE_X11Y110_A2 = LIOB33_X0Y111_IOB_X0Y111_I;
  assign CLBLM_L_X8Y110_SLICE_X11Y110_A3 = RIOB33_X105Y101_IOB_X1Y101_I;
  assign CLBLM_L_X8Y110_SLICE_X11Y110_A4 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLM_L_X8Y110_SLICE_X11Y110_A5 = 1'b1;
  assign CLBLM_L_X8Y110_SLICE_X11Y110_A6 = 1'b1;
  assign CLBLM_L_X8Y110_SLICE_X11Y110_B1 = CLBLM_L_X10Y109_SLICE_X12Y109_AO6;
  assign CLBLM_L_X8Y110_SLICE_X11Y110_B2 = LIOB33_X0Y109_IOB_X0Y109_I;
  assign CLBLM_L_X8Y110_SLICE_X11Y110_B3 = LIOB33_X0Y109_IOB_X0Y110_I;
  assign CLBLM_L_X8Y110_SLICE_X11Y110_B4 = RIOB33_X105Y101_IOB_X1Y101_I;
  assign CLBLM_L_X8Y110_SLICE_X11Y110_B5 = CLBLM_R_X11Y109_SLICE_X14Y109_BO6;
  assign CLBLM_L_X8Y110_SLICE_X11Y110_B6 = CLBLM_L_X10Y110_SLICE_X12Y110_AO6;
  assign CLBLL_L_X4Y116_SLICE_X4Y116_A1 = 1'b1;
  assign CLBLL_L_X4Y116_SLICE_X4Y116_A2 = 1'b1;
  assign CLBLL_L_X4Y116_SLICE_X4Y116_A3 = CLBLL_L_X4Y115_SLICE_X4Y115_AO6;
  assign CLBLL_L_X4Y116_SLICE_X4Y116_A4 = 1'b1;
  assign CLBLL_L_X4Y116_SLICE_X4Y116_A5 = 1'b1;
  assign CLBLL_L_X4Y116_SLICE_X4Y116_A6 = CLBLL_L_X4Y114_SLICE_X4Y114_CO6;
  assign CLBLM_L_X8Y110_SLICE_X11Y110_C3 = CLBLM_L_X10Y109_SLICE_X12Y109_AO6;
  assign CLBLM_L_X8Y110_SLICE_X11Y110_C1 = CLBLM_R_X11Y109_SLICE_X14Y109_BO6;
  assign CLBLM_L_X8Y110_SLICE_X11Y110_C6 = LIOB33_X0Y109_IOB_X0Y109_I;
  assign CLBLM_L_X8Y110_SLICE_X11Y110_C2 = CLBLM_L_X10Y110_SLICE_X12Y110_AO6;
  assign CLBLL_L_X4Y116_SLICE_X4Y116_B1 = 1'b1;
  assign CLBLL_L_X4Y116_SLICE_X4Y116_B2 = 1'b1;
  assign CLBLL_L_X4Y116_SLICE_X4Y116_B3 = 1'b1;
  assign CLBLL_L_X4Y116_SLICE_X4Y116_B4 = 1'b1;
  assign CLBLL_L_X4Y116_SLICE_X4Y116_B5 = 1'b1;
  assign CLBLL_L_X4Y116_SLICE_X4Y116_B6 = 1'b1;
  assign CLBLL_L_X4Y116_SLICE_X4Y116_C1 = 1'b1;
  assign CLBLL_L_X4Y116_SLICE_X4Y116_C2 = 1'b1;
  assign CLBLL_L_X4Y116_SLICE_X4Y116_C3 = 1'b1;
  assign CLBLL_L_X4Y116_SLICE_X4Y116_C4 = 1'b1;
  assign CLBLL_L_X4Y116_SLICE_X4Y116_C5 = 1'b1;
  assign CLBLL_L_X4Y116_SLICE_X4Y116_C6 = 1'b1;
  assign CLBLM_L_X8Y110_SLICE_X11Y110_D1 = 1'b1;
  assign CLBLM_L_X8Y110_SLICE_X11Y110_D2 = 1'b1;
  assign CLBLM_L_X8Y110_SLICE_X11Y110_D3 = 1'b1;
  assign CLBLM_L_X8Y110_SLICE_X11Y110_D4 = 1'b1;
  assign CLBLM_L_X8Y110_SLICE_X11Y110_D5 = 1'b1;
  assign CLBLM_L_X8Y110_SLICE_X11Y110_D6 = 1'b1;
  assign CLBLM_L_X8Y110_SLICE_X10Y110_A1 = CLBLM_L_X8Y110_SLICE_X11Y110_AO5;
  assign CLBLM_L_X8Y110_SLICE_X10Y110_A3 = CLBLM_L_X8Y110_SLICE_X11Y110_AO6;
  assign CLBLM_L_X8Y110_SLICE_X10Y110_A4 = CLBLM_L_X8Y110_SLICE_X11Y110_CO6;
  assign CLBLM_L_X8Y110_SLICE_X10Y110_A5 = CLBLM_L_X8Y108_SLICE_X11Y108_AO6;
  assign CLBLM_L_X8Y110_SLICE_X10Y110_A2 = CLBLM_L_X8Y110_SLICE_X11Y110_BO6;
  assign CLBLL_L_X4Y116_SLICE_X4Y116_D1 = 1'b1;
  assign CLBLL_L_X4Y116_SLICE_X4Y116_D2 = 1'b1;
  assign CLBLL_L_X4Y116_SLICE_X4Y116_D3 = 1'b1;
  assign CLBLL_L_X4Y116_SLICE_X4Y116_D4 = 1'b1;
  assign CLBLL_L_X4Y116_SLICE_X4Y116_D5 = 1'b1;
  assign CLBLL_L_X4Y116_SLICE_X4Y116_D6 = 1'b1;
  assign CLBLM_L_X8Y110_SLICE_X10Y110_A6 = CLBLM_L_X10Y112_SLICE_X12Y112_AO6;
  assign CLBLM_L_X8Y110_SLICE_X10Y110_B1 = CLBLM_L_X8Y110_SLICE_X11Y110_AO5;
  assign CLBLM_L_X8Y110_SLICE_X10Y110_B2 = CLBLM_L_X8Y110_SLICE_X11Y110_BO6;
  assign CLBLM_L_X8Y110_SLICE_X10Y110_B3 = CLBLM_L_X8Y110_SLICE_X11Y110_AO6;
  assign CLBLM_L_X8Y110_SLICE_X10Y110_B4 = CLBLM_L_X8Y112_SLICE_X10Y112_AO6;
  assign CLBLM_L_X8Y110_SLICE_X10Y110_B5 = CLBLM_L_X8Y108_SLICE_X11Y108_AO6;
  assign CLBLM_L_X8Y110_SLICE_X10Y110_B6 = CLBLM_L_X10Y110_SLICE_X13Y110_BO6;
  assign CLBLM_L_X8Y110_SLICE_X10Y110_C1 = CLBLM_L_X8Y108_SLICE_X11Y108_AO6;
  assign CLBLM_L_X8Y110_SLICE_X10Y110_C2 = CLBLM_L_X8Y110_SLICE_X11Y110_CO6;
  assign CLBLM_L_X8Y110_SLICE_X10Y110_C3 = CLBLM_L_X8Y110_SLICE_X11Y110_BO6;
  assign CLBLM_L_X8Y110_SLICE_X10Y110_C4 = CLBLM_L_X10Y112_SLICE_X12Y112_AO6;
  assign CLBLM_L_X8Y110_SLICE_X10Y110_C5 = CLBLM_L_X8Y110_SLICE_X11Y110_AO5;
  assign CLBLM_L_X8Y110_SLICE_X10Y110_C6 = CLBLM_L_X8Y110_SLICE_X11Y110_AO6;
  assign CLBLM_L_X8Y110_SLICE_X10Y110_D1 = 1'b1;
  assign CLBLM_L_X8Y110_SLICE_X10Y110_D2 = 1'b1;
  assign CLBLM_L_X8Y110_SLICE_X10Y110_D3 = 1'b1;
  assign CLBLL_L_X4Y116_SLICE_X5Y116_A4 = 1'b1;
  assign CLBLL_L_X4Y116_SLICE_X5Y116_A5 = 1'b1;
  assign CLBLL_L_X4Y116_SLICE_X5Y116_A6 = 1'b1;
  assign CLBLM_L_X8Y110_SLICE_X10Y110_D4 = 1'b1;
  assign CLBLM_L_X8Y110_SLICE_X10Y110_D5 = 1'b1;
  assign CLBLL_L_X4Y116_SLICE_X5Y116_A1 = 1'b1;
  assign CLBLL_L_X4Y116_SLICE_X5Y116_A2 = 1'b1;
  assign CLBLL_L_X4Y116_SLICE_X5Y116_A3 = 1'b1;
  assign CLBLM_L_X8Y110_SLICE_X10Y110_D6 = 1'b1;
  assign CLBLL_L_X4Y116_SLICE_X5Y116_B1 = 1'b1;
  assign CLBLL_L_X4Y116_SLICE_X5Y116_B2 = 1'b1;
  assign CLBLL_L_X4Y116_SLICE_X5Y116_B3 = 1'b1;
  assign CLBLL_L_X4Y116_SLICE_X5Y116_B4 = 1'b1;
  assign CLBLL_L_X4Y116_SLICE_X5Y116_B5 = 1'b1;
  assign CLBLL_L_X4Y116_SLICE_X5Y116_B6 = 1'b1;
  assign CLBLL_L_X4Y116_SLICE_X5Y116_C1 = 1'b1;
  assign CLBLL_L_X4Y116_SLICE_X5Y116_C2 = 1'b1;
  assign CLBLL_L_X4Y116_SLICE_X5Y116_C3 = 1'b1;
  assign CLBLL_L_X4Y116_SLICE_X5Y116_C4 = 1'b1;
  assign CLBLL_L_X4Y116_SLICE_X5Y116_C5 = 1'b1;
  assign CLBLL_L_X4Y116_SLICE_X5Y116_C6 = 1'b1;
  assign CLBLL_L_X4Y116_SLICE_X5Y116_D1 = 1'b1;
  assign CLBLL_L_X4Y116_SLICE_X5Y116_D2 = 1'b1;
  assign CLBLL_L_X4Y116_SLICE_X5Y116_D3 = 1'b1;
  assign CLBLL_L_X4Y116_SLICE_X5Y116_D4 = 1'b1;
  assign CLBLL_L_X4Y116_SLICE_X5Y116_D5 = 1'b1;
  assign CLBLL_L_X4Y116_SLICE_X5Y116_D6 = 1'b1;
  assign CLBLM_R_X7Y104_SLICE_X9Y104_A1 = LIOB33_X0Y105_IOB_X0Y105_I;
  assign CLBLM_R_X7Y104_SLICE_X9Y104_A2 = LIOB33_X0Y103_IOB_X0Y104_I;
  assign CLBLM_R_X7Y104_SLICE_X9Y104_A3 = 1'b1;
  assign CLBLM_R_X7Y104_SLICE_X9Y104_A4 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLM_R_X7Y104_SLICE_X9Y104_A5 = 1'b1;
  assign CLBLM_R_X7Y104_SLICE_X9Y104_A6 = 1'b1;
  assign CLBLM_R_X7Y104_SLICE_X9Y104_B1 = CLBLM_L_X8Y104_SLICE_X10Y104_CO6;
  assign CLBLM_R_X7Y104_SLICE_X9Y104_B2 = CLBLM_L_X10Y102_SLICE_X12Y102_BO6;
  assign CLBLM_R_X7Y104_SLICE_X9Y104_B3 = CLBLM_L_X8Y105_SLICE_X11Y105_AO6;
  assign CLBLM_R_X7Y104_SLICE_X9Y104_B4 = CLBLM_R_X7Y104_SLICE_X8Y104_DO6;
  assign CLBLM_R_X7Y104_SLICE_X9Y104_B5 = CLBLM_R_X7Y104_SLICE_X9Y104_AO6;
  assign CLBLM_R_X7Y104_SLICE_X9Y104_B6 = CLBLM_L_X8Y104_SLICE_X10Y104_BO6;
  assign CLBLM_R_X7Y104_SLICE_X9Y104_C1 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLM_R_X7Y104_SLICE_X9Y104_C2 = LIOB33_X0Y103_IOB_X0Y104_I;
  assign CLBLM_R_X7Y104_SLICE_X9Y104_C3 = CLBLM_R_X7Y104_SLICE_X8Y104_DO6;
  assign CLBLM_R_X7Y104_SLICE_X9Y104_C4 = CLBLM_L_X8Y104_SLICE_X10Y104_DO6;
  assign CLBLM_R_X7Y104_SLICE_X9Y104_C5 = RIOB33_X105Y101_IOB_X1Y101_I;
  assign CLBLM_R_X7Y104_SLICE_X9Y104_C6 = LIOB33_X0Y101_IOB_X0Y102_I;
  assign CLBLM_R_X7Y104_SLICE_X9Y104_D1 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLM_R_X7Y104_SLICE_X9Y104_D2 = CLBLM_L_X8Y104_SLICE_X10Y104_DO6;
  assign CLBLM_R_X7Y104_SLICE_X9Y104_D3 = CLBLM_R_X7Y104_SLICE_X8Y104_BO5;
  assign CLBLM_R_X7Y104_SLICE_X9Y104_D4 = CLBLM_L_X8Y103_SLICE_X10Y103_AO6;
  assign CLBLM_R_X7Y104_SLICE_X9Y104_D5 = RIOB33_X105Y101_IOB_X1Y101_I;
  assign CLBLM_R_X7Y104_SLICE_X9Y104_D6 = LIOB33_X0Y101_IOB_X0Y102_I;
  assign CLBLM_R_X7Y104_SLICE_X8Y104_A1 = 1'b1;
  assign CLBLM_R_X7Y104_SLICE_X8Y104_A2 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLM_R_X7Y104_SLICE_X8Y104_A3 = LIOB33_X0Y101_IOB_X0Y101_I;
  assign CLBLM_R_X7Y104_SLICE_X8Y104_A4 = LIOB33_X0Y101_IOB_X0Y102_I;
  assign CLBLM_R_X7Y104_SLICE_X8Y104_A5 = 1'b1;
  assign CLBLM_R_X7Y104_SLICE_X8Y104_A6 = 1'b1;
  assign CLBLM_R_X7Y104_SLICE_X8Y104_B1 = 1'b1;
  assign CLBLM_R_X7Y104_SLICE_X8Y104_B2 = CLBLM_R_X7Y103_SLICE_X8Y103_CO6;
  assign CLBLM_R_X7Y104_SLICE_X8Y104_B3 = CLBLM_R_X7Y103_SLICE_X8Y103_AO6;
  assign CLBLM_R_X7Y104_SLICE_X8Y104_B4 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLM_R_X7Y104_SLICE_X8Y104_B5 = LIOB33_X0Y101_IOB_X0Y101_I;
  assign CLBLM_R_X7Y104_SLICE_X8Y104_B6 = 1'b1;
  assign LIOI3_X0Y115_ILOGIC_X0Y116_D = LIOB33_X0Y115_IOB_X0Y116_I;
  assign LIOI3_X0Y115_ILOGIC_X0Y115_D = LIOB33_X0Y115_IOB_X0Y115_I;
  assign CLBLM_R_X7Y104_SLICE_X8Y104_C1 = CLBLM_R_X7Y104_SLICE_X8Y104_AO6;
  assign CLBLM_R_X7Y104_SLICE_X8Y104_C2 = CLBLM_R_X7Y103_SLICE_X8Y103_CO6;
  assign CLBLM_R_X7Y104_SLICE_X8Y104_C3 = CLBLM_R_X7Y103_SLICE_X8Y103_AO6;
  assign CLBLM_R_X7Y104_SLICE_X8Y104_C4 = CLBLM_R_X7Y104_SLICE_X8Y104_AO5;
  assign CLBLM_R_X7Y104_SLICE_X8Y104_C5 = CLBLM_L_X8Y104_SLICE_X10Y104_AO6;
  assign CLBLM_R_X7Y104_SLICE_X8Y104_C6 = CLBLM_R_X7Y103_SLICE_X8Y103_BO6;
  assign CLBLM_R_X7Y104_SLICE_X8Y104_D1 = CLBLM_R_X7Y104_SLICE_X8Y104_AO6;
  assign CLBLM_R_X7Y104_SLICE_X8Y104_D2 = CLBLM_R_X7Y103_SLICE_X8Y103_CO6;
  assign CLBLM_R_X7Y104_SLICE_X8Y104_D3 = CLBLM_R_X7Y103_SLICE_X8Y103_AO6;
  assign CLBLM_R_X7Y104_SLICE_X8Y104_D4 = CLBLM_R_X7Y104_SLICE_X8Y104_AO5;
  assign CLBLM_R_X7Y104_SLICE_X8Y104_D5 = CLBLM_L_X8Y104_SLICE_X10Y104_AO6;
  assign CLBLM_R_X7Y104_SLICE_X8Y104_D6 = CLBLM_R_X7Y103_SLICE_X8Y103_BO6;
  assign CLBLM_L_X8Y111_SLICE_X11Y111_A1 = CLBLM_L_X10Y112_SLICE_X13Y112_CO6;
  assign CLBLM_L_X8Y111_SLICE_X11Y111_A2 = LIOB33_X0Y109_IOB_X0Y110_I;
  assign CLBLM_L_X8Y111_SLICE_X11Y111_A3 = 1'b1;
  assign CLBLM_L_X8Y111_SLICE_X11Y111_A4 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X8Y111_SLICE_X11Y111_A5 = CLBLM_L_X10Y111_SLICE_X12Y111_DO6;
  assign CLBLM_L_X8Y111_SLICE_X11Y111_A6 = 1'b1;
  assign CLBLM_L_X8Y111_SLICE_X11Y111_B1 = CLBLM_L_X8Y111_SLICE_X11Y111_DO6;
  assign CLBLM_L_X8Y111_SLICE_X11Y111_B2 = CLBLM_L_X10Y111_SLICE_X12Y111_BO6;
  assign CLBLM_L_X8Y111_SLICE_X11Y111_B3 = CLBLM_L_X10Y111_SLICE_X13Y111_AO5;
  assign CLBLM_L_X8Y111_SLICE_X11Y111_B4 = CLBLM_R_X11Y111_SLICE_X14Y111_AO5;
  assign CLBLM_L_X8Y111_SLICE_X11Y111_B5 = CLBLM_L_X10Y111_SLICE_X12Y111_DO6;
  assign CLBLM_L_X8Y111_SLICE_X11Y111_B6 = CLBLM_L_X10Y112_SLICE_X13Y112_CO6;
  assign CLBLM_L_X8Y111_SLICE_X11Y111_C1 = CLBLM_L_X8Y111_SLICE_X11Y111_AO6;
  assign CLBLM_L_X8Y111_SLICE_X11Y111_C2 = CLBLM_L_X10Y111_SLICE_X12Y111_BO6;
  assign CLBLM_L_X8Y111_SLICE_X11Y111_C3 = RIOB33_X105Y103_IOB_X1Y104_I;
  assign CLBLM_L_X8Y111_SLICE_X11Y111_C4 = LIOB33_X0Y109_IOB_X0Y110_I;
  assign CLBLM_L_X8Y111_SLICE_X11Y111_C5 = LIOB33_X0Y111_IOB_X0Y111_I;
  assign CLBLM_L_X8Y111_SLICE_X11Y111_C6 = CLBLM_R_X11Y111_SLICE_X14Y111_AO5;
  assign CLBLM_L_X8Y111_SLICE_X11Y111_D1 = 1'b1;
  assign CLBLM_L_X8Y111_SLICE_X11Y111_D2 = LIOB33_X0Y109_IOB_X0Y110_I;
  assign CLBLM_L_X8Y111_SLICE_X11Y111_D3 = 1'b1;
  assign CLBLM_L_X8Y111_SLICE_X11Y111_D4 = 1'b1;
  assign CLBLM_L_X8Y111_SLICE_X11Y111_D5 = 1'b1;
  assign CLBLM_L_X8Y111_SLICE_X11Y111_D6 = RIOB33_X105Y103_IOB_X1Y104_I;
  assign CLBLM_L_X8Y111_SLICE_X10Y111_A1 = CLBLM_L_X10Y111_SLICE_X12Y111_CO6;
  assign CLBLM_L_X8Y111_SLICE_X10Y111_A2 = RIOB33_X105Y103_IOB_X1Y104_I;
  assign CLBLM_L_X8Y111_SLICE_X10Y111_A3 = LIOB33_X0Y109_IOB_X0Y110_I;
  assign CLBLM_L_X8Y111_SLICE_X10Y111_A4 = CLBLM_R_X11Y111_SLICE_X14Y111_AO5;
  assign CLBLM_L_X8Y111_SLICE_X10Y111_A5 = CLBLM_L_X10Y111_SLICE_X12Y111_BO6;
  assign CLBLM_L_X8Y111_SLICE_X10Y111_A6 = 1'b1;
  assign CLBLM_L_X8Y111_SLICE_X10Y111_B1 = LIOB33_X0Y111_IOB_X0Y111_I;
  assign CLBLM_L_X8Y111_SLICE_X10Y111_B2 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLM_L_X8Y111_SLICE_X10Y111_B3 = CLBLM_L_X8Y108_SLICE_X11Y108_AO6;
  assign CLBLM_L_X8Y111_SLICE_X10Y111_B4 = CLBLM_L_X10Y110_SLICE_X12Y110_BO6;
  assign CLBLM_L_X8Y111_SLICE_X10Y111_B5 = LIOB33_X0Y109_IOB_X0Y110_I;
  assign CLBLM_L_X8Y111_SLICE_X10Y111_B6 = RIOB33_X105Y101_IOB_X1Y101_I;
  assign CLBLM_L_X8Y111_SLICE_X10Y111_C1 = CLBLM_L_X8Y108_SLICE_X11Y108_AO6;
  assign CLBLM_L_X8Y111_SLICE_X10Y111_C2 = RIOB33_X105Y101_IOB_X1Y101_I;
  assign CLBLM_L_X8Y111_SLICE_X10Y111_C3 = LIOB33_X0Y111_IOB_X0Y111_I;
  assign CLBLM_L_X8Y111_SLICE_X10Y111_C4 = CLBLM_L_X10Y110_SLICE_X12Y110_BO6;
  assign CLBLM_L_X8Y111_SLICE_X10Y111_C5 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLM_L_X8Y111_SLICE_X10Y111_C6 = LIOB33_X0Y109_IOB_X0Y110_I;
  assign CLBLM_L_X8Y111_SLICE_X10Y111_D1 = 1'b1;
  assign CLBLM_L_X8Y111_SLICE_X10Y111_D2 = 1'b1;
  assign CLBLM_L_X8Y111_SLICE_X10Y111_D3 = 1'b1;
  assign CLBLM_L_X8Y111_SLICE_X10Y111_D4 = 1'b1;
  assign CLBLM_L_X8Y111_SLICE_X10Y111_D5 = 1'b1;
  assign CLBLM_L_X8Y111_SLICE_X10Y111_D6 = 1'b1;
  assign CLBLL_L_X4Y112_SLICE_X4Y112_B3 = RIOB33_X105Y101_IOB_X1Y101_I;
  assign CLBLL_L_X4Y112_SLICE_X4Y112_B4 = CLBLM_R_X7Y112_SLICE_X9Y112_CO6;
  assign CLBLL_L_X4Y112_SLICE_X4Y112_B5 = LIOB33_X0Y115_IOB_X0Y115_I;
  assign CLBLL_L_X4Y112_SLICE_X4Y112_B6 = LIOB33_X0Y113_IOB_X0Y113_I;
  assign CLBLM_R_X7Y105_SLICE_X9Y105_A1 = CLBLM_R_X5Y104_SLICE_X7Y104_BO6;
  assign CLBLM_R_X7Y105_SLICE_X9Y105_A2 = CLBLM_R_X5Y106_SLICE_X7Y106_AO6;
  assign CLBLM_R_X7Y105_SLICE_X9Y105_A3 = CLBLM_R_X7Y104_SLICE_X9Y104_BO6;
  assign CLBLM_R_X7Y105_SLICE_X9Y105_A4 = CLBLM_L_X8Y105_SLICE_X10Y105_AO6;
  assign CLBLM_R_X7Y105_SLICE_X9Y105_A5 = CLBLM_R_X7Y104_SLICE_X9Y104_CO6;
  assign CLBLM_R_X7Y105_SLICE_X9Y105_A6 = CLBLM_R_X7Y104_SLICE_X9Y104_AO5;
  assign CLBLM_R_X7Y105_SLICE_X9Y105_B1 = CLBLM_R_X5Y104_SLICE_X7Y104_BO6;
  assign CLBLM_R_X7Y105_SLICE_X9Y105_B2 = CLBLM_L_X8Y105_SLICE_X10Y105_AO6;
  assign CLBLM_R_X7Y105_SLICE_X9Y105_B3 = CLBLM_R_X7Y104_SLICE_X9Y104_BO6;
  assign CLBLM_R_X7Y105_SLICE_X9Y105_B4 = CLBLM_R_X5Y106_SLICE_X7Y106_AO6;
  assign CLBLM_R_X7Y105_SLICE_X9Y105_B5 = CLBLM_R_X7Y104_SLICE_X9Y104_CO6;
  assign CLBLM_R_X7Y105_SLICE_X9Y105_B6 = CLBLM_R_X7Y104_SLICE_X9Y104_AO5;
  assign CLBLM_R_X7Y105_SLICE_X9Y105_C1 = LIOB33_X0Y115_IOB_X0Y116_I;
  assign CLBLM_R_X7Y105_SLICE_X9Y105_C2 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLM_R_X7Y105_SLICE_X9Y105_C3 = LIOB33_X0Y105_IOB_X0Y105_I;
  assign CLBLM_R_X7Y105_SLICE_X9Y105_C4 = CLBLM_R_X7Y104_SLICE_X9Y104_BO6;
  assign CLBLM_R_X7Y105_SLICE_X9Y105_C5 = CLBLM_R_X5Y104_SLICE_X7Y104_BO6;
  assign CLBLM_R_X7Y105_SLICE_X9Y105_C6 = CLBLM_R_X7Y104_SLICE_X9Y104_CO6;
  assign CLBLM_R_X7Y105_SLICE_X9Y105_D1 = LIOB33_X0Y115_IOB_X0Y116_I;
  assign CLBLM_R_X7Y105_SLICE_X9Y105_D2 = LIOB33_X0Y103_IOB_X0Y104_I;
  assign CLBLM_R_X7Y105_SLICE_X9Y105_D3 = LIOB33_X0Y105_IOB_X0Y105_I;
  assign CLBLM_R_X7Y105_SLICE_X9Y105_D4 = CLBLM_R_X5Y104_SLICE_X7Y104_BO6;
  assign CLBLM_R_X7Y105_SLICE_X9Y105_D5 = CLBLM_R_X7Y104_SLICE_X9Y104_DO6;
  assign CLBLM_R_X7Y105_SLICE_X9Y105_D6 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLM_R_X7Y105_SLICE_X8Y105_A1 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLM_R_X7Y105_SLICE_X8Y105_A2 = CLBLM_R_X7Y105_SLICE_X9Y105_BO6;
  assign CLBLM_R_X7Y105_SLICE_X8Y105_A3 = CLBLM_L_X8Y106_SLICE_X11Y106_AO6;
  assign CLBLM_R_X7Y105_SLICE_X8Y105_A4 = CLBLM_L_X8Y104_SLICE_X11Y104_CO6;
  assign CLBLM_R_X7Y105_SLICE_X8Y105_A5 = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLM_R_X7Y105_SLICE_X8Y105_A6 = 1'b1;
  assign CLBLM_R_X7Y105_SLICE_X8Y105_B1 = CLBLM_R_X7Y105_SLICE_X9Y105_CO6;
  assign CLBLM_R_X7Y105_SLICE_X8Y105_B2 = LIOB33_X0Y107_IOB_X0Y107_I;
  assign CLBLM_R_X7Y105_SLICE_X8Y105_B3 = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLM_R_X7Y105_SLICE_X8Y105_B4 = CLBLM_R_X5Y105_SLICE_X7Y105_CO6;
  assign CLBLM_R_X7Y105_SLICE_X8Y105_B5 = LIOB33_X0Y115_IOB_X0Y116_I;
  assign CLBLM_R_X7Y105_SLICE_X8Y105_B6 = LIOB33_X0Y113_IOB_X0Y114_I;
  assign CLBLM_R_X7Y105_SLICE_X8Y105_C1 = LIOB33_X0Y115_IOB_X0Y116_I;
  assign CLBLM_R_X7Y105_SLICE_X8Y105_C2 = LIOB33_X0Y113_IOB_X0Y114_I;
  assign CLBLM_R_X7Y105_SLICE_X8Y105_C3 = LIOB33_X0Y107_IOB_X0Y108_I;
  assign CLBLM_R_X7Y105_SLICE_X8Y105_C4 = CLBLM_R_X7Y105_SLICE_X8Y105_AO5;
  assign CLBLM_R_X7Y105_SLICE_X8Y105_C5 = LIOB33_X0Y107_IOB_X0Y107_I;
  assign CLBLM_R_X7Y105_SLICE_X8Y105_C6 = CLBLM_R_X7Y105_SLICE_X8Y105_BO6;
  assign CLBLM_R_X7Y105_SLICE_X8Y105_D1 = LIOB33_X0Y115_IOB_X0Y116_I;
  assign CLBLM_R_X7Y105_SLICE_X8Y105_D2 = LIOB33_X0Y113_IOB_X0Y114_I;
  assign CLBLM_R_X7Y105_SLICE_X8Y105_D3 = LIOB33_X0Y107_IOB_X0Y108_I;
  assign CLBLM_R_X7Y105_SLICE_X8Y105_D4 = CLBLM_R_X7Y105_SLICE_X8Y105_AO5;
  assign CLBLM_R_X7Y105_SLICE_X8Y105_D5 = LIOB33_X0Y107_IOB_X0Y107_I;
  assign CLBLM_R_X7Y105_SLICE_X8Y105_D6 = CLBLM_R_X7Y105_SLICE_X8Y105_BO6;
  assign CLBLM_R_X5Y113_SLICE_X7Y113_C4 = CLBLM_R_X5Y111_SLICE_X7Y111_DO6;
  assign CLBLM_R_X5Y113_SLICE_X7Y113_C5 = LIOB33_X0Y113_IOB_X0Y113_I;
  assign CLBLM_R_X5Y113_SLICE_X7Y113_C6 = CLBLM_R_X5Y112_SLICE_X7Y112_CO6;
  assign CLBLM_L_X8Y112_SLICE_X11Y112_A1 = RIOB33_X105Y101_IOB_X1Y102_I;
  assign CLBLM_L_X8Y112_SLICE_X11Y112_A2 = LIOB33_X0Y111_IOB_X0Y111_I;
  assign CLBLM_L_X8Y112_SLICE_X11Y112_A3 = CLBLM_L_X10Y110_SLICE_X12Y110_DO6;
  assign CLBLM_L_X8Y112_SLICE_X11Y112_A4 = RIOB33_X105Y101_IOB_X1Y101_I;
  assign CLBLM_L_X8Y112_SLICE_X11Y112_A5 = LIOB33_X0Y109_IOB_X0Y110_I;
  assign CLBLM_L_X8Y112_SLICE_X11Y112_A6 = CLBLM_L_X8Y110_SLICE_X11Y110_CO6;
  assign CLBLM_L_X8Y112_SLICE_X11Y112_B1 = LIOB33_X0Y111_IOB_X0Y111_I;
  assign CLBLM_L_X8Y112_SLICE_X11Y112_B2 = CLBLM_L_X10Y112_SLICE_X12Y112_BO6;
  assign CLBLM_L_X8Y112_SLICE_X11Y112_B3 = LIOB33_X0Y109_IOB_X0Y110_I;
  assign CLBLM_L_X8Y112_SLICE_X11Y112_B4 = RIOB33_X105Y103_IOB_X1Y103_I;
  assign CLBLM_L_X8Y112_SLICE_X11Y112_B5 = CLBLM_L_X10Y111_SLICE_X13Y111_CO6;
  assign CLBLM_L_X8Y112_SLICE_X11Y112_B6 = RIOB33_X105Y101_IOB_X1Y102_I;
  assign CLBLM_L_X8Y112_SLICE_X11Y112_C1 = LIOB33_X0Y109_IOB_X0Y110_I;
  assign CLBLM_L_X8Y112_SLICE_X11Y112_C2 = CLBLM_L_X8Y110_SLICE_X11Y110_CO6;
  assign CLBLM_L_X8Y112_SLICE_X11Y112_C3 = LIOB33_X0Y111_IOB_X0Y111_I;
  assign CLBLM_L_X8Y112_SLICE_X11Y112_C4 = RIOB33_X105Y101_IOB_X1Y102_I;
  assign CLBLM_L_X8Y112_SLICE_X11Y112_C5 = CLBLM_L_X10Y110_SLICE_X12Y110_DO6;
  assign CLBLM_L_X8Y112_SLICE_X11Y112_C6 = RIOB33_X105Y101_IOB_X1Y101_I;
  assign CLBLM_L_X8Y112_SLICE_X11Y112_D1 = LIOB33_X0Y109_IOB_X0Y110_I;
  assign CLBLM_L_X8Y112_SLICE_X11Y112_D2 = CLBLM_L_X10Y112_SLICE_X12Y112_BO6;
  assign CLBLM_L_X8Y112_SLICE_X11Y112_D3 = LIOB33_X0Y111_IOB_X0Y111_I;
  assign CLBLM_L_X8Y112_SLICE_X11Y112_D4 = RIOB33_X105Y101_IOB_X1Y102_I;
  assign CLBLM_L_X8Y112_SLICE_X11Y112_D5 = CLBLM_L_X10Y111_SLICE_X13Y111_CO6;
  assign CLBLM_L_X8Y112_SLICE_X11Y112_D6 = RIOB33_X105Y103_IOB_X1Y103_I;
  assign CLBLM_L_X8Y112_SLICE_X10Y112_A1 = CLBLM_L_X8Y111_SLICE_X10Y111_CO6;
  assign CLBLM_L_X8Y112_SLICE_X10Y112_A2 = 1'b1;
  assign CLBLM_L_X8Y112_SLICE_X10Y112_A3 = CLBLM_L_X8Y112_SLICE_X11Y112_AO6;
  assign CLBLM_L_X8Y112_SLICE_X10Y112_A4 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLM_L_X8Y112_SLICE_X10Y112_A5 = LIOB33_X0Y111_IOB_X0Y112_I;
  assign CLBLM_L_X8Y112_SLICE_X10Y112_A6 = 1'b1;
  assign CLBLM_L_X8Y112_SLICE_X10Y112_B1 = CLBLM_L_X8Y110_SLICE_X11Y110_CO6;
  assign CLBLM_L_X8Y112_SLICE_X10Y112_B2 = CLBLM_L_X10Y111_SLICE_X12Y111_AO6;
  assign CLBLM_L_X8Y112_SLICE_X10Y112_B3 = CLBLM_L_X10Y112_SLICE_X12Y112_AO6;
  assign CLBLM_L_X8Y112_SLICE_X10Y112_B4 = CLBLM_R_X5Y112_SLICE_X7Y112_AO6;
  assign CLBLM_L_X8Y112_SLICE_X10Y112_B5 = CLBLM_L_X8Y110_SLICE_X11Y110_AO5;
  assign CLBLM_L_X8Y112_SLICE_X10Y112_B6 = CLBLM_L_X10Y112_SLICE_X12Y112_BO6;
  assign CLBLM_L_X8Y112_SLICE_X10Y112_C1 = CLBLM_L_X8Y110_SLICE_X11Y110_AO5;
  assign CLBLM_L_X8Y112_SLICE_X10Y112_C2 = CLBLM_L_X10Y112_SLICE_X12Y112_AO6;
  assign CLBLM_L_X8Y112_SLICE_X10Y112_C3 = CLBLM_L_X10Y110_SLICE_X13Y110_CO6;
  assign CLBLM_L_X8Y112_SLICE_X10Y112_C4 = CLBLM_L_X8Y110_SLICE_X11Y110_CO6;
  assign CLBLM_L_X8Y112_SLICE_X10Y112_C5 = CLBLM_R_X7Y112_SLICE_X8Y112_AO6;
  assign CLBLM_L_X8Y112_SLICE_X10Y112_C6 = CLBLM_R_X5Y112_SLICE_X7Y112_AO6;
  assign CLBLL_L_X2Y104_SLICE_X0Y104_A1 = RIOB33_SING_X105Y100_IOB_X1Y100_I;
  assign CLBLL_L_X2Y104_SLICE_X0Y104_A2 = CLBLL_L_X2Y104_SLICE_X1Y104_BO6;
  assign CLBLL_L_X2Y104_SLICE_X0Y104_A3 = LIOB33_X0Y103_IOB_X0Y104_I;
  assign CLBLL_L_X2Y104_SLICE_X0Y104_A4 = 1'b1;
  assign CLBLL_L_X2Y104_SLICE_X0Y104_A5 = LIOB33_X0Y103_IOB_X0Y103_I;
  assign CLBLL_L_X2Y104_SLICE_X0Y104_A6 = 1'b1;
  assign CLBLM_L_X8Y112_SLICE_X10Y112_D1 = LIOB33_X0Y111_IOB_X0Y112_I;
  assign CLBLM_L_X8Y112_SLICE_X10Y112_D2 = CLBLM_L_X8Y111_SLICE_X10Y111_CO6;
  assign CLBLL_L_X2Y104_SLICE_X0Y104_B1 = RIOB33_X105Y111_IOB_X1Y112_I;
  assign CLBLL_L_X2Y104_SLICE_X0Y104_B2 = RIOB33_X105Y105_IOB_X1Y106_I;
  assign CLBLL_L_X2Y104_SLICE_X0Y104_B3 = RIOB33_X105Y113_IOB_X1Y113_I;
  assign CLBLL_L_X2Y104_SLICE_X0Y104_B4 = LIOB33_SING_X0Y100_IOB_X0Y100_I;
  assign CLBLL_L_X2Y104_SLICE_X0Y104_B5 = LIOB33_X0Y103_IOB_X0Y103_I;
  assign CLBLL_L_X2Y104_SLICE_X0Y104_B6 = LIOB33_X0Y113_IOB_X0Y114_I;
  assign CLBLL_L_X2Y104_SLICE_X0Y104_C1 = LIOB33_X0Y103_IOB_X0Y103_I;
  assign CLBLL_L_X2Y104_SLICE_X0Y104_C2 = RIOB33_X105Y105_IOB_X1Y106_I;
  assign CLBLL_L_X2Y104_SLICE_X0Y104_C3 = RIOB33_X105Y111_IOB_X1Y112_I;
  assign CLBLL_L_X2Y104_SLICE_X0Y104_C4 = LIOB33_SING_X0Y100_IOB_X0Y100_I;
  assign CLBLL_L_X2Y104_SLICE_X0Y104_C5 = RIOB33_X105Y113_IOB_X1Y113_I;
  assign CLBLL_L_X2Y104_SLICE_X0Y104_C6 = LIOB33_X0Y113_IOB_X0Y114_I;
  assign LIOI3_X0Y117_OLOGIC_X0Y118_D1 = CLBLL_L_X2Y109_SLICE_X0Y109_AO5;
  assign CLBLL_L_X2Y104_SLICE_X0Y104_D1 = 1'b1;
  assign CLBLL_L_X2Y104_SLICE_X0Y104_D2 = 1'b1;
  assign CLBLL_L_X2Y104_SLICE_X0Y104_D3 = 1'b1;
  assign CLBLL_L_X2Y104_SLICE_X0Y104_D4 = 1'b1;
  assign CLBLL_L_X2Y104_SLICE_X0Y104_D5 = 1'b1;
  assign CLBLL_L_X2Y104_SLICE_X0Y104_D6 = 1'b1;
  assign LIOI3_X0Y117_OLOGIC_X0Y118_T1 = 1'b1;
  assign CLBLM_R_X7Y106_SLICE_X9Y106_A1 = CLBLM_R_X7Y106_SLICE_X8Y106_AO6;
  assign CLBLM_R_X7Y106_SLICE_X9Y106_A2 = CLBLM_R_X7Y105_SLICE_X8Y105_BO6;
  assign CLBLM_R_X7Y106_SLICE_X9Y106_A3 = CLBLM_R_X7Y106_SLICE_X8Y106_CO6;
  assign CLBLM_R_X7Y106_SLICE_X9Y106_A4 = CLBLM_R_X7Y106_SLICE_X8Y106_AO5;
  assign CLBLM_R_X7Y106_SLICE_X9Y106_A5 = CLBLM_L_X8Y105_SLICE_X10Y105_BO6;
  assign CLBLM_R_X7Y106_SLICE_X9Y106_A6 = CLBLM_L_X8Y106_SLICE_X10Y106_BO6;
  assign CLBLL_L_X2Y104_SLICE_X1Y104_A1 = RIOB33_X105Y105_IOB_X1Y106_I;
  assign CLBLL_L_X2Y104_SLICE_X1Y104_A2 = CLBLL_L_X2Y104_SLICE_X0Y104_BO6;
  assign CLBLL_L_X2Y104_SLICE_X1Y104_A3 = CLBLL_L_X2Y104_SLICE_X0Y104_CO6;
  assign CLBLM_R_X7Y106_SLICE_X9Y106_B4 = CLBLM_R_X7Y106_SLICE_X8Y106_AO5;
  assign CLBLM_R_X7Y106_SLICE_X9Y106_B5 = CLBLM_L_X8Y106_SLICE_X10Y106_DO6;
  assign CLBLM_R_X7Y106_SLICE_X9Y106_B6 = CLBLM_R_X5Y106_SLICE_X6Y106_AO5;
  assign CLBLL_L_X2Y104_SLICE_X1Y104_A4 = 1'b1;
  assign CLBLL_L_X2Y104_SLICE_X1Y104_A5 = LIOB33_X0Y101_IOB_X0Y101_I;
  assign CLBLL_L_X2Y104_SLICE_X1Y104_A6 = 1'b1;
  assign CLBLM_R_X7Y106_SLICE_X9Y106_B1 = CLBLM_R_X7Y106_SLICE_X8Y106_AO6;
  assign CLBLM_R_X7Y106_SLICE_X9Y106_B2 = CLBLM_R_X7Y105_SLICE_X8Y105_BO6;
  assign CLBLM_R_X7Y106_SLICE_X9Y106_C3 = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLM_R_X7Y106_SLICE_X9Y106_C4 = CLBLM_L_X8Y104_SLICE_X11Y104_CO6;
  assign CLBLM_R_X7Y106_SLICE_X9Y106_C5 = CLBLM_L_X8Y105_SLICE_X11Y105_DO6;
  assign CLBLM_R_X7Y106_SLICE_X9Y106_C6 = RIOB33_X105Y101_IOB_X1Y101_I;
  assign CLBLL_L_X2Y104_SLICE_X1Y104_B1 = CLBLL_L_X2Y106_SLICE_X1Y106_AO5;
  assign CLBLL_L_X2Y104_SLICE_X1Y104_B2 = CLBLL_L_X2Y104_SLICE_X1Y104_CO6;
  assign CLBLL_L_X2Y104_SLICE_X1Y104_B3 = LIOB33_X0Y101_IOB_X0Y102_I;
  assign CLBLL_L_X2Y104_SLICE_X1Y104_B4 = RIOB33_X105Y105_IOB_X1Y106_I;
  assign CLBLL_L_X2Y104_SLICE_X1Y104_B5 = RIOB33_SING_X105Y100_IOB_X1Y100_I;
  assign CLBLL_L_X2Y104_SLICE_X1Y104_B6 = CLBLL_L_X2Y104_SLICE_X1Y104_AO5;
  assign CLBLL_L_X2Y104_SLICE_X1Y104_C1 = LIOB33_X0Y101_IOB_X0Y101_I;
  assign CLBLL_L_X2Y104_SLICE_X1Y104_C2 = CLBLL_L_X2Y104_SLICE_X0Y104_CO6;
  assign CLBLL_L_X2Y104_SLICE_X1Y104_C3 = CLBLL_L_X2Y104_SLICE_X0Y104_BO6;
  assign CLBLM_R_X7Y106_SLICE_X9Y106_D2 = CLBLM_R_X7Y106_SLICE_X8Y106_CO6;
  assign CLBLM_R_X7Y106_SLICE_X9Y106_D3 = CLBLM_L_X8Y106_SLICE_X10Y106_DO6;
  assign CLBLM_R_X7Y106_SLICE_X9Y106_D4 = CLBLM_R_X5Y106_SLICE_X6Y106_AO5;
  assign CLBLM_R_X7Y106_SLICE_X9Y106_D5 = CLBLM_R_X7Y106_SLICE_X8Y106_AO6;
  assign CLBLM_R_X7Y106_SLICE_X9Y106_D6 = CLBLM_R_X7Y106_SLICE_X8Y106_AO5;
  assign CLBLL_L_X2Y104_SLICE_X1Y104_C4 = LIOB33_X0Y103_IOB_X0Y103_I;
  assign CLBLL_L_X2Y104_SLICE_X1Y104_C5 = CLBLM_R_X3Y105_SLICE_X2Y105_AO6;
  assign CLBLL_L_X2Y104_SLICE_X1Y104_C6 = RIOB33_X105Y105_IOB_X1Y106_I;
  assign CLBLL_L_X2Y104_SLICE_X1Y104_D1 = CLBLL_L_X2Y104_SLICE_X1Y104_AO6;
  assign CLBLL_L_X2Y104_SLICE_X1Y104_D2 = CLBLM_R_X3Y104_SLICE_X2Y104_BO6;
  assign CLBLM_R_X7Y106_SLICE_X8Y106_A1 = LIOB33_X0Y107_IOB_X0Y108_I;
  assign CLBLM_R_X7Y106_SLICE_X8Y106_A2 = 1'b1;
  assign CLBLM_R_X7Y106_SLICE_X8Y106_A3 = LIOB33_X0Y113_IOB_X0Y114_I;
  assign CLBLM_R_X7Y106_SLICE_X8Y106_A4 = 1'b1;
  assign CLBLM_R_X7Y106_SLICE_X8Y106_A5 = LIOB33_X0Y115_IOB_X0Y116_I;
  assign CLBLM_R_X7Y106_SLICE_X8Y106_A6 = 1'b1;
  assign CLBLL_L_X2Y104_SLICE_X1Y104_D3 = LIOB33_X0Y103_IOB_X0Y103_I;
  assign CLBLL_L_X2Y104_SLICE_X1Y104_D4 = RIOB33_X105Y105_IOB_X1Y106_I;
  assign CLBLL_L_X2Y104_SLICE_X1Y104_D5 = LIOB33_X0Y101_IOB_X0Y102_I;
  assign CLBLL_L_X2Y104_SLICE_X1Y104_D6 = CLBLM_R_X3Y104_SLICE_X2Y104_AO6;
  assign CLBLM_R_X7Y106_SLICE_X8Y106_B1 = CLBLM_L_X8Y106_SLICE_X10Y106_AO6;
  assign CLBLM_R_X7Y106_SLICE_X8Y106_B3 = CLBLM_R_X7Y105_SLICE_X9Y105_AO6;
  assign CLBLM_R_X7Y106_SLICE_X8Y106_B4 = CLBLM_R_X5Y106_SLICE_X7Y106_BO6;
  assign CLBLM_R_X7Y106_SLICE_X8Y106_B5 = CLBLM_R_X7Y105_SLICE_X9Y105_BO6;
  assign CLBLM_R_X7Y106_SLICE_X8Y106_B6 = CLBLM_R_X5Y105_SLICE_X7Y105_CO6;
  assign CLBLM_R_X7Y106_SLICE_X8Y106_B2 = CLBLM_L_X8Y104_SLICE_X11Y104_AO6;
  assign CLBLM_R_X7Y106_SLICE_X8Y106_C1 = CLBLM_R_X7Y105_SLICE_X9Y105_BO6;
  assign CLBLM_R_X7Y106_SLICE_X8Y106_C2 = CLBLM_L_X8Y104_SLICE_X11Y104_CO6;
  assign CLBLM_R_X7Y106_SLICE_X8Y106_C3 = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLM_R_X7Y106_SLICE_X8Y106_C4 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLM_R_X7Y106_SLICE_X8Y106_C5 = CLBLM_L_X8Y106_SLICE_X10Y106_AO6;
  assign CLBLM_R_X7Y106_SLICE_X8Y106_C6 = CLBLM_L_X8Y106_SLICE_X11Y106_AO6;
  assign CLBLM_R_X7Y106_SLICE_X8Y106_D1 = CLBLM_R_X3Y106_SLICE_X2Y106_AO6;
  assign CLBLM_R_X7Y106_SLICE_X8Y106_D2 = CLBLM_L_X8Y104_SLICE_X11Y104_CO6;
  assign CLBLM_R_X7Y106_SLICE_X8Y106_D3 = RIOB33_X105Y107_IOB_X1Y108_I;
  assign CLBLM_R_X7Y106_SLICE_X8Y106_D4 = LIOB33_X0Y103_IOB_X0Y104_I;
  assign CLBLM_R_X7Y106_SLICE_X8Y106_D5 = CLBLM_L_X8Y106_SLICE_X11Y106_AO6;
  assign CLBLM_R_X7Y106_SLICE_X8Y106_D6 = CLBLM_L_X12Y107_SLICE_X17Y107_AO5;
  assign CLBLM_L_X8Y113_SLICE_X11Y113_A1 = 1'b1;
  assign CLBLM_L_X8Y113_SLICE_X11Y113_A2 = 1'b1;
  assign CLBLM_L_X8Y113_SLICE_X11Y113_A3 = 1'b1;
  assign CLBLM_L_X8Y113_SLICE_X11Y113_A4 = 1'b1;
  assign CLBLM_L_X8Y113_SLICE_X11Y113_A5 = 1'b1;
  assign CLBLM_L_X8Y113_SLICE_X11Y113_A6 = 1'b1;
  assign CLBLM_L_X8Y113_SLICE_X11Y113_B1 = 1'b1;
  assign CLBLM_L_X8Y113_SLICE_X11Y113_B2 = 1'b1;
  assign CLBLM_L_X8Y113_SLICE_X11Y113_B3 = 1'b1;
  assign CLBLM_L_X8Y113_SLICE_X11Y113_B4 = 1'b1;
  assign CLBLM_L_X8Y113_SLICE_X11Y113_B5 = 1'b1;
  assign CLBLM_L_X8Y113_SLICE_X11Y113_B6 = 1'b1;
  assign LIOI3_X0Y117_ILOGIC_X0Y117_D = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLM_L_X8Y113_SLICE_X11Y113_C1 = 1'b1;
  assign CLBLM_L_X8Y113_SLICE_X11Y113_C2 = 1'b1;
  assign CLBLM_L_X8Y113_SLICE_X11Y113_C3 = 1'b1;
  assign CLBLM_L_X8Y113_SLICE_X11Y113_C4 = 1'b1;
  assign CLBLM_L_X8Y113_SLICE_X11Y113_C5 = 1'b1;
  assign CLBLM_L_X8Y113_SLICE_X11Y113_C6 = 1'b1;
  assign CLBLM_R_X5Y113_SLICE_X7Y113_D5 = 1'b1;
  assign CLBLM_L_X8Y113_SLICE_X11Y113_D1 = 1'b1;
  assign CLBLM_L_X8Y113_SLICE_X11Y113_D2 = 1'b1;
  assign CLBLM_L_X8Y113_SLICE_X11Y113_D3 = 1'b1;
  assign CLBLM_L_X8Y113_SLICE_X11Y113_D4 = 1'b1;
  assign CLBLM_L_X8Y113_SLICE_X11Y113_D5 = 1'b1;
  assign CLBLM_L_X8Y113_SLICE_X11Y113_D6 = 1'b1;
  assign RIOI3_X105Y101_ILOGIC_X1Y102_D = RIOB33_X105Y101_IOB_X1Y102_I;
  assign RIOI3_X105Y101_ILOGIC_X1Y101_D = RIOB33_X105Y101_IOB_X1Y101_I;
  assign CLBLM_L_X8Y113_SLICE_X10Y113_A1 = RIOB33_X105Y107_IOB_X1Y107_I;
  assign CLBLM_L_X8Y113_SLICE_X10Y113_A2 = CLBLM_R_X7Y110_SLICE_X9Y110_BO5;
  assign CLBLM_L_X8Y113_SLICE_X10Y113_A3 = CLBLM_L_X10Y112_SLICE_X13Y112_BO6;
  assign CLBLM_L_X8Y113_SLICE_X10Y113_A4 = CLBLM_L_X8Y111_SLICE_X11Y111_AO5;
  assign CLBLM_L_X8Y113_SLICE_X10Y113_A5 = LIOB33_X0Y109_IOB_X0Y110_I;
  assign CLBLM_L_X8Y113_SLICE_X10Y113_A6 = 1'b1;
  assign CLBLM_L_X8Y113_SLICE_X10Y113_B1 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X8Y113_SLICE_X10Y113_B2 = RIOB33_X105Y103_IOB_X1Y104_I;
  assign CLBLM_L_X8Y113_SLICE_X10Y113_B3 = LIOB33_X0Y111_IOB_X0Y112_I;
  assign CLBLM_L_X8Y113_SLICE_X10Y113_B4 = LIOB33_X0Y111_IOB_X0Y111_I;
  assign CLBLM_L_X8Y113_SLICE_X10Y113_B5 = CLBLM_L_X8Y113_SLICE_X10Y113_AO6;
  assign CLBLM_L_X8Y113_SLICE_X10Y113_B6 = CLBLM_L_X8Y111_SLICE_X11Y111_CO6;
  assign CLBLM_L_X8Y113_SLICE_X10Y113_C1 = LIOB33_X0Y111_IOB_X0Y112_I;
  assign CLBLM_L_X8Y113_SLICE_X10Y113_C2 = CLBLM_L_X8Y113_SLICE_X10Y113_AO6;
  assign CLBLM_L_X8Y113_SLICE_X10Y113_C3 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X8Y113_SLICE_X10Y113_C4 = CLBLM_L_X8Y111_SLICE_X11Y111_CO6;
  assign CLBLM_L_X8Y113_SLICE_X10Y113_C5 = RIOB33_X105Y103_IOB_X1Y104_I;
  assign CLBLM_L_X8Y113_SLICE_X10Y113_C6 = LIOB33_X0Y111_IOB_X0Y111_I;
  assign CLBLM_L_X8Y113_SLICE_X10Y113_D1 = 1'b1;
  assign CLBLM_L_X8Y113_SLICE_X10Y113_D2 = 1'b1;
  assign CLBLM_L_X8Y113_SLICE_X10Y113_D3 = 1'b1;
  assign CLBLM_L_X8Y113_SLICE_X10Y113_D4 = 1'b1;
  assign CLBLM_L_X8Y113_SLICE_X10Y113_D5 = 1'b1;
  assign CLBLM_L_X8Y113_SLICE_X10Y113_D6 = 1'b1;
  assign CLBLM_R_X7Y107_SLICE_X9Y107_A1 = LIOB33_X0Y107_IOB_X0Y108_I;
  assign CLBLM_R_X7Y107_SLICE_X9Y107_A2 = LIOB33_X0Y107_IOB_X0Y107_I;
  assign CLBLM_R_X7Y107_SLICE_X9Y107_A3 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLM_R_X7Y107_SLICE_X9Y107_A4 = CLBLM_L_X8Y105_SLICE_X10Y105_BO6;
  assign CLBLM_R_X7Y107_SLICE_X9Y107_A5 = LIOB33_X0Y115_IOB_X0Y116_I;
  assign CLBLM_R_X7Y107_SLICE_X9Y107_A6 = CLBLM_R_X7Y106_SLICE_X9Y106_CO6;
  assign CLBLM_R_X7Y107_SLICE_X9Y107_B1 = CLBLM_R_X7Y105_SLICE_X8Y105_DO6;
  assign CLBLM_R_X7Y107_SLICE_X9Y107_B2 = LIOB33_X0Y115_IOB_X0Y116_I;
  assign CLBLM_R_X7Y107_SLICE_X9Y107_B3 = LIOB33_X0Y113_IOB_X0Y114_I;
  assign CLBLM_R_X7Y107_SLICE_X9Y107_B4 = CLBLM_L_X8Y107_SLICE_X10Y107_AO6;
  assign CLBLM_R_X7Y107_SLICE_X9Y107_B5 = CLBLM_R_X7Y107_SLICE_X9Y107_AO6;
  assign CLBLM_R_X7Y107_SLICE_X9Y107_B6 = LIOB33_X0Y109_IOB_X0Y109_I;
  assign CLBLM_R_X7Y107_SLICE_X9Y107_C1 = CLBLM_R_X7Y107_SLICE_X9Y107_AO6;
  assign CLBLM_R_X7Y107_SLICE_X9Y107_C2 = LIOB33_X0Y109_IOB_X0Y110_I;
  assign CLBLM_R_X7Y107_SLICE_X9Y107_C3 = CLBLM_R_X7Y105_SLICE_X8Y105_DO6;
  assign CLBLM_R_X7Y107_SLICE_X9Y107_C4 = LIOB33_X0Y109_IOB_X0Y109_I;
  assign CLBLM_R_X7Y107_SLICE_X9Y107_C5 = LIOB33_X0Y113_IOB_X0Y114_I;
  assign CLBLM_R_X7Y107_SLICE_X9Y107_C6 = CLBLM_L_X8Y106_SLICE_X11Y106_BO6;
  assign CLBLM_R_X7Y107_SLICE_X9Y107_D1 = CLBLM_R_X7Y107_SLICE_X9Y107_AO6;
  assign CLBLM_R_X7Y107_SLICE_X9Y107_D2 = LIOB33_X0Y109_IOB_X0Y109_I;
  assign CLBLM_R_X7Y107_SLICE_X9Y107_D3 = LIOB33_X0Y109_IOB_X0Y110_I;
  assign CLBLM_R_X7Y107_SLICE_X9Y107_D4 = CLBLM_R_X7Y105_SLICE_X8Y105_DO6;
  assign CLBLM_R_X7Y107_SLICE_X9Y107_D5 = LIOB33_X0Y113_IOB_X0Y114_I;
  assign CLBLM_R_X7Y107_SLICE_X9Y107_D6 = CLBLM_L_X8Y106_SLICE_X11Y106_BO6;
  assign CLBLM_R_X7Y107_SLICE_X8Y107_A1 = LIOB33_X0Y103_IOB_X0Y103_I;
  assign CLBLM_R_X7Y107_SLICE_X8Y107_A2 = CLBLM_R_X7Y107_SLICE_X9Y107_BO6;
  assign CLBLM_R_X7Y107_SLICE_X8Y107_A3 = LIOB33_X0Y113_IOB_X0Y114_I;
  assign CLBLM_R_X7Y107_SLICE_X8Y107_A4 = LIOB33_X0Y111_IOB_X0Y111_I;
  assign CLBLM_R_X7Y107_SLICE_X8Y107_A5 = LIOB33_X0Y109_IOB_X0Y110_I;
  assign CLBLM_R_X7Y107_SLICE_X8Y107_A6 = CLBLM_R_X5Y107_SLICE_X7Y107_CO6;
  assign CLBLM_R_X7Y107_SLICE_X8Y107_B1 = CLBLM_R_X7Y108_SLICE_X9Y108_BO6;
  assign CLBLM_R_X7Y107_SLICE_X8Y107_B2 = CLBLM_R_X5Y108_SLICE_X7Y108_AO5;
  assign CLBLM_R_X7Y107_SLICE_X8Y107_B3 = CLBLM_R_X7Y107_SLICE_X9Y107_CO6;
  assign CLBLM_R_X7Y107_SLICE_X8Y107_B4 = CLBLM_R_X7Y108_SLICE_X8Y108_AO6;
  assign CLBLM_R_X7Y107_SLICE_X8Y107_B5 = CLBLM_R_X7Y107_SLICE_X9Y107_DO6;
  assign CLBLM_R_X7Y107_SLICE_X8Y107_B6 = CLBLM_R_X5Y107_SLICE_X7Y107_CO6;
  assign CLBLM_R_X7Y107_SLICE_X8Y107_C1 = LIOB33_X0Y113_IOB_X0Y114_I;
  assign CLBLM_R_X7Y107_SLICE_X8Y107_C2 = LIOB33_X0Y109_IOB_X0Y110_I;
  assign CLBLM_R_X7Y107_SLICE_X8Y107_C3 = CLBLM_R_X7Y107_SLICE_X9Y107_BO6;
  assign CLBLM_R_X7Y107_SLICE_X8Y107_C4 = CLBLM_R_X5Y107_SLICE_X7Y107_CO6;
  assign CLBLM_R_X7Y107_SLICE_X8Y107_C5 = LIOB33_X0Y103_IOB_X0Y103_I;
  assign CLBLM_R_X7Y107_SLICE_X8Y107_C6 = LIOB33_X0Y111_IOB_X0Y111_I;
  assign CLBLM_R_X7Y107_SLICE_X8Y107_D1 = CLBLM_L_X8Y107_SLICE_X10Y107_BO6;
  assign CLBLM_R_X7Y107_SLICE_X8Y107_D2 = CLBLM_R_X7Y107_SLICE_X9Y107_CO6;
  assign CLBLM_R_X7Y107_SLICE_X8Y107_D3 = CLBLM_R_X5Y110_SLICE_X7Y110_BO6;
  assign CLBLM_R_X7Y107_SLICE_X8Y107_D4 = CLBLM_R_X5Y107_SLICE_X7Y107_CO6;
  assign CLBLM_R_X7Y107_SLICE_X8Y107_D5 = CLBLM_R_X7Y108_SLICE_X8Y108_AO6;
  assign CLBLM_R_X7Y107_SLICE_X8Y107_D6 = CLBLM_R_X5Y108_SLICE_X7Y108_AO5;
  assign CLBLL_L_X2Y106_SLICE_X0Y106_A1 = 1'b1;
  assign CLBLL_L_X2Y106_SLICE_X0Y106_A2 = RIOB33_SING_X105Y100_IOB_X1Y100_I;
  assign CLBLL_L_X2Y106_SLICE_X0Y106_A3 = CLBLL_L_X2Y106_SLICE_X1Y106_CO6;
  assign CLBLL_L_X2Y106_SLICE_X0Y106_A4 = LIOB33_X0Y101_IOB_X0Y102_I;
  assign CLBLL_L_X2Y106_SLICE_X0Y106_A5 = 1'b1;
  assign CLBLL_L_X2Y106_SLICE_X0Y106_A6 = 1'b1;
  assign CLBLL_L_X2Y106_SLICE_X0Y106_B1 = RIOB33_X105Y105_IOB_X1Y106_I;
  assign CLBLL_L_X2Y106_SLICE_X0Y106_B2 = CLBLL_L_X2Y106_SLICE_X1Y106_DO6;
  assign CLBLL_L_X2Y106_SLICE_X0Y106_B3 = LIOB33_X0Y103_IOB_X0Y104_I;
  assign CLBLL_L_X2Y106_SLICE_X0Y106_B4 = CLBLL_L_X2Y104_SLICE_X1Y104_CO6;
  assign CLBLL_L_X2Y106_SLICE_X0Y106_B5 = RIOB33_SING_X105Y100_IOB_X1Y100_I;
  assign CLBLL_L_X2Y106_SLICE_X0Y106_B6 = LIOB33_X0Y101_IOB_X0Y102_I;
  assign CLBLL_L_X2Y106_SLICE_X0Y106_C1 = 1'b1;
  assign CLBLL_L_X2Y106_SLICE_X0Y106_C2 = 1'b1;
  assign CLBLL_L_X2Y106_SLICE_X0Y106_C3 = 1'b1;
  assign CLBLL_L_X2Y106_SLICE_X0Y106_C4 = 1'b1;
  assign CLBLL_L_X2Y106_SLICE_X0Y106_C5 = 1'b1;
  assign CLBLL_L_X2Y106_SLICE_X0Y106_C6 = 1'b1;
  assign CLBLL_L_X2Y106_SLICE_X0Y106_D1 = 1'b1;
  assign CLBLL_L_X2Y106_SLICE_X0Y106_D2 = 1'b1;
  assign CLBLL_L_X2Y106_SLICE_X0Y106_D3 = 1'b1;
  assign CLBLL_L_X2Y106_SLICE_X0Y106_D4 = 1'b1;
  assign CLBLL_L_X2Y106_SLICE_X0Y106_D5 = 1'b1;
  assign CLBLL_L_X2Y106_SLICE_X0Y106_D6 = 1'b1;
  assign CLBLL_L_X2Y106_SLICE_X1Y106_A1 = RIOB33_SING_X105Y100_IOB_X1Y100_I;
  assign CLBLL_L_X2Y106_SLICE_X1Y106_A2 = CLBLM_R_X3Y106_SLICE_X2Y106_CO6;
  assign CLBLL_L_X2Y106_SLICE_X1Y106_A3 = LIOB33_X0Y101_IOB_X0Y101_I;
  assign CLBLM_R_X7Y108_SLICE_X9Y108_A4 = CLBLM_R_X7Y106_SLICE_X9Y106_CO6;
  assign CLBLM_R_X7Y108_SLICE_X9Y108_A5 = LIOB33_X0Y115_IOB_X0Y116_I;
  assign CLBLM_R_X7Y108_SLICE_X9Y108_A6 = LIOB33_X0Y107_IOB_X0Y107_I;
  assign CLBLL_L_X2Y106_SLICE_X1Y106_A4 = CLBLL_L_X2Y106_SLICE_X1Y106_BO6;
  assign CLBLL_L_X2Y106_SLICE_X1Y106_A5 = 1'b1;
  assign CLBLL_L_X2Y106_SLICE_X1Y106_A6 = 1'b1;
  assign CLBLM_R_X7Y108_SLICE_X9Y108_A1 = LIOB33_X0Y107_IOB_X0Y108_I;
  assign CLBLM_R_X7Y108_SLICE_X9Y108_A2 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLM_R_X7Y108_SLICE_X9Y108_B3 = LIOB33_X0Y109_IOB_X0Y110_I;
  assign CLBLM_R_X7Y108_SLICE_X9Y108_B4 = LIOB33_X0Y115_IOB_X0Y116_I;
  assign CLBLM_R_X7Y108_SLICE_X9Y108_B5 = CLBLM_L_X8Y108_SLICE_X10Y108_BO6;
  assign CLBLM_R_X7Y108_SLICE_X9Y108_B6 = LIOB33_X0Y109_IOB_X0Y109_I;
  assign CLBLL_L_X2Y106_SLICE_X1Y106_B1 = RIOB33_X105Y105_IOB_X1Y106_I;
  assign CLBLL_L_X2Y106_SLICE_X1Y106_B2 = RIOB33_X105Y111_IOB_X1Y112_I;
  assign CLBLL_L_X2Y106_SLICE_X1Y106_B3 = LIOB33_SING_X0Y100_IOB_X0Y100_I;
  assign CLBLL_L_X2Y106_SLICE_X1Y106_B4 = LIOB33_X0Y103_IOB_X0Y103_I;
  assign CLBLL_L_X2Y106_SLICE_X1Y106_B5 = RIOB33_X105Y113_IOB_X1Y113_I;
  assign CLBLM_R_X7Y108_SLICE_X9Y108_C3 = CLBLM_L_X8Y107_SLICE_X11Y107_CO6;
  assign CLBLM_R_X7Y108_SLICE_X9Y108_C4 = LIOB33_X0Y109_IOB_X0Y110_I;
  assign CLBLM_R_X7Y108_SLICE_X9Y108_C5 = CLBLM_R_X7Y108_SLICE_X9Y108_AO6;
  assign CLBLL_L_X2Y106_SLICE_X1Y106_C1 = LIOB33_X0Y101_IOB_X0Y101_I;
  assign CLBLL_L_X2Y106_SLICE_X1Y106_C2 = CLBLM_R_X3Y106_SLICE_X2Y106_CO6;
  assign CLBLL_L_X2Y106_SLICE_X1Y106_C3 = RIOB33_X105Y105_IOB_X1Y106_I;
  assign CLBLL_L_X2Y106_SLICE_X1Y106_C4 = RIOB33_SING_X105Y100_IOB_X1Y100_I;
  assign CLBLL_L_X2Y106_SLICE_X1Y106_C5 = CLBLL_L_X2Y104_SLICE_X0Y104_BO6;
  assign CLBLL_L_X2Y106_SLICE_X1Y106_C6 = CLBLL_L_X2Y106_SLICE_X1Y106_BO6;
  assign CLBLM_L_X8Y107_SLICE_X11Y107_D2 = CLBLM_L_X10Y106_SLICE_X12Y106_AO6;
  assign CLBLM_L_X8Y107_SLICE_X11Y107_D3 = CLBLM_L_X10Y107_SLICE_X12Y107_AO6;
  assign CLBLL_L_X2Y106_SLICE_X1Y106_D1 = CLBLL_L_X2Y106_SLICE_X1Y106_AO6;
  assign CLBLL_L_X2Y106_SLICE_X1Y106_D2 = CLBLM_R_X13Y106_SLICE_X18Y106_AO5;
  assign CLBLL_L_X2Y106_SLICE_X1Y106_D3 = CLBLM_R_X3Y106_SLICE_X2Y106_CO6;
  assign CLBLL_L_X2Y106_SLICE_X1Y106_D4 = CLBLL_L_X2Y104_SLICE_X0Y104_BO6;
  assign CLBLL_L_X2Y106_SLICE_X1Y106_D5 = CLBLL_L_X2Y106_SLICE_X0Y106_AO6;
  assign CLBLL_L_X2Y106_SLICE_X1Y106_D6 = CLBLL_L_X2Y106_SLICE_X1Y106_BO6;
  assign CLBLM_R_X7Y108_SLICE_X9Y108_D1 = CLBLM_L_X8Y108_SLICE_X10Y108_BO6;
  assign CLBLM_R_X7Y108_SLICE_X9Y108_D2 = CLBLM_L_X8Y107_SLICE_X10Y107_CO6;
  assign CLBLM_R_X7Y108_SLICE_X9Y108_D3 = LIOB33_X0Y115_IOB_X0Y116_I;
  assign CLBLM_R_X7Y108_SLICE_X9Y108_D4 = LIOB33_X0Y109_IOB_X0Y109_I;
  assign CLBLM_L_X8Y107_SLICE_X11Y107_D6 = CLBLM_L_X8Y107_SLICE_X11Y107_BO6;
  assign CLBLM_R_X7Y108_SLICE_X8Y108_A1 = 1'b1;
  assign CLBLM_R_X7Y108_SLICE_X8Y108_A2 = 1'b1;
  assign CLBLM_R_X7Y108_SLICE_X8Y108_A3 = LIOB33_X0Y115_IOB_X0Y116_I;
  assign CLBLM_R_X7Y108_SLICE_X8Y108_A4 = LIOB33_X0Y111_IOB_X0Y111_I;
  assign CLBLM_R_X7Y108_SLICE_X8Y108_A5 = LIOB33_X0Y113_IOB_X0Y114_I;
  assign CLBLM_R_X7Y108_SLICE_X8Y108_A6 = 1'b1;
  assign CLBLM_R_X7Y108_SLICE_X8Y108_B1 = CLBLM_R_X7Y107_SLICE_X9Y107_DO6;
  assign CLBLM_R_X7Y108_SLICE_X8Y108_B2 = CLBLM_R_X7Y108_SLICE_X9Y108_BO6;
  assign CLBLM_R_X7Y108_SLICE_X8Y108_B3 = CLBLM_R_X7Y109_SLICE_X8Y109_AO6;
  assign CLBLM_R_X7Y108_SLICE_X8Y108_B4 = CLBLM_L_X8Y108_SLICE_X10Y108_CO6;
  assign CLBLM_R_X7Y108_SLICE_X8Y108_B5 = CLBLM_R_X7Y108_SLICE_X8Y108_AO6;
  assign CLBLM_R_X7Y108_SLICE_X8Y108_B6 = CLBLM_R_X7Y108_SLICE_X8Y108_AO5;
  assign CLBLM_R_X7Y108_SLICE_X8Y108_C1 = CLBLM_R_X7Y108_SLICE_X8Y108_AO6;
  assign CLBLM_R_X7Y108_SLICE_X8Y108_C2 = CLBLM_R_X7Y108_SLICE_X9Y108_CO6;
  assign CLBLM_R_X7Y108_SLICE_X8Y108_C3 = CLBLM_R_X7Y108_SLICE_X9Y108_BO6;
  assign CLBLM_R_X7Y108_SLICE_X8Y108_C4 = CLBLM_R_X7Y108_SLICE_X8Y108_AO5;
  assign CLBLM_R_X7Y108_SLICE_X8Y108_C5 = CLBLM_L_X8Y108_SLICE_X11Y108_BO6;
  assign CLBLM_R_X7Y108_SLICE_X8Y108_C6 = CLBLM_R_X7Y107_SLICE_X9Y107_DO6;
  assign CLBLM_R_X7Y108_SLICE_X8Y108_D1 = 1'b1;
  assign CLBLM_R_X7Y108_SLICE_X8Y108_D2 = 1'b1;
  assign CLBLM_R_X7Y108_SLICE_X8Y108_D3 = 1'b1;
  assign CLBLM_R_X7Y108_SLICE_X8Y108_D4 = 1'b1;
  assign CLBLM_R_X7Y108_SLICE_X8Y108_D5 = 1'b1;
  assign CLBLM_R_X7Y108_SLICE_X8Y108_D6 = 1'b1;
  assign LIOI3_X0Y121_OLOGIC_X0Y122_D1 = CLBLL_L_X2Y104_SLICE_X0Y104_AO6;
  assign LIOI3_X0Y121_OLOGIC_X0Y122_T1 = 1'b1;
  assign LIOI3_X0Y121_OLOGIC_X0Y121_D1 = CLBLL_L_X2Y106_SLICE_X0Y106_AO5;
  assign LIOI3_X0Y121_OLOGIC_X0Y121_T1 = 1'b1;
  assign CLBLM_L_X8Y107_SLICE_X10Y107_B4 = CLBLM_R_X5Y107_SLICE_X7Y107_AO5;
  assign CLBLL_L_X2Y107_SLICE_X0Y107_A1 = RIOB33_X105Y105_IOB_X1Y106_I;
  assign CLBLL_L_X2Y107_SLICE_X0Y107_A2 = CLBLL_L_X2Y106_SLICE_X0Y106_BO6;
  assign CLBLL_L_X2Y107_SLICE_X0Y107_A3 = LIOB33_X0Y103_IOB_X0Y104_I;
  assign CLBLL_L_X2Y107_SLICE_X0Y107_A4 = RIOB33_SING_X105Y100_IOB_X1Y100_I;
  assign CLBLL_L_X2Y107_SLICE_X0Y107_A5 = LIOB33_X0Y105_IOB_X0Y105_I;
  assign CLBLL_L_X2Y107_SLICE_X0Y107_A6 = CLBLL_L_X2Y104_SLICE_X1Y104_DO6;
  assign CLBLL_L_X2Y107_SLICE_X0Y107_B1 = CLBLL_L_X2Y106_SLICE_X0Y106_BO6;
  assign CLBLL_L_X2Y107_SLICE_X0Y107_B2 = RIOB33_SING_X105Y100_IOB_X1Y100_I;
  assign CLBLL_L_X2Y107_SLICE_X0Y107_B3 = LIOB33_X0Y105_IOB_X0Y105_I;
  assign CLBLL_L_X2Y107_SLICE_X0Y107_B4 = CLBLL_L_X2Y104_SLICE_X1Y104_DO6;
  assign CLBLL_L_X2Y107_SLICE_X0Y107_B5 = LIOB33_X0Y103_IOB_X0Y104_I;
  assign CLBLL_L_X2Y107_SLICE_X0Y107_B6 = RIOB33_X105Y105_IOB_X1Y106_I;
  assign CLBLL_L_X2Y107_SLICE_X0Y107_C1 = 1'b1;
  assign CLBLL_L_X2Y107_SLICE_X0Y107_C2 = 1'b1;
  assign CLBLL_L_X2Y107_SLICE_X0Y107_C3 = 1'b1;
  assign CLBLL_L_X2Y107_SLICE_X0Y107_C4 = 1'b1;
  assign CLBLL_L_X2Y107_SLICE_X0Y107_C5 = 1'b1;
  assign CLBLL_L_X2Y107_SLICE_X0Y107_C6 = 1'b1;
  assign CLBLL_L_X2Y107_SLICE_X0Y107_D1 = 1'b1;
  assign CLBLL_L_X2Y107_SLICE_X0Y107_D2 = 1'b1;
  assign CLBLL_L_X2Y107_SLICE_X0Y107_D3 = 1'b1;
  assign CLBLL_L_X2Y107_SLICE_X0Y107_D4 = 1'b1;
  assign CLBLL_L_X2Y107_SLICE_X0Y107_D5 = 1'b1;
  assign CLBLL_L_X2Y107_SLICE_X0Y107_D6 = 1'b1;
  assign CLBLL_L_X2Y107_SLICE_X1Y107_A1 = 1'b1;
  assign CLBLL_L_X2Y107_SLICE_X1Y107_A2 = 1'b1;
  assign CLBLL_L_X2Y107_SLICE_X1Y107_A3 = 1'b1;
  assign CLBLL_L_X2Y107_SLICE_X1Y107_A4 = 1'b1;
  assign CLBLL_L_X2Y107_SLICE_X1Y107_A5 = 1'b1;
  assign CLBLL_L_X2Y107_SLICE_X1Y107_A6 = 1'b1;
  assign CLBLM_R_X7Y109_SLICE_X9Y109_A1 = LIOB33_X0Y107_IOB_X0Y107_I;
  assign CLBLM_R_X7Y109_SLICE_X9Y109_A2 = CLBLM_L_X10Y109_SLICE_X12Y109_CO6;
  assign CLBLM_R_X7Y109_SLICE_X9Y109_A3 = RIOB33_SING_X105Y100_IOB_X1Y100_I;
  assign CLBLL_L_X2Y107_SLICE_X1Y107_B1 = 1'b1;
  assign CLBLL_L_X2Y107_SLICE_X1Y107_B2 = 1'b1;
  assign CLBLL_L_X2Y107_SLICE_X1Y107_B3 = 1'b1;
  assign CLBLL_L_X2Y107_SLICE_X1Y107_B4 = 1'b1;
  assign CLBLM_R_X7Y109_SLICE_X9Y109_B1 = CLBLM_L_X8Y109_SLICE_X10Y109_AO6;
  assign CLBLM_R_X7Y109_SLICE_X9Y109_B2 = RIOB33_X105Y109_IOB_X1Y110_I;
  assign CLBLM_R_X7Y109_SLICE_X9Y109_B3 = LIOB33_X0Y109_IOB_X0Y110_I;
  assign CLBLM_R_X7Y109_SLICE_X9Y109_B4 = LIOB33_X0Y109_IOB_X0Y109_I;
  assign CLBLM_R_X7Y109_SLICE_X9Y109_B5 = RIOB33_X105Y109_IOB_X1Y109_I;
  assign CLBLM_R_X7Y109_SLICE_X9Y109_B6 = CLBLM_R_X7Y109_SLICE_X9Y109_CO6;
  assign CLBLL_L_X2Y107_SLICE_X1Y107_B5 = 1'b1;
  assign CLBLL_L_X2Y107_SLICE_X1Y107_B6 = 1'b1;
  assign CLBLL_L_X2Y107_SLICE_X1Y107_C1 = 1'b1;
  assign CLBLL_L_X2Y107_SLICE_X1Y107_C2 = 1'b1;
  assign CLBLL_L_X2Y107_SLICE_X1Y107_C3 = 1'b1;
  assign CLBLL_L_X2Y107_SLICE_X1Y107_C4 = 1'b1;
  assign CLBLL_L_X2Y107_SLICE_X1Y107_C5 = 1'b1;
  assign CLBLL_L_X2Y107_SLICE_X1Y107_C6 = 1'b1;
  assign CLBLM_R_X7Y109_SLICE_X9Y109_C1 = RIOB33_X105Y111_IOB_X1Y111_I;
  assign CLBLM_R_X7Y109_SLICE_X9Y109_C2 = LIOB33_X0Y107_IOB_X0Y108_I;
  assign CLBLM_R_X7Y109_SLICE_X9Y109_C3 = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLM_R_X7Y109_SLICE_X9Y109_C4 = CLBLM_L_X10Y109_SLICE_X12Y109_DO6;
  assign CLBLM_R_X7Y109_SLICE_X9Y109_C5 = LIOB33_X0Y107_IOB_X0Y107_I;
  assign CLBLM_R_X7Y109_SLICE_X9Y109_C6 = RIOB33_X105Y109_IOB_X1Y110_I;
  assign CLBLL_L_X2Y107_SLICE_X1Y107_D1 = 1'b1;
  assign CLBLL_L_X2Y107_SLICE_X1Y107_D2 = 1'b1;
  assign CLBLL_L_X2Y107_SLICE_X1Y107_D3 = 1'b1;
  assign CLBLL_L_X2Y107_SLICE_X1Y107_D4 = 1'b1;
  assign CLBLL_L_X2Y107_SLICE_X1Y107_D5 = 1'b1;
  assign CLBLL_L_X2Y107_SLICE_X1Y107_D6 = 1'b1;
  assign CLBLM_R_X7Y109_SLICE_X9Y109_D1 = LIOB33_X0Y109_IOB_X0Y110_I;
  assign CLBLM_R_X7Y109_SLICE_X9Y109_D2 = RIOB33_X105Y109_IOB_X1Y109_I;
  assign CLBLM_R_X7Y109_SLICE_X9Y109_D3 = LIOB33_X0Y109_IOB_X0Y109_I;
  assign CLBLM_R_X7Y109_SLICE_X9Y109_D4 = CLBLM_R_X7Y109_SLICE_X9Y109_CO6;
  assign CLBLM_R_X7Y109_SLICE_X9Y109_D5 = CLBLM_L_X8Y109_SLICE_X10Y109_AO6;
  assign CLBLM_R_X7Y109_SLICE_X9Y109_D6 = RIOB33_X105Y109_IOB_X1Y110_I;
  assign CLBLM_R_X7Y109_SLICE_X8Y109_A1 = 1'b1;
  assign CLBLM_R_X7Y109_SLICE_X8Y109_A2 = 1'b1;
  assign CLBLM_R_X7Y109_SLICE_X8Y109_A3 = LIOB33_X0Y115_IOB_X0Y116_I;
  assign CLBLM_R_X7Y109_SLICE_X8Y109_A4 = LIOB33_X0Y111_IOB_X0Y112_I;
  assign CLBLM_R_X7Y109_SLICE_X8Y109_A5 = LIOB33_X0Y113_IOB_X0Y114_I;
  assign CLBLM_R_X7Y109_SLICE_X8Y109_A6 = 1'b1;
  assign CLBLM_R_X7Y109_SLICE_X8Y109_B1 = CLBLM_L_X8Y110_SLICE_X11Y110_BO6;
  assign CLBLM_R_X7Y109_SLICE_X8Y109_B2 = CLBLM_L_X8Y108_SLICE_X11Y108_BO6;
  assign CLBLM_R_X7Y109_SLICE_X8Y109_B3 = CLBLM_L_X8Y110_SLICE_X11Y110_AO6;
  assign CLBLM_R_X7Y109_SLICE_X8Y109_B4 = CLBLM_R_X7Y108_SLICE_X9Y108_CO6;
  assign CLBLM_R_X7Y109_SLICE_X8Y109_B5 = CLBLM_L_X8Y108_SLICE_X11Y108_AO6;
  assign CLBLM_R_X7Y109_SLICE_X8Y109_B6 = CLBLM_R_X7Y108_SLICE_X8Y108_AO5;
  assign CLBLM_R_X7Y109_SLICE_X8Y109_C1 = LIOB33_X0Y111_IOB_X0Y111_I;
  assign CLBLM_R_X7Y109_SLICE_X8Y109_C2 = LIOB33_X0Y115_IOB_X0Y116_I;
  assign CLBLM_R_X7Y109_SLICE_X8Y109_C3 = CLBLM_R_X7Y108_SLICE_X9Y108_CO6;
  assign CLBLM_R_X7Y109_SLICE_X8Y109_C4 = CLBLM_L_X8Y108_SLICE_X11Y108_CO6;
  assign CLBLM_R_X7Y109_SLICE_X8Y109_C5 = LIOB33_X0Y109_IOB_X0Y110_I;
  assign CLBLM_R_X7Y109_SLICE_X8Y109_C6 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLM_R_X7Y109_SLICE_X8Y109_D1 = CLBLM_L_X8Y108_SLICE_X10Y108_DO6;
  assign CLBLM_R_X7Y109_SLICE_X8Y109_D2 = CLBLM_R_X7Y108_SLICE_X8Y108_AO5;
  assign CLBLM_R_X7Y109_SLICE_X8Y109_D3 = CLBLM_R_X7Y108_SLICE_X9Y108_CO6;
  assign CLBLM_R_X7Y109_SLICE_X8Y109_D4 = CLBLM_R_X7Y109_SLICE_X8Y109_AO5;
  assign CLBLM_R_X7Y109_SLICE_X8Y109_D5 = CLBLM_L_X8Y110_SLICE_X11Y110_AO6;
  assign CLBLM_R_X7Y109_SLICE_X8Y109_D6 = CLBLM_L_X8Y108_SLICE_X11Y108_BO6;
  assign CLBLM_R_X7Y110_SLICE_X9Y110_A1 = 1'b1;
  assign CLBLM_R_X7Y110_SLICE_X9Y110_A2 = CLBLM_R_X7Y109_SLICE_X9Y109_BO6;
  assign CLBLM_R_X7Y110_SLICE_X9Y110_A3 = LIOB33_X0Y111_IOB_X0Y111_I;
  assign CLBLM_R_X7Y110_SLICE_X9Y110_A4 = RIOB33_X105Y107_IOB_X1Y108_I;
  assign CLBLM_R_X7Y110_SLICE_X9Y110_A5 = CLBLM_R_X7Y110_SLICE_X9Y110_CO6;
  assign CLBLM_R_X7Y110_SLICE_X9Y110_A6 = 1'b1;
  assign CLBLM_R_X7Y110_SLICE_X9Y110_B1 = CLBLM_L_X10Y110_SLICE_X13Y110_DO6;
  assign CLBLM_R_X7Y110_SLICE_X9Y110_B2 = CLBLM_L_X8Y109_SLICE_X10Y109_CO6;
  assign CLBLM_R_X7Y110_SLICE_X9Y110_B3 = LIOB33_X0Y109_IOB_X0Y109_I;
  assign CLBLM_R_X7Y110_SLICE_X9Y110_B4 = RIOB33_X105Y107_IOB_X1Y108_I;
  assign CLBLM_R_X7Y110_SLICE_X9Y110_B5 = CLBLM_L_X8Y109_SLICE_X10Y109_BO6;
  assign CLBLM_R_X7Y110_SLICE_X9Y110_B6 = 1'b1;
  assign CLBLM_R_X7Y110_SLICE_X9Y110_C1 = LIOB33_X0Y109_IOB_X0Y110_I;
  assign CLBLM_R_X7Y110_SLICE_X9Y110_C2 = CLBLM_L_X8Y109_SLICE_X10Y109_CO6;
  assign CLBLM_R_X7Y110_SLICE_X9Y110_C3 = RIOB33_X105Y107_IOB_X1Y108_I;
  assign CLBLM_R_X7Y110_SLICE_X9Y110_C4 = LIOB33_X0Y109_IOB_X0Y109_I;
  assign CLBLM_R_X7Y110_SLICE_X9Y110_C5 = CLBLM_L_X10Y110_SLICE_X13Y110_DO6;
  assign CLBLM_R_X7Y110_SLICE_X9Y110_C6 = CLBLM_L_X8Y109_SLICE_X10Y109_BO6;
  assign CLBLM_R_X7Y110_SLICE_X9Y110_D1 = LIOB33_X0Y109_IOB_X0Y110_I;
  assign CLBLM_R_X7Y110_SLICE_X9Y110_D2 = CLBLM_L_X8Y109_SLICE_X10Y109_CO6;
  assign CLBLM_R_X7Y110_SLICE_X9Y110_D3 = RIOB33_X105Y107_IOB_X1Y108_I;
  assign CLBLM_R_X7Y110_SLICE_X9Y110_D4 = CLBLM_L_X10Y110_SLICE_X13Y110_DO6;
  assign CLBLM_R_X7Y110_SLICE_X9Y110_D5 = LIOB33_X0Y109_IOB_X0Y109_I;
  assign CLBLM_R_X7Y110_SLICE_X9Y110_D6 = CLBLM_L_X8Y109_SLICE_X10Y109_BO6;
  assign CLBLM_R_X7Y110_SLICE_X8Y110_A1 = CLBLM_R_X7Y110_SLICE_X8Y110_BO6;
  assign CLBLM_R_X7Y110_SLICE_X8Y110_A2 = CLBLM_L_X8Y110_SLICE_X10Y110_AO6;
  assign CLBLM_R_X7Y110_SLICE_X8Y110_A3 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLM_R_X7Y110_SLICE_X8Y110_A4 = LIOB33_X0Y115_IOB_X0Y116_I;
  assign CLBLM_R_X7Y110_SLICE_X8Y110_A5 = LIOB33_X0Y111_IOB_X0Y112_I;
  assign CLBLM_R_X7Y110_SLICE_X8Y110_A6 = CLBLM_L_X8Y111_SLICE_X10Y111_BO6;
  assign CLBLM_R_X7Y110_SLICE_X8Y110_B1 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLM_R_X7Y110_SLICE_X8Y110_B2 = LIOB33_X0Y115_IOB_X0Y116_I;
  assign CLBLM_R_X7Y110_SLICE_X8Y110_B3 = CLBLM_L_X8Y108_SLICE_X11Y108_CO6;
  assign CLBLM_R_X7Y110_SLICE_X8Y110_B4 = LIOB33_X0Y109_IOB_X0Y110_I;
  assign CLBLM_R_X7Y110_SLICE_X8Y110_B5 = LIOB33_X0Y111_IOB_X0Y111_I;
  assign CLBLM_R_X7Y110_SLICE_X8Y110_B6 = CLBLM_R_X7Y108_SLICE_X9Y108_CO6;
  assign CLBLM_R_X7Y110_SLICE_X8Y110_C1 = CLBLM_L_X8Y107_SLICE_X10Y107_DO6;
  assign CLBLM_R_X7Y110_SLICE_X8Y110_C2 = CLBLM_R_X7Y107_SLICE_X8Y107_AO6;
  assign CLBLM_R_X7Y110_SLICE_X8Y110_C3 = CLBLM_R_X7Y110_SLICE_X9Y110_BO6;
  assign CLBLM_R_X7Y110_SLICE_X8Y110_C4 = CLBLM_L_X8Y109_SLICE_X10Y109_CO6;
  assign CLBLM_R_X7Y110_SLICE_X8Y110_C5 = CLBLM_R_X5Y112_SLICE_X7Y112_DO6;
  assign CLBLM_R_X7Y110_SLICE_X8Y110_C6 = CLBLM_R_X7Y106_SLICE_X8Y106_DO6;
  assign CLBLM_R_X7Y110_SLICE_X8Y110_D1 = 1'b1;
  assign CLBLM_R_X7Y110_SLICE_X8Y110_D2 = 1'b1;
  assign CLBLM_R_X7Y110_SLICE_X8Y110_D3 = 1'b1;
  assign CLBLM_R_X7Y110_SLICE_X8Y110_D4 = 1'b1;
  assign CLBLM_R_X7Y110_SLICE_X8Y110_D5 = 1'b1;
  assign CLBLM_R_X7Y110_SLICE_X8Y110_D6 = 1'b1;
  assign LIOI3_X0Y123_OLOGIC_X0Y124_D1 = CLBLM_R_X3Y107_SLICE_X2Y107_AO6;
  assign LIOI3_X0Y123_OLOGIC_X0Y124_T1 = 1'b1;
  assign LIOI3_X0Y123_OLOGIC_X0Y123_D1 = CLBLL_L_X2Y107_SLICE_X0Y107_AO6;
  assign CLBLL_L_X2Y109_SLICE_X0Y109_A1 = RIOB33_X105Y113_IOB_X1Y113_I;
  assign CLBLL_L_X2Y109_SLICE_X0Y109_A2 = RIOB33_X105Y105_IOB_X1Y106_I;
  assign CLBLL_L_X2Y109_SLICE_X0Y109_A3 = RIOB33_X105Y111_IOB_X1Y112_I;
  assign CLBLL_L_X2Y109_SLICE_X0Y109_A4 = RIOB33_SING_X105Y100_IOB_X1Y100_I;
  assign CLBLL_L_X2Y109_SLICE_X0Y109_A5 = LIOB33_SING_X0Y100_IOB_X0Y100_I;
  assign CLBLL_L_X2Y109_SLICE_X0Y109_A6 = 1'b1;
  assign LIOI3_X0Y123_OLOGIC_X0Y123_T1 = 1'b1;
  assign CLBLL_L_X2Y109_SLICE_X0Y109_B1 = 1'b1;
  assign CLBLL_L_X2Y109_SLICE_X0Y109_B2 = 1'b1;
  assign CLBLL_L_X2Y109_SLICE_X0Y109_B3 = 1'b1;
  assign CLBLL_L_X2Y109_SLICE_X0Y109_B4 = 1'b1;
  assign CLBLL_L_X2Y109_SLICE_X0Y109_B5 = 1'b1;
  assign CLBLL_L_X2Y109_SLICE_X0Y109_B6 = 1'b1;
  assign CLBLL_L_X2Y109_SLICE_X0Y109_C1 = 1'b1;
  assign CLBLL_L_X2Y109_SLICE_X0Y109_C2 = 1'b1;
  assign CLBLL_L_X2Y109_SLICE_X0Y109_C3 = 1'b1;
  assign CLBLL_L_X2Y109_SLICE_X0Y109_C4 = 1'b1;
  assign CLBLL_L_X2Y109_SLICE_X0Y109_C5 = 1'b1;
  assign CLBLL_L_X2Y109_SLICE_X0Y109_C6 = 1'b1;
  assign CLBLL_L_X2Y109_SLICE_X0Y109_D1 = 1'b1;
  assign CLBLL_L_X2Y109_SLICE_X0Y109_D2 = 1'b1;
  assign CLBLL_L_X2Y109_SLICE_X0Y109_D3 = 1'b1;
  assign CLBLL_L_X2Y109_SLICE_X0Y109_D4 = 1'b1;
  assign CLBLL_L_X2Y109_SLICE_X0Y109_D5 = 1'b1;
  assign CLBLL_L_X2Y109_SLICE_X0Y109_D6 = 1'b1;
  assign CLBLL_L_X2Y109_SLICE_X1Y109_A1 = 1'b1;
  assign CLBLL_L_X2Y109_SLICE_X1Y109_A2 = 1'b1;
  assign CLBLL_L_X2Y109_SLICE_X1Y109_A3 = 1'b1;
  assign CLBLL_L_X2Y109_SLICE_X1Y109_A4 = 1'b1;
  assign CLBLL_L_X2Y109_SLICE_X1Y109_A5 = 1'b1;
  assign CLBLL_L_X2Y109_SLICE_X1Y109_A6 = 1'b1;
  assign CLBLL_L_X2Y109_SLICE_X1Y109_B1 = 1'b1;
  assign CLBLL_L_X2Y109_SLICE_X1Y109_B2 = 1'b1;
  assign CLBLL_L_X2Y109_SLICE_X1Y109_B3 = 1'b1;
  assign CLBLL_L_X2Y109_SLICE_X1Y109_B4 = 1'b1;
  assign CLBLL_L_X2Y109_SLICE_X1Y109_B5 = 1'b1;
  assign CLBLL_L_X2Y109_SLICE_X1Y109_B6 = 1'b1;
  assign CLBLM_R_X7Y111_SLICE_X9Y111_A1 = 1'b1;
  assign CLBLM_R_X7Y111_SLICE_X9Y111_A2 = RIOB33_X105Y109_IOB_X1Y109_I;
  assign CLBLM_R_X7Y111_SLICE_X9Y111_A3 = LIOB33_X0Y111_IOB_X0Y111_I;
  assign CLBLL_L_X2Y109_SLICE_X1Y109_C1 = 1'b1;
  assign CLBLL_L_X2Y109_SLICE_X1Y109_C2 = 1'b1;
  assign CLBLL_L_X2Y109_SLICE_X1Y109_C3 = 1'b1;
  assign CLBLL_L_X2Y109_SLICE_X1Y109_C4 = 1'b1;
  assign CLBLL_L_X2Y109_SLICE_X1Y109_C5 = 1'b1;
  assign CLBLL_L_X2Y109_SLICE_X1Y109_C6 = 1'b1;
  assign CLBLM_R_X7Y111_SLICE_X9Y111_A4 = CLBLM_R_X7Y111_SLICE_X9Y111_BO6;
  assign CLBLM_R_X7Y111_SLICE_X9Y111_A5 = CLBLM_R_X7Y109_SLICE_X9Y109_DO6;
  assign CLBLM_R_X7Y111_SLICE_X9Y111_A6 = 1'b1;
  assign CLBLM_R_X7Y111_SLICE_X9Y111_B5 = LIOB33_X0Y109_IOB_X0Y109_I;
  assign CLBLM_R_X7Y111_SLICE_X9Y111_B6 = CLBLM_R_X7Y111_SLICE_X9Y111_CO6;
  assign CLBLM_R_X7Y111_SLICE_X9Y111_B1 = RIOB33_X105Y111_IOB_X1Y111_I;
  assign CLBLM_R_X7Y111_SLICE_X9Y111_B2 = RIOB33_X105Y109_IOB_X1Y110_I;
  assign CLBLM_R_X7Y111_SLICE_X9Y111_B3 = LIOB33_X0Y109_IOB_X0Y110_I;
  assign CLBLM_R_X7Y111_SLICE_X9Y111_B4 = LIOB33_X0Y107_IOB_X0Y108_I;
  assign CLBLL_L_X2Y109_SLICE_X1Y109_D1 = 1'b1;
  assign CLBLL_L_X2Y109_SLICE_X1Y109_D2 = 1'b1;
  assign CLBLL_L_X2Y109_SLICE_X1Y109_D3 = 1'b1;
  assign CLBLL_L_X2Y109_SLICE_X1Y109_D4 = 1'b1;
  assign CLBLL_L_X2Y109_SLICE_X1Y109_D5 = 1'b1;
  assign CLBLL_L_X2Y109_SLICE_X1Y109_D6 = 1'b1;
  assign CLBLM_R_X7Y111_SLICE_X9Y111_C1 = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLM_R_X7Y111_SLICE_X9Y111_C2 = LIOB33_X0Y107_IOB_X0Y108_I;
  assign CLBLM_R_X7Y111_SLICE_X9Y111_C3 = CLBLM_L_X10Y109_SLICE_X12Y109_DO6;
  assign CLBLM_R_X7Y111_SLICE_X9Y111_C4 = RIOB33_X105Y109_IOB_X1Y110_I;
  assign CLBLM_R_X7Y111_SLICE_X9Y111_C5 = RIOB33_X105Y111_IOB_X1Y111_I;
  assign CLBLM_R_X7Y111_SLICE_X9Y111_D1 = 1'b1;
  assign CLBLM_R_X7Y111_SLICE_X9Y111_D2 = 1'b1;
  assign CLBLM_R_X7Y111_SLICE_X9Y111_D3 = 1'b1;
  assign CLBLM_R_X7Y111_SLICE_X9Y111_D4 = 1'b1;
  assign CLBLM_R_X7Y111_SLICE_X9Y111_D5 = 1'b1;
  assign CLBLM_R_X7Y111_SLICE_X9Y111_D6 = 1'b1;
  assign CLBLM_R_X7Y111_SLICE_X8Y111_A1 = CLBLM_L_X8Y111_SLICE_X10Y111_AO5;
  assign CLBLM_R_X7Y111_SLICE_X8Y111_A2 = CLBLM_L_X8Y111_SLICE_X10Y111_AO6;
  assign CLBLM_R_X7Y111_SLICE_X8Y111_A3 = RIOB33_X105Y103_IOB_X1Y103_I;
  assign CLBLM_R_X7Y111_SLICE_X8Y111_A4 = CLBLM_L_X10Y111_SLICE_X12Y111_CO6;
  assign CLBLM_R_X7Y111_SLICE_X8Y111_A5 = LIOB33_X0Y111_IOB_X0Y111_I;
  assign CLBLM_R_X7Y111_SLICE_X8Y111_A6 = 1'b1;
  assign CLBLM_R_X7Y111_SLICE_X8Y111_B1 = RIOB33_X105Y103_IOB_X1Y103_I;
  assign CLBLM_R_X7Y111_SLICE_X8Y111_B2 = CLBLM_L_X8Y111_SLICE_X10Y111_AO6;
  assign CLBLM_R_X7Y111_SLICE_X8Y111_B3 = LIOB33_X0Y111_IOB_X0Y111_I;
  assign CLBLM_R_X7Y111_SLICE_X8Y111_B4 = CLBLM_L_X10Y111_SLICE_X12Y111_CO6;
  assign CLBLM_R_X7Y111_SLICE_X8Y111_B5 = RIOB33_X105Y103_IOB_X1Y104_I;
  assign CLBLM_R_X7Y111_SLICE_X8Y111_B6 = CLBLM_L_X8Y111_SLICE_X11Y111_BO6;
  assign CLBLM_R_X7Y111_SLICE_X8Y111_C1 = 1'b1;
  assign CLBLM_R_X7Y111_SLICE_X8Y111_C2 = 1'b1;
  assign CLBLM_R_X7Y111_SLICE_X8Y111_C3 = 1'b1;
  assign CLBLM_R_X7Y111_SLICE_X8Y111_C4 = 1'b1;
  assign CLBLM_R_X7Y111_SLICE_X8Y111_C5 = 1'b1;
  assign CLBLM_R_X7Y111_SLICE_X8Y111_C6 = 1'b1;
  assign CLBLM_R_X7Y111_SLICE_X8Y111_D1 = 1'b1;
  assign CLBLM_R_X7Y111_SLICE_X8Y111_D2 = 1'b1;
  assign CLBLM_R_X7Y111_SLICE_X8Y111_D3 = 1'b1;
  assign CLBLM_R_X7Y111_SLICE_X8Y111_D4 = 1'b1;
  assign CLBLM_R_X7Y111_SLICE_X8Y111_D5 = 1'b1;
  assign CLBLM_R_X7Y111_SLICE_X8Y111_D6 = 1'b1;
  assign RIOI3_X105Y105_ILOGIC_X1Y106_D = RIOB33_X105Y105_IOB_X1Y106_I;
  assign RIOI3_X105Y105_ILOGIC_X1Y105_D = RIOB33_X105Y105_IOB_X1Y105_I;
  assign LIOI3_TBYTESRC_X0Y107_ILOGIC_X0Y108_D = LIOB33_X0Y107_IOB_X0Y108_I;
  assign LIOI3_TBYTESRC_X0Y107_ILOGIC_X0Y107_D = LIOB33_X0Y107_IOB_X0Y107_I;
  assign RIOI3_TBYTETERM_X105Y113_ILOGIC_X1Y113_D = RIOB33_X105Y113_IOB_X1Y113_I;
  assign CLBLL_L_X2Y110_SLICE_X0Y110_A1 = 1'b1;
  assign CLBLL_L_X2Y110_SLICE_X0Y110_A2 = RIOB33_X105Y111_IOB_X1Y112_I;
  assign CLBLL_L_X2Y110_SLICE_X0Y110_A3 = LIOB33_X0Y113_IOB_X0Y113_I;
  assign CLBLL_L_X2Y110_SLICE_X0Y110_A4 = CLBLL_L_X4Y108_SLICE_X4Y108_CO6;
  assign CLBLL_L_X2Y110_SLICE_X0Y110_A5 = RIOB33_SING_X105Y100_IOB_X1Y100_I;
  assign CLBLL_L_X2Y110_SLICE_X0Y110_A6 = 1'b1;
  assign CLBLL_L_X2Y110_SLICE_X0Y110_B1 = 1'b1;
  assign CLBLL_L_X2Y110_SLICE_X0Y110_B2 = 1'b1;
  assign CLBLL_L_X2Y110_SLICE_X0Y110_B3 = 1'b1;
  assign CLBLL_L_X2Y110_SLICE_X0Y110_B4 = 1'b1;
  assign CLBLL_L_X2Y110_SLICE_X0Y110_B5 = 1'b1;
  assign CLBLL_L_X2Y110_SLICE_X0Y110_B6 = 1'b1;
  assign RIOI3_SING_X105Y100_ILOGIC_X1Y100_D = RIOB33_SING_X105Y100_IOB_X1Y100_I;
  assign CLBLL_L_X2Y110_SLICE_X0Y110_C1 = 1'b1;
  assign CLBLL_L_X2Y110_SLICE_X0Y110_C2 = 1'b1;
  assign CLBLL_L_X2Y110_SLICE_X0Y110_C3 = 1'b1;
  assign CLBLL_L_X2Y110_SLICE_X0Y110_C4 = 1'b1;
  assign CLBLL_L_X2Y110_SLICE_X0Y110_C5 = 1'b1;
  assign CLBLL_L_X2Y110_SLICE_X0Y110_C6 = 1'b1;
  assign CLBLL_L_X2Y110_SLICE_X0Y110_D1 = 1'b1;
  assign CLBLL_L_X2Y110_SLICE_X0Y110_D2 = 1'b1;
  assign CLBLL_L_X2Y110_SLICE_X0Y110_D3 = 1'b1;
  assign CLBLL_L_X2Y110_SLICE_X0Y110_D4 = 1'b1;
  assign CLBLL_L_X2Y110_SLICE_X0Y110_D5 = 1'b1;
  assign CLBLL_L_X2Y110_SLICE_X0Y110_D6 = 1'b1;
  assign CLBLL_L_X2Y110_SLICE_X1Y110_A1 = 1'b1;
  assign CLBLL_L_X2Y110_SLICE_X1Y110_A2 = 1'b1;
  assign CLBLL_L_X2Y110_SLICE_X1Y110_A3 = 1'b1;
  assign CLBLL_L_X2Y110_SLICE_X1Y110_A4 = 1'b1;
  assign CLBLL_L_X2Y110_SLICE_X1Y110_A5 = 1'b1;
  assign CLBLL_L_X2Y110_SLICE_X1Y110_A6 = 1'b1;
  assign CLBLL_L_X2Y110_SLICE_X1Y110_B1 = 1'b1;
  assign CLBLL_L_X2Y110_SLICE_X1Y110_B2 = 1'b1;
  assign CLBLL_L_X2Y110_SLICE_X1Y110_B3 = 1'b1;
  assign CLBLL_L_X2Y110_SLICE_X1Y110_B4 = 1'b1;
  assign CLBLL_L_X2Y110_SLICE_X1Y110_B5 = 1'b1;
  assign CLBLL_L_X2Y110_SLICE_X1Y110_B6 = 1'b1;
  assign CLBLL_L_X2Y110_SLICE_X1Y110_C1 = 1'b1;
  assign CLBLL_L_X2Y110_SLICE_X1Y110_C2 = 1'b1;
  assign CLBLL_L_X2Y110_SLICE_X1Y110_C3 = 1'b1;
  assign CLBLL_L_X2Y110_SLICE_X1Y110_C4 = 1'b1;
  assign CLBLL_L_X2Y110_SLICE_X1Y110_C5 = 1'b1;
  assign CLBLL_L_X2Y110_SLICE_X1Y110_C6 = 1'b1;
  assign CLBLM_R_X7Y112_SLICE_X9Y112_A1 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLM_R_X7Y112_SLICE_X9Y112_A2 = CLBLM_L_X8Y112_SLICE_X11Y112_AO6;
  assign CLBLM_R_X7Y112_SLICE_X9Y112_A3 = RIOB33_X105Y101_IOB_X1Y101_I;
  assign CLBLM_R_X7Y112_SLICE_X9Y112_A4 = LIOB33_X0Y111_IOB_X0Y112_I;
  assign CLBLM_R_X7Y112_SLICE_X9Y112_A5 = CLBLM_L_X8Y112_SLICE_X10Y112_BO6;
  assign CLBLM_R_X7Y112_SLICE_X9Y112_B2 = LIOB33_X0Y115_IOB_X0Y116_I;
  assign CLBLM_R_X7Y112_SLICE_X9Y112_A6 = CLBLM_L_X8Y111_SLICE_X10Y111_CO6;
  assign CLBLM_R_X7Y112_SLICE_X9Y112_B5 = CLBLM_R_X7Y110_SLICE_X8Y110_BO6;
  assign CLBLM_R_X7Y112_SLICE_X9Y112_B1 = LIOB33_X0Y113_IOB_X0Y113_I;
  assign CLBLL_L_X2Y110_SLICE_X1Y110_D1 = 1'b1;
  assign CLBLL_L_X2Y110_SLICE_X1Y110_D2 = 1'b1;
  assign CLBLL_L_X2Y110_SLICE_X1Y110_D3 = 1'b1;
  assign CLBLL_L_X2Y110_SLICE_X1Y110_D4 = 1'b1;
  assign CLBLL_L_X2Y110_SLICE_X1Y110_D5 = 1'b1;
  assign CLBLL_L_X2Y110_SLICE_X1Y110_D6 = 1'b1;
  assign CLBLM_R_X7Y112_SLICE_X9Y112_B6 = LIOB33_X0Y111_IOB_X0Y112_I;
  assign CLBLM_R_X7Y112_SLICE_X9Y112_C1 = CLBLM_L_X8Y112_SLICE_X10Y112_BO6;
  assign CLBLM_R_X7Y112_SLICE_X9Y112_C2 = CLBLM_L_X8Y112_SLICE_X10Y112_AO5;
  assign CLBLM_R_X7Y112_SLICE_X9Y112_C3 = LIOB33_X0Y111_IOB_X0Y112_I;
  assign CLBLM_R_X7Y112_SLICE_X9Y112_C4 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLM_R_X7Y112_SLICE_X9Y112_C5 = LIOB33_X0Y113_IOB_X0Y113_I;
  assign CLBLM_R_X7Y112_SLICE_X9Y112_C6 = RIOB33_X105Y101_IOB_X1Y101_I;
  assign CLBLM_R_X7Y112_SLICE_X9Y112_D1 = CLBLM_R_X7Y110_SLICE_X8Y110_BO6;
  assign CLBLM_R_X7Y112_SLICE_X9Y112_D2 = LIOB33_X0Y115_IOB_X0Y116_I;
  assign CLBLM_R_X7Y112_SLICE_X9Y112_D3 = LIOB33_X0Y113_IOB_X0Y113_I;
  assign CLBLM_R_X7Y112_SLICE_X9Y112_D4 = CLBLM_L_X8Y111_SLICE_X10Y111_BO6;
  assign CLBLM_R_X7Y112_SLICE_X9Y112_D5 = CLBLM_L_X8Y110_SLICE_X10Y110_BO6;
  assign CLBLM_R_X7Y112_SLICE_X9Y112_D6 = LIOB33_X0Y111_IOB_X0Y112_I;
  assign CLBLM_R_X7Y112_SLICE_X8Y112_A1 = CLBLM_L_X8Y112_SLICE_X11Y112_CO6;
  assign CLBLM_R_X7Y112_SLICE_X8Y112_A2 = LIOB33_X0Y111_IOB_X0Y112_I;
  assign CLBLM_R_X7Y112_SLICE_X8Y112_A3 = RIOB33_X105Y101_IOB_X1Y101_I;
  assign CLBLM_R_X7Y112_SLICE_X8Y112_A4 = CLBLM_R_X7Y112_SLICE_X8Y112_BO6;
  assign CLBLM_R_X7Y112_SLICE_X8Y112_A5 = CLBLM_L_X8Y112_SLICE_X11Y112_BO6;
  assign CLBLM_R_X7Y112_SLICE_X8Y112_A6 = 1'b1;
  assign CLBLM_R_X7Y112_SLICE_X8Y112_B1 = RIOB33_X105Y101_IOB_X1Y102_I;
  assign CLBLM_R_X7Y112_SLICE_X8Y112_B2 = CLBLM_L_X8Y112_SLICE_X11Y112_DO6;
  assign CLBLM_R_X7Y112_SLICE_X8Y112_B3 = LIOB33_X0Y111_IOB_X0Y111_I;
  assign CLBLM_R_X7Y112_SLICE_X8Y112_B4 = LIOB33_X0Y111_IOB_X0Y112_I;
  assign CLBLM_R_X7Y112_SLICE_X8Y112_B5 = RIOB33_X105Y103_IOB_X1Y103_I;
  assign CLBLM_R_X7Y112_SLICE_X8Y112_B6 = CLBLM_L_X8Y111_SLICE_X10Y111_AO5;
  assign CLBLM_R_X7Y112_SLICE_X8Y112_C1 = RIOB33_X105Y101_IOB_X1Y101_I;
  assign CLBLM_R_X7Y112_SLICE_X8Y112_C2 = LIOB33_X0Y111_IOB_X0Y112_I;
  assign CLBLM_R_X7Y112_SLICE_X8Y112_C3 = CLBLM_L_X8Y112_SLICE_X11Y112_CO6;
  assign CLBLM_R_X7Y112_SLICE_X8Y112_C4 = CLBLM_L_X8Y112_SLICE_X11Y112_BO6;
  assign CLBLM_R_X7Y112_SLICE_X8Y112_C5 = LIOB33_X0Y113_IOB_X0Y113_I;
  assign CLBLM_R_X7Y112_SLICE_X8Y112_C6 = CLBLM_R_X7Y112_SLICE_X8Y112_BO6;
  assign CLBLM_R_X7Y114_SLICE_X9Y114_C4 = 1'b1;
  assign CLBLM_R_X7Y114_SLICE_X9Y114_C5 = 1'b1;
  assign CLBLM_R_X7Y114_SLICE_X9Y114_C6 = 1'b1;
  assign CLBLM_R_X7Y112_SLICE_X8Y112_D1 = 1'b1;
  assign CLBLM_R_X7Y112_SLICE_X8Y112_D2 = 1'b1;
  assign CLBLM_R_X7Y112_SLICE_X8Y112_D3 = 1'b1;
  assign CLBLM_R_X7Y112_SLICE_X8Y112_D4 = 1'b1;
  assign CLBLM_R_X7Y112_SLICE_X8Y112_D5 = 1'b1;
  assign CLBLM_R_X7Y112_SLICE_X8Y112_D6 = 1'b1;
  assign CLBLM_R_X7Y114_SLICE_X9Y114_D5 = 1'b1;
  assign CLBLM_R_X7Y114_SLICE_X9Y114_D6 = 1'b1;
  assign CLBLM_R_X7Y114_SLICE_X8Y114_C1 = CLBLM_R_X7Y113_SLICE_X8Y113_BO6;
  assign CLBLM_R_X7Y113_SLICE_X9Y113_A1 = CLBLM_L_X8Y111_SLICE_X11Y111_AO5;
  assign CLBLM_R_X7Y113_SLICE_X9Y113_A2 = CLBLM_L_X8Y113_SLICE_X10Y113_AO5;
  assign CLBLM_R_X7Y113_SLICE_X9Y113_A3 = LIOB33_X0Y111_IOB_X0Y112_I;
  assign CLBLM_R_X7Y113_SLICE_X9Y113_A4 = LIOB33_X0Y111_IOB_X0Y111_I;
  assign CLBLM_R_X7Y113_SLICE_X9Y113_A5 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X7Y113_SLICE_X9Y113_A6 = CLBLM_R_X7Y113_SLICE_X9Y113_CO6;
  assign LIOI3_X0Y125_OLOGIC_X0Y126_D1 = CLBLM_R_X3Y107_SLICE_X2Y107_CO6;
  assign CLBLM_R_X7Y113_SLICE_X9Y113_B1 = CLBLM_R_X7Y110_SLICE_X9Y110_DO6;
  assign CLBLM_R_X7Y113_SLICE_X9Y113_B2 = CLBLM_R_X7Y110_SLICE_X9Y110_BO5;
  assign CLBLM_R_X7Y113_SLICE_X9Y113_B3 = RIOB33_X105Y107_IOB_X1Y107_I;
  assign CLBLM_R_X7Y113_SLICE_X9Y113_B4 = LIOB33_X0Y111_IOB_X0Y111_I;
  assign CLBLM_R_X7Y113_SLICE_X9Y113_B5 = LIOB33_X0Y109_IOB_X0Y110_I;
  assign CLBLM_R_X7Y113_SLICE_X9Y113_B6 = CLBLM_L_X10Y112_SLICE_X13Y112_BO6;
  assign LIOI3_X0Y125_OLOGIC_X0Y126_T1 = 1'b1;
  assign CLBLM_R_X7Y113_SLICE_X9Y113_C1 = RIOB33_X105Y107_IOB_X1Y107_I;
  assign CLBLM_R_X7Y113_SLICE_X9Y113_C2 = CLBLM_R_X7Y110_SLICE_X9Y110_BO5;
  assign CLBLM_R_X7Y113_SLICE_X9Y113_C3 = CLBLM_R_X7Y110_SLICE_X9Y110_DO6;
  assign CLBLM_R_X7Y113_SLICE_X9Y113_C4 = CLBLM_L_X10Y112_SLICE_X13Y112_BO6;
  assign CLBLM_R_X7Y113_SLICE_X9Y113_C5 = LIOB33_X0Y111_IOB_X0Y111_I;
  assign CLBLM_R_X7Y113_SLICE_X9Y113_C6 = LIOB33_X0Y109_IOB_X0Y110_I;
  assign LIOI3_X0Y125_OLOGIC_X0Y125_D1 = CLBLM_R_X7Y109_SLICE_X9Y109_AO5;
  assign CLBLM_R_X7Y113_SLICE_X9Y113_D1 = LIOB33_X0Y111_IOB_X0Y112_I;
  assign CLBLM_R_X7Y113_SLICE_X9Y113_D2 = LIOB33_X0Y111_IOB_X0Y111_I;
  assign CLBLM_R_X7Y113_SLICE_X9Y113_D3 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X7Y113_SLICE_X9Y113_D4 = CLBLM_R_X7Y113_SLICE_X9Y113_CO6;
  assign CLBLM_R_X7Y113_SLICE_X9Y113_D5 = CLBLM_L_X8Y111_SLICE_X11Y111_AO5;
  assign CLBLM_R_X7Y113_SLICE_X9Y113_D6 = CLBLM_L_X8Y113_SLICE_X10Y113_AO5;
  assign CLBLM_L_X8Y108_SLICE_X11Y108_D2 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign LIOI3_X0Y125_OLOGIC_X0Y125_T1 = 1'b1;
  assign CLBLM_R_X7Y113_SLICE_X8Y113_A1 = LIOB33_X0Y113_IOB_X0Y113_I;
  assign CLBLM_R_X7Y113_SLICE_X8Y113_A2 = CLBLM_R_X7Y113_SLICE_X8Y113_BO5;
  assign CLBLM_R_X7Y113_SLICE_X8Y113_A3 = RIOB33_X105Y103_IOB_X1Y104_I;
  assign CLBLM_R_X7Y113_SLICE_X8Y113_A4 = RIOB33_X105Y107_IOB_X1Y107_I;
  assign CLBLM_R_X7Y113_SLICE_X8Y113_A5 = CLBLM_R_X5Y110_SLICE_X7Y110_AO5;
  assign CLBLM_R_X7Y113_SLICE_X8Y113_A6 = 1'b1;
  assign LIOI3_TBYTESRC_X0Y119_OLOGIC_X0Y120_D1 = CLBLM_R_X3Y106_SLICE_X2Y106_AO5;
  assign CLBLM_R_X7Y113_SLICE_X8Y113_B1 = 1'b1;
  assign CLBLM_R_X7Y113_SLICE_X8Y113_B2 = CLBLM_R_X7Y113_SLICE_X9Y113_BO6;
  assign CLBLM_R_X7Y113_SLICE_X8Y113_B3 = CLBLM_R_X7Y110_SLICE_X9Y110_AO6;
  assign CLBLM_R_X7Y113_SLICE_X8Y113_B4 = RIOB33_X105Y107_IOB_X1Y107_I;
  assign CLBLM_R_X7Y113_SLICE_X8Y113_B5 = LIOB33_X0Y111_IOB_X0Y112_I;
  assign CLBLM_R_X7Y113_SLICE_X8Y113_B6 = 1'b1;
  assign LIOI3_TBYTESRC_X0Y119_OLOGIC_X0Y120_T1 = 1'b1;
  assign CLBLM_R_X7Y113_SLICE_X8Y113_C1 = CLBLM_R_X5Y111_SLICE_X7Y111_BO6;
  assign CLBLM_R_X7Y113_SLICE_X8Y113_C2 = CLBLM_R_X5Y110_SLICE_X7Y110_AO5;
  assign CLBLM_R_X7Y113_SLICE_X8Y113_C3 = LIOB33_X0Y113_IOB_X0Y113_I;
  assign CLBLM_R_X7Y113_SLICE_X8Y113_C4 = RIOB33_X105Y107_IOB_X1Y107_I;
  assign CLBLM_R_X7Y113_SLICE_X8Y113_C5 = CLBLM_R_X7Y113_SLICE_X8Y113_BO5;
  assign CLBLM_R_X7Y113_SLICE_X8Y113_C6 = LIOB33_X0Y115_IOB_X0Y115_I;
  assign LIOI3_TBYTESRC_X0Y119_OLOGIC_X0Y119_D1 = CLBLL_L_X2Y109_SLICE_X0Y109_AO6;
  assign LIOI3_TBYTESRC_X0Y119_OLOGIC_X0Y119_T1 = 1'b1;
  assign CLBLM_R_X7Y113_SLICE_X8Y113_D1 = CLBLM_R_X5Y111_SLICE_X7Y111_BO6;
  assign CLBLM_R_X7Y113_SLICE_X8Y113_D2 = CLBLM_R_X5Y110_SLICE_X7Y110_AO5;
  assign CLBLM_R_X7Y113_SLICE_X8Y113_D3 = LIOB33_X0Y113_IOB_X0Y113_I;
  assign CLBLM_R_X7Y113_SLICE_X8Y113_D4 = RIOB33_X105Y107_IOB_X1Y107_I;
  assign CLBLM_R_X7Y113_SLICE_X8Y113_D5 = CLBLM_R_X7Y113_SLICE_X8Y113_BO5;
  assign CLBLM_R_X7Y113_SLICE_X8Y113_D6 = LIOB33_X0Y115_IOB_X0Y115_I;
  assign RIOI3_X105Y109_ILOGIC_X1Y110_D = RIOB33_X105Y109_IOB_X1Y110_I;
  assign RIOI3_X105Y109_ILOGIC_X1Y109_D = RIOB33_X105Y109_IOB_X1Y109_I;
  assign CLBLM_R_X7Y114_SLICE_X9Y114_A1 = 1'b1;
  assign CLBLM_R_X7Y114_SLICE_X9Y114_A2 = 1'b1;
  assign CLBLM_R_X7Y114_SLICE_X9Y114_A3 = 1'b1;
  assign CLBLM_R_X7Y114_SLICE_X9Y114_A4 = 1'b1;
  assign CLBLM_R_X7Y114_SLICE_X9Y114_A5 = 1'b1;
  assign CLBLM_R_X7Y114_SLICE_X9Y114_A6 = 1'b1;
  assign CLBLM_R_X7Y114_SLICE_X9Y114_B1 = 1'b1;
  assign CLBLM_R_X7Y114_SLICE_X9Y114_B2 = 1'b1;
  assign CLBLM_R_X7Y114_SLICE_X9Y114_B3 = 1'b1;
  assign CLBLM_R_X7Y114_SLICE_X9Y114_B4 = 1'b1;
  assign CLBLM_R_X7Y114_SLICE_X9Y114_B5 = 1'b1;
  assign CLBLM_R_X7Y114_SLICE_X9Y114_B6 = 1'b1;
  assign CLBLM_R_X5Y104_SLICE_X7Y104_A1 = CLBLM_R_X7Y104_SLICE_X8Y104_CO6;
  assign CLBLM_R_X5Y104_SLICE_X7Y104_A2 = CLBLM_L_X8Y104_SLICE_X10Y104_BO6;
  assign CLBLM_R_X5Y104_SLICE_X7Y104_A3 = CLBLM_R_X5Y104_SLICE_X6Y104_AO5;
  assign CLBLM_R_X5Y104_SLICE_X7Y104_A4 = CLBLM_R_X7Y104_SLICE_X9Y104_AO6;
  assign CLBLM_R_X5Y104_SLICE_X7Y104_A5 = CLBLM_R_X7Y104_SLICE_X8Y104_DO6;
  assign CLBLM_R_X5Y104_SLICE_X7Y104_A6 = CLBLL_L_X4Y103_SLICE_X5Y103_CO6;
  assign CLBLM_R_X7Y114_SLICE_X9Y114_C1 = 1'b1;
  assign CLBLM_R_X7Y114_SLICE_X9Y114_C2 = 1'b1;
  assign CLBLM_R_X7Y114_SLICE_X9Y114_C3 = 1'b1;
  assign CLBLM_R_X5Y104_SLICE_X7Y104_B1 = LIOB33_X0Y115_IOB_X0Y116_I;
  assign CLBLM_R_X5Y104_SLICE_X7Y104_B2 = LIOB33_X0Y103_IOB_X0Y104_I;
  assign CLBLM_R_X5Y104_SLICE_X7Y104_B3 = CLBLM_R_X7Y103_SLICE_X8Y103_DO6;
  assign CLBLM_R_X5Y104_SLICE_X7Y104_B4 = LIOB33_X0Y101_IOB_X0Y102_I;
  assign CLBLM_R_X5Y104_SLICE_X7Y104_B5 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLM_R_X5Y104_SLICE_X7Y104_B6 = CLBLL_L_X4Y103_SLICE_X5Y103_CO6;
  assign CLBLM_R_X7Y114_SLICE_X9Y114_D1 = 1'b1;
  assign CLBLM_R_X7Y114_SLICE_X9Y114_D2 = 1'b1;
  assign CLBLM_R_X5Y104_SLICE_X7Y104_C1 = 1'b1;
  assign CLBLM_R_X5Y104_SLICE_X7Y104_C2 = 1'b1;
  assign CLBLM_R_X5Y104_SLICE_X7Y104_C3 = 1'b1;
  assign CLBLM_R_X5Y104_SLICE_X7Y104_C4 = 1'b1;
  assign CLBLM_R_X5Y104_SLICE_X7Y104_C5 = 1'b1;
  assign CLBLM_R_X5Y104_SLICE_X7Y104_C6 = 1'b1;
  assign CLBLM_R_X7Y114_SLICE_X9Y114_D3 = 1'b1;
  assign CLBLM_R_X7Y114_SLICE_X9Y114_D4 = 1'b1;
  assign CLBLM_R_X7Y114_SLICE_X8Y114_A1 = LIOB33_X0Y113_IOB_X0Y113_I;
  assign CLBLM_R_X7Y114_SLICE_X8Y114_A2 = 1'b1;
  assign CLBLM_R_X7Y114_SLICE_X8Y114_A3 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X7Y114_SLICE_X8Y114_A4 = CLBLM_R_X7Y113_SLICE_X9Y113_DO6;
  assign CLBLM_R_X7Y114_SLICE_X8Y114_A5 = CLBLM_R_X7Y113_SLICE_X8Y113_BO6;
  assign CLBLM_R_X7Y114_SLICE_X8Y114_A6 = 1'b1;
  assign CLBLM_R_X5Y104_SLICE_X7Y104_D1 = 1'b1;
  assign CLBLM_R_X5Y104_SLICE_X7Y104_D2 = 1'b1;
  assign CLBLM_R_X5Y104_SLICE_X7Y104_D3 = 1'b1;
  assign CLBLM_R_X5Y104_SLICE_X7Y104_D4 = 1'b1;
  assign CLBLM_R_X5Y104_SLICE_X7Y104_D5 = 1'b1;
  assign CLBLM_R_X5Y104_SLICE_X7Y104_D6 = 1'b1;
  assign CLBLM_R_X7Y114_SLICE_X8Y114_B1 = CLBLM_R_X7Y113_SLICE_X8Y113_BO6;
  assign CLBLM_R_X7Y114_SLICE_X8Y114_B6 = CLBLM_R_X7Y113_SLICE_X9Y113_DO6;
  assign CLBLM_R_X7Y114_SLICE_X8Y114_B2 = CLBLM_R_X7Y113_SLICE_X9Y113_AO6;
  assign CLBLM_R_X7Y114_SLICE_X8Y114_B3 = CLBLM_R_X7Y113_SLICE_X8Y113_AO6;
  assign CLBLM_R_X7Y114_SLICE_X8Y114_B4 = CLBLM_L_X8Y113_SLICE_X10Y113_CO6;
  assign CLBLM_R_X7Y114_SLICE_X8Y114_B5 = CLBLM_R_X7Y114_SLICE_X8Y114_AO6;
  assign CLBLM_R_X5Y104_SLICE_X6Y104_A1 = 1'b1;
  assign CLBLM_R_X5Y104_SLICE_X6Y104_A2 = 1'b1;
  assign CLBLM_R_X7Y114_SLICE_X8Y114_C2 = CLBLM_R_X7Y113_SLICE_X8Y113_AO5;
  assign CLBLM_R_X7Y114_SLICE_X8Y114_C3 = LIOB33_X0Y113_IOB_X0Y113_I;
  assign CLBLM_R_X7Y114_SLICE_X8Y114_C4 = CLBLM_R_X7Y113_SLICE_X9Y113_DO6;
  assign CLBLM_R_X7Y114_SLICE_X8Y114_C5 = LIOB33_X0Y115_IOB_X0Y115_I;
  assign CLBLM_R_X7Y114_SLICE_X8Y114_C6 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X5Y104_SLICE_X6Y104_A3 = LIOB33_X0Y115_IOB_X0Y116_I;
  assign CLBLM_R_X5Y104_SLICE_X6Y104_A4 = LIOB33_X0Y103_IOB_X0Y104_I;
  assign CLBLM_R_X5Y104_SLICE_X6Y104_A5 = LIOB33_X0Y113_IOB_X0Y114_I;
  assign CLBLM_R_X5Y104_SLICE_X6Y104_A6 = 1'b1;
  assign CLBLM_R_X5Y104_SLICE_X6Y104_B1 = LIOB33_SING_X0Y100_IOB_X0Y100_I;
  assign CLBLM_R_X5Y104_SLICE_X6Y104_B2 = RIOB33_X105Y111_IOB_X1Y112_I;
  assign CLBLM_R_X5Y104_SLICE_X6Y104_B3 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLM_R_X5Y104_SLICE_X6Y104_B4 = LIOB33_X0Y115_IOB_X0Y116_I;
  assign CLBLM_R_X5Y104_SLICE_X6Y104_B5 = RIOB33_X105Y113_IOB_X1Y113_I;
  assign CLBLM_R_X5Y104_SLICE_X6Y104_B6 = RIOB33_X105Y101_IOB_X1Y101_I;
  assign CLBLM_R_X7Y114_SLICE_X8Y114_D1 = CLBLM_R_X7Y113_SLICE_X8Y113_BO6;
  assign CLBLM_R_X7Y114_SLICE_X8Y114_D2 = CLBLM_R_X7Y113_SLICE_X8Y113_AO5;
  assign CLBLM_R_X7Y114_SLICE_X8Y114_D3 = LIOB33_X0Y113_IOB_X0Y113_I;
  assign CLBLM_R_X5Y104_SLICE_X6Y104_C1 = CLBLM_R_X7Y103_SLICE_X8Y103_DO6;
  assign CLBLM_R_X5Y104_SLICE_X6Y104_C2 = LIOB33_X0Y115_IOB_X0Y116_I;
  assign CLBLM_R_X5Y104_SLICE_X6Y104_C3 = LIOB33_X0Y103_IOB_X0Y104_I;
  assign CLBLM_R_X5Y104_SLICE_X6Y104_C4 = CLBLL_L_X4Y103_SLICE_X5Y103_CO6;
  assign CLBLM_R_X5Y104_SLICE_X6Y104_C5 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLM_R_X5Y104_SLICE_X6Y104_C6 = LIOB33_X0Y101_IOB_X0Y102_I;
  assign CLBLM_R_X7Y114_SLICE_X8Y114_D4 = CLBLM_R_X7Y113_SLICE_X9Y113_DO6;
  assign CLBLM_R_X7Y114_SLICE_X8Y114_D5 = LIOB33_X0Y115_IOB_X0Y115_I;
  assign CLBLM_R_X7Y114_SLICE_X8Y114_D6 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X5Y104_SLICE_X6Y104_D1 = CLBLM_R_X7Y103_SLICE_X8Y103_DO6;
  assign CLBLM_R_X5Y104_SLICE_X6Y104_D2 = LIOB33_X0Y115_IOB_X0Y116_I;
  assign CLBLM_R_X5Y104_SLICE_X6Y104_D3 = CLBLL_L_X4Y104_SLICE_X5Y104_AO5;
  assign CLBLM_R_X5Y104_SLICE_X6Y104_D4 = CLBLM_R_X7Y104_SLICE_X8Y104_BO6;
  assign CLBLM_R_X5Y104_SLICE_X6Y104_D5 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLM_R_X5Y104_SLICE_X6Y104_D6 = LIOB33_X0Y101_IOB_X0Y102_I;
  assign CLBLM_R_X5Y105_SLICE_X7Y105_A1 = LIOB33_X0Y113_IOB_X0Y114_I;
  assign CLBLM_R_X5Y105_SLICE_X7Y105_A2 = 1'b1;
  assign CLBLM_R_X5Y105_SLICE_X7Y105_A3 = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLM_R_X5Y105_SLICE_X7Y105_A4 = 1'b1;
  assign CLBLM_R_X5Y105_SLICE_X7Y105_A5 = LIOB33_X0Y103_IOB_X0Y103_I;
  assign CLBLM_R_X5Y105_SLICE_X7Y105_A6 = 1'b1;
  assign CLBLM_R_X5Y105_SLICE_X7Y105_B1 = CLBLM_R_X5Y104_SLICE_X6Y104_CO6;
  assign CLBLM_R_X5Y105_SLICE_X7Y105_B2 = CLBLM_R_X5Y106_SLICE_X7Y106_AO6;
  assign CLBLM_R_X5Y105_SLICE_X7Y105_B3 = CLBLM_R_X5Y104_SLICE_X7Y104_AO6;
  assign CLBLM_R_X5Y105_SLICE_X7Y105_B4 = CLBLL_L_X4Y105_SLICE_X5Y105_AO6;
  assign CLBLM_R_X5Y105_SLICE_X7Y105_B5 = CLBLM_R_X5Y105_SLICE_X7Y105_AO6;
  assign CLBLM_R_X5Y105_SLICE_X7Y105_B6 = CLBLM_R_X5Y106_SLICE_X7Y106_AO5;
  assign CLBLM_R_X5Y105_SLICE_X7Y105_C1 = CLBLM_R_X5Y105_SLICE_X7Y105_AO6;
  assign CLBLM_R_X5Y105_SLICE_X7Y105_C2 = CLBLM_R_X5Y106_SLICE_X7Y106_AO6;
  assign CLBLM_R_X5Y105_SLICE_X7Y105_C3 = CLBLM_R_X5Y106_SLICE_X7Y106_AO5;
  assign CLBLM_R_X5Y105_SLICE_X7Y105_C4 = CLBLM_R_X5Y104_SLICE_X7Y104_AO6;
  assign CLBLM_R_X5Y105_SLICE_X7Y105_C5 = CLBLM_R_X5Y104_SLICE_X6Y104_CO6;
  assign CLBLM_R_X5Y105_SLICE_X7Y105_C6 = CLBLL_L_X4Y105_SLICE_X5Y105_AO6;
  assign CLBLM_R_X5Y105_SLICE_X7Y105_D1 = 1'b1;
  assign CLBLM_R_X5Y105_SLICE_X7Y105_D2 = 1'b1;
  assign CLBLM_R_X5Y105_SLICE_X7Y105_D3 = 1'b1;
  assign CLBLM_R_X5Y105_SLICE_X7Y105_D4 = 1'b1;
  assign CLBLM_R_X5Y105_SLICE_X7Y105_D5 = 1'b1;
  assign CLBLM_R_X5Y105_SLICE_X7Y105_D6 = 1'b1;
  assign CLBLM_R_X5Y105_SLICE_X6Y105_A1 = LIOB33_X0Y105_IOB_X0Y105_I;
  assign CLBLM_R_X5Y105_SLICE_X6Y105_A2 = CLBLM_R_X5Y104_SLICE_X6Y104_CO6;
  assign CLBLM_R_X5Y105_SLICE_X6Y105_A3 = CLBLM_R_X5Y104_SLICE_X7Y104_AO6;
  assign CLBLM_R_X5Y105_SLICE_X6Y105_A4 = LIOB33_X0Y115_IOB_X0Y116_I;
  assign CLBLM_R_X5Y105_SLICE_X6Y105_A5 = LIOB33_X0Y113_IOB_X0Y114_I;
  assign CLBLM_R_X5Y105_SLICE_X6Y105_A6 = CLBLL_L_X4Y105_SLICE_X5Y105_AO6;
  assign CLBLM_R_X5Y105_SLICE_X6Y105_B1 = LIOB33_X0Y105_IOB_X0Y105_I;
  assign CLBLM_R_X5Y105_SLICE_X6Y105_B2 = LIOB33_X0Y115_IOB_X0Y116_I;
  assign CLBLM_R_X5Y105_SLICE_X6Y105_B3 = LIOB33_X0Y103_IOB_X0Y104_I;
  assign CLBLM_R_X5Y105_SLICE_X6Y105_B4 = CLBLM_R_X5Y104_SLICE_X6Y104_DO6;
  assign CLBLM_R_X5Y105_SLICE_X6Y105_B5 = LIOB33_X0Y113_IOB_X0Y114_I;
  assign CLBLM_R_X5Y105_SLICE_X6Y105_B6 = CLBLL_L_X4Y105_SLICE_X5Y105_AO6;
  assign CLBLM_R_X5Y105_SLICE_X6Y105_C1 = LIOB33_X0Y113_IOB_X0Y114_I;
  assign CLBLM_R_X5Y105_SLICE_X6Y105_C2 = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLM_R_X5Y105_SLICE_X6Y105_C3 = CLBLM_R_X7Y105_SLICE_X9Y105_CO6;
  assign CLBLM_R_X5Y105_SLICE_X6Y105_C4 = CLBLM_R_X7Y105_SLICE_X9Y105_DO6;
  assign CLBLM_R_X5Y105_SLICE_X6Y105_C5 = CLBLM_R_X5Y105_SLICE_X6Y105_DO6;
  assign CLBLM_R_X5Y105_SLICE_X6Y105_C6 = LIOB33_X0Y115_IOB_X0Y116_I;
  assign CLBLM_R_X5Y105_SLICE_X6Y105_D1 = LIOB33_X0Y103_IOB_X0Y104_I;
  assign CLBLM_R_X5Y105_SLICE_X6Y105_D2 = LIOB33_X0Y113_IOB_X0Y114_I;
  assign CLBLM_R_X5Y105_SLICE_X6Y105_D3 = LIOB33_X0Y105_IOB_X0Y105_I;
  assign CLBLM_R_X5Y105_SLICE_X6Y105_D4 = CLBLM_R_X5Y104_SLICE_X6Y104_DO6;
  assign CLBLM_R_X5Y105_SLICE_X6Y105_D5 = LIOB33_X0Y115_IOB_X0Y116_I;
  assign CLBLM_R_X5Y105_SLICE_X6Y105_D6 = CLBLL_L_X4Y105_SLICE_X5Y105_AO6;
  assign LIOI3_X0Y127_OLOGIC_X0Y128_D1 = CLBLM_R_X3Y107_SLICE_X3Y107_BO6;
  assign LIOI3_X0Y127_OLOGIC_X0Y128_T1 = 1'b1;
  assign LIOI3_X0Y127_OLOGIC_X0Y127_D1 = CLBLM_R_X3Y107_SLICE_X3Y107_AO6;
  assign LIOI3_X0Y127_OLOGIC_X0Y127_T1 = 1'b1;
  assign LIOI3_TBYTESRC_X0Y131_OLOGIC_X0Y132_D1 = CLBLL_L_X2Y110_SLICE_X0Y110_AO5;
  assign LIOI3_TBYTESRC_X0Y131_OLOGIC_X0Y132_T1 = 1'b1;
  assign LIOI3_TBYTESRC_X0Y131_OLOGIC_X0Y131_D1 = CLBLL_L_X4Y108_SLICE_X4Y108_AO6;
  assign LIOI3_TBYTESRC_X0Y131_OLOGIC_X0Y131_T1 = 1'b1;
  assign CLBLM_R_X5Y106_SLICE_X7Y106_A1 = LIOB33_X0Y113_IOB_X0Y114_I;
  assign CLBLM_R_X5Y106_SLICE_X7Y106_A2 = 1'b1;
  assign CLBLM_R_X5Y106_SLICE_X7Y106_A3 = LIOB33_X0Y105_IOB_X0Y105_I;
  assign CLBLM_R_X5Y106_SLICE_X7Y106_A4 = LIOB33_X0Y115_IOB_X0Y116_I;
  assign CLBLM_R_X5Y106_SLICE_X7Y106_A5 = 1'b1;
  assign CLBLM_R_X5Y106_SLICE_X7Y106_A6 = 1'b1;
  assign RIOI3_X105Y103_ILOGIC_X1Y104_D = RIOB33_X105Y103_IOB_X1Y104_I;
  assign CLBLM_R_X5Y106_SLICE_X7Y106_B1 = LIOB33_X0Y113_IOB_X0Y114_I;
  assign CLBLM_R_X5Y106_SLICE_X7Y106_B2 = 1'b1;
  assign CLBLM_R_X5Y106_SLICE_X7Y106_B3 = LIOB33_X0Y103_IOB_X0Y103_I;
  assign CLBLM_R_X5Y106_SLICE_X7Y106_B4 = 1'b1;
  assign CLBLM_R_X5Y106_SLICE_X7Y106_B5 = LIOB33_X0Y107_IOB_X0Y107_I;
  assign CLBLM_R_X5Y106_SLICE_X7Y106_B6 = 1'b1;
  assign RIOI3_X105Y111_ILOGIC_X1Y112_D = RIOB33_X105Y111_IOB_X1Y112_I;
  assign RIOI3_X105Y111_ILOGIC_X1Y111_D = RIOB33_X105Y111_IOB_X1Y111_I;
  assign CLBLM_R_X5Y106_SLICE_X7Y106_C1 = CLBLL_L_X4Y105_SLICE_X5Y105_BO6;
  assign CLBLM_R_X5Y106_SLICE_X7Y106_C2 = CLBLM_R_X7Y105_SLICE_X9Y105_AO6;
  assign CLBLM_R_X5Y106_SLICE_X7Y106_C3 = CLBLM_R_X5Y105_SLICE_X7Y105_BO6;
  assign CLBLM_R_X5Y106_SLICE_X7Y106_C4 = CLBLM_R_X5Y105_SLICE_X7Y105_CO6;
  assign CLBLM_R_X5Y106_SLICE_X7Y106_C5 = CLBLM_R_X5Y106_SLICE_X7Y106_BO5;
  assign CLBLM_R_X5Y106_SLICE_X7Y106_C6 = CLBLM_R_X5Y106_SLICE_X7Y106_BO6;
  assign RIOI3_X105Y103_ILOGIC_X1Y103_D = RIOB33_X105Y103_IOB_X1Y103_I;
  assign CLBLM_R_X5Y106_SLICE_X7Y106_D1 = LIOB33_X0Y107_IOB_X0Y107_I;
  assign CLBLM_R_X5Y106_SLICE_X7Y106_D2 = CLBLM_R_X7Y105_SLICE_X9Y105_CO6;
  assign CLBLM_R_X5Y106_SLICE_X7Y106_D3 = LIOB33_X0Y113_IOB_X0Y114_I;
  assign CLBLM_R_X5Y106_SLICE_X7Y106_D4 = CLBLM_R_X5Y105_SLICE_X7Y105_CO6;
  assign CLBLM_R_X5Y106_SLICE_X7Y106_D5 = LIOB33_X0Y115_IOB_X0Y116_I;
  assign CLBLM_R_X5Y106_SLICE_X7Y106_D6 = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLM_R_X5Y106_SLICE_X6Y106_A1 = 1'b1;
  assign CLBLM_R_X5Y106_SLICE_X6Y106_A2 = 1'b1;
  assign CLBLM_R_X5Y106_SLICE_X6Y106_A3 = LIOB33_X0Y113_IOB_X0Y114_I;
  assign CLBLM_R_X5Y106_SLICE_X6Y106_A4 = LIOB33_X0Y109_IOB_X0Y109_I;
  assign CLBLM_R_X5Y106_SLICE_X6Y106_A5 = LIOB33_X0Y103_IOB_X0Y103_I;
  assign CLBLM_R_X5Y106_SLICE_X6Y106_A6 = 1'b1;
  assign CLBLM_R_X5Y106_SLICE_X6Y106_B1 = LIOB33_X0Y107_IOB_X0Y108_I;
  assign CLBLM_R_X5Y106_SLICE_X6Y106_B2 = CLBLM_R_X5Y106_SLICE_X7Y106_DO6;
  assign CLBLM_R_X5Y106_SLICE_X6Y106_B3 = LIOB33_X0Y113_IOB_X0Y114_I;
  assign CLBLM_R_X5Y106_SLICE_X6Y106_B4 = CLBLM_R_X7Y106_SLICE_X8Y106_BO6;
  assign CLBLM_R_X5Y106_SLICE_X6Y106_B5 = CLBLL_L_X4Y106_SLICE_X5Y106_BO6;
  assign CLBLM_R_X5Y106_SLICE_X6Y106_B6 = LIOB33_X0Y103_IOB_X0Y103_I;
  assign CLBLM_R_X5Y106_SLICE_X6Y106_C1 = CLBLM_R_X5Y106_SLICE_X6Y106_AO6;
  assign CLBLM_R_X5Y106_SLICE_X6Y106_C2 = CLBLL_L_X4Y107_SLICE_X5Y107_AO6;
  assign CLBLM_R_X5Y106_SLICE_X6Y106_C3 = CLBLM_R_X5Y106_SLICE_X7Y106_DO6;
  assign CLBLM_R_X5Y106_SLICE_X6Y106_C4 = CLBLL_L_X4Y106_SLICE_X5Y106_BO6;
  assign CLBLM_R_X5Y106_SLICE_X6Y106_C5 = CLBLM_R_X7Y106_SLICE_X8Y106_AO5;
  assign CLBLM_R_X5Y106_SLICE_X6Y106_C6 = CLBLM_R_X7Y106_SLICE_X8Y106_BO6;
  assign CLBLM_R_X5Y106_SLICE_X6Y106_D1 = CLBLM_R_X5Y106_SLICE_X6Y106_AO6;
  assign CLBLM_R_X5Y106_SLICE_X6Y106_D2 = CLBLL_L_X4Y107_SLICE_X5Y107_AO6;
  assign CLBLM_R_X5Y106_SLICE_X6Y106_D3 = CLBLM_R_X5Y106_SLICE_X7Y106_DO6;
  assign CLBLM_R_X5Y106_SLICE_X6Y106_D4 = CLBLL_L_X4Y106_SLICE_X5Y106_BO6;
  assign CLBLM_R_X5Y106_SLICE_X6Y106_D5 = CLBLM_R_X7Y106_SLICE_X8Y106_AO5;
  assign CLBLM_R_X5Y106_SLICE_X6Y106_D6 = CLBLM_R_X7Y106_SLICE_X8Y106_BO6;
  assign CLBLM_R_X5Y107_SLICE_X7Y107_A1 = LIOB33_X0Y109_IOB_X0Y110_I;
  assign CLBLM_R_X5Y107_SLICE_X7Y107_A2 = 1'b1;
  assign CLBLM_R_X5Y107_SLICE_X7Y107_A3 = LIOB33_X0Y113_IOB_X0Y114_I;
  assign CLBLM_R_X5Y107_SLICE_X7Y107_A4 = 1'b1;
  assign CLBLM_R_X5Y107_SLICE_X7Y107_A5 = LIOB33_X0Y103_IOB_X0Y103_I;
  assign CLBLM_R_X5Y107_SLICE_X7Y107_A6 = 1'b1;
  assign CLBLM_R_X5Y107_SLICE_X7Y107_B1 = LIOB33_X0Y103_IOB_X0Y103_I;
  assign CLBLM_R_X5Y107_SLICE_X7Y107_B2 = CLBLM_R_X7Y105_SLICE_X8Y105_CO6;
  assign CLBLM_R_X5Y107_SLICE_X7Y107_B3 = LIOB33_X0Y109_IOB_X0Y109_I;
  assign CLBLM_R_X5Y107_SLICE_X7Y107_B4 = CLBLM_R_X7Y106_SLICE_X9Y106_AO6;
  assign CLBLM_R_X5Y107_SLICE_X7Y107_B5 = CLBLL_L_X4Y106_SLICE_X5Y106_DO6;
  assign CLBLM_R_X5Y107_SLICE_X7Y107_B6 = LIOB33_X0Y113_IOB_X0Y114_I;
  assign CLBLM_R_X5Y107_SLICE_X7Y107_C1 = CLBLL_L_X4Y106_SLICE_X5Y106_DO6;
  assign CLBLM_R_X5Y107_SLICE_X7Y107_C2 = CLBLM_R_X7Y105_SLICE_X8Y105_CO6;
  assign CLBLM_R_X5Y107_SLICE_X7Y107_C3 = LIOB33_X0Y103_IOB_X0Y103_I;
  assign CLBLM_R_X5Y107_SLICE_X7Y107_C4 = LIOB33_X0Y109_IOB_X0Y110_I;
  assign CLBLM_R_X5Y107_SLICE_X7Y107_C5 = LIOB33_X0Y109_IOB_X0Y109_I;
  assign CLBLM_R_X5Y107_SLICE_X7Y107_C6 = CLBLM_R_X7Y106_SLICE_X9Y106_BO6;
  assign CLBLM_R_X5Y107_SLICE_X7Y107_D1 = 1'b1;
  assign CLBLM_R_X5Y107_SLICE_X7Y107_D2 = 1'b1;
  assign CLBLM_R_X5Y107_SLICE_X7Y107_D3 = 1'b1;
  assign CLBLM_R_X5Y107_SLICE_X7Y107_D4 = 1'b1;
  assign CLBLM_R_X5Y107_SLICE_X7Y107_D5 = 1'b1;
  assign CLBLM_R_X5Y107_SLICE_X7Y107_D6 = 1'b1;
  assign CLBLM_R_X5Y107_SLICE_X6Y107_A1 = RIOB33_X105Y105_IOB_X1Y106_I;
  assign CLBLM_R_X5Y107_SLICE_X6Y107_A2 = CLBLM_R_X5Y106_SLICE_X6Y106_BO6;
  assign CLBLM_R_X5Y107_SLICE_X6Y107_A3 = LIOB33_X0Y109_IOB_X0Y109_I;
  assign CLBLM_R_X5Y107_SLICE_X6Y107_A4 = CLBLL_L_X4Y107_SLICE_X4Y107_CO6;
  assign CLBLM_R_X5Y107_SLICE_X6Y107_A5 = LIOB33_X0Y103_IOB_X0Y103_I;
  assign CLBLM_R_X5Y107_SLICE_X6Y107_A6 = CLBLL_L_X4Y106_SLICE_X5Y106_CO6;
  assign CLBLM_R_X5Y107_SLICE_X6Y107_B1 = RIOB33_X105Y105_IOB_X1Y106_I;
  assign CLBLM_R_X5Y107_SLICE_X6Y107_B2 = CLBLL_L_X4Y107_SLICE_X4Y107_CO6;
  assign CLBLM_R_X5Y107_SLICE_X6Y107_B3 = LIOB33_X0Y109_IOB_X0Y110_I;
  assign CLBLM_R_X5Y107_SLICE_X6Y107_B4 = CLBLL_L_X4Y106_SLICE_X5Y106_CO6;
  assign CLBLM_R_X5Y107_SLICE_X6Y107_B5 = LIOB33_X0Y109_IOB_X0Y109_I;
  assign CLBLM_R_X5Y107_SLICE_X6Y107_B6 = CLBLM_R_X5Y106_SLICE_X6Y106_CO6;
  assign CLBLM_R_X5Y107_SLICE_X6Y107_C1 = CLBLM_R_X7Y106_SLICE_X9Y106_BO6;
  assign CLBLM_R_X5Y107_SLICE_X6Y107_C2 = CLBLM_R_X5Y107_SLICE_X7Y107_AO6;
  assign CLBLM_R_X5Y107_SLICE_X6Y107_C3 = CLBLM_R_X5Y106_SLICE_X6Y106_DO6;
  assign CLBLM_R_X5Y107_SLICE_X6Y107_C4 = CLBLM_R_X5Y106_SLICE_X6Y106_CO6;
  assign CLBLM_R_X5Y107_SLICE_X6Y107_C5 = CLBLM_R_X3Y107_SLICE_X3Y107_BO5;
  assign CLBLM_R_X5Y107_SLICE_X6Y107_C6 = CLBLL_L_X4Y107_SLICE_X5Y107_DO6;
  assign CLBLM_R_X5Y107_SLICE_X6Y107_D1 = LIOB33_X0Y109_IOB_X0Y110_I;
  assign CLBLM_R_X5Y107_SLICE_X6Y107_D2 = CLBLL_L_X4Y107_SLICE_X4Y107_CO6;
  assign CLBLM_R_X5Y107_SLICE_X6Y107_D3 = RIOB33_X105Y105_IOB_X1Y106_I;
  assign CLBLM_R_X5Y107_SLICE_X6Y107_D4 = CLBLM_R_X5Y106_SLICE_X6Y106_CO6;
  assign CLBLM_R_X5Y107_SLICE_X6Y107_D5 = LIOB33_X0Y109_IOB_X0Y109_I;
  assign CLBLM_R_X5Y107_SLICE_X6Y107_D6 = CLBLL_L_X4Y106_SLICE_X5Y106_CO6;
  assign LIOI3_X0Y129_OLOGIC_X0Y130_D1 = CLBLL_L_X2Y110_SLICE_X0Y110_AO6;
  assign LIOI3_X0Y129_OLOGIC_X0Y130_T1 = 1'b1;
  assign LIOI3_X0Y129_OLOGIC_X0Y129_D1 = CLBLM_R_X3Y108_SLICE_X3Y108_AO6;
  assign LIOI3_X0Y129_OLOGIC_X0Y129_T1 = 1'b1;
  assign LIOI3_TBYTESRC_X0Y143_OLOGIC_X0Y144_D1 = CLBLL_L_X4Y116_SLICE_X4Y116_AO6;
  assign LIOI3_TBYTESRC_X0Y143_OLOGIC_X0Y144_T1 = 1'b1;
  assign LIOI3_TBYTESRC_X0Y143_OLOGIC_X0Y143_D1 = CLBLL_L_X4Y115_SLICE_X4Y115_DO6;
  assign LIOI3_TBYTESRC_X0Y143_OLOGIC_X0Y143_T1 = 1'b1;
  assign CLBLM_R_X5Y108_SLICE_X7Y108_A1 = RIOB33_X105Y105_IOB_X1Y106_I;
  assign CLBLM_R_X5Y108_SLICE_X7Y108_A2 = 1'b1;
  assign CLBLM_R_X5Y108_SLICE_X7Y108_A3 = 1'b1;
  assign CLBLM_R_X5Y108_SLICE_X7Y108_A4 = LIOB33_X0Y111_IOB_X0Y111_I;
  assign CLBLM_R_X5Y108_SLICE_X7Y108_A5 = LIOB33_X0Y103_IOB_X0Y103_I;
  assign CLBLM_R_X5Y108_SLICE_X7Y108_A6 = 1'b1;
  assign CLBLM_R_X5Y108_SLICE_X7Y108_B1 = LIOB33_X0Y111_IOB_X0Y111_I;
  assign CLBLM_R_X5Y108_SLICE_X7Y108_B2 = CLBLM_R_X7Y107_SLICE_X9Y107_DO6;
  assign CLBLM_R_X5Y108_SLICE_X7Y108_B3 = LIOB33_X0Y109_IOB_X0Y110_I;
  assign CLBLM_R_X5Y108_SLICE_X7Y108_B4 = CLBLM_R_X7Y108_SLICE_X9Y108_DO6;
  assign CLBLM_R_X5Y108_SLICE_X7Y108_B5 = LIOB33_X0Y115_IOB_X0Y116_I;
  assign CLBLM_R_X5Y108_SLICE_X7Y108_B6 = LIOB33_X0Y113_IOB_X0Y114_I;
  assign CLBLM_R_X5Y108_SLICE_X7Y108_C1 = LIOB33_X0Y109_IOB_X0Y110_I;
  assign CLBLM_R_X5Y108_SLICE_X7Y108_C2 = LIOB33_X0Y111_IOB_X0Y111_I;
  assign CLBLM_R_X5Y108_SLICE_X7Y108_C3 = CLBLM_R_X7Y108_SLICE_X9Y108_DO6;
  assign CLBLM_R_X5Y108_SLICE_X7Y108_C4 = LIOB33_X0Y113_IOB_X0Y114_I;
  assign CLBLM_R_X5Y108_SLICE_X7Y108_C5 = LIOB33_X0Y115_IOB_X0Y116_I;
  assign CLBLM_R_X5Y108_SLICE_X7Y108_C6 = CLBLM_R_X7Y107_SLICE_X9Y107_DO6;
  assign CLBLM_L_X8Y109_SLICE_X11Y109_D2 = 1'b1;
  assign CLBLM_R_X5Y108_SLICE_X7Y108_D1 = 1'b1;
  assign CLBLM_R_X5Y108_SLICE_X7Y108_D2 = 1'b1;
  assign CLBLM_R_X5Y108_SLICE_X7Y108_D3 = 1'b1;
  assign CLBLM_R_X5Y108_SLICE_X7Y108_D4 = 1'b1;
  assign CLBLM_R_X5Y108_SLICE_X7Y108_D5 = 1'b1;
  assign CLBLM_R_X5Y108_SLICE_X7Y108_D6 = 1'b1;
  assign CLBLM_L_X8Y109_SLICE_X11Y109_D4 = 1'b1;
  assign CLBLM_R_X5Y108_SLICE_X6Y108_A1 = RIOB33_X105Y105_IOB_X1Y106_I;
  assign CLBLM_R_X5Y108_SLICE_X6Y108_A2 = LIOB33_X0Y111_IOB_X0Y111_I;
  assign CLBLM_R_X5Y108_SLICE_X6Y108_A3 = LIOB33_X0Y109_IOB_X0Y110_I;
  assign CLBLM_R_X5Y108_SLICE_X6Y108_A4 = CLBLM_R_X5Y107_SLICE_X6Y107_BO6;
  assign CLBLM_R_X5Y108_SLICE_X6Y108_A5 = CLBLM_R_X5Y107_SLICE_X7Y107_BO6;
  assign CLBLM_R_X5Y108_SLICE_X6Y108_A6 = LIOB33_X0Y103_IOB_X0Y103_I;
  assign CLBLM_R_X5Y108_SLICE_X6Y108_B1 = RIOB33_X105Y105_IOB_X1Y106_I;
  assign CLBLM_R_X5Y108_SLICE_X6Y108_B2 = CLBLM_R_X5Y107_SLICE_X6Y107_BO6;
  assign CLBLM_R_X5Y108_SLICE_X6Y108_B3 = LIOB33_X0Y109_IOB_X0Y110_I;
  assign CLBLM_R_X5Y108_SLICE_X6Y108_B4 = LIOB33_X0Y103_IOB_X0Y103_I;
  assign CLBLM_R_X5Y108_SLICE_X6Y108_B5 = CLBLM_R_X5Y107_SLICE_X7Y107_BO6;
  assign CLBLM_R_X5Y108_SLICE_X6Y108_B6 = LIOB33_X0Y111_IOB_X0Y111_I;
  assign CLBLM_R_X5Y108_SLICE_X6Y108_C1 = CLBLL_L_X4Y107_SLICE_X4Y107_BO6;
  assign CLBLM_R_X5Y108_SLICE_X6Y108_C2 = CLBLM_R_X5Y107_SLICE_X6Y107_CO6;
  assign CLBLM_R_X5Y108_SLICE_X6Y108_C3 = CLBLM_R_X5Y108_SLICE_X7Y108_AO6;
  assign CLBLM_R_X5Y108_SLICE_X6Y108_C4 = CLBLM_R_X5Y110_SLICE_X6Y110_AO6;
  assign CLBLM_R_X5Y108_SLICE_X6Y108_C5 = CLBLM_R_X5Y110_SLICE_X7Y110_AO6;
  assign CLBLM_R_X5Y108_SLICE_X6Y108_C6 = CLBLM_R_X5Y107_SLICE_X6Y107_DO6;
  assign CLBLM_R_X5Y108_SLICE_X6Y108_D1 = 1'b1;
  assign CLBLM_R_X5Y108_SLICE_X6Y108_D2 = 1'b1;
  assign CLBLM_R_X5Y108_SLICE_X6Y108_D3 = 1'b1;
  assign CLBLM_R_X5Y108_SLICE_X6Y108_D4 = 1'b1;
  assign CLBLM_R_X5Y108_SLICE_X6Y108_D5 = 1'b1;
  assign CLBLM_R_X5Y108_SLICE_X6Y108_D6 = 1'b1;
  assign CLBLM_R_X5Y109_SLICE_X7Y109_A1 = CLBLM_R_X7Y109_SLICE_X8Y109_CO6;
  assign CLBLM_R_X5Y109_SLICE_X7Y109_A2 = CLBLM_R_X7Y109_SLICE_X8Y109_BO6;
  assign CLBLM_R_X5Y109_SLICE_X7Y109_A3 = LIOB33_X0Y115_IOB_X0Y116_I;
  assign CLBLM_R_X5Y109_SLICE_X7Y109_A4 = CLBLM_R_X5Y108_SLICE_X7Y108_BO6;
  assign CLBLM_R_X5Y109_SLICE_X7Y109_A5 = LIOB33_X0Y111_IOB_X0Y112_I;
  assign CLBLM_R_X5Y109_SLICE_X7Y109_A6 = LIOB33_X0Y113_IOB_X0Y114_I;
  assign CLBLM_R_X5Y109_SLICE_X7Y109_B1 = CLBLM_R_X7Y109_SLICE_X8Y109_CO6;
  assign CLBLM_R_X5Y109_SLICE_X7Y109_B2 = CLBLM_R_X5Y108_SLICE_X7Y108_BO6;
  assign CLBLM_R_X5Y109_SLICE_X7Y109_B3 = LIOB33_X0Y113_IOB_X0Y114_I;
  assign CLBLM_R_X5Y109_SLICE_X7Y109_B4 = CLBLM_R_X7Y109_SLICE_X8Y109_DO6;
  assign CLBLM_R_X5Y109_SLICE_X7Y109_B5 = LIOB33_X0Y111_IOB_X0Y112_I;
  assign CLBLM_R_X5Y109_SLICE_X7Y109_B6 = LIOB33_X0Y113_IOB_X0Y113_I;
  assign CLBLM_R_X5Y109_SLICE_X7Y109_C1 = 1'b1;
  assign CLBLM_R_X5Y109_SLICE_X7Y109_C2 = 1'b1;
  assign CLBLM_R_X5Y109_SLICE_X7Y109_C3 = 1'b1;
  assign CLBLM_R_X5Y109_SLICE_X7Y109_C4 = 1'b1;
  assign CLBLM_R_X5Y109_SLICE_X7Y109_C5 = 1'b1;
  assign CLBLM_R_X5Y109_SLICE_X7Y109_C6 = 1'b1;
  assign CLBLM_R_X5Y109_SLICE_X7Y109_D1 = 1'b1;
  assign CLBLM_R_X5Y109_SLICE_X7Y109_D2 = 1'b1;
  assign CLBLM_R_X5Y109_SLICE_X7Y109_D3 = 1'b1;
  assign CLBLM_R_X5Y109_SLICE_X7Y109_D4 = 1'b1;
  assign CLBLM_R_X5Y109_SLICE_X7Y109_D5 = 1'b1;
  assign CLBLM_R_X5Y109_SLICE_X7Y109_D6 = 1'b1;
  assign CLBLM_R_X5Y109_SLICE_X6Y109_A1 = 1'b1;
  assign CLBLM_R_X5Y109_SLICE_X6Y109_A2 = 1'b1;
  assign CLBLM_R_X5Y109_SLICE_X6Y109_A3 = 1'b1;
  assign CLBLM_R_X5Y109_SLICE_X6Y109_A4 = 1'b1;
  assign CLBLM_R_X5Y109_SLICE_X6Y109_A5 = 1'b1;
  assign CLBLM_R_X5Y109_SLICE_X6Y109_A6 = 1'b1;
  assign CLBLM_R_X5Y109_SLICE_X6Y109_B1 = 1'b1;
  assign CLBLM_R_X5Y109_SLICE_X6Y109_B2 = 1'b1;
  assign CLBLM_R_X5Y109_SLICE_X6Y109_B3 = 1'b1;
  assign CLBLM_R_X5Y109_SLICE_X6Y109_B4 = 1'b1;
  assign CLBLM_R_X5Y109_SLICE_X6Y109_B5 = 1'b1;
  assign CLBLM_R_X5Y109_SLICE_X6Y109_B6 = 1'b1;
  assign CLBLM_R_X5Y109_SLICE_X6Y109_C1 = 1'b1;
  assign CLBLM_R_X5Y109_SLICE_X6Y109_C2 = 1'b1;
  assign CLBLM_R_X5Y109_SLICE_X6Y109_C3 = 1'b1;
  assign CLBLM_R_X5Y109_SLICE_X6Y109_C4 = 1'b1;
  assign CLBLM_R_X5Y109_SLICE_X6Y109_C5 = 1'b1;
  assign CLBLM_R_X5Y109_SLICE_X6Y109_C6 = 1'b1;
  assign CLBLM_R_X5Y109_SLICE_X6Y109_D1 = 1'b1;
  assign CLBLM_R_X5Y109_SLICE_X6Y109_D2 = 1'b1;
  assign CLBLM_R_X5Y109_SLICE_X6Y109_D3 = 1'b1;
  assign CLBLM_R_X5Y109_SLICE_X6Y109_D4 = 1'b1;
  assign CLBLM_R_X5Y109_SLICE_X6Y109_D5 = 1'b1;
  assign CLBLM_R_X5Y109_SLICE_X6Y109_D6 = 1'b1;
  assign CLBLM_R_X5Y110_SLICE_X7Y110_A1 = CLBLM_R_X7Y110_SLICE_X9Y110_AO5;
  assign CLBLM_R_X5Y110_SLICE_X7Y110_A2 = CLBLM_R_X7Y111_SLICE_X9Y111_AO6;
  assign CLBLM_R_X5Y110_SLICE_X7Y110_A3 = LIOB33_X0Y111_IOB_X0Y112_I;
  assign CLBLM_R_X5Y110_SLICE_X7Y110_A4 = RIOB33_SING_X105Y100_IOB_X1Y100_I;
  assign CLBLM_R_X5Y110_SLICE_X7Y110_A5 = RIOB33_X105Y107_IOB_X1Y108_I;
  assign CLBLM_R_X5Y110_SLICE_X7Y110_A6 = 1'b1;
  assign LIOI3_X0Y133_OLOGIC_X0Y134_D1 = 1'b0;
  assign CLBLM_R_X5Y110_SLICE_X7Y110_B1 = 1'b1;
  assign CLBLM_R_X5Y110_SLICE_X7Y110_B2 = RIOB33_X105Y103_IOB_X1Y103_I;
  assign CLBLM_R_X5Y110_SLICE_X7Y110_B3 = LIOB33_X0Y103_IOB_X0Y103_I;
  assign CLBLM_R_X5Y110_SLICE_X7Y110_B4 = LIOB33_X0Y111_IOB_X0Y112_I;
  assign CLBLM_R_X5Y110_SLICE_X7Y110_B5 = CLBLM_R_X7Y111_SLICE_X8Y111_BO6;
  assign CLBLM_R_X5Y110_SLICE_X7Y110_B6 = 1'b1;
  assign CLBLM_R_X5Y110_SLICE_X7Y110_C1 = CLBLM_R_X7Y111_SLICE_X8Y111_BO6;
  assign CLBLM_R_X5Y110_SLICE_X7Y110_C2 = LIOB33_X0Y111_IOB_X0Y112_I;
  assign CLBLM_R_X5Y110_SLICE_X7Y110_C3 = CLBLM_L_X8Y112_SLICE_X11Y112_DO6;
  assign CLBLM_R_X5Y110_SLICE_X7Y110_C4 = CLBLM_R_X7Y111_SLICE_X8Y111_AO6;
  assign CLBLM_R_X5Y110_SLICE_X7Y110_C5 = RIOB33_X105Y101_IOB_X1Y102_I;
  assign CLBLM_R_X5Y110_SLICE_X7Y110_C6 = RIOB33_X105Y103_IOB_X1Y103_I;
  assign LIOI3_X0Y133_OLOGIC_X0Y134_T1 = 1'b1;
  assign LIOI3_X0Y133_OLOGIC_X0Y133_D1 = CLBLM_R_X3Y109_SLICE_X3Y109_AO6;
  assign CLBLM_R_X5Y110_SLICE_X7Y110_D1 = RIOB33_X105Y101_IOB_X1Y102_I;
  assign CLBLM_R_X5Y110_SLICE_X7Y110_D2 = CLBLM_R_X7Y111_SLICE_X8Y111_AO6;
  assign CLBLM_R_X5Y110_SLICE_X7Y110_D3 = CLBLM_L_X8Y112_SLICE_X11Y112_DO6;
  assign CLBLM_R_X5Y110_SLICE_X7Y110_D4 = LIOB33_X0Y113_IOB_X0Y113_I;
  assign CLBLM_R_X5Y110_SLICE_X7Y110_D5 = CLBLM_R_X5Y110_SLICE_X7Y110_BO5;
  assign CLBLM_R_X5Y110_SLICE_X7Y110_D6 = LIOB33_X0Y111_IOB_X0Y112_I;
  assign LIOI3_X0Y133_OLOGIC_X0Y133_T1 = 1'b1;
  assign CLBLM_R_X5Y110_SLICE_X6Y110_A1 = CLBLM_L_X8Y111_SLICE_X11Y111_BO6;
  assign CLBLM_R_X5Y110_SLICE_X6Y110_A2 = RIOB33_SING_X105Y100_IOB_X1Y100_I;
  assign CLBLM_R_X5Y110_SLICE_X6Y110_A3 = RIOB33_X105Y103_IOB_X1Y104_I;
  assign CLBLM_R_X5Y110_SLICE_X6Y110_A4 = 1'b1;
  assign CLBLM_R_X5Y110_SLICE_X6Y110_A5 = LIOB33_X0Y111_IOB_X0Y111_I;
  assign CLBLM_R_X5Y110_SLICE_X6Y110_A6 = 1'b1;
  assign CLBLM_R_X5Y110_SLICE_X6Y110_B1 = CLBLM_R_X5Y112_SLICE_X7Y112_DO6;
  assign CLBLM_R_X5Y110_SLICE_X6Y110_B2 = RIOB33_X105Y109_IOB_X1Y110_I;
  assign CLBLM_R_X5Y110_SLICE_X6Y110_B3 = LIOB33_X0Y111_IOB_X0Y111_I;
  assign CLBLM_R_X5Y110_SLICE_X6Y110_B4 = LIOB33_X0Y111_IOB_X0Y112_I;
  assign CLBLM_R_X5Y110_SLICE_X6Y110_B5 = RIOB33_X105Y111_IOB_X1Y111_I;
  assign CLBLM_R_X5Y110_SLICE_X6Y110_B6 = 1'b1;
  assign CLBLM_R_X5Y110_SLICE_X6Y110_C1 = CLBLM_L_X8Y110_SLICE_X10Y110_CO6;
  assign CLBLM_R_X5Y110_SLICE_X6Y110_C2 = CLBLM_R_X7Y110_SLICE_X8Y110_CO6;
  assign CLBLM_R_X5Y110_SLICE_X6Y110_C3 = CLBLM_R_X5Y112_SLICE_X6Y112_AO5;
  assign CLBLM_R_X5Y110_SLICE_X6Y110_C4 = CLBLM_R_X5Y111_SLICE_X6Y111_CO6;
  assign CLBLM_R_X5Y110_SLICE_X6Y110_C5 = CLBLM_R_X5Y110_SLICE_X6Y110_DO6;
  assign CLBLM_R_X5Y110_SLICE_X6Y110_C6 = CLBLM_R_X5Y110_SLICE_X6Y110_BO6;
  assign CLBLM_R_X5Y110_SLICE_X6Y110_D1 = 1'b1;
  assign CLBLM_R_X5Y110_SLICE_X6Y110_D2 = 1'b1;
  assign CLBLM_R_X5Y110_SLICE_X6Y110_D3 = CLBLM_R_X5Y108_SLICE_X6Y108_BO6;
  assign CLBLM_R_X5Y110_SLICE_X6Y110_D4 = 1'b1;
  assign CLBLM_R_X5Y110_SLICE_X6Y110_D5 = 1'b1;
  assign CLBLM_R_X5Y110_SLICE_X6Y110_D6 = CLBLM_R_X7Y107_SLICE_X8Y107_AO6;
  assign CLBLM_R_X5Y111_SLICE_X7Y111_A1 = RIOB33_X105Y109_IOB_X1Y109_I;
  assign CLBLM_R_X5Y111_SLICE_X7Y111_A2 = RIOB33_X105Y109_IOB_X1Y110_I;
  assign CLBLM_R_X5Y111_SLICE_X7Y111_A3 = LIOB33_X0Y111_IOB_X0Y111_I;
  assign CLBLM_R_X5Y111_SLICE_X7Y111_A4 = CLBLM_R_X7Y111_SLICE_X9Y111_AO5;
  assign CLBLM_R_X5Y111_SLICE_X7Y111_A5 = LIOB33_X0Y111_IOB_X0Y112_I;
  assign CLBLM_R_X5Y111_SLICE_X7Y111_A6 = CLBLM_R_X5Y111_SLICE_X7Y111_CO6;
  assign CLBLM_R_X5Y111_SLICE_X7Y111_B1 = LIOB33_X0Y113_IOB_X0Y113_I;
  assign CLBLM_R_X5Y111_SLICE_X7Y111_B2 = CLBLM_R_X7Y110_SLICE_X9Y110_AO5;
  assign CLBLM_R_X5Y111_SLICE_X7Y111_B3 = RIOB33_X105Y107_IOB_X1Y108_I;
  assign CLBLM_R_X5Y111_SLICE_X7Y111_B4 = LIOB33_X0Y111_IOB_X0Y112_I;
  assign CLBLM_R_X5Y111_SLICE_X7Y111_B5 = CLBLM_R_X7Y111_SLICE_X9Y111_AO6;
  assign CLBLM_R_X5Y111_SLICE_X7Y111_B6 = CLBLM_R_X5Y111_SLICE_X7Y111_AO6;
  assign CLBLM_R_X5Y111_SLICE_X7Y111_C1 = LIOB33_X0Y109_IOB_X0Y109_I;
  assign CLBLM_R_X5Y111_SLICE_X7Y111_C2 = CLBLM_R_X7Y111_SLICE_X9Y111_CO6;
  assign CLBLM_R_X5Y111_SLICE_X7Y111_C3 = LIOB33_X0Y109_IOB_X0Y110_I;
  assign CLBLM_R_X5Y111_SLICE_X7Y111_C4 = LIOB33_X0Y107_IOB_X0Y108_I;
  assign CLBLM_R_X5Y111_SLICE_X7Y111_C5 = RIOB33_X105Y109_IOB_X1Y110_I;
  assign CLBLM_R_X5Y111_SLICE_X7Y111_C6 = RIOB33_X105Y111_IOB_X1Y111_I;
  assign CLBLM_R_X5Y111_SLICE_X7Y111_D1 = CLBLM_R_X7Y111_SLICE_X9Y111_AO5;
  assign CLBLM_R_X5Y111_SLICE_X7Y111_D2 = LIOB33_X0Y111_IOB_X0Y111_I;
  assign CLBLM_R_X5Y111_SLICE_X7Y111_D3 = RIOB33_X105Y109_IOB_X1Y110_I;
  assign CLBLM_R_X5Y111_SLICE_X7Y111_D4 = CLBLM_R_X5Y111_SLICE_X7Y111_CO6;
  assign CLBLM_R_X5Y111_SLICE_X7Y111_D5 = RIOB33_X105Y109_IOB_X1Y109_I;
  assign CLBLM_R_X5Y111_SLICE_X7Y111_D6 = LIOB33_X0Y111_IOB_X0Y112_I;
  assign CLBLM_R_X5Y111_SLICE_X6Y111_A1 = LIOB33_X0Y113_IOB_X0Y113_I;
  assign CLBLM_R_X5Y111_SLICE_X6Y111_A2 = RIOB33_X105Y101_IOB_X1Y101_I;
  assign CLBLM_R_X5Y111_SLICE_X6Y111_A3 = CLBLM_R_X5Y110_SLICE_X7Y110_CO6;
  assign CLBLM_R_X5Y111_SLICE_X6Y111_A4 = RIOB33_X105Y101_IOB_X1Y102_I;
  assign CLBLM_R_X5Y111_SLICE_X6Y111_A5 = LIOB33_X0Y115_IOB_X0Y115_I;
  assign CLBLM_R_X5Y111_SLICE_X6Y111_A6 = CLBLM_R_X7Y112_SLICE_X8Y112_CO6;
  assign CLBLM_R_X5Y111_SLICE_X6Y111_B1 = LIOB33_X0Y113_IOB_X0Y113_I;
  assign CLBLM_R_X5Y111_SLICE_X6Y111_B2 = RIOB33_X105Y103_IOB_X1Y103_I;
  assign CLBLM_R_X5Y111_SLICE_X6Y111_B3 = CLBLM_R_X7Y111_SLICE_X8Y111_AO5;
  assign CLBLM_R_X5Y111_SLICE_X6Y111_B4 = CLBLM_L_X8Y113_SLICE_X10Y113_BO6;
  assign CLBLM_R_X5Y111_SLICE_X6Y111_B5 = LIOB33_X0Y111_IOB_X0Y112_I;
  assign CLBLM_R_X5Y111_SLICE_X6Y111_B6 = CLBLM_R_X5Y110_SLICE_X6Y110_AO5;
  assign CLBLM_R_X5Y111_SLICE_X6Y111_C1 = RIOB33_X105Y107_IOB_X1Y108_I;
  assign CLBLM_R_X5Y111_SLICE_X6Y111_C2 = CLBLM_R_X7Y111_SLICE_X9Y111_AO6;
  assign CLBLM_R_X5Y111_SLICE_X6Y111_C3 = CLBLM_R_X5Y111_SLICE_X7Y111_AO6;
  assign CLBLM_R_X5Y111_SLICE_X6Y111_C4 = CLBLM_R_X7Y110_SLICE_X9Y110_AO5;
  assign CLBLM_R_X5Y111_SLICE_X6Y111_C5 = LIOB33_X0Y113_IOB_X0Y113_I;
  assign CLBLM_R_X5Y111_SLICE_X6Y111_C6 = LIOB33_X0Y111_IOB_X0Y112_I;
  assign CLBLM_R_X5Y111_SLICE_X6Y111_D1 = LIOB33_X0Y111_IOB_X0Y112_I;
  assign CLBLM_R_X5Y111_SLICE_X6Y111_D2 = 1'b1;
  assign CLBLM_R_X5Y111_SLICE_X6Y111_D3 = CLBLM_R_X7Y111_SLICE_X8Y111_AO5;
  assign CLBLM_R_X5Y111_SLICE_X6Y111_D4 = CLBLM_R_X5Y110_SLICE_X6Y110_AO5;
  assign CLBLM_R_X5Y111_SLICE_X6Y111_D5 = RIOB33_X105Y103_IOB_X1Y103_I;
  assign CLBLM_R_X5Y111_SLICE_X6Y111_D6 = CLBLM_L_X8Y113_SLICE_X10Y113_BO6;
  assign CLBLM_R_X5Y112_SLICE_X7Y112_A1 = 1'b1;
  assign CLBLM_R_X5Y112_SLICE_X7Y112_A2 = LIOB33_X0Y115_IOB_X0Y115_I;
  assign CLBLM_R_X5Y112_SLICE_X7Y112_A3 = LIOB33_X0Y111_IOB_X0Y111_I;
  assign CLBLM_R_X5Y112_SLICE_X7Y112_A4 = RIOB33_X105Y101_IOB_X1Y102_I;
  assign CLBLM_R_X5Y112_SLICE_X7Y112_A5 = 1'b1;
  assign CLBLM_R_X5Y112_SLICE_X7Y112_A6 = 1'b1;
  assign CLBLM_R_X5Y112_SLICE_X7Y112_B1 = RIOB33_X105Y111_IOB_X1Y111_I;
  assign CLBLM_R_X5Y112_SLICE_X7Y112_B2 = LIOB33_X0Y109_IOB_X0Y109_I;
  assign CLBLM_R_X5Y112_SLICE_X7Y112_B3 = LIOB33_X0Y107_IOB_X0Y108_I;
  assign CLBLM_R_X5Y112_SLICE_X7Y112_B4 = RIOB33_X105Y109_IOB_X1Y110_I;
  assign CLBLM_R_X5Y112_SLICE_X7Y112_B5 = CLBLM_R_X7Y111_SLICE_X9Y111_CO6;
  assign CLBLM_R_X5Y112_SLICE_X7Y112_B6 = LIOB33_X0Y109_IOB_X0Y110_I;
  assign CLBLM_R_X5Y112_SLICE_X7Y112_C1 = LIOB33_X0Y111_IOB_X0Y111_I;
  assign CLBLM_R_X5Y112_SLICE_X7Y112_C2 = RIOB33_X105Y109_IOB_X1Y110_I;
  assign CLBLM_R_X5Y112_SLICE_X7Y112_C3 = LIOB33_X0Y113_IOB_X0Y113_I;
  assign CLBLM_R_X5Y112_SLICE_X7Y112_C4 = RIOB33_X105Y111_IOB_X1Y111_I;
  assign CLBLM_R_X5Y112_SLICE_X7Y112_C5 = CLBLM_R_X5Y112_SLICE_X7Y112_DO6;
  assign CLBLM_R_X5Y112_SLICE_X7Y112_C6 = LIOB33_X0Y111_IOB_X0Y112_I;
  assign CLBLM_R_X5Y112_SLICE_X7Y112_D1 = LIOB33_X0Y111_IOB_X0Y111_I;
  assign CLBLM_R_X5Y112_SLICE_X7Y112_D2 = LIOB33_X0Y109_IOB_X0Y110_I;
  assign CLBLM_R_X5Y112_SLICE_X7Y112_D3 = 1'b1;
  assign CLBLM_R_X5Y112_SLICE_X7Y112_D4 = RIOB33_X105Y109_IOB_X1Y110_I;
  assign CLBLM_R_X5Y112_SLICE_X7Y112_D5 = RIOB33_X105Y111_IOB_X1Y111_I;
  assign CLBLM_R_X5Y112_SLICE_X7Y112_D6 = CLBLM_R_X5Y112_SLICE_X7Y112_BO6;
  assign CLBLM_R_X5Y112_SLICE_X6Y112_A1 = CLBLM_R_X5Y111_SLICE_X6Y111_DO6;
  assign CLBLM_R_X5Y112_SLICE_X6Y112_A2 = RIOB33_X105Y103_IOB_X1Y103_I;
  assign CLBLM_R_X5Y112_SLICE_X6Y112_A3 = RIOB33_X105Y109_IOB_X1Y109_I;
  assign CLBLM_R_X5Y112_SLICE_X6Y112_A4 = LIOB33_X0Y113_IOB_X0Y113_I;
  assign CLBLM_R_X5Y112_SLICE_X6Y112_A5 = CLBLM_R_X5Y112_SLICE_X6Y112_CO6;
  assign CLBLM_R_X5Y112_SLICE_X6Y112_A6 = 1'b1;
  assign CLBLM_R_X5Y112_SLICE_X6Y112_B1 = CLBLM_R_X5Y111_SLICE_X6Y111_DO6;
  assign CLBLM_R_X5Y112_SLICE_X6Y112_B2 = LIOB33_X0Y113_IOB_X0Y113_I;
  assign CLBLM_R_X5Y112_SLICE_X6Y112_B3 = RIOB33_X105Y101_IOB_X1Y102_I;
  assign CLBLM_R_X5Y112_SLICE_X6Y112_B4 = LIOB33_X0Y115_IOB_X0Y115_I;
  assign CLBLM_R_X5Y112_SLICE_X6Y112_B5 = RIOB33_X105Y103_IOB_X1Y103_I;
  assign CLBLM_R_X5Y112_SLICE_X6Y112_B6 = CLBLM_R_X5Y110_SLICE_X7Y110_DO6;
  assign CLBLM_R_X5Y112_SLICE_X6Y112_C1 = LIOB33_X0Y111_IOB_X0Y111_I;
  assign CLBLM_R_X5Y112_SLICE_X6Y112_C2 = RIOB33_X105Y111_IOB_X1Y111_I;
  assign CLBLM_R_X5Y112_SLICE_X6Y112_C3 = CLBLM_R_X5Y112_SLICE_X7Y112_DO6;
  assign CLBLM_R_X5Y112_SLICE_X6Y112_C4 = CLBLM_R_X5Y111_SLICE_X7Y111_DO6;
  assign CLBLM_R_X5Y112_SLICE_X6Y112_C5 = RIOB33_X105Y109_IOB_X1Y110_I;
  assign CLBLM_R_X5Y112_SLICE_X6Y112_C6 = LIOB33_X0Y111_IOB_X0Y112_I;
  assign CLBLM_R_X5Y112_SLICE_X6Y112_D1 = 1'b1;
  assign CLBLM_R_X5Y112_SLICE_X6Y112_D2 = CLBLM_R_X5Y111_SLICE_X6Y111_CO6;
  assign CLBLM_R_X5Y112_SLICE_X6Y112_D3 = 1'b1;
  assign CLBLM_R_X5Y112_SLICE_X6Y112_D4 = CLBLM_R_X5Y112_SLICE_X6Y112_AO5;
  assign CLBLM_R_X5Y112_SLICE_X6Y112_D5 = 1'b1;
  assign CLBLM_R_X5Y112_SLICE_X6Y112_D6 = 1'b1;
  assign LIOI3_X0Y135_OLOGIC_X0Y136_D1 = CLBLL_L_X4Y110_SLICE_X5Y110_AO5;
  assign LIOI3_X0Y135_OLOGIC_X0Y136_T1 = 1'b1;
  assign LIOI3_X0Y135_OLOGIC_X0Y135_D1 = CLBLL_L_X4Y110_SLICE_X5Y110_AO6;
  assign LIOI3_X0Y135_OLOGIC_X0Y135_T1 = 1'b1;
  assign CLBLM_L_X8Y110_SLICE_X11Y110_C4 = RIOB33_X105Y101_IOB_X1Y101_I;
  assign CLBLM_L_X8Y110_SLICE_X11Y110_C5 = LIOB33_X0Y109_IOB_X0Y110_I;
  assign CLBLM_R_X5Y113_SLICE_X7Y113_A1 = RIOB33_X105Y103_IOB_X1Y104_I;
  assign CLBLM_R_X5Y113_SLICE_X7Y113_A2 = 1'b1;
  assign CLBLM_R_X5Y113_SLICE_X7Y113_A3 = LIOB33_X0Y113_IOB_X0Y113_I;
  assign CLBLM_R_X5Y113_SLICE_X7Y113_A4 = CLBLM_R_X7Y113_SLICE_X9Y113_AO6;
  assign CLBLM_R_X5Y113_SLICE_X7Y113_A5 = CLBLM_L_X8Y113_SLICE_X10Y113_CO6;
  assign CLBLM_R_X5Y113_SLICE_X7Y113_A6 = 1'b1;
  assign CLBLM_R_X5Y113_SLICE_X7Y113_B1 = CLBLM_R_X5Y110_SLICE_X6Y110_BO5;
  assign CLBLM_R_X5Y113_SLICE_X7Y113_B2 = LIOB33_X0Y115_IOB_X0Y115_I;
  assign CLBLM_R_X5Y113_SLICE_X7Y113_B3 = LIOB33_X0Y113_IOB_X0Y113_I;
  assign CLBLM_R_X5Y113_SLICE_X7Y113_B4 = CLBLM_R_X5Y112_SLICE_X7Y112_CO6;
  assign CLBLM_R_X5Y113_SLICE_X7Y113_B5 = RIOB33_X105Y109_IOB_X1Y109_I;
  assign CLBLM_R_X5Y113_SLICE_X7Y113_B6 = CLBLM_R_X5Y111_SLICE_X7Y111_DO6;
  assign CLBLM_R_X3Y103_SLICE_X3Y103_A1 = LIOB33_X0Y113_IOB_X0Y114_I;
  assign CLBLM_R_X3Y103_SLICE_X3Y103_A2 = CLBLM_R_X3Y103_SLICE_X2Y103_BO6;
  assign CLBLM_R_X3Y103_SLICE_X3Y103_A3 = CLBLM_R_X3Y103_SLICE_X2Y103_AO6;
  assign CLBLM_R_X3Y103_SLICE_X3Y103_A4 = CLBLM_R_X3Y103_SLICE_X3Y103_BO6;
  assign CLBLM_R_X3Y103_SLICE_X3Y103_A5 = LIOB33_X0Y101_IOB_X0Y101_I;
  assign CLBLM_R_X3Y103_SLICE_X3Y103_A6 = 1'b1;
  assign CLBLM_R_X5Y113_SLICE_X7Y113_C1 = RIOB33_X105Y109_IOB_X1Y109_I;
  assign CLBLM_R_X5Y113_SLICE_X7Y113_C2 = LIOB33_X0Y115_IOB_X0Y115_I;
  assign CLBLM_R_X5Y113_SLICE_X7Y113_C3 = CLBLM_R_X5Y110_SLICE_X6Y110_BO5;
  assign CLBLM_R_X3Y103_SLICE_X3Y103_B1 = LIOB33_SING_X0Y100_IOB_X0Y100_I;
  assign CLBLM_R_X3Y103_SLICE_X3Y103_B2 = 1'b1;
  assign CLBLM_R_X3Y103_SLICE_X3Y103_B3 = LIOB33_X0Y115_IOB_X0Y116_I;
  assign CLBLM_R_X3Y103_SLICE_X3Y103_B4 = LIOB33_X0Y113_IOB_X0Y114_I;
  assign CLBLM_R_X3Y103_SLICE_X3Y103_B5 = RIOB33_X105Y113_IOB_X1Y113_I;
  assign CLBLM_R_X3Y103_SLICE_X3Y103_B6 = RIOB33_X105Y111_IOB_X1Y112_I;
  assign CLBLM_R_X5Y113_SLICE_X7Y113_D1 = 1'b1;
  assign CLBLM_R_X5Y113_SLICE_X7Y113_D2 = 1'b1;
  assign CLBLM_R_X3Y103_SLICE_X3Y103_C1 = 1'b1;
  assign CLBLM_R_X3Y103_SLICE_X3Y103_C2 = 1'b1;
  assign CLBLM_R_X3Y103_SLICE_X3Y103_C3 = 1'b1;
  assign CLBLM_R_X3Y103_SLICE_X3Y103_C4 = 1'b1;
  assign CLBLM_R_X3Y103_SLICE_X3Y103_C5 = 1'b1;
  assign CLBLM_R_X3Y103_SLICE_X3Y103_C6 = 1'b1;
  assign CLBLM_R_X5Y113_SLICE_X7Y113_D3 = 1'b1;
  assign CLBLM_R_X5Y113_SLICE_X7Y113_D4 = 1'b1;
  assign CLBLM_R_X5Y113_SLICE_X6Y113_A1 = 1'b1;
  assign CLBLM_R_X5Y113_SLICE_X6Y113_A2 = 1'b1;
  assign CLBLM_R_X5Y113_SLICE_X6Y113_A3 = 1'b1;
  assign CLBLM_R_X5Y113_SLICE_X6Y113_A4 = 1'b1;
  assign CLBLM_R_X5Y113_SLICE_X6Y113_A5 = 1'b1;
  assign CLBLM_R_X5Y113_SLICE_X6Y113_A6 = 1'b1;
  assign CLBLM_R_X3Y103_SLICE_X3Y103_D1 = 1'b1;
  assign CLBLM_R_X3Y103_SLICE_X3Y103_D2 = 1'b1;
  assign CLBLM_R_X3Y103_SLICE_X3Y103_D3 = 1'b1;
  assign CLBLM_R_X3Y103_SLICE_X3Y103_D4 = 1'b1;
  assign CLBLM_R_X3Y103_SLICE_X3Y103_D5 = 1'b1;
  assign CLBLM_R_X3Y103_SLICE_X3Y103_D6 = 1'b1;
  assign CLBLM_R_X5Y113_SLICE_X6Y113_B1 = 1'b1;
  assign CLBLM_R_X5Y113_SLICE_X6Y113_B2 = 1'b1;
  assign CLBLM_R_X5Y113_SLICE_X6Y113_B3 = 1'b1;
  assign CLBLM_R_X11Y104_SLICE_X15Y104_B4 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X5Y113_SLICE_X6Y113_B4 = 1'b1;
  assign CLBLM_R_X5Y113_SLICE_X6Y113_B5 = 1'b1;
  assign CLBLM_R_X3Y103_SLICE_X2Y103_A1 = LIOB33_SING_X0Y100_IOB_X0Y100_I;
  assign CLBLM_R_X3Y103_SLICE_X2Y103_A2 = LIOB33_X0Y115_IOB_X0Y116_I;
  assign CLBLM_R_X3Y103_SLICE_X2Y103_A3 = RIOB33_X105Y113_IOB_X1Y113_I;
  assign CLBLM_R_X3Y103_SLICE_X2Y103_A4 = LIOB33_X0Y113_IOB_X0Y114_I;
  assign CLBLM_R_X3Y103_SLICE_X2Y103_A5 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLM_R_X3Y103_SLICE_X2Y103_A6 = RIOB33_X105Y111_IOB_X1Y112_I;
  assign CLBLM_R_X5Y113_SLICE_X6Y113_C1 = 1'b1;
  assign CLBLM_R_X5Y113_SLICE_X6Y113_C2 = 1'b1;
  assign CLBLM_R_X5Y113_SLICE_X6Y113_C3 = 1'b1;
  assign CLBLM_R_X3Y103_SLICE_X2Y103_B1 = LIOB33_SING_X0Y100_IOB_X0Y100_I;
  assign CLBLM_R_X3Y103_SLICE_X2Y103_B2 = RIOB33_X105Y113_IOB_X1Y113_I;
  assign CLBLM_R_X3Y103_SLICE_X2Y103_B3 = LIOB33_X0Y115_IOB_X0Y116_I;
  assign CLBLM_R_X3Y103_SLICE_X2Y103_B4 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLM_R_X3Y103_SLICE_X2Y103_B5 = 1'b1;
  assign CLBLM_R_X3Y103_SLICE_X2Y103_B6 = RIOB33_X105Y111_IOB_X1Y112_I;
  assign CLBLM_R_X5Y113_SLICE_X6Y113_D1 = 1'b1;
  assign CLBLM_R_X5Y113_SLICE_X6Y113_D2 = 1'b1;
  assign CLBLM_R_X5Y113_SLICE_X6Y113_D3 = 1'b1;
  assign CLBLM_R_X3Y103_SLICE_X2Y103_C1 = 1'b1;
  assign CLBLM_R_X3Y103_SLICE_X2Y103_C2 = 1'b1;
  assign CLBLM_R_X3Y103_SLICE_X2Y103_C3 = 1'b1;
  assign CLBLM_R_X3Y103_SLICE_X2Y103_C4 = 1'b1;
  assign CLBLM_R_X3Y103_SLICE_X2Y103_C5 = 1'b1;
  assign CLBLM_R_X3Y103_SLICE_X2Y103_C6 = 1'b1;
  assign CLBLM_R_X5Y113_SLICE_X6Y113_D4 = 1'b1;
  assign CLBLM_R_X5Y113_SLICE_X6Y113_D5 = 1'b1;
  assign CLBLM_R_X5Y113_SLICE_X6Y113_D6 = 1'b1;
  assign CLBLM_R_X3Y103_SLICE_X2Y103_D1 = 1'b1;
  assign CLBLM_R_X3Y103_SLICE_X2Y103_D2 = 1'b1;
  assign CLBLM_R_X3Y103_SLICE_X2Y103_D3 = 1'b1;
  assign CLBLM_R_X3Y103_SLICE_X2Y103_D4 = 1'b1;
  assign CLBLM_R_X3Y103_SLICE_X2Y103_D5 = 1'b1;
  assign CLBLM_R_X3Y103_SLICE_X2Y103_D6 = 1'b1;
  assign CLBLM_R_X11Y104_SLICE_X15Y104_C3 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X11Y104_SLICE_X15Y104_C4 = RIOB33_X105Y107_IOB_X1Y107_I;
  assign CLBLM_R_X11Y104_SLICE_X15Y104_C5 = RIOB33_X105Y111_IOB_X1Y112_I;
  assign CLBLM_R_X11Y104_SLICE_X15Y104_C6 = RIOB33_X105Y107_IOB_X1Y108_I;
  assign CLBLM_R_X7Y106_SLICE_X9Y106_B3 = CLBLM_R_X7Y106_SLICE_X8Y106_CO6;
  assign CLBLM_R_X7Y106_SLICE_X9Y106_C1 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLM_R_X7Y106_SLICE_X9Y106_C2 = CLBLM_L_X8Y106_SLICE_X11Y106_AO6;
  assign CLBLM_R_X3Y104_SLICE_X3Y104_A1 = 1'b1;
  assign CLBLM_R_X3Y104_SLICE_X3Y104_A2 = RIOB33_X105Y105_IOB_X1Y106_I;
  assign CLBLM_R_X3Y104_SLICE_X3Y104_A3 = LIOB33_X0Y101_IOB_X0Y102_I;
  assign CLBLM_R_X3Y104_SLICE_X3Y104_A4 = 1'b1;
  assign CLBLM_R_X3Y104_SLICE_X3Y104_A5 = LIOB33_X0Y103_IOB_X0Y103_I;
  assign CLBLM_R_X3Y104_SLICE_X3Y104_A6 = 1'b1;
  assign CLBLM_R_X3Y104_SLICE_X3Y104_B1 = LIOB33_X0Y101_IOB_X0Y102_I;
  assign CLBLM_R_X3Y104_SLICE_X3Y104_B2 = CLBLM_R_X3Y104_SLICE_X2Y104_BO6;
  assign CLBLM_R_X3Y104_SLICE_X3Y104_B3 = LIOB33_X0Y103_IOB_X0Y103_I;
  assign CLBLM_R_X3Y104_SLICE_X3Y104_B4 = RIOB33_X105Y105_IOB_X1Y106_I;
  assign CLBLM_R_X3Y104_SLICE_X3Y104_B5 = LIOB33_X0Y103_IOB_X0Y104_I;
  assign CLBLM_R_X3Y104_SLICE_X3Y104_B6 = CLBLM_R_X3Y104_SLICE_X3Y104_CO6;
  assign CLBLM_R_X7Y106_SLICE_X9Y106_D1 = CLBLM_R_X7Y105_SLICE_X8Y105_BO6;
  assign CLBLM_R_X3Y104_SLICE_X3Y104_C1 = CLBLM_R_X3Y105_SLICE_X2Y105_AO6;
  assign CLBLM_R_X3Y104_SLICE_X3Y104_C2 = CLBLL_L_X2Y104_SLICE_X0Y104_BO6;
  assign CLBLM_R_X3Y104_SLICE_X3Y104_C3 = CLBLL_L_X2Y104_SLICE_X0Y104_CO6;
  assign CLBLM_R_X3Y104_SLICE_X3Y104_C4 = CLBLM_R_X3Y104_SLICE_X3Y104_AO5;
  assign CLBLM_R_X3Y104_SLICE_X3Y104_C5 = CLBLL_L_X4Y103_SLICE_X4Y103_AO6;
  assign CLBLM_R_X3Y104_SLICE_X3Y104_C6 = CLBLM_R_X13Y106_SLICE_X18Y106_AO5;
  assign CLBLM_R_X3Y104_SLICE_X3Y104_D1 = CLBLM_R_X3Y104_SLICE_X3Y104_AO6;
  assign CLBLM_R_X3Y104_SLICE_X3Y104_D2 = CLBLM_R_X3Y104_SLICE_X2Y104_CO6;
  assign CLBLM_R_X3Y104_SLICE_X3Y104_D3 = CLBLM_R_X3Y106_SLICE_X2Y106_BO5;
  assign CLBLM_R_X3Y104_SLICE_X3Y104_D4 = CLBLM_R_X3Y105_SLICE_X2Y105_AO6;
  assign CLBLM_R_X3Y104_SLICE_X3Y104_D5 = CLBLL_L_X4Y103_SLICE_X4Y103_AO6;
  assign CLBLM_R_X3Y104_SLICE_X3Y104_D6 = CLBLM_R_X3Y103_SLICE_X2Y103_AO6;
  assign CLBLM_R_X3Y104_SLICE_X2Y104_A1 = LIOB33_X0Y103_IOB_X0Y103_I;
  assign CLBLM_R_X3Y104_SLICE_X2Y104_A2 = CLBLM_R_X3Y104_SLICE_X2Y104_CO6;
  assign CLBLM_R_X3Y104_SLICE_X2Y104_A3 = CLBLM_R_X3Y105_SLICE_X2Y105_AO6;
  assign CLBLM_R_X3Y104_SLICE_X2Y104_A4 = 1'b1;
  assign CLBLM_R_X3Y104_SLICE_X2Y104_A5 = LIOB33_X0Y101_IOB_X0Y101_I;
  assign CLBLM_R_X3Y104_SLICE_X2Y104_A6 = 1'b1;
  assign CLBLM_R_X3Y104_SLICE_X2Y104_B1 = LIOB33_X0Y103_IOB_X0Y103_I;
  assign CLBLM_R_X3Y104_SLICE_X2Y104_B2 = CLBLM_R_X3Y103_SLICE_X2Y103_AO6;
  assign CLBLM_R_X3Y104_SLICE_X2Y104_B3 = LIOB33_X0Y101_IOB_X0Y101_I;
  assign CLBLM_R_X3Y104_SLICE_X2Y104_B4 = LIOB33_X0Y113_IOB_X0Y114_I;
  assign CLBLM_R_X3Y104_SLICE_X2Y104_B5 = CLBLM_R_X3Y105_SLICE_X2Y105_AO6;
  assign CLBLM_R_X3Y104_SLICE_X2Y104_B6 = CLBLM_R_X3Y104_SLICE_X2Y104_CO6;
  assign CLBLM_R_X3Y104_SLICE_X2Y104_C1 = LIOB33_X0Y103_IOB_X0Y103_I;
  assign CLBLM_R_X3Y104_SLICE_X2Y104_C2 = RIOB33_X105Y113_IOB_X1Y113_I;
  assign CLBLM_R_X3Y104_SLICE_X2Y104_C3 = LIOB33_SING_X0Y100_IOB_X0Y100_I;
  assign CLBLM_R_X3Y104_SLICE_X2Y104_C4 = LIOB33_X0Y113_IOB_X0Y114_I;
  assign CLBLM_R_X3Y104_SLICE_X2Y104_C5 = LIOB33_X0Y115_IOB_X0Y116_I;
  assign CLBLM_R_X3Y104_SLICE_X2Y104_C6 = RIOB33_X105Y111_IOB_X1Y112_I;
  assign CLBLM_R_X3Y104_SLICE_X2Y104_D1 = CLBLM_R_X3Y103_SLICE_X3Y103_AO6;
  assign CLBLM_R_X3Y104_SLICE_X2Y104_D2 = LIOB33_X0Y103_IOB_X0Y103_I;
  assign CLBLM_R_X3Y104_SLICE_X2Y104_D3 = LIOB33_X0Y101_IOB_X0Y102_I;
  assign CLBLM_R_X3Y104_SLICE_X2Y104_D4 = CLBLM_R_X3Y104_SLICE_X2Y104_AO5;
  assign CLBLM_R_X3Y104_SLICE_X2Y104_D5 = CLBLL_L_X4Y103_SLICE_X4Y103_BO6;
  assign CLBLM_R_X3Y104_SLICE_X2Y104_D6 = LIOB33_X0Y113_IOB_X0Y114_I;
  assign LIOB33_SING_X0Y149_IOB_X0Y149_O = CLBLM_R_X3Y112_SLICE_X2Y112_DO6;
  assign LIOI3_X0Y139_OLOGIC_X0Y140_D1 = CLBLL_L_X4Y112_SLICE_X4Y112_AO5;
  assign LIOI3_X0Y139_OLOGIC_X0Y140_T1 = 1'b1;
  assign LIOI3_X0Y139_OLOGIC_X0Y139_D1 = CLBLL_L_X4Y112_SLICE_X4Y112_AO6;
  assign LIOI3_X0Y139_OLOGIC_X0Y139_T1 = 1'b1;
  assign CLBLM_R_X3Y105_SLICE_X3Y105_A1 = 1'b1;
  assign CLBLM_R_X3Y105_SLICE_X3Y105_A2 = 1'b1;
  assign CLBLM_R_X3Y105_SLICE_X3Y105_A3 = 1'b1;
  assign CLBLM_R_X3Y105_SLICE_X3Y105_A4 = 1'b1;
  assign CLBLM_R_X3Y105_SLICE_X3Y105_A5 = 1'b1;
  assign CLBLM_R_X3Y105_SLICE_X3Y105_A6 = 1'b1;
  assign CLBLM_R_X3Y105_SLICE_X3Y105_B1 = 1'b1;
  assign CLBLM_R_X3Y105_SLICE_X3Y105_B2 = 1'b1;
  assign CLBLM_R_X3Y105_SLICE_X3Y105_B3 = 1'b1;
  assign CLBLM_R_X3Y105_SLICE_X3Y105_B4 = 1'b1;
  assign CLBLM_R_X3Y105_SLICE_X3Y105_B5 = 1'b1;
  assign CLBLM_R_X3Y105_SLICE_X3Y105_B6 = 1'b1;
  assign CLBLM_R_X3Y105_SLICE_X3Y105_C1 = 1'b1;
  assign CLBLM_R_X3Y105_SLICE_X3Y105_C2 = 1'b1;
  assign CLBLM_R_X3Y105_SLICE_X3Y105_C3 = 1'b1;
  assign CLBLM_R_X3Y105_SLICE_X3Y105_C4 = 1'b1;
  assign CLBLM_R_X3Y105_SLICE_X3Y105_C5 = 1'b1;
  assign CLBLM_R_X3Y105_SLICE_X3Y105_C6 = 1'b1;
  assign CLBLM_R_X3Y105_SLICE_X3Y105_D1 = 1'b1;
  assign CLBLM_R_X3Y105_SLICE_X3Y105_D2 = 1'b1;
  assign CLBLM_R_X3Y105_SLICE_X3Y105_D3 = 1'b1;
  assign CLBLM_R_X3Y105_SLICE_X3Y105_D4 = 1'b1;
  assign CLBLM_R_X3Y105_SLICE_X3Y105_D5 = 1'b1;
  assign CLBLM_R_X3Y105_SLICE_X3Y105_D6 = 1'b1;
  assign LIOB33_X0Y117_IOB_X0Y118_O = CLBLL_L_X2Y109_SLICE_X0Y109_AO5;
  assign CLBLM_R_X3Y105_SLICE_X2Y105_A1 = LIOB33_SING_X0Y100_IOB_X0Y100_I;
  assign CLBLM_R_X3Y105_SLICE_X2Y105_A2 = LIOB33_X0Y113_IOB_X0Y114_I;
  assign CLBLM_R_X3Y105_SLICE_X2Y105_A3 = LIOB33_X0Y103_IOB_X0Y103_I;
  assign CLBLM_R_X3Y105_SLICE_X2Y105_A4 = RIOB33_X105Y113_IOB_X1Y113_I;
  assign CLBLM_R_X3Y105_SLICE_X2Y105_A5 = LIOB33_X0Y115_IOB_X0Y116_I;
  assign CLBLM_R_X3Y105_SLICE_X2Y105_A6 = RIOB33_X105Y111_IOB_X1Y112_I;
  assign CLBLM_R_X3Y105_SLICE_X2Y105_B1 = RIOB33_X105Y105_IOB_X1Y106_I;
  assign CLBLM_R_X3Y105_SLICE_X2Y105_B2 = LIOB33_X0Y103_IOB_X0Y104_I;
  assign CLBLM_R_X3Y105_SLICE_X2Y105_B3 = LIOB33_X0Y103_IOB_X0Y103_I;
  assign CLBLM_R_X3Y105_SLICE_X2Y105_B4 = CLBLM_R_X3Y104_SLICE_X2Y104_DO6;
  assign CLBLM_R_X3Y105_SLICE_X2Y105_B5 = CLBLM_R_X3Y104_SLICE_X3Y104_BO6;
  assign CLBLM_R_X3Y105_SLICE_X2Y105_B6 = LIOB33_X0Y105_IOB_X0Y105_I;
  assign CLBLM_R_X3Y105_SLICE_X2Y105_C1 = LIOB33_X0Y103_IOB_X0Y103_I;
  assign CLBLM_R_X3Y105_SLICE_X2Y105_C2 = RIOB33_X105Y105_IOB_X1Y106_I;
  assign CLBLM_R_X3Y105_SLICE_X2Y105_C3 = LIOB33_X0Y103_IOB_X0Y104_I;
  assign CLBLM_R_X3Y105_SLICE_X2Y105_C4 = CLBLM_R_X3Y104_SLICE_X2Y104_DO6;
  assign CLBLM_R_X3Y105_SLICE_X2Y105_C5 = CLBLM_R_X3Y104_SLICE_X3Y104_BO6;
  assign CLBLM_R_X3Y105_SLICE_X2Y105_C6 = LIOB33_X0Y105_IOB_X0Y105_I;
  assign CLBLM_R_X3Y105_SLICE_X2Y105_D1 = 1'b1;
  assign CLBLM_R_X3Y105_SLICE_X2Y105_D2 = 1'b1;
  assign CLBLM_R_X3Y105_SLICE_X2Y105_D3 = 1'b1;
  assign CLBLM_R_X3Y105_SLICE_X2Y105_D4 = 1'b1;
  assign CLBLM_R_X3Y105_SLICE_X2Y105_D5 = 1'b1;
  assign CLBLM_R_X3Y105_SLICE_X2Y105_D6 = 1'b1;
  assign RIOI3_TBYTESRC_X105Y107_ILOGIC_X1Y108_D = RIOB33_X105Y107_IOB_X1Y108_I;
  assign RIOI3_TBYTESRC_X105Y107_ILOGIC_X1Y107_D = RIOB33_X105Y107_IOB_X1Y107_I;
  assign CLBLM_R_X3Y106_SLICE_X3Y106_A1 = 1'b1;
  assign CLBLM_R_X3Y106_SLICE_X3Y106_A2 = RIOB33_X105Y105_IOB_X1Y106_I;
  assign CLBLM_R_X3Y106_SLICE_X3Y106_A3 = LIOB33_X0Y103_IOB_X0Y103_I;
  assign CLBLM_R_X3Y106_SLICE_X3Y106_A4 = LIOB33_X0Y105_IOB_X0Y105_I;
  assign CLBLM_R_X3Y106_SLICE_X3Y106_A5 = 1'b1;
  assign CLBLM_R_X3Y106_SLICE_X3Y106_A6 = 1'b1;
  assign LIOB33_X0Y119_IOB_X0Y119_O = CLBLL_L_X2Y109_SLICE_X0Y109_AO6;
  assign LIOB33_X0Y119_IOB_X0Y120_O = CLBLM_R_X3Y106_SLICE_X2Y106_AO5;
  assign CLBLM_R_X3Y106_SLICE_X3Y106_B1 = CLBLL_L_X4Y105_SLICE_X4Y105_AO6;
  assign CLBLM_R_X3Y106_SLICE_X3Y106_B2 = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLM_R_X3Y106_SLICE_X3Y106_B3 = LIOB33_X0Y103_IOB_X0Y103_I;
  assign CLBLM_R_X3Y106_SLICE_X3Y106_B4 = CLBLL_L_X4Y106_SLICE_X4Y106_AO6;
  assign CLBLM_R_X3Y106_SLICE_X3Y106_B5 = RIOB33_X105Y105_IOB_X1Y106_I;
  assign CLBLM_R_X3Y106_SLICE_X3Y106_B6 = CLBLM_R_X3Y105_SLICE_X2Y105_CO6;
  assign CLBLM_R_X3Y106_SLICE_X3Y106_C1 = CLBLM_R_X3Y106_SLICE_X3Y106_AO6;
  assign CLBLM_R_X3Y106_SLICE_X3Y106_C2 = CLBLL_L_X4Y104_SLICE_X4Y104_BO6;
  assign CLBLM_R_X3Y106_SLICE_X3Y106_C3 = CLBLM_R_X3Y107_SLICE_X2Y107_AO5;
  assign CLBLM_R_X3Y106_SLICE_X3Y106_C4 = CLBLM_R_X3Y106_SLICE_X3Y106_AO5;
  assign CLBLM_R_X3Y106_SLICE_X3Y106_C5 = CLBLL_L_X4Y104_SLICE_X4Y104_AO6;
  assign CLBLM_R_X3Y106_SLICE_X3Y106_C6 = CLBLM_R_X3Y104_SLICE_X3Y104_BO6;
  assign CLBLM_R_X3Y106_SLICE_X3Y106_D1 = CLBLM_R_X3Y106_SLICE_X3Y106_AO6;
  assign CLBLM_R_X3Y106_SLICE_X3Y106_D2 = CLBLL_L_X4Y104_SLICE_X4Y104_BO6;
  assign CLBLM_R_X3Y106_SLICE_X3Y106_D3 = CLBLM_R_X3Y107_SLICE_X2Y107_AO5;
  assign CLBLM_R_X3Y106_SLICE_X3Y106_D4 = CLBLM_R_X3Y106_SLICE_X3Y106_AO5;
  assign CLBLM_R_X3Y106_SLICE_X3Y106_D5 = CLBLL_L_X4Y104_SLICE_X4Y104_AO6;
  assign CLBLM_R_X3Y106_SLICE_X3Y106_D6 = CLBLM_R_X3Y104_SLICE_X3Y104_BO6;
  assign CLBLM_R_X3Y106_SLICE_X2Y106_A1 = RIOB33_SING_X105Y100_IOB_X1Y100_I;
  assign CLBLM_R_X3Y106_SLICE_X2Y106_A2 = CLBLL_L_X2Y106_SLICE_X1Y106_BO6;
  assign CLBLM_R_X3Y106_SLICE_X2Y106_A3 = CLBLM_R_X3Y103_SLICE_X2Y103_BO6;
  assign CLBLM_R_X3Y106_SLICE_X2Y106_A4 = CLBLM_R_X3Y106_SLICE_X2Y106_BO6;
  assign CLBLM_R_X3Y106_SLICE_X2Y106_A5 = LIOB33_X0Y101_IOB_X0Y101_I;
  assign CLBLM_R_X3Y106_SLICE_X2Y106_A6 = 1'b1;
  assign CLBLM_R_X3Y106_SLICE_X2Y106_B1 = RIOB33_X105Y113_IOB_X1Y113_I;
  assign CLBLM_R_X3Y106_SLICE_X2Y106_B2 = LIOB33_X0Y113_IOB_X0Y114_I;
  assign CLBLM_R_X3Y106_SLICE_X2Y106_B3 = LIOB33_X0Y103_IOB_X0Y103_I;
  assign CLBLM_R_X3Y106_SLICE_X2Y106_B4 = RIOB33_X105Y111_IOB_X1Y112_I;
  assign CLBLM_R_X3Y106_SLICE_X2Y106_B5 = LIOB33_X0Y101_IOB_X0Y101_I;
  assign CLBLM_R_X3Y106_SLICE_X2Y106_B6 = 1'b1;
  assign CLBLM_R_X3Y106_SLICE_X2Y106_C1 = LIOB33_X0Y103_IOB_X0Y103_I;
  assign CLBLM_R_X3Y106_SLICE_X2Y106_C2 = RIOB33_X105Y113_IOB_X1Y113_I;
  assign CLBLM_R_X3Y106_SLICE_X2Y106_C3 = LIOB33_SING_X0Y100_IOB_X0Y100_I;
  assign CLBLM_R_X3Y106_SLICE_X2Y106_C4 = RIOB33_X105Y111_IOB_X1Y112_I;
  assign CLBLM_R_X3Y106_SLICE_X2Y106_C5 = RIOB33_SING_X105Y100_IOB_X1Y100_I;
  assign CLBLM_R_X3Y106_SLICE_X2Y106_C6 = RIOB33_X105Y105_IOB_X1Y106_I;
  assign CLBLM_R_X3Y106_SLICE_X2Y106_D1 = LIOB33_X0Y103_IOB_X0Y103_I;
  assign CLBLM_R_X3Y106_SLICE_X2Y106_D2 = CLBLL_L_X4Y104_SLICE_X4Y104_AO6;
  assign CLBLM_R_X3Y106_SLICE_X2Y106_D3 = CLBLL_L_X4Y104_SLICE_X4Y104_BO6;
  assign CLBLM_R_X3Y106_SLICE_X2Y106_D4 = RIOB33_X105Y105_IOB_X1Y106_I;
  assign CLBLM_R_X3Y106_SLICE_X2Y106_D5 = CLBLM_R_X3Y104_SLICE_X3Y104_BO6;
  assign CLBLM_R_X3Y106_SLICE_X2Y106_D6 = LIOB33_X0Y105_IOB_X0Y105_I;
  assign LIOB33_X0Y121_IOB_X0Y122_O = CLBLL_L_X2Y104_SLICE_X0Y104_AO6;
  assign LIOB33_X0Y121_IOB_X0Y121_O = CLBLL_L_X2Y106_SLICE_X0Y106_AO5;
  assign CLBLM_R_X3Y107_SLICE_X3Y107_A1 = RIOB33_SING_X105Y100_IOB_X1Y100_I;
  assign CLBLM_R_X3Y107_SLICE_X3Y107_A2 = CLBLL_L_X4Y107_SLICE_X4Y107_AO6;
  assign CLBLM_R_X3Y107_SLICE_X3Y107_A3 = RIOB33_X105Y105_IOB_X1Y106_I;
  assign CLBLM_R_X3Y107_SLICE_X3Y107_A4 = LIOB33_X0Y109_IOB_X0Y109_I;
  assign CLBLM_R_X3Y107_SLICE_X3Y107_A5 = CLBLM_R_X3Y107_SLICE_X3Y107_CO6;
  assign CLBLM_R_X3Y107_SLICE_X3Y107_A6 = 1'b1;
  assign CLBLM_R_X3Y107_SLICE_X3Y107_B1 = CLBLM_R_X3Y107_SLICE_X3Y107_DO6;
  assign CLBLM_R_X3Y107_SLICE_X3Y107_B2 = RIOB33_X105Y105_IOB_X1Y106_I;
  assign CLBLM_R_X3Y107_SLICE_X3Y107_B3 = RIOB33_SING_X105Y100_IOB_X1Y100_I;
  assign CLBLM_R_X3Y107_SLICE_X3Y107_B4 = 1'b1;
  assign CLBLM_R_X3Y107_SLICE_X3Y107_B5 = LIOB33_X0Y109_IOB_X0Y110_I;
  assign CLBLM_R_X3Y107_SLICE_X3Y107_B6 = 1'b1;
  assign LIOI3_X0Y141_OLOGIC_X0Y142_D1 = CLBLL_L_X4Y114_SLICE_X4Y114_DO6;
  assign LIOI3_X0Y103_ILOGIC_X0Y104_D = LIOB33_X0Y103_IOB_X0Y104_I;
  assign CLBLM_R_X3Y107_SLICE_X3Y107_C1 = RIOB33_X105Y105_IOB_X1Y106_I;
  assign CLBLM_R_X3Y107_SLICE_X3Y107_C2 = LIOB33_X0Y107_IOB_X0Y107_I;
  assign CLBLM_R_X3Y107_SLICE_X3Y107_C3 = CLBLM_R_X3Y107_SLICE_X2Y107_DO6;
  assign CLBLM_R_X3Y107_SLICE_X3Y107_C4 = RIOB33_SING_X105Y100_IOB_X1Y100_I;
  assign CLBLM_R_X3Y107_SLICE_X3Y107_C5 = LIOB33_X0Y107_IOB_X0Y108_I;
  assign CLBLM_R_X3Y107_SLICE_X3Y107_C6 = CLBLM_R_X3Y106_SLICE_X3Y106_BO6;
  assign LIOI3_X0Y141_OLOGIC_X0Y142_T1 = 1'b1;
  assign CLBLM_R_X3Y107_SLICE_X3Y107_D1 = LIOB33_X0Y109_IOB_X0Y109_I;
  assign CLBLM_R_X3Y107_SLICE_X3Y107_D2 = CLBLL_L_X4Y107_SLICE_X5Y107_BO6;
  assign CLBLM_R_X3Y107_SLICE_X3Y107_D3 = RIOB33_X105Y105_IOB_X1Y106_I;
  assign CLBLM_R_X3Y107_SLICE_X3Y107_D4 = CLBLM_R_X3Y107_SLICE_X3Y107_CO6;
  assign CLBLM_R_X3Y107_SLICE_X3Y107_D5 = RIOB33_SING_X105Y100_IOB_X1Y100_I;
  assign CLBLM_R_X3Y107_SLICE_X3Y107_D6 = CLBLL_L_X4Y107_SLICE_X4Y107_AO6;
  assign LIOI3_X0Y103_ILOGIC_X0Y103_D = LIOB33_X0Y103_IOB_X0Y103_I;
  assign LIOI3_X0Y141_OLOGIC_X0Y141_D1 = CLBLL_L_X4Y112_SLICE_X5Y112_DO6;
  assign CLBLM_R_X3Y107_SLICE_X2Y107_A1 = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLM_R_X3Y107_SLICE_X2Y107_A2 = CLBLM_R_X3Y105_SLICE_X2Y105_BO6;
  assign CLBLM_R_X3Y107_SLICE_X2Y107_A3 = CLBLL_L_X2Y107_SLICE_X0Y107_BO6;
  assign CLBLM_R_X3Y107_SLICE_X2Y107_A4 = RIOB33_X105Y105_IOB_X1Y106_I;
  assign CLBLM_R_X3Y107_SLICE_X2Y107_A5 = RIOB33_SING_X105Y100_IOB_X1Y100_I;
  assign CLBLM_R_X3Y107_SLICE_X2Y107_A6 = 1'b1;
  assign LIOI3_X0Y141_OLOGIC_X0Y141_T1 = 1'b1;
  assign CLBLM_R_X3Y107_SLICE_X2Y107_B1 = RIOB33_SING_X105Y100_IOB_X1Y100_I;
  assign CLBLM_R_X3Y107_SLICE_X2Y107_B2 = CLBLM_R_X3Y105_SLICE_X2Y105_BO6;
  assign CLBLM_R_X3Y107_SLICE_X2Y107_B3 = CLBLL_L_X2Y107_SLICE_X0Y107_BO6;
  assign CLBLM_R_X3Y107_SLICE_X2Y107_B4 = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLM_R_X3Y107_SLICE_X2Y107_B5 = RIOB33_X105Y105_IOB_X1Y106_I;
  assign CLBLM_R_X3Y107_SLICE_X2Y107_B6 = CLBLM_R_X3Y106_SLICE_X2Y106_DO6;
  assign CLBLM_R_X3Y107_SLICE_X2Y107_C1 = RIOB33_X105Y105_IOB_X1Y106_I;
  assign CLBLM_R_X3Y107_SLICE_X2Y107_C2 = RIOB33_SING_X105Y100_IOB_X1Y100_I;
  assign CLBLM_R_X3Y107_SLICE_X2Y107_C3 = LIOB33_X0Y107_IOB_X0Y108_I;
  assign CLBLM_R_X3Y107_SLICE_X2Y107_C4 = CLBLM_R_X3Y106_SLICE_X3Y106_BO6;
  assign CLBLM_R_X3Y107_SLICE_X2Y107_C5 = CLBLM_R_X3Y107_SLICE_X2Y107_DO6;
  assign CLBLM_R_X3Y107_SLICE_X2Y107_C6 = LIOB33_X0Y107_IOB_X0Y107_I;
  assign CLBLM_R_X3Y107_SLICE_X2Y107_D1 = CLBLL_L_X2Y107_SLICE_X0Y107_BO6;
  assign CLBLM_R_X3Y107_SLICE_X2Y107_D2 = CLBLM_R_X3Y106_SLICE_X3Y106_CO6;
  assign CLBLM_R_X3Y107_SLICE_X2Y107_D3 = RIOB33_SING_X105Y100_IOB_X1Y100_I;
  assign CLBLM_R_X3Y107_SLICE_X2Y107_D4 = CLBLM_R_X3Y105_SLICE_X2Y105_BO6;
  assign CLBLM_R_X3Y107_SLICE_X2Y107_D5 = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLM_R_X3Y107_SLICE_X2Y107_D6 = LIOB33_X0Y107_IOB_X0Y107_I;
  assign LIOB33_X0Y123_IOB_X0Y124_O = CLBLM_R_X3Y107_SLICE_X2Y107_AO6;
  assign LIOB33_X0Y123_IOB_X0Y123_O = CLBLL_L_X2Y107_SLICE_X0Y107_AO6;
  assign CLBLM_R_X3Y108_SLICE_X3Y108_A1 = LIOB33_X0Y111_IOB_X0Y111_I;
  assign CLBLM_R_X3Y108_SLICE_X3Y108_A2 = CLBLM_R_X5Y107_SLICE_X6Y107_AO6;
  assign CLBLM_R_X3Y108_SLICE_X3Y108_A3 = RIOB33_X105Y105_IOB_X1Y106_I;
  assign CLBLM_R_X3Y108_SLICE_X3Y108_A4 = LIOB33_X0Y109_IOB_X0Y110_I;
  assign CLBLM_R_X3Y108_SLICE_X3Y108_A5 = RIOB33_SING_X105Y100_IOB_X1Y100_I;
  assign CLBLM_R_X3Y108_SLICE_X3Y108_A6 = CLBLL_L_X4Y107_SLICE_X4Y107_BO6;
  assign CLBLM_R_X3Y108_SLICE_X3Y108_B1 = 1'b1;
  assign CLBLM_R_X3Y108_SLICE_X3Y108_B2 = 1'b1;
  assign CLBLM_R_X3Y108_SLICE_X3Y108_B3 = 1'b1;
  assign CLBLM_R_X3Y108_SLICE_X3Y108_B4 = 1'b1;
  assign CLBLM_R_X3Y108_SLICE_X3Y108_B5 = 1'b1;
  assign CLBLM_R_X3Y108_SLICE_X3Y108_B6 = 1'b1;
  assign CLBLM_R_X3Y108_SLICE_X3Y108_C1 = 1'b1;
  assign CLBLM_R_X3Y108_SLICE_X3Y108_C2 = 1'b1;
  assign CLBLM_R_X3Y108_SLICE_X3Y108_C3 = 1'b1;
  assign CLBLM_R_X3Y108_SLICE_X3Y108_C4 = 1'b1;
  assign CLBLM_R_X3Y108_SLICE_X3Y108_C5 = 1'b1;
  assign CLBLM_R_X3Y108_SLICE_X3Y108_C6 = 1'b1;
  assign CLBLM_R_X3Y108_SLICE_X3Y108_D1 = 1'b1;
  assign CLBLM_R_X3Y108_SLICE_X3Y108_D2 = 1'b1;
  assign CLBLM_R_X3Y108_SLICE_X3Y108_D3 = 1'b1;
  assign CLBLM_R_X3Y108_SLICE_X3Y108_D4 = 1'b1;
  assign CLBLM_R_X3Y108_SLICE_X3Y108_D5 = 1'b1;
  assign CLBLM_R_X3Y108_SLICE_X3Y108_D6 = 1'b1;
  assign CLBLM_R_X11Y105_SLICE_X15Y105_B1 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X11Y105_SLICE_X15Y105_B2 = CLBLM_L_X12Y105_SLICE_X16Y105_CO6;
  assign CLBLM_R_X3Y108_SLICE_X2Y108_A1 = 1'b1;
  assign CLBLM_R_X3Y108_SLICE_X2Y108_A2 = 1'b1;
  assign CLBLM_R_X3Y108_SLICE_X2Y108_A3 = 1'b1;
  assign CLBLM_R_X3Y108_SLICE_X2Y108_A4 = 1'b1;
  assign CLBLM_R_X3Y108_SLICE_X2Y108_A5 = 1'b1;
  assign CLBLM_R_X3Y108_SLICE_X2Y108_A6 = 1'b1;
  assign CLBLM_R_X3Y108_SLICE_X2Y108_B1 = 1'b1;
  assign CLBLM_R_X3Y108_SLICE_X2Y108_B2 = 1'b1;
  assign CLBLM_R_X3Y108_SLICE_X2Y108_B3 = 1'b1;
  assign CLBLM_R_X3Y108_SLICE_X2Y108_B4 = 1'b1;
  assign CLBLM_R_X3Y108_SLICE_X2Y108_B5 = 1'b1;
  assign CLBLM_R_X3Y108_SLICE_X2Y108_B6 = 1'b1;
  assign CLBLM_R_X11Y105_SLICE_X15Y105_B5 = CLBLM_R_X11Y104_SLICE_X14Y104_CO6;
  assign CLBLM_R_X3Y108_SLICE_X2Y108_C1 = 1'b1;
  assign CLBLM_R_X3Y108_SLICE_X2Y108_C2 = 1'b1;
  assign CLBLM_R_X3Y108_SLICE_X2Y108_C3 = 1'b1;
  assign CLBLM_R_X3Y108_SLICE_X2Y108_C4 = 1'b1;
  assign CLBLM_R_X3Y108_SLICE_X2Y108_C5 = 1'b1;
  assign CLBLM_R_X3Y108_SLICE_X2Y108_C6 = 1'b1;
  assign CLBLM_R_X3Y108_SLICE_X2Y108_D1 = 1'b1;
  assign CLBLM_R_X3Y108_SLICE_X2Y108_D2 = 1'b1;
  assign CLBLM_R_X3Y108_SLICE_X2Y108_D3 = 1'b1;
  assign CLBLM_R_X3Y108_SLICE_X2Y108_D4 = 1'b1;
  assign CLBLM_R_X3Y108_SLICE_X2Y108_D5 = 1'b1;
  assign CLBLM_R_X3Y108_SLICE_X2Y108_D6 = 1'b1;
  assign CLBLM_R_X11Y105_SLICE_X15Y105_C1 = CLBLM_R_X11Y104_SLICE_X14Y104_CO6;
  assign CLBLM_R_X11Y105_SLICE_X15Y105_C2 = LIOB33_X0Y103_IOB_X0Y104_I;
  assign CLBLM_R_X11Y105_SLICE_X15Y105_D6 = CLBLM_L_X12Y105_SLICE_X16Y105_CO6;
  assign LIOB33_X0Y125_IOB_X0Y126_O = CLBLM_R_X3Y107_SLICE_X2Y107_CO6;
  assign LIOB33_X0Y125_IOB_X0Y125_O = CLBLM_R_X7Y109_SLICE_X9Y109_AO5;
  assign CLBLM_R_X3Y109_SLICE_X3Y109_A1 = LIOB33_X0Y113_IOB_X0Y113_I;
  assign CLBLM_R_X3Y109_SLICE_X3Y109_A2 = LIOB33_X0Y115_IOB_X0Y115_I;
  assign CLBLM_R_X3Y109_SLICE_X3Y109_A3 = CLBLL_L_X4Y108_SLICE_X5Y108_AO6;
  assign CLBLM_R_X3Y109_SLICE_X3Y109_A4 = RIOB33_X105Y105_IOB_X1Y106_I;
  assign CLBLM_R_X3Y109_SLICE_X3Y109_A5 = CLBLL_L_X4Y108_SLICE_X4Y108_DO6;
  assign CLBLM_R_X3Y109_SLICE_X3Y109_A6 = RIOB33_SING_X105Y100_IOB_X1Y100_I;
  assign CLBLM_R_X3Y109_SLICE_X3Y109_B1 = 1'b1;
  assign CLBLM_R_X3Y109_SLICE_X3Y109_B2 = 1'b1;
  assign CLBLM_R_X3Y109_SLICE_X3Y109_B3 = 1'b1;
  assign CLBLM_R_X3Y109_SLICE_X3Y109_B4 = 1'b1;
  assign CLBLM_R_X3Y109_SLICE_X3Y109_B5 = 1'b1;
  assign CLBLM_R_X3Y109_SLICE_X3Y109_B6 = 1'b1;
  assign CLBLM_R_X3Y109_SLICE_X3Y109_C1 = 1'b1;
  assign CLBLM_R_X3Y109_SLICE_X3Y109_C2 = 1'b1;
  assign CLBLM_R_X3Y109_SLICE_X3Y109_C3 = 1'b1;
  assign CLBLM_R_X3Y109_SLICE_X3Y109_C4 = 1'b1;
  assign CLBLM_R_X3Y109_SLICE_X3Y109_C5 = 1'b1;
  assign CLBLM_R_X3Y109_SLICE_X3Y109_C6 = 1'b1;
  assign CLBLM_R_X3Y109_SLICE_X3Y109_D1 = 1'b1;
  assign CLBLM_R_X3Y109_SLICE_X3Y109_D2 = 1'b1;
  assign CLBLM_R_X3Y109_SLICE_X3Y109_D3 = 1'b1;
  assign CLBLM_R_X3Y109_SLICE_X3Y109_D4 = 1'b1;
  assign CLBLM_R_X3Y109_SLICE_X3Y109_D5 = 1'b1;
  assign CLBLM_R_X3Y109_SLICE_X3Y109_D6 = 1'b1;
  assign CLBLM_R_X3Y109_SLICE_X2Y109_A1 = 1'b1;
  assign CLBLM_R_X3Y109_SLICE_X2Y109_A2 = 1'b1;
  assign CLBLM_R_X3Y109_SLICE_X2Y109_A3 = 1'b1;
  assign CLBLM_R_X3Y109_SLICE_X2Y109_A4 = 1'b1;
  assign CLBLM_R_X3Y109_SLICE_X2Y109_A5 = 1'b1;
  assign CLBLM_R_X3Y109_SLICE_X2Y109_A6 = 1'b1;
  assign CLBLM_R_X3Y109_SLICE_X2Y109_B1 = 1'b1;
  assign CLBLM_R_X3Y109_SLICE_X2Y109_B2 = 1'b1;
  assign CLBLM_R_X3Y109_SLICE_X2Y109_B3 = 1'b1;
  assign CLBLM_R_X3Y109_SLICE_X2Y109_B4 = 1'b1;
  assign CLBLM_R_X3Y109_SLICE_X2Y109_B5 = 1'b1;
  assign CLBLM_R_X3Y109_SLICE_X2Y109_B6 = 1'b1;
  assign CLBLM_R_X3Y109_SLICE_X2Y109_C1 = 1'b1;
  assign CLBLM_R_X3Y109_SLICE_X2Y109_C2 = 1'b1;
  assign CLBLM_R_X3Y109_SLICE_X2Y109_C3 = 1'b1;
  assign CLBLM_R_X3Y109_SLICE_X2Y109_C4 = 1'b1;
  assign CLBLM_R_X3Y109_SLICE_X2Y109_C5 = 1'b1;
  assign CLBLM_R_X3Y109_SLICE_X2Y109_C6 = 1'b1;
  assign CLBLM_R_X3Y109_SLICE_X2Y109_D1 = 1'b1;
  assign CLBLM_R_X3Y109_SLICE_X2Y109_D2 = 1'b1;
  assign CLBLM_R_X3Y109_SLICE_X2Y109_D3 = 1'b1;
  assign CLBLM_R_X3Y109_SLICE_X2Y109_D4 = 1'b1;
  assign CLBLM_R_X3Y109_SLICE_X2Y109_D5 = 1'b1;
  assign CLBLM_R_X3Y109_SLICE_X2Y109_D6 = 1'b1;
  assign CLBLM_L_X12Y104_SLICE_X17Y104_A1 = 1'b1;
  assign CLBLM_L_X12Y104_SLICE_X17Y104_A2 = 1'b1;
  assign CLBLM_L_X12Y104_SLICE_X17Y104_A3 = 1'b1;
  assign CLBLM_L_X12Y104_SLICE_X17Y104_A4 = 1'b1;
  assign CLBLM_L_X12Y104_SLICE_X17Y104_A5 = 1'b1;
  assign CLBLM_L_X12Y104_SLICE_X17Y104_A6 = 1'b1;
  assign CLBLM_L_X12Y104_SLICE_X17Y104_B1 = 1'b1;
  assign CLBLM_L_X12Y104_SLICE_X17Y104_B2 = 1'b1;
  assign CLBLM_L_X12Y104_SLICE_X17Y104_B3 = 1'b1;
  assign CLBLM_L_X12Y104_SLICE_X17Y104_B4 = 1'b1;
  assign CLBLM_L_X12Y104_SLICE_X17Y104_B5 = 1'b1;
  assign CLBLM_L_X12Y104_SLICE_X17Y104_B6 = 1'b1;
  assign CLBLM_L_X12Y104_SLICE_X17Y104_C1 = 1'b1;
  assign CLBLM_L_X12Y104_SLICE_X17Y104_C2 = 1'b1;
  assign CLBLM_L_X12Y104_SLICE_X17Y104_C3 = 1'b1;
  assign CLBLM_L_X12Y104_SLICE_X17Y104_C4 = 1'b1;
  assign CLBLM_L_X12Y104_SLICE_X17Y104_C5 = 1'b1;
  assign CLBLM_L_X12Y104_SLICE_X17Y104_C6 = 1'b1;
  assign CLBLM_L_X12Y104_SLICE_X17Y104_D1 = 1'b1;
  assign CLBLM_L_X12Y104_SLICE_X17Y104_D2 = 1'b1;
  assign CLBLM_L_X12Y104_SLICE_X17Y104_D3 = 1'b1;
  assign CLBLM_L_X12Y104_SLICE_X17Y104_D4 = 1'b1;
  assign CLBLM_L_X12Y104_SLICE_X17Y104_D5 = 1'b1;
  assign CLBLM_L_X12Y104_SLICE_X17Y104_D6 = 1'b1;
  assign LIOI3_X0Y145_OLOGIC_X0Y146_D1 = CLBLL_L_X4Y115_SLICE_X4Y115_CO6;
  assign CLBLM_L_X12Y104_SLICE_X16Y104_A1 = 1'b1;
  assign CLBLM_L_X12Y104_SLICE_X16Y104_A2 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X12Y104_SLICE_X16Y104_A3 = LIOB33_X0Y101_IOB_X0Y102_I;
  assign CLBLM_L_X12Y104_SLICE_X16Y104_A4 = LIOB33_X0Y101_IOB_X0Y101_I;
  assign CLBLM_L_X12Y104_SLICE_X16Y104_A5 = 1'b1;
  assign CLBLM_L_X12Y104_SLICE_X16Y104_A6 = 1'b1;
  assign LIOI3_X0Y145_OLOGIC_X0Y146_T1 = 1'b1;
  assign CLBLM_L_X12Y104_SLICE_X16Y104_B1 = CLBLM_R_X11Y104_SLICE_X15Y104_CO6;
  assign CLBLM_L_X12Y104_SLICE_X16Y104_B2 = CLBLM_L_X12Y106_SLICE_X17Y106_AO6;
  assign CLBLM_L_X12Y104_SLICE_X16Y104_B3 = CLBLM_L_X12Y105_SLICE_X16Y105_BO6;
  assign CLBLM_L_X12Y104_SLICE_X16Y104_B4 = CLBLM_L_X12Y104_SLICE_X16Y104_CO6;
  assign CLBLM_L_X12Y104_SLICE_X16Y104_B5 = CLBLM_L_X12Y104_SLICE_X16Y104_AO6;
  assign CLBLM_L_X12Y104_SLICE_X16Y104_B6 = CLBLM_L_X12Y104_SLICE_X16Y104_AO5;
  assign LIOI3_X0Y145_OLOGIC_X0Y145_D1 = CLBLL_L_X4Y115_SLICE_X4Y115_AO5;
  assign CLBLM_L_X12Y104_SLICE_X16Y104_C1 = RIOB33_X105Y113_IOB_X1Y113_I;
  assign CLBLM_L_X12Y104_SLICE_X16Y104_C2 = LIOB33_SING_X0Y100_IOB_X0Y100_I;
  assign CLBLM_L_X12Y104_SLICE_X16Y104_C3 = RIOB33_X105Y111_IOB_X1Y112_I;
  assign CLBLM_L_X12Y104_SLICE_X16Y104_C4 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X12Y104_SLICE_X16Y104_C5 = RIOB33_X105Y107_IOB_X1Y107_I;
  assign CLBLM_L_X12Y104_SLICE_X16Y104_C6 = RIOB33_X105Y107_IOB_X1Y108_I;
  assign LIOI3_X0Y145_OLOGIC_X0Y145_T1 = 1'b1;
  assign CLBLM_L_X12Y104_SLICE_X16Y104_D1 = CLBLM_L_X12Y106_SLICE_X17Y106_AO6;
  assign CLBLM_L_X12Y104_SLICE_X16Y104_D2 = CLBLM_L_X12Y104_SLICE_X16Y104_AO6;
  assign CLBLM_L_X12Y104_SLICE_X16Y104_D3 = CLBLM_L_X12Y104_SLICE_X16Y104_CO6;
  assign CLBLM_L_X12Y104_SLICE_X16Y104_D4 = CLBLM_L_X12Y104_SLICE_X16Y104_AO5;
  assign CLBLM_L_X12Y104_SLICE_X16Y104_D5 = CLBLM_R_X11Y104_SLICE_X15Y104_CO6;
  assign CLBLM_L_X12Y104_SLICE_X16Y104_D6 = CLBLM_L_X12Y105_SLICE_X16Y105_BO6;
  assign LIOB33_X0Y127_IOB_X0Y128_O = CLBLM_R_X3Y107_SLICE_X3Y107_BO6;
  assign LIOB33_X0Y127_IOB_X0Y127_O = CLBLM_R_X3Y107_SLICE_X3Y107_AO6;
  assign CLBLM_R_X11Y104_SLICE_X15Y104_B5 = RIOB33_X105Y113_IOB_X1Y113_I;
  assign CLBLM_R_X11Y104_SLICE_X15Y104_B6 = LIOB33_SING_X0Y100_IOB_X0Y100_I;
  assign CLBLM_L_X12Y105_SLICE_X17Y105_A1 = CLBLM_L_X12Y105_SLICE_X17Y105_DO6;
  assign CLBLM_L_X12Y105_SLICE_X17Y105_A2 = CLBLM_R_X13Y105_SLICE_X18Y105_AO6;
  assign CLBLM_L_X12Y105_SLICE_X17Y105_A3 = LIOB33_X0Y101_IOB_X0Y102_I;
  assign CLBLM_L_X12Y105_SLICE_X17Y105_A4 = LIOB33_X0Y101_IOB_X0Y101_I;
  assign CLBLM_L_X12Y105_SLICE_X17Y105_A5 = RIOB33_X105Y109_IOB_X1Y109_I;
  assign CLBLM_L_X12Y105_SLICE_X17Y105_A6 = CLBLM_L_X12Y105_SLICE_X17Y105_CO6;
  assign CLBLM_L_X12Y105_SLICE_X17Y105_B1 = CLBLM_L_X12Y105_SLICE_X17Y105_DO6;
  assign CLBLM_L_X12Y105_SLICE_X17Y105_B2 = LIOB33_X0Y101_IOB_X0Y101_I;
  assign CLBLM_L_X12Y105_SLICE_X17Y105_B3 = LIOB33_X0Y101_IOB_X0Y102_I;
  assign CLBLM_L_X12Y105_SLICE_X17Y105_B4 = RIOB33_X105Y109_IOB_X1Y109_I;
  assign CLBLM_L_X12Y105_SLICE_X17Y105_B5 = CLBLM_R_X13Y105_SLICE_X18Y105_AO6;
  assign CLBLM_L_X12Y105_SLICE_X17Y105_B6 = CLBLM_L_X12Y105_SLICE_X17Y105_CO6;
  assign CLBLM_L_X12Y105_SLICE_X17Y105_C1 = RIOB33_X105Y113_IOB_X1Y113_I;
  assign CLBLM_L_X12Y105_SLICE_X17Y105_C2 = RIOB33_X105Y111_IOB_X1Y112_I;
  assign CLBLM_L_X12Y105_SLICE_X17Y105_C3 = RIOB33_X105Y109_IOB_X1Y110_I;
  assign CLBLM_L_X12Y105_SLICE_X17Y105_C4 = LIOB33_SING_X0Y100_IOB_X0Y100_I;
  assign CLBLM_L_X12Y105_SLICE_X17Y105_C5 = RIOB33_X105Y111_IOB_X1Y111_I;
  assign CLBLM_L_X12Y105_SLICE_X17Y105_C6 = LIOB33_X0Y101_IOB_X0Y101_I;
  assign CLBLM_L_X12Y105_SLICE_X17Y105_D1 = RIOB33_X105Y113_IOB_X1Y113_I;
  assign CLBLM_L_X12Y105_SLICE_X17Y105_D2 = LIOB33_SING_X0Y100_IOB_X0Y100_I;
  assign CLBLM_L_X12Y105_SLICE_X17Y105_D3 = RIOB33_X105Y111_IOB_X1Y111_I;
  assign CLBLM_L_X12Y105_SLICE_X17Y105_D4 = RIOB33_X105Y111_IOB_X1Y112_I;
  assign CLBLM_L_X12Y105_SLICE_X17Y105_D5 = RIOB33_X105Y109_IOB_X1Y110_I;
  assign CLBLM_L_X12Y105_SLICE_X17Y105_D6 = RIOB33_X105Y109_IOB_X1Y109_I;
  assign CLBLM_L_X12Y105_SLICE_X16Y105_A1 = 1'b1;
  assign CLBLM_L_X12Y105_SLICE_X16Y105_A2 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X12Y105_SLICE_X16Y105_A3 = CLBLM_L_X12Y104_SLICE_X16Y104_CO6;
  assign CLBLM_L_X12Y105_SLICE_X16Y105_A4 = LIOB33_X0Y101_IOB_X0Y101_I;
  assign CLBLM_L_X12Y105_SLICE_X16Y105_A5 = CLBLM_R_X11Y104_SLICE_X15Y104_CO6;
  assign CLBLM_L_X12Y105_SLICE_X16Y105_A6 = 1'b1;
  assign CLBLM_L_X12Y105_SLICE_X16Y105_B1 = RIOB33_X105Y109_IOB_X1Y109_I;
  assign CLBLM_L_X12Y105_SLICE_X16Y105_B2 = RIOB33_X105Y107_IOB_X1Y107_I;
  assign CLBLM_L_X12Y105_SLICE_X16Y105_B3 = RIOB33_X105Y111_IOB_X1Y112_I;
  assign CLBLM_L_X12Y105_SLICE_X16Y105_B4 = LIOB33_SING_X0Y100_IOB_X0Y100_I;
  assign CLBLM_L_X12Y105_SLICE_X16Y105_B5 = RIOB33_X105Y113_IOB_X1Y113_I;
  assign CLBLM_L_X12Y105_SLICE_X16Y105_B6 = RIOB33_X105Y107_IOB_X1Y108_I;
  assign CLBLM_L_X12Y105_SLICE_X16Y105_C1 = CLBLM_L_X12Y104_SLICE_X16Y104_CO6;
  assign CLBLM_L_X12Y105_SLICE_X16Y105_C2 = RIOB33_X105Y107_IOB_X1Y107_I;
  assign CLBLM_L_X12Y105_SLICE_X16Y105_C3 = CLBLM_R_X11Y104_SLICE_X15Y104_CO6;
  assign CLBLM_L_X12Y105_SLICE_X16Y105_C4 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X12Y105_SLICE_X16Y105_C5 = LIOB33_X0Y101_IOB_X0Y101_I;
  assign CLBLM_L_X12Y105_SLICE_X16Y105_C6 = CLBLM_L_X12Y105_SLICE_X16Y105_BO6;
  assign LIOB33_X0Y129_IOB_X0Y129_O = CLBLM_R_X3Y108_SLICE_X3Y108_AO6;
  assign LIOB33_X0Y129_IOB_X0Y130_O = CLBLL_L_X2Y110_SLICE_X0Y110_AO6;
  assign CLBLM_L_X12Y105_SLICE_X16Y105_D1 = RIOB33_X105Y113_IOB_X1Y113_I;
  assign CLBLM_L_X12Y105_SLICE_X16Y105_D2 = RIOB33_X105Y111_IOB_X1Y112_I;
  assign CLBLM_L_X12Y105_SLICE_X16Y105_D3 = RIOB33_X105Y107_IOB_X1Y107_I;
  assign CLBLM_L_X12Y105_SLICE_X16Y105_D4 = LIOB33_SING_X0Y100_IOB_X0Y100_I;
  assign CLBLM_L_X12Y105_SLICE_X16Y105_D5 = RIOB33_X105Y109_IOB_X1Y109_I;
  assign CLBLM_L_X12Y105_SLICE_X16Y105_D6 = RIOB33_X105Y107_IOB_X1Y108_I;
  assign CLBLM_L_X12Y106_SLICE_X17Y106_A1 = LIOB33_X0Y101_IOB_X0Y102_I;
  assign CLBLM_L_X12Y106_SLICE_X17Y106_A2 = RIOB33_X105Y107_IOB_X1Y107_I;
  assign CLBLM_L_X12Y106_SLICE_X17Y106_A3 = LIOB33_X0Y101_IOB_X0Y101_I;
  assign CLBLM_L_X12Y106_SLICE_X17Y106_A4 = 1'b1;
  assign CLBLM_L_X12Y106_SLICE_X17Y106_A5 = 1'b1;
  assign CLBLM_L_X12Y106_SLICE_X17Y106_A6 = 1'b1;
  assign CLBLM_L_X12Y106_SLICE_X17Y106_B1 = CLBLM_R_X13Y106_SLICE_X19Y106_CO6;
  assign CLBLM_L_X12Y106_SLICE_X17Y106_B2 = CLBLM_L_X12Y105_SLICE_X16Y105_DO6;
  assign CLBLM_L_X12Y106_SLICE_X17Y106_B3 = CLBLM_L_X12Y106_SLICE_X16Y106_AO6;
  assign CLBLM_L_X12Y106_SLICE_X17Y106_B4 = CLBLM_L_X12Y105_SLICE_X16Y105_BO6;
  assign CLBLM_L_X12Y106_SLICE_X17Y106_B5 = CLBLM_L_X12Y106_SLICE_X17Y106_AO6;
  assign CLBLM_L_X12Y106_SLICE_X17Y106_B6 = CLBLM_L_X12Y106_SLICE_X17Y106_AO5;
  assign CLBLM_L_X12Y106_SLICE_X17Y106_C1 = RIOB33_X105Y107_IOB_X1Y108_I;
  assign CLBLM_L_X12Y106_SLICE_X17Y106_C2 = RIOB33_X105Y107_IOB_X1Y107_I;
  assign CLBLM_L_X12Y106_SLICE_X17Y106_C3 = CLBLM_L_X12Y106_SLICE_X16Y106_BO5;
  assign CLBLM_L_X12Y106_SLICE_X17Y106_C4 = CLBLM_R_X13Y106_SLICE_X18Y106_DO6;
  assign CLBLM_L_X12Y106_SLICE_X17Y106_C5 = LIOB33_X0Y101_IOB_X0Y102_I;
  assign CLBLM_L_X12Y106_SLICE_X17Y106_C6 = CLBLM_R_X13Y106_SLICE_X19Y106_AO6;
  assign CLBLM_L_X12Y106_SLICE_X17Y106_D1 = CLBLM_L_X12Y106_SLICE_X17Y106_AO6;
  assign CLBLM_L_X12Y106_SLICE_X17Y106_D2 = CLBLM_L_X12Y106_SLICE_X16Y106_AO6;
  assign CLBLM_L_X12Y106_SLICE_X17Y106_D3 = CLBLM_L_X12Y105_SLICE_X16Y105_DO6;
  assign CLBLM_L_X12Y106_SLICE_X17Y106_D4 = CLBLM_L_X12Y106_SLICE_X17Y106_AO5;
  assign CLBLM_L_X12Y106_SLICE_X17Y106_D5 = CLBLM_R_X13Y106_SLICE_X19Y106_CO6;
  assign CLBLM_L_X12Y106_SLICE_X17Y106_D6 = CLBLM_L_X12Y105_SLICE_X16Y105_BO6;
  assign LIOB33_X0Y131_IOB_X0Y131_O = CLBLL_L_X4Y108_SLICE_X4Y108_AO6;
  assign LIOB33_X0Y131_IOB_X0Y132_O = CLBLL_L_X2Y110_SLICE_X0Y110_AO5;
  assign CLBLM_L_X12Y106_SLICE_X16Y106_A1 = 1'b1;
  assign CLBLM_L_X12Y106_SLICE_X16Y106_A2 = RIOB33_X105Y107_IOB_X1Y108_I;
  assign CLBLM_L_X12Y106_SLICE_X16Y106_A3 = LIOB33_X0Y103_IOB_X0Y104_I;
  assign CLBLM_L_X12Y106_SLICE_X16Y106_A4 = 1'b1;
  assign CLBLM_L_X12Y106_SLICE_X16Y106_A5 = LIOB33_X0Y101_IOB_X0Y101_I;
  assign CLBLM_L_X12Y106_SLICE_X16Y106_A6 = 1'b1;
  assign CLBLM_L_X12Y106_SLICE_X16Y106_B1 = CLBLM_L_X12Y105_SLICE_X16Y105_DO6;
  assign CLBLM_L_X12Y106_SLICE_X16Y106_B2 = CLBLM_L_X12Y105_SLICE_X16Y105_BO6;
  assign CLBLM_L_X12Y106_SLICE_X16Y106_B3 = 1'b1;
  assign CLBLM_L_X12Y106_SLICE_X16Y106_B4 = RIOB33_X105Y107_IOB_X1Y107_I;
  assign CLBLM_L_X12Y106_SLICE_X16Y106_B5 = LIOB33_X0Y101_IOB_X0Y101_I;
  assign CLBLM_L_X12Y106_SLICE_X16Y106_B6 = 1'b1;
  assign CLBLM_L_X12Y106_SLICE_X16Y106_C1 = CLBLM_L_X12Y105_SLICE_X16Y105_AO6;
  assign CLBLM_L_X12Y106_SLICE_X16Y106_C2 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X12Y106_SLICE_X16Y106_C3 = LIOB33_X0Y101_IOB_X0Y102_I;
  assign CLBLM_L_X12Y106_SLICE_X16Y106_C4 = RIOB33_X105Y107_IOB_X1Y107_I;
  assign CLBLM_L_X12Y106_SLICE_X16Y106_C5 = CLBLM_L_X12Y106_SLICE_X16Y106_DO6;
  assign CLBLM_L_X12Y106_SLICE_X16Y106_C6 = CLBLM_L_X12Y106_SLICE_X16Y106_BO6;
  assign CLBLM_L_X12Y106_SLICE_X16Y106_D1 = RIOB33_X105Y107_IOB_X1Y108_I;
  assign CLBLM_L_X12Y106_SLICE_X16Y106_D2 = LIOB33_X0Y101_IOB_X0Y101_I;
  assign CLBLM_L_X12Y106_SLICE_X16Y106_D3 = CLBLM_R_X13Y106_SLICE_X19Y106_CO6;
  assign CLBLM_L_X12Y106_SLICE_X16Y106_D4 = RIOB33_X105Y107_IOB_X1Y107_I;
  assign CLBLM_L_X12Y106_SLICE_X16Y106_D5 = CLBLM_L_X12Y105_SLICE_X16Y105_DO6;
  assign CLBLM_L_X12Y106_SLICE_X16Y106_D6 = CLBLM_L_X12Y105_SLICE_X16Y105_BO6;
  assign LIOI3_X0Y147_OLOGIC_X0Y148_D1 = CLBLM_R_X3Y112_SLICE_X2Y112_CO6;
  assign LIOI3_X0Y147_OLOGIC_X0Y148_T1 = 1'b1;
  assign LIOI3_X0Y147_OLOGIC_X0Y147_D1 = CLBLM_R_X3Y112_SLICE_X2Y112_AO5;
  assign LIOI3_X0Y147_OLOGIC_X0Y147_T1 = 1'b1;
  assign CLBLM_R_X3Y112_SLICE_X3Y112_A1 = LIOB33_X0Y113_IOB_X0Y113_I;
  assign CLBLM_R_X3Y112_SLICE_X3Y112_A2 = LIOB33_X0Y115_IOB_X0Y115_I;
  assign CLBLM_R_X3Y112_SLICE_X3Y112_A3 = RIOB33_X105Y111_IOB_X1Y111_I;
  assign CLBLM_R_X3Y112_SLICE_X3Y112_A4 = CLBLM_R_X3Y112_SLICE_X3Y112_BO6;
  assign CLBLM_R_X3Y112_SLICE_X3Y112_A5 = RIOB33_X105Y109_IOB_X1Y110_I;
  assign CLBLM_R_X3Y112_SLICE_X3Y112_A6 = 1'b1;
  assign CLBLM_R_X3Y112_SLICE_X3Y112_B1 = LIOB33_X0Y113_IOB_X0Y113_I;
  assign CLBLM_R_X3Y112_SLICE_X3Y112_B2 = LIOB33_X0Y111_IOB_X0Y112_I;
  assign CLBLM_R_X3Y112_SLICE_X3Y112_B3 = LIOB33_X0Y111_IOB_X0Y111_I;
  assign CLBLM_R_X3Y112_SLICE_X3Y112_B4 = RIOB33_X105Y109_IOB_X1Y110_I;
  assign CLBLM_R_X3Y112_SLICE_X3Y112_B5 = RIOB33_X105Y111_IOB_X1Y111_I;
  assign CLBLM_R_X3Y112_SLICE_X3Y112_B6 = CLBLM_R_X5Y112_SLICE_X7Y112_DO6;
  assign CLBLM_R_X3Y112_SLICE_X3Y112_C1 = 1'b1;
  assign CLBLM_R_X3Y112_SLICE_X3Y112_C2 = 1'b1;
  assign CLBLM_R_X3Y112_SLICE_X3Y112_C3 = 1'b1;
  assign CLBLM_R_X3Y112_SLICE_X3Y112_C4 = 1'b1;
  assign CLBLM_R_X3Y112_SLICE_X3Y112_C5 = 1'b1;
  assign CLBLM_R_X3Y112_SLICE_X3Y112_C6 = 1'b1;
  assign CLBLM_R_X3Y112_SLICE_X3Y112_D1 = 1'b1;
  assign CLBLM_R_X3Y112_SLICE_X3Y112_D2 = 1'b1;
  assign CLBLM_R_X3Y112_SLICE_X3Y112_D3 = 1'b1;
  assign CLBLM_R_X3Y112_SLICE_X3Y112_D4 = 1'b1;
  assign CLBLM_R_X3Y112_SLICE_X3Y112_D5 = 1'b1;
  assign CLBLM_R_X3Y112_SLICE_X3Y112_D6 = 1'b1;
  assign CLBLM_R_X3Y112_SLICE_X2Y112_A1 = CLBLM_R_X3Y112_SLICE_X2Y112_BO6;
  assign CLBLM_R_X3Y112_SLICE_X2Y112_A2 = CLBLM_R_X5Y113_SLICE_X7Y113_CO6;
  assign CLBLM_R_X3Y112_SLICE_X2Y112_A3 = LIOB33_X0Y115_IOB_X0Y115_I;
  assign CLBLM_R_X3Y112_SLICE_X2Y112_A4 = CLBLL_L_X4Y113_SLICE_X4Y113_BO6;
  assign CLBLM_R_X3Y112_SLICE_X2Y112_A5 = RIOB33_X105Y109_IOB_X1Y110_I;
  assign CLBLM_R_X3Y112_SLICE_X2Y112_A6 = 1'b1;
  assign CLBLM_R_X3Y112_SLICE_X2Y112_B1 = LIOB33_X0Y113_IOB_X0Y113_I;
  assign CLBLM_R_X3Y112_SLICE_X2Y112_B2 = RIOB33_X105Y109_IOB_X1Y110_I;
  assign CLBLM_R_X3Y112_SLICE_X2Y112_B3 = RIOB33_X105Y111_IOB_X1Y111_I;
  assign CLBLM_R_X3Y112_SLICE_X2Y112_B4 = CLBLM_R_X5Y112_SLICE_X7Y112_DO6;
  assign CLBLM_R_X3Y112_SLICE_X2Y112_B5 = LIOB33_X0Y111_IOB_X0Y111_I;
  assign CLBLM_R_X3Y112_SLICE_X2Y112_B6 = LIOB33_X0Y111_IOB_X0Y112_I;
  assign CLBLM_R_X3Y112_SLICE_X2Y112_C1 = CLBLM_R_X3Y112_SLICE_X2Y112_AO6;
  assign CLBLM_R_X3Y112_SLICE_X2Y112_C2 = CLBLM_R_X3Y112_SLICE_X3Y112_AO5;
  assign CLBLM_R_X3Y112_SLICE_X2Y112_C3 = CLBLM_R_X5Y113_SLICE_X7Y113_CO6;
  assign CLBLM_R_X3Y112_SLICE_X2Y112_C4 = RIOB33_X105Y111_IOB_X1Y111_I;
  assign CLBLM_R_X3Y112_SLICE_X2Y112_C5 = LIOB33_X0Y115_IOB_X0Y115_I;
  assign CLBLM_R_X3Y112_SLICE_X2Y112_C6 = CLBLL_L_X4Y113_SLICE_X4Y113_BO6;
  assign CLBLM_R_X3Y112_SLICE_X2Y112_D1 = RIOB33_X105Y109_IOB_X1Y110_I;
  assign CLBLM_R_X3Y112_SLICE_X2Y112_D2 = CLBLM_R_X3Y112_SLICE_X3Y112_AO6;
  assign CLBLM_R_X3Y112_SLICE_X2Y112_D3 = CLBLM_R_X5Y113_SLICE_X7Y113_CO6;
  assign CLBLM_R_X3Y112_SLICE_X2Y112_D4 = LIOB33_X0Y115_IOB_X0Y115_I;
  assign CLBLM_R_X3Y112_SLICE_X2Y112_D5 = CLBLM_R_X3Y112_SLICE_X2Y112_BO6;
  assign CLBLM_R_X3Y112_SLICE_X2Y112_D6 = CLBLL_L_X4Y113_SLICE_X4Y113_BO6;
  assign CLBLM_L_X12Y107_SLICE_X17Y107_A1 = RIOB33_X105Y107_IOB_X1Y108_I;
  assign CLBLM_L_X12Y107_SLICE_X17Y107_A2 = CLBLM_R_X13Y106_SLICE_X19Y106_AO5;
  assign CLBLM_L_X12Y107_SLICE_X17Y107_A3 = CLBLM_R_X13Y106_SLICE_X18Y106_AO6;
  assign CLBLM_L_X12Y107_SLICE_X17Y107_A4 = CLBLM_L_X12Y105_SLICE_X17Y105_BO6;
  assign CLBLM_L_X12Y107_SLICE_X17Y107_A5 = LIOB33_X0Y101_IOB_X0Y102_I;
  assign CLBLM_L_X12Y107_SLICE_X17Y107_A6 = 1'b1;
  assign LIOB33_X0Y133_IOB_X0Y134_O = 1'b0;
  assign CLBLM_L_X12Y107_SLICE_X17Y107_B1 = CLBLM_R_X13Y106_SLICE_X18Y106_AO6;
  assign CLBLM_L_X12Y107_SLICE_X17Y107_B2 = CLBLM_R_X13Y106_SLICE_X19Y106_AO5;
  assign CLBLM_L_X12Y107_SLICE_X17Y107_B3 = LIOB33_X0Y103_IOB_X0Y104_I;
  assign CLBLM_L_X12Y107_SLICE_X17Y107_B4 = CLBLM_L_X12Y105_SLICE_X17Y105_BO6;
  assign CLBLM_L_X12Y107_SLICE_X17Y107_B5 = LIOB33_X0Y101_IOB_X0Y102_I;
  assign CLBLM_L_X12Y107_SLICE_X17Y107_B6 = RIOB33_X105Y107_IOB_X1Y108_I;
  assign LIOB33_X0Y133_IOB_X0Y133_O = CLBLM_R_X3Y109_SLICE_X3Y109_AO6;
  assign CLBLM_L_X12Y107_SLICE_X17Y107_C1 = LIOB33_X0Y103_IOB_X0Y104_I;
  assign CLBLM_L_X12Y107_SLICE_X17Y107_C2 = CLBLM_R_X13Y106_SLICE_X19Y106_AO5;
  assign CLBLM_L_X12Y107_SLICE_X17Y107_C3 = RIOB33_X105Y107_IOB_X1Y108_I;
  assign CLBLM_L_X12Y107_SLICE_X17Y107_C4 = CLBLM_L_X12Y105_SLICE_X17Y105_BO6;
  assign CLBLM_L_X12Y107_SLICE_X17Y107_C5 = CLBLM_R_X13Y106_SLICE_X18Y106_AO6;
  assign CLBLM_L_X12Y107_SLICE_X17Y107_C6 = LIOB33_X0Y101_IOB_X0Y102_I;
  assign CLBLM_L_X12Y107_SLICE_X17Y107_D1 = LIOB33_X0Y103_IOB_X0Y104_I;
  assign CLBLM_L_X12Y107_SLICE_X17Y107_D2 = CLBLM_L_X12Y106_SLICE_X17Y106_DO6;
  assign CLBLM_L_X12Y107_SLICE_X17Y107_D3 = RIOB33_X105Y107_IOB_X1Y107_I;
  assign CLBLM_L_X12Y107_SLICE_X17Y107_D4 = CLBLM_R_X13Y106_SLICE_X18Y106_DO6;
  assign CLBLM_L_X12Y107_SLICE_X17Y107_D5 = RIOB33_X105Y107_IOB_X1Y108_I;
  assign CLBLM_L_X12Y107_SLICE_X17Y107_D6 = LIOB33_X0Y101_IOB_X0Y102_I;
  assign CLBLM_L_X12Y107_SLICE_X16Y107_A1 = CLBLM_R_X13Y106_SLICE_X18Y106_CO6;
  assign CLBLM_L_X12Y107_SLICE_X16Y107_A2 = CLBLM_L_X12Y105_SLICE_X17Y105_BO6;
  assign CLBLM_L_X12Y107_SLICE_X16Y107_A3 = CLBLM_L_X12Y108_SLICE_X16Y108_AO5;
  assign CLBLM_L_X12Y107_SLICE_X16Y107_A4 = CLBLM_L_X12Y106_SLICE_X17Y106_DO6;
  assign CLBLM_L_X12Y107_SLICE_X16Y107_A5 = CLBLM_R_X13Y106_SLICE_X18Y106_BO6;
  assign CLBLM_L_X12Y107_SLICE_X16Y107_A6 = CLBLM_L_X12Y106_SLICE_X16Y106_AO5;
  assign CLBLM_L_X12Y107_SLICE_X16Y107_B1 = CLBLM_L_X12Y106_SLICE_X16Y106_DO6;
  assign CLBLM_L_X12Y107_SLICE_X16Y107_B2 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X12Y107_SLICE_X16Y107_B3 = LIOB33_X0Y103_IOB_X0Y104_I;
  assign CLBLM_L_X12Y107_SLICE_X16Y107_B4 = RIOB33_X105Y107_IOB_X1Y107_I;
  assign CLBLM_L_X12Y107_SLICE_X16Y107_B5 = LIOB33_X0Y101_IOB_X0Y102_I;
  assign CLBLM_L_X12Y107_SLICE_X16Y107_B6 = CLBLM_L_X12Y104_SLICE_X16Y104_DO6;
  assign CLBLM_L_X12Y107_SLICE_X16Y107_C1 = CLBLM_L_X12Y106_SLICE_X17Y106_BO6;
  assign CLBLM_L_X12Y107_SLICE_X16Y107_C2 = CLBLM_R_X11Y107_SLICE_X14Y107_AO6;
  assign CLBLM_L_X12Y107_SLICE_X16Y107_C3 = CLBLM_R_X13Y106_SLICE_X18Y106_CO6;
  assign CLBLM_L_X12Y107_SLICE_X16Y107_C4 = CLBLM_L_X12Y106_SLICE_X17Y106_DO6;
  assign CLBLM_L_X12Y107_SLICE_X16Y107_C5 = CLBLM_L_X12Y108_SLICE_X16Y108_AO5;
  assign CLBLM_L_X12Y107_SLICE_X16Y107_C6 = CLBLM_L_X12Y104_SLICE_X16Y104_DO6;
  assign CLBLM_L_X12Y107_SLICE_X16Y107_D1 = CLBLM_L_X12Y105_SLICE_X17Y105_AO6;
  assign CLBLM_L_X12Y107_SLICE_X16Y107_D2 = CLBLM_L_X12Y105_SLICE_X17Y105_BO6;
  assign CLBLM_L_X12Y107_SLICE_X16Y107_D3 = CLBLM_R_X13Y106_SLICE_X18Y106_BO6;
  assign CLBLM_L_X12Y107_SLICE_X16Y107_D4 = CLBLM_L_X12Y106_SLICE_X16Y106_AO5;
  assign CLBLM_L_X12Y107_SLICE_X16Y107_D5 = CLBLM_R_X11Y107_SLICE_X15Y107_AO6;
  assign CLBLM_L_X12Y107_SLICE_X16Y107_D6 = CLBLM_R_X11Y107_SLICE_X14Y107_BO5;
  assign CLBLM_R_X11Y106_SLICE_X15Y106_A4 = CLBLM_L_X10Y108_SLICE_X13Y108_DO6;
  assign CLBLM_R_X11Y106_SLICE_X15Y106_A5 = LIOB33_X0Y101_IOB_X0Y101_I;
  assign CLBLM_R_X11Y106_SLICE_X15Y106_A6 = 1'b1;
  assign CLBLM_R_X11Y106_SLICE_X15Y106_B3 = CLBLM_L_X12Y105_SLICE_X17Y105_AO6;
  assign CLBLM_R_X11Y106_SLICE_X15Y106_B4 = RIOB33_X105Y109_IOB_X1Y109_I;
  assign CLBLM_R_X11Y106_SLICE_X15Y106_B5 = LIOB33_X0Y101_IOB_X0Y102_I;
  assign LIOB33_X0Y135_IOB_X0Y135_O = CLBLL_L_X4Y110_SLICE_X5Y110_AO6;
  assign LIOB33_X0Y135_IOB_X0Y136_O = CLBLL_L_X4Y110_SLICE_X5Y110_AO5;
  assign CLBLM_R_X11Y106_SLICE_X15Y106_B6 = CLBLM_L_X10Y107_SLICE_X13Y107_DO6;
  assign CLBLM_L_X12Y108_SLICE_X17Y108_A1 = RIOB33_X105Y107_IOB_X1Y107_I;
  assign CLBLM_L_X12Y108_SLICE_X17Y108_A2 = CLBLM_L_X12Y107_SLICE_X16Y107_BO6;
  assign CLBLM_L_X12Y108_SLICE_X17Y108_A3 = CLBLM_R_X13Y107_SLICE_X18Y107_AO6;
  assign CLBLM_L_X12Y108_SLICE_X17Y108_A4 = LIOB33_X0Y105_IOB_X0Y105_I;
  assign CLBLM_L_X12Y108_SLICE_X17Y108_A5 = CLBLM_L_X12Y107_SLICE_X16Y107_AO6;
  assign CLBLM_L_X12Y108_SLICE_X17Y108_A6 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X12Y108_SLICE_X17Y108_B1 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X12Y108_SLICE_X17Y108_B2 = LIOB33_X0Y103_IOB_X0Y104_I;
  assign CLBLM_L_X12Y108_SLICE_X17Y108_B3 = LIOB33_X0Y105_IOB_X0Y105_I;
  assign CLBLM_L_X12Y108_SLICE_X17Y108_B4 = CLBLM_L_X12Y107_SLICE_X16Y107_BO6;
  assign CLBLM_L_X12Y108_SLICE_X17Y108_B5 = RIOB33_X105Y107_IOB_X1Y107_I;
  assign CLBLM_L_X12Y108_SLICE_X17Y108_B6 = CLBLM_L_X12Y106_SLICE_X17Y106_CO6;
  assign CLBLM_L_X12Y108_SLICE_X17Y108_C1 = RIOB33_X105Y103_IOB_X1Y104_I;
  assign CLBLM_L_X12Y108_SLICE_X17Y108_C2 = CLBLM_L_X12Y106_SLICE_X16Y106_CO6;
  assign CLBLM_L_X12Y108_SLICE_X17Y108_C3 = LIOB33_X0Y103_IOB_X0Y104_I;
  assign CLBLM_L_X12Y108_SLICE_X17Y108_C4 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X12Y108_SLICE_X17Y108_C5 = CLBLM_R_X11Y105_SLICE_X15Y105_CO6;
  assign CLBLM_L_X12Y108_SLICE_X17Y108_C6 = LIOB33_X0Y105_IOB_X0Y105_I;
  assign CLBLM_L_X10Y110_SLICE_X12Y110_D4 = CLBLM_L_X10Y110_SLICE_X12Y110_CO6;
  assign CLBLM_L_X12Y108_SLICE_X17Y108_D1 = LIOB33_X0Y105_IOB_X0Y105_I;
  assign CLBLM_L_X12Y108_SLICE_X17Y108_D2 = CLBLM_L_X12Y106_SLICE_X17Y106_CO6;
  assign CLBLM_L_X12Y108_SLICE_X17Y108_D3 = LIOB33_X0Y103_IOB_X0Y104_I;
  assign CLBLM_L_X12Y108_SLICE_X17Y108_D4 = RIOB33_X105Y107_IOB_X1Y107_I;
  assign CLBLM_L_X10Y110_SLICE_X12Y110_D5 = RIOB33_X105Y103_IOB_X1Y103_I;
  assign CLBLM_L_X12Y108_SLICE_X17Y108_D5 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X12Y108_SLICE_X17Y108_D6 = CLBLM_L_X12Y107_SLICE_X16Y107_BO6;
  assign CLBLM_L_X10Y110_SLICE_X12Y110_D6 = CLBLM_L_X12Y110_SLICE_X16Y110_BO6;
  assign CLBLM_L_X12Y108_SLICE_X16Y108_A1 = 1'b1;
  assign CLBLM_L_X12Y108_SLICE_X16Y108_A2 = LIOB33_X0Y105_IOB_X0Y105_I;
  assign CLBLM_L_X12Y108_SLICE_X16Y108_A3 = 1'b1;
  assign CLBLM_L_X12Y108_SLICE_X16Y108_A4 = LIOB33_X0Y103_IOB_X0Y104_I;
  assign CLBLM_L_X12Y108_SLICE_X16Y108_A5 = RIOB33_X105Y107_IOB_X1Y107_I;
  assign CLBLM_L_X12Y108_SLICE_X16Y108_A6 = 1'b1;
  assign CLBLM_L_X12Y108_SLICE_X16Y108_B1 = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLM_L_X12Y108_SLICE_X16Y108_B2 = CLBLM_R_X11Y106_SLICE_X15Y106_BO6;
  assign CLBLM_L_X12Y108_SLICE_X16Y108_B3 = RIOB33_X105Y107_IOB_X1Y108_I;
  assign CLBLM_L_X12Y108_SLICE_X16Y108_B4 = LIOB33_X0Y105_IOB_X0Y105_I;
  assign CLBLM_L_X12Y108_SLICE_X16Y108_B5 = CLBLM_R_X11Y107_SLICE_X15Y107_DO6;
  assign CLBLM_L_X12Y108_SLICE_X16Y108_B6 = CLBLM_L_X12Y107_SLICE_X17Y107_CO6;
  assign CLBLM_L_X12Y108_SLICE_X16Y108_C1 = CLBLM_R_X11Y107_SLICE_X15Y107_DO6;
  assign CLBLM_L_X12Y108_SLICE_X16Y108_C2 = CLBLM_R_X11Y106_SLICE_X15Y106_BO6;
  assign CLBLM_L_X12Y108_SLICE_X16Y108_C3 = RIOB33_X105Y107_IOB_X1Y108_I;
  assign CLBLM_L_X12Y108_SLICE_X16Y108_C4 = CLBLM_L_X12Y107_SLICE_X17Y107_CO6;
  assign CLBLM_L_X12Y108_SLICE_X16Y108_C5 = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLM_L_X12Y108_SLICE_X16Y108_C6 = LIOB33_X0Y105_IOB_X0Y105_I;
  assign CLBLM_L_X12Y108_SLICE_X16Y108_D1 = LIOB33_X0Y105_IOB_X0Y105_I;
  assign CLBLM_L_X12Y108_SLICE_X16Y108_D2 = CLBLM_L_X12Y107_SLICE_X17Y107_AO5;
  assign CLBLM_L_X12Y108_SLICE_X16Y108_D3 = RIOB33_X105Y107_IOB_X1Y107_I;
  assign CLBLM_L_X12Y108_SLICE_X16Y108_D4 = RIOB33_X105Y107_IOB_X1Y108_I;
  assign CLBLM_L_X12Y108_SLICE_X16Y108_D5 = CLBLM_L_X12Y107_SLICE_X17Y107_DO6;
  assign CLBLM_L_X12Y108_SLICE_X16Y108_D6 = LIOB33_X0Y103_IOB_X0Y104_I;
  assign CLBLM_R_X7Y108_SLICE_X9Y108_A3 = CLBLM_L_X8Y105_SLICE_X10Y105_BO6;
  assign CLBLM_R_X7Y108_SLICE_X9Y108_B1 = CLBLM_R_X7Y108_SLICE_X9Y108_AO6;
  assign CLBLM_R_X7Y108_SLICE_X9Y108_B2 = CLBLM_L_X8Y107_SLICE_X11Y107_CO6;
  assign CLBLM_R_X7Y108_SLICE_X9Y108_C1 = CLBLM_L_X8Y108_SLICE_X10Y108_BO6;
  assign CLBLM_R_X7Y108_SLICE_X9Y108_C2 = LIOB33_X0Y109_IOB_X0Y109_I;
  assign CLBLM_L_X8Y112_SLICE_X10Y112_D3 = CLBLM_L_X8Y112_SLICE_X11Y112_AO6;
  assign CLBLM_R_X7Y108_SLICE_X9Y108_C6 = LIOB33_X0Y115_IOB_X0Y116_I;
  assign CLBLM_L_X8Y112_SLICE_X10Y112_D4 = CLBLM_L_X8Y112_SLICE_X10Y112_CO6;
  assign CLBLM_L_X8Y112_SLICE_X10Y112_D5 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLM_L_X8Y112_SLICE_X10Y112_D6 = LIOB33_X0Y113_IOB_X0Y113_I;
  assign LIOB33_X0Y137_IOB_X0Y138_O = CLBLL_L_X4Y111_SLICE_X4Y111_AO5;
  assign LIOB33_X0Y137_IOB_X0Y137_O = CLBLL_L_X4Y111_SLICE_X4Y111_AO6;
  assign CLBLM_R_X7Y108_SLICE_X9Y108_D5 = CLBLM_R_X7Y108_SLICE_X9Y108_AO6;
  assign CLBLM_R_X7Y108_SLICE_X9Y108_D6 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLM_L_X12Y109_SLICE_X17Y109_A1 = CLBLM_L_X12Y108_SLICE_X17Y108_CO6;
  assign CLBLM_L_X12Y109_SLICE_X17Y109_A2 = CLBLM_L_X12Y108_SLICE_X17Y108_AO6;
  assign CLBLM_L_X12Y109_SLICE_X17Y109_A3 = CLBLM_L_X12Y108_SLICE_X17Y108_BO6;
  assign CLBLM_L_X12Y109_SLICE_X17Y109_A4 = RIOB33_X105Y103_IOB_X1Y104_I;
  assign CLBLM_L_X12Y109_SLICE_X17Y109_A5 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X12Y109_SLICE_X17Y109_A6 = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLM_L_X12Y109_SLICE_X17Y109_B1 = CLBLM_L_X12Y107_SLICE_X16Y107_DO6;
  assign CLBLM_L_X12Y109_SLICE_X17Y109_B2 = LIOB33_X0Y105_IOB_X0Y105_I;
  assign CLBLM_L_X12Y109_SLICE_X17Y109_B3 = RIOB33_X105Y107_IOB_X1Y107_I;
  assign CLBLM_L_X12Y109_SLICE_X17Y109_B4 = RIOB33_X105Y107_IOB_X1Y108_I;
  assign CLBLM_L_X12Y109_SLICE_X17Y109_B5 = CLBLM_L_X12Y107_SLICE_X17Y107_BO6;
  assign CLBLM_L_X12Y109_SLICE_X17Y109_B6 = CLBLM_L_X12Y107_SLICE_X17Y107_DO6;
  assign CLBLM_L_X12Y109_SLICE_X17Y109_C1 = 1'b1;
  assign CLBLM_L_X12Y109_SLICE_X17Y109_C2 = 1'b1;
  assign CLBLM_L_X12Y109_SLICE_X17Y109_C3 = 1'b1;
  assign CLBLM_L_X12Y109_SLICE_X17Y109_C4 = 1'b1;
  assign CLBLM_L_X12Y109_SLICE_X17Y109_C5 = 1'b1;
  assign CLBLM_L_X12Y109_SLICE_X17Y109_C6 = 1'b1;
  assign CLBLM_L_X12Y109_SLICE_X17Y109_D1 = 1'b1;
  assign CLBLM_L_X12Y109_SLICE_X17Y109_D2 = 1'b1;
  assign CLBLM_L_X12Y109_SLICE_X17Y109_D3 = 1'b1;
  assign CLBLM_L_X12Y109_SLICE_X17Y109_D4 = 1'b1;
  assign CLBLM_L_X12Y109_SLICE_X17Y109_D5 = 1'b1;
  assign CLBLM_L_X12Y109_SLICE_X17Y109_D6 = 1'b1;
  assign CLBLM_L_X12Y109_SLICE_X16Y109_A1 = LIOB33_X0Y105_IOB_X0Y105_I;
  assign CLBLM_L_X12Y109_SLICE_X16Y109_A2 = RIOB33_X105Y107_IOB_X1Y108_I;
  assign CLBLM_L_X12Y109_SLICE_X16Y109_A3 = CLBLM_L_X12Y107_SLICE_X17Y107_CO6;
  assign CLBLM_L_X12Y109_SLICE_X16Y109_A4 = CLBLM_R_X11Y106_SLICE_X15Y106_BO6;
  assign CLBLM_L_X12Y109_SLICE_X16Y109_A5 = 1'b1;
  assign CLBLM_L_X12Y109_SLICE_X16Y109_A6 = 1'b1;
  assign CLBLM_L_X12Y109_SLICE_X16Y109_B1 = CLBLM_L_X12Y107_SLICE_X16Y107_DO6;
  assign CLBLM_L_X12Y109_SLICE_X16Y109_B2 = CLBLM_L_X12Y107_SLICE_X17Y107_BO6;
  assign CLBLM_L_X12Y109_SLICE_X16Y109_B3 = CLBLM_L_X12Y108_SLICE_X16Y108_AO6;
  assign CLBLM_L_X12Y109_SLICE_X16Y109_B4 = CLBLM_L_X12Y110_SLICE_X16Y110_AO6;
  assign CLBLM_L_X12Y109_SLICE_X16Y109_B5 = CLBLM_L_X12Y109_SLICE_X16Y109_AO6;
  assign CLBLM_L_X12Y109_SLICE_X16Y109_B6 = CLBLM_L_X12Y107_SLICE_X17Y107_DO6;
  assign CLBLM_L_X12Y109_SLICE_X16Y109_C1 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X12Y109_SLICE_X16Y109_C2 = CLBLM_R_X11Y108_SLICE_X15Y108_DO6;
  assign CLBLM_L_X12Y109_SLICE_X16Y109_C3 = CLBLM_L_X12Y109_SLICE_X17Y109_BO6;
  assign CLBLM_L_X12Y109_SLICE_X16Y109_C4 = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLM_L_X12Y109_SLICE_X16Y109_C5 = RIOB33_X105Y107_IOB_X1Y107_I;
  assign CLBLM_L_X12Y109_SLICE_X16Y109_C6 = CLBLM_L_X12Y108_SLICE_X17Y108_DO6;
  assign CLBLM_L_X12Y109_SLICE_X16Y109_D1 = CLBLM_L_X12Y109_SLICE_X16Y109_AO6;
  assign CLBLM_L_X12Y109_SLICE_X16Y109_D2 = CLBLM_L_X12Y107_SLICE_X16Y107_DO6;
  assign CLBLM_L_X12Y109_SLICE_X16Y109_D3 = CLBLM_L_X12Y107_SLICE_X17Y107_BO6;
  assign CLBLM_L_X12Y109_SLICE_X16Y109_D4 = CLBLM_L_X12Y110_SLICE_X16Y110_AO6;
  assign CLBLM_L_X12Y109_SLICE_X16Y109_D5 = CLBLM_L_X12Y108_SLICE_X16Y108_AO6;
  assign CLBLM_L_X12Y109_SLICE_X16Y109_D6 = CLBLM_L_X12Y107_SLICE_X17Y107_DO6;
  assign LIOB33_X0Y139_IOB_X0Y140_O = CLBLL_L_X4Y112_SLICE_X4Y112_AO5;
  assign LIOB33_X0Y139_IOB_X0Y139_O = CLBLL_L_X4Y112_SLICE_X4Y112_AO6;
  assign CLBLM_L_X12Y110_SLICE_X17Y110_A1 = 1'b1;
  assign CLBLM_L_X12Y110_SLICE_X17Y110_A2 = 1'b1;
  assign CLBLM_L_X12Y110_SLICE_X17Y110_A3 = 1'b1;
  assign CLBLM_L_X12Y110_SLICE_X17Y110_A4 = 1'b1;
  assign CLBLM_L_X12Y110_SLICE_X17Y110_A5 = 1'b1;
  assign CLBLM_L_X12Y110_SLICE_X17Y110_A6 = 1'b1;
  assign CLBLM_L_X12Y110_SLICE_X17Y110_B1 = 1'b1;
  assign CLBLM_L_X12Y110_SLICE_X17Y110_B2 = 1'b1;
  assign CLBLM_L_X12Y110_SLICE_X17Y110_B3 = 1'b1;
  assign CLBLM_L_X12Y110_SLICE_X17Y110_B4 = 1'b1;
  assign CLBLM_L_X12Y110_SLICE_X17Y110_B5 = 1'b1;
  assign CLBLM_L_X12Y110_SLICE_X17Y110_B6 = 1'b1;
  assign CLBLM_L_X12Y110_SLICE_X17Y110_C1 = 1'b1;
  assign CLBLM_L_X12Y110_SLICE_X17Y110_C2 = 1'b1;
  assign CLBLM_L_X12Y110_SLICE_X17Y110_C3 = 1'b1;
  assign CLBLM_L_X12Y110_SLICE_X17Y110_C4 = 1'b1;
  assign CLBLM_L_X12Y110_SLICE_X17Y110_C5 = 1'b1;
  assign CLBLM_L_X12Y110_SLICE_X17Y110_C6 = 1'b1;
  assign CLBLM_L_X12Y110_SLICE_X17Y110_D1 = 1'b1;
  assign CLBLM_L_X12Y110_SLICE_X17Y110_D2 = 1'b1;
  assign CLBLM_L_X12Y110_SLICE_X17Y110_D3 = 1'b1;
  assign CLBLM_L_X12Y110_SLICE_X17Y110_D4 = 1'b1;
  assign CLBLM_L_X12Y110_SLICE_X17Y110_D5 = 1'b1;
  assign CLBLM_L_X12Y110_SLICE_X17Y110_D6 = 1'b1;
  assign CLBLM_L_X12Y110_SLICE_X16Y110_A1 = 1'b1;
  assign CLBLM_L_X12Y110_SLICE_X16Y110_A2 = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLM_L_X12Y110_SLICE_X16Y110_A3 = LIOB33_X0Y107_IOB_X0Y107_I;
  assign CLBLM_L_X12Y110_SLICE_X16Y110_A4 = RIOB33_X105Y107_IOB_X1Y107_I;
  assign CLBLM_L_X12Y110_SLICE_X16Y110_A5 = 1'b1;
  assign CLBLM_L_X12Y110_SLICE_X16Y110_A6 = 1'b1;
  assign CLBLM_L_X12Y110_SLICE_X16Y110_B1 = LIOB33_X0Y107_IOB_X0Y108_I;
  assign CLBLM_L_X12Y110_SLICE_X16Y110_B2 = CLBLM_R_X11Y109_SLICE_X15Y109_BO6;
  assign CLBLM_L_X12Y110_SLICE_X16Y110_B3 = LIOB33_X0Y107_IOB_X0Y107_I;
  assign CLBLM_L_X12Y110_SLICE_X16Y110_B4 = RIOB33_X105Y103_IOB_X1Y104_I;
  assign CLBLM_L_X12Y110_SLICE_X16Y110_B5 = CLBLM_L_X12Y109_SLICE_X17Y109_AO6;
  assign CLBLM_L_X12Y110_SLICE_X16Y110_B6 = RIOB33_X105Y103_IOB_X1Y103_I;
  assign CLBLM_L_X12Y110_SLICE_X16Y110_C1 = CLBLM_L_X12Y109_SLICE_X17Y109_AO6;
  assign CLBLM_L_X12Y110_SLICE_X16Y110_C2 = LIOB33_X0Y107_IOB_X0Y107_I;
  assign CLBLM_L_X12Y110_SLICE_X16Y110_C3 = RIOB33_X105Y103_IOB_X1Y103_I;
  assign CLBLM_L_X12Y110_SLICE_X16Y110_C4 = RIOB33_X105Y103_IOB_X1Y104_I;
  assign CLBLM_L_X12Y110_SLICE_X16Y110_C5 = LIOB33_X0Y107_IOB_X0Y108_I;
  assign CLBLM_L_X12Y110_SLICE_X16Y110_C6 = CLBLM_R_X11Y109_SLICE_X15Y109_BO6;
  assign CLBLM_L_X12Y110_SLICE_X16Y110_D1 = CLBLM_R_X11Y107_SLICE_X15Y107_CO6;
  assign CLBLM_L_X12Y110_SLICE_X16Y110_D2 = CLBLM_L_X12Y108_SLICE_X16Y108_CO6;
  assign CLBLM_L_X12Y110_SLICE_X16Y110_D3 = CLBLM_L_X12Y109_SLICE_X16Y109_DO6;
  assign CLBLM_L_X12Y110_SLICE_X16Y110_D4 = CLBLM_L_X12Y110_SLICE_X16Y110_AO5;
  assign CLBLM_L_X12Y110_SLICE_X16Y110_D5 = CLBLM_R_X11Y111_SLICE_X15Y111_BO5;
  assign CLBLM_L_X12Y110_SLICE_X16Y110_D6 = CLBLM_L_X12Y109_SLICE_X16Y109_BO6;
  assign LIOB33_X0Y141_IOB_X0Y142_O = CLBLL_L_X4Y114_SLICE_X4Y114_DO6;
  assign LIOB33_X0Y141_IOB_X0Y141_O = CLBLL_L_X4Y112_SLICE_X5Y112_DO6;
  assign LIOI3_SING_X0Y100_ILOGIC_X0Y100_D = LIOB33_SING_X0Y100_IOB_X0Y100_I;
  assign CLBLM_R_X13Y105_SLICE_X19Y105_A1 = 1'b1;
  assign CLBLM_R_X13Y105_SLICE_X19Y105_A2 = 1'b1;
  assign CLBLM_R_X13Y105_SLICE_X19Y105_A3 = 1'b1;
  assign CLBLM_R_X13Y105_SLICE_X19Y105_A4 = 1'b1;
  assign CLBLM_R_X13Y105_SLICE_X19Y105_A5 = 1'b1;
  assign CLBLM_R_X13Y105_SLICE_X19Y105_A6 = 1'b1;
  assign CLBLM_R_X13Y105_SLICE_X19Y105_B1 = 1'b1;
  assign CLBLM_R_X13Y105_SLICE_X19Y105_B2 = 1'b1;
  assign CLBLM_R_X13Y105_SLICE_X19Y105_B3 = 1'b1;
  assign CLBLM_R_X13Y105_SLICE_X19Y105_B4 = 1'b1;
  assign CLBLM_R_X13Y105_SLICE_X19Y105_B5 = 1'b1;
  assign CLBLM_R_X13Y105_SLICE_X19Y105_B6 = 1'b1;
  assign CLBLM_R_X13Y105_SLICE_X19Y105_C1 = 1'b1;
  assign CLBLM_R_X13Y105_SLICE_X19Y105_C2 = 1'b1;
  assign CLBLM_R_X13Y105_SLICE_X19Y105_C3 = 1'b1;
  assign CLBLM_R_X13Y105_SLICE_X19Y105_C4 = 1'b1;
  assign CLBLM_R_X13Y105_SLICE_X19Y105_C5 = 1'b1;
  assign CLBLM_R_X13Y105_SLICE_X19Y105_C6 = 1'b1;
  assign LIOB33_X0Y143_IOB_X0Y143_O = CLBLL_L_X4Y115_SLICE_X4Y115_DO6;
  assign CLBLM_R_X13Y105_SLICE_X19Y105_D1 = 1'b1;
  assign CLBLM_R_X13Y105_SLICE_X19Y105_D2 = 1'b1;
  assign CLBLM_R_X13Y105_SLICE_X19Y105_D3 = 1'b1;
  assign CLBLM_R_X13Y105_SLICE_X19Y105_D4 = 1'b1;
  assign CLBLM_R_X13Y105_SLICE_X19Y105_D5 = 1'b1;
  assign CLBLM_R_X13Y105_SLICE_X19Y105_D6 = 1'b1;
  assign CLBLM_R_X13Y105_SLICE_X18Y105_A1 = RIOB33_X105Y111_IOB_X1Y111_I;
  assign CLBLM_R_X13Y105_SLICE_X18Y105_A2 = LIOB33_SING_X0Y100_IOB_X0Y100_I;
  assign CLBLM_R_X13Y105_SLICE_X18Y105_A3 = RIOB33_X105Y109_IOB_X1Y109_I;
  assign CLBLM_R_X13Y105_SLICE_X18Y105_A4 = RIOB33_X105Y113_IOB_X1Y113_I;
  assign CLBLM_R_X13Y105_SLICE_X18Y105_A5 = RIOB33_X105Y111_IOB_X1Y112_I;
  assign CLBLM_R_X13Y105_SLICE_X18Y105_A6 = RIOB33_X105Y109_IOB_X1Y110_I;
  assign CLBLM_R_X13Y105_SLICE_X18Y105_B1 = 1'b1;
  assign CLBLM_R_X13Y105_SLICE_X18Y105_B2 = 1'b1;
  assign CLBLM_R_X13Y105_SLICE_X18Y105_B3 = 1'b1;
  assign CLBLM_R_X13Y105_SLICE_X18Y105_B4 = 1'b1;
  assign CLBLM_R_X13Y105_SLICE_X18Y105_B5 = 1'b1;
  assign CLBLM_R_X13Y105_SLICE_X18Y105_B6 = 1'b1;
  assign CLBLM_R_X13Y105_SLICE_X18Y105_C1 = 1'b1;
  assign CLBLM_R_X13Y105_SLICE_X18Y105_C2 = 1'b1;
  assign CLBLM_R_X13Y105_SLICE_X18Y105_C3 = 1'b1;
  assign CLBLM_R_X13Y105_SLICE_X18Y105_C4 = 1'b1;
  assign CLBLM_R_X13Y105_SLICE_X18Y105_C5 = 1'b1;
  assign CLBLM_R_X13Y105_SLICE_X18Y105_C6 = 1'b1;
  assign CLBLM_R_X13Y105_SLICE_X18Y105_D1 = 1'b1;
  assign CLBLM_R_X13Y105_SLICE_X18Y105_D2 = 1'b1;
  assign CLBLM_R_X13Y105_SLICE_X18Y105_D3 = 1'b1;
  assign CLBLM_R_X13Y105_SLICE_X18Y105_D4 = 1'b1;
  assign CLBLM_R_X13Y105_SLICE_X18Y105_D5 = 1'b1;
  assign CLBLM_R_X13Y105_SLICE_X18Y105_D6 = 1'b1;
  assign LIOI3_SING_X0Y149_OLOGIC_X0Y149_D1 = CLBLM_R_X3Y112_SLICE_X2Y112_DO6;
  assign LIOI3_SING_X0Y149_OLOGIC_X0Y149_T1 = 1'b1;
  assign CLBLM_L_X10Y102_SLICE_X13Y102_A1 = 1'b1;
  assign CLBLM_L_X10Y102_SLICE_X13Y102_A2 = 1'b1;
  assign CLBLM_L_X10Y102_SLICE_X13Y102_A3 = 1'b1;
  assign CLBLM_L_X10Y102_SLICE_X13Y102_A4 = 1'b1;
  assign CLBLM_L_X10Y102_SLICE_X13Y102_A5 = 1'b1;
  assign CLBLM_L_X10Y102_SLICE_X13Y102_A6 = 1'b1;
  assign CLBLM_L_X10Y102_SLICE_X13Y102_B1 = 1'b1;
  assign CLBLM_L_X10Y102_SLICE_X13Y102_B2 = 1'b1;
  assign CLBLM_L_X10Y102_SLICE_X13Y102_B3 = 1'b1;
  assign CLBLM_L_X10Y102_SLICE_X13Y102_B4 = 1'b1;
  assign CLBLM_L_X10Y102_SLICE_X13Y102_B5 = 1'b1;
  assign CLBLM_L_X10Y102_SLICE_X13Y102_B6 = 1'b1;
  assign CLBLM_L_X10Y102_SLICE_X13Y102_C1 = 1'b1;
  assign CLBLM_L_X10Y102_SLICE_X13Y102_C2 = 1'b1;
  assign CLBLM_L_X10Y102_SLICE_X13Y102_C3 = 1'b1;
  assign CLBLM_L_X10Y102_SLICE_X13Y102_C4 = 1'b1;
  assign CLBLM_L_X10Y102_SLICE_X13Y102_C5 = 1'b1;
  assign CLBLM_L_X10Y102_SLICE_X13Y102_C6 = 1'b1;
  assign CLBLM_L_X10Y102_SLICE_X13Y102_D1 = 1'b1;
  assign CLBLM_L_X10Y102_SLICE_X13Y102_D2 = 1'b1;
  assign CLBLM_L_X10Y102_SLICE_X13Y102_D3 = 1'b1;
  assign CLBLM_L_X10Y102_SLICE_X13Y102_D4 = 1'b1;
  assign CLBLM_L_X10Y102_SLICE_X13Y102_D5 = 1'b1;
  assign CLBLM_L_X10Y102_SLICE_X13Y102_D6 = 1'b1;
  assign CLBLM_L_X10Y102_SLICE_X12Y102_A1 = LIOB33_X0Y101_IOB_X0Y101_I;
  assign CLBLM_L_X10Y102_SLICE_X12Y102_A2 = RIOB33_X105Y101_IOB_X1Y102_I;
  assign CLBLM_L_X10Y102_SLICE_X12Y102_A3 = 1'b1;
  assign CLBLM_L_X10Y102_SLICE_X12Y102_A4 = LIOB33_X0Y101_IOB_X0Y102_I;
  assign CLBLM_L_X10Y102_SLICE_X12Y102_A5 = 1'b1;
  assign CLBLM_L_X10Y102_SLICE_X12Y102_A6 = 1'b1;
  assign CLBLM_L_X10Y102_SLICE_X12Y102_B1 = CLBLM_L_X10Y104_SLICE_X12Y104_BO6;
  assign CLBLM_L_X10Y102_SLICE_X12Y102_B2 = CLBLM_L_X10Y104_SLICE_X13Y104_AO6;
  assign CLBLM_L_X10Y102_SLICE_X12Y102_B3 = CLBLM_L_X10Y104_SLICE_X12Y104_AO6;
  assign CLBLM_L_X10Y102_SLICE_X12Y102_B4 = CLBLM_L_X10Y103_SLICE_X12Y103_BO6;
  assign CLBLM_L_X10Y102_SLICE_X12Y102_B5 = CLBLM_L_X10Y102_SLICE_X12Y102_AO6;
  assign CLBLM_L_X10Y102_SLICE_X12Y102_B6 = CLBLM_L_X10Y102_SLICE_X12Y102_AO5;
  assign CLBLM_L_X10Y102_SLICE_X12Y102_C1 = CLBLM_L_X10Y104_SLICE_X13Y104_AO6;
  assign CLBLM_L_X10Y102_SLICE_X12Y102_C2 = CLBLM_L_X10Y102_SLICE_X12Y102_AO6;
  assign CLBLM_L_X10Y102_SLICE_X12Y102_C3 = CLBLM_L_X10Y104_SLICE_X12Y104_AO6;
  assign CLBLM_L_X10Y102_SLICE_X12Y102_C4 = CLBLM_L_X10Y102_SLICE_X12Y102_AO5;
  assign CLBLM_L_X10Y102_SLICE_X12Y102_C5 = CLBLM_L_X10Y104_SLICE_X12Y104_BO6;
  assign CLBLM_L_X10Y102_SLICE_X12Y102_C6 = CLBLM_L_X10Y103_SLICE_X12Y103_BO6;
  assign CLBLM_L_X10Y102_SLICE_X12Y102_D1 = 1'b1;
  assign CLBLM_L_X10Y102_SLICE_X12Y102_D2 = 1'b1;
  assign CLBLM_L_X10Y102_SLICE_X12Y102_D3 = 1'b1;
  assign CLBLM_L_X10Y102_SLICE_X12Y102_D4 = 1'b1;
  assign CLBLM_L_X10Y102_SLICE_X12Y102_D5 = 1'b1;
  assign CLBLM_L_X10Y102_SLICE_X12Y102_D6 = 1'b1;
  assign LIOB33_X0Y145_IOB_X0Y146_O = CLBLL_L_X4Y115_SLICE_X4Y115_CO6;
  assign LIOB33_X0Y145_IOB_X0Y145_O = CLBLL_L_X4Y115_SLICE_X4Y115_AO5;
  assign CLBLM_R_X13Y106_SLICE_X19Y106_A1 = CLBLM_R_X13Y106_SLICE_X19Y106_BO6;
  assign CLBLM_R_X13Y106_SLICE_X19Y106_A2 = RIOB33_X105Y107_IOB_X1Y108_I;
  assign CLBLM_R_X13Y106_SLICE_X19Y106_A3 = 1'b1;
  assign CLBLM_R_X13Y106_SLICE_X19Y106_A4 = LIOB33_X0Y101_IOB_X0Y101_I;
  assign CLBLM_R_X13Y106_SLICE_X19Y106_A5 = CLBLM_R_X13Y106_SLICE_X19Y106_CO6;
  assign CLBLM_R_X13Y106_SLICE_X19Y106_A6 = 1'b1;
  assign CLBLM_R_X13Y106_SLICE_X19Y106_B1 = RIOB33_X105Y109_IOB_X1Y109_I;
  assign CLBLM_R_X13Y106_SLICE_X19Y106_B2 = RIOB33_X105Y107_IOB_X1Y108_I;
  assign CLBLM_R_X13Y106_SLICE_X19Y106_B3 = RIOB33_X105Y111_IOB_X1Y112_I;
  assign CLBLM_R_X13Y106_SLICE_X19Y106_B4 = RIOB33_X105Y113_IOB_X1Y113_I;
  assign CLBLM_R_X13Y106_SLICE_X19Y106_B5 = RIOB33_X105Y109_IOB_X1Y110_I;
  assign CLBLM_R_X13Y106_SLICE_X19Y106_B6 = LIOB33_SING_X0Y100_IOB_X0Y100_I;
  assign CLBLM_R_X13Y106_SLICE_X19Y106_C1 = RIOB33_X105Y111_IOB_X1Y112_I;
  assign CLBLM_R_X13Y106_SLICE_X19Y106_C2 = RIOB33_X105Y107_IOB_X1Y108_I;
  assign CLBLM_R_X13Y106_SLICE_X19Y106_C3 = RIOB33_X105Y109_IOB_X1Y109_I;
  assign CLBLM_R_X13Y106_SLICE_X19Y106_C4 = LIOB33_SING_X0Y100_IOB_X0Y100_I;
  assign CLBLM_R_X13Y106_SLICE_X19Y106_C5 = RIOB33_X105Y113_IOB_X1Y113_I;
  assign CLBLM_R_X13Y106_SLICE_X19Y106_C6 = RIOB33_X105Y109_IOB_X1Y110_I;
  assign CLBLM_R_X13Y106_SLICE_X19Y106_D1 = 1'b1;
  assign CLBLM_R_X13Y106_SLICE_X19Y106_D2 = 1'b1;
  assign CLBLM_R_X13Y106_SLICE_X19Y106_D3 = 1'b1;
  assign CLBLM_R_X13Y106_SLICE_X19Y106_D4 = 1'b1;
  assign CLBLM_R_X13Y106_SLICE_X19Y106_D5 = 1'b1;
  assign CLBLM_R_X13Y106_SLICE_X19Y106_D6 = 1'b1;
  assign CLBLM_R_X13Y106_SLICE_X18Y106_A1 = 1'b1;
  assign CLBLM_R_X13Y106_SLICE_X18Y106_A2 = LIOB33_X0Y101_IOB_X0Y101_I;
  assign CLBLM_R_X13Y106_SLICE_X18Y106_A3 = CLBLM_R_X13Y105_SLICE_X18Y105_AO6;
  assign CLBLM_R_X13Y106_SLICE_X18Y106_A4 = RIOB33_X105Y109_IOB_X1Y109_I;
  assign CLBLM_R_X13Y106_SLICE_X18Y106_A5 = RIOB33_X105Y105_IOB_X1Y106_I;
  assign CLBLM_R_X13Y106_SLICE_X18Y106_A6 = 1'b1;
  assign CLBLM_R_X13Y106_SLICE_X18Y106_B1 = CLBLM_L_X12Y107_SLICE_X17Y107_AO6;
  assign CLBLM_R_X13Y106_SLICE_X18Y106_B2 = CLBLM_R_X13Y106_SLICE_X19Y106_BO6;
  assign CLBLM_R_X13Y106_SLICE_X18Y106_B3 = CLBLM_R_X13Y106_SLICE_X19Y106_CO6;
  assign CLBLM_R_X13Y106_SLICE_X18Y106_B4 = CLBLM_R_X11Y106_SLICE_X15Y106_AO6;
  assign CLBLM_R_X13Y106_SLICE_X18Y106_B5 = CLBLM_R_X13Y105_SLICE_X18Y105_AO6;
  assign CLBLM_R_X13Y106_SLICE_X18Y106_B6 = CLBLM_L_X12Y106_SLICE_X16Y106_AO6;
  assign CLBLM_R_X13Y106_SLICE_X18Y106_C1 = CLBLM_R_X13Y105_SLICE_X18Y105_AO6;
  assign CLBLM_R_X13Y106_SLICE_X18Y106_C2 = CLBLM_R_X13Y106_SLICE_X19Y106_CO6;
  assign CLBLM_R_X13Y106_SLICE_X18Y106_C3 = CLBLM_R_X13Y106_SLICE_X19Y106_BO6;
  assign CLBLM_R_X13Y106_SLICE_X18Y106_C4 = CLBLM_R_X11Y106_SLICE_X15Y106_AO6;
  assign CLBLM_R_X13Y106_SLICE_X18Y106_C5 = CLBLM_L_X12Y107_SLICE_X17Y107_AO6;
  assign CLBLM_R_X13Y106_SLICE_X18Y106_C6 = CLBLM_L_X12Y106_SLICE_X16Y106_AO6;
  assign CLBLM_R_X13Y106_SLICE_X18Y106_D1 = CLBLM_R_X13Y105_SLICE_X18Y105_AO6;
  assign CLBLM_R_X13Y106_SLICE_X18Y106_D2 = CLBLM_R_X13Y106_SLICE_X19Y106_CO6;
  assign CLBLM_R_X13Y106_SLICE_X18Y106_D3 = CLBLM_R_X13Y106_SLICE_X19Y106_BO6;
  assign CLBLM_R_X13Y106_SLICE_X18Y106_D4 = LIOB33_X0Y101_IOB_X0Y101_I;
  assign CLBLM_R_X13Y106_SLICE_X18Y106_D5 = RIOB33_X105Y109_IOB_X1Y109_I;
  assign CLBLM_R_X13Y106_SLICE_X18Y106_D6 = RIOB33_X105Y107_IOB_X1Y108_I;
  assign CLBLM_R_X11Y107_SLICE_X15Y107_A2 = CLBLM_R_X11Y107_SLICE_X14Y107_DO6;
  assign CLBLM_R_X11Y107_SLICE_X15Y107_B1 = CLBLM_R_X11Y107_SLICE_X14Y107_AO5;
  assign CLBLM_R_X11Y107_SLICE_X15Y107_B2 = CLBLM_R_X11Y111_SLICE_X15Y111_BO6;
  assign CLBLM_R_X11Y107_SLICE_X15Y107_B3 = CLBLM_L_X12Y107_SLICE_X16Y107_AO6;
  assign CLBLM_R_X11Y107_SLICE_X15Y107_B4 = CLBLM_L_X12Y108_SLICE_X16Y108_AO6;
  assign CLBLM_R_X11Y107_SLICE_X15Y107_B5 = CLBLM_L_X12Y107_SLICE_X16Y107_BO6;
  assign CLBLM_L_X10Y103_SLICE_X13Y103_A1 = 1'b1;
  assign CLBLM_L_X10Y103_SLICE_X13Y103_A2 = 1'b1;
  assign CLBLM_L_X10Y103_SLICE_X13Y103_A3 = 1'b1;
  assign CLBLM_L_X10Y103_SLICE_X13Y103_A4 = 1'b1;
  assign CLBLM_L_X10Y103_SLICE_X13Y103_A5 = 1'b1;
  assign CLBLM_L_X10Y103_SLICE_X13Y103_A6 = 1'b1;
  assign CLBLM_L_X10Y103_SLICE_X13Y103_B1 = 1'b1;
  assign CLBLM_L_X10Y103_SLICE_X13Y103_B2 = 1'b1;
  assign CLBLM_L_X10Y103_SLICE_X13Y103_B3 = 1'b1;
  assign CLBLM_L_X10Y103_SLICE_X13Y103_B4 = 1'b1;
  assign CLBLM_L_X10Y103_SLICE_X13Y103_B5 = 1'b1;
  assign CLBLM_L_X10Y111_SLICE_X12Y111_D2 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X10Y103_SLICE_X13Y103_B6 = 1'b1;
  assign CLBLM_L_X10Y103_SLICE_X13Y103_C1 = 1'b1;
  assign CLBLM_L_X10Y103_SLICE_X13Y103_C2 = 1'b1;
  assign CLBLM_L_X10Y103_SLICE_X13Y103_C3 = 1'b1;
  assign CLBLM_L_X10Y103_SLICE_X13Y103_C4 = 1'b1;
  assign CLBLM_L_X10Y103_SLICE_X13Y103_C5 = 1'b1;
  assign CLBLM_L_X10Y103_SLICE_X13Y103_C6 = 1'b1;
  assign CLBLM_L_X10Y103_SLICE_X13Y103_D1 = 1'b1;
  assign CLBLM_L_X10Y103_SLICE_X13Y103_D2 = 1'b1;
  assign CLBLM_L_X10Y103_SLICE_X13Y103_D3 = 1'b1;
  assign CLBLM_L_X10Y103_SLICE_X13Y103_D4 = 1'b1;
  assign CLBLM_L_X10Y103_SLICE_X13Y103_D5 = 1'b1;
  assign CLBLM_L_X10Y103_SLICE_X13Y103_D6 = 1'b1;
  assign CLBLM_L_X10Y103_SLICE_X12Y103_A1 = LIOB33_X0Y101_IOB_X0Y101_I;
  assign CLBLM_L_X10Y103_SLICE_X12Y103_A2 = 1'b1;
  assign CLBLM_L_X10Y103_SLICE_X12Y103_A3 = CLBLM_L_X10Y104_SLICE_X12Y104_AO6;
  assign CLBLM_L_X10Y103_SLICE_X12Y103_A4 = CLBLM_L_X10Y103_SLICE_X12Y103_BO6;
  assign CLBLM_L_X10Y103_SLICE_X12Y103_A5 = RIOB33_X105Y101_IOB_X1Y102_I;
  assign CLBLM_L_X10Y103_SLICE_X12Y103_A6 = 1'b1;
  assign CLBLM_L_X10Y103_SLICE_X12Y103_B1 = RIOB33_X105Y101_IOB_X1Y102_I;
  assign CLBLM_L_X10Y103_SLICE_X12Y103_B2 = RIOB33_X105Y103_IOB_X1Y103_I;
  assign CLBLM_L_X10Y103_SLICE_X12Y103_B3 = RIOB33_X105Y111_IOB_X1Y112_I;
  assign CLBLM_L_X10Y103_SLICE_X12Y103_B4 = RIOB33_X105Y103_IOB_X1Y104_I;
  assign CLBLM_L_X10Y103_SLICE_X12Y103_B5 = LIOB33_SING_X0Y100_IOB_X0Y100_I;
  assign CLBLM_L_X10Y103_SLICE_X12Y103_B6 = RIOB33_X105Y113_IOB_X1Y113_I;
  assign CLBLM_L_X10Y103_SLICE_X12Y103_C1 = RIOB33_X105Y103_IOB_X1Y103_I;
  assign CLBLM_L_X10Y103_SLICE_X12Y103_C2 = CLBLM_L_X10Y104_SLICE_X12Y104_BO6;
  assign CLBLM_L_X10Y103_SLICE_X12Y103_C3 = LIOB33_X0Y101_IOB_X0Y101_I;
  assign CLBLM_L_X10Y103_SLICE_X12Y103_C4 = CLBLM_L_X10Y104_SLICE_X12Y104_AO6;
  assign CLBLM_L_X10Y103_SLICE_X12Y103_C5 = RIOB33_X105Y101_IOB_X1Y102_I;
endmodule
