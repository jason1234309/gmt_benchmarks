module top(
  input LIOB33_SING_X0Y50_IOB_X0Y50_IPAD,
  input LIOB33_X0Y51_IOB_X0Y51_IPAD,
  input LIOB33_X0Y51_IOB_X0Y52_IPAD,
  input LIOB33_X0Y53_IOB_X0Y53_IPAD,
  input LIOB33_X0Y53_IOB_X0Y54_IPAD,
  input LIOB33_X0Y55_IOB_X0Y55_IPAD,
  input LIOB33_X0Y55_IOB_X0Y56_IPAD,
  input LIOB33_X0Y57_IOB_X0Y57_IPAD,
  input LIOB33_X0Y57_IOB_X0Y58_IPAD,
  input LIOB33_X0Y59_IOB_X0Y59_IPAD,
  input LIOB33_X0Y59_IOB_X0Y60_IPAD,
  input LIOB33_X0Y61_IOB_X0Y61_IPAD,
  input LIOB33_X0Y61_IOB_X0Y62_IPAD,
  input LIOB33_X0Y63_IOB_X0Y63_IPAD,
  input LIOB33_X0Y77_IOB_X0Y78_IPAD,
  input RIOB33_SING_X105Y100_IOB_X1Y100_IPAD,
  input RIOB33_SING_X105Y149_IOB_X1Y149_IPAD,
  input RIOB33_X105Y101_IOB_X1Y101_IPAD,
  input RIOB33_X105Y101_IOB_X1Y102_IPAD,
  input RIOB33_X105Y103_IOB_X1Y103_IPAD,
  input RIOB33_X105Y103_IOB_X1Y104_IPAD,
  input RIOB33_X105Y105_IOB_X1Y105_IPAD,
  input RIOB33_X105Y105_IOB_X1Y106_IPAD,
  input RIOB33_X105Y107_IOB_X1Y107_IPAD,
  input RIOB33_X105Y107_IOB_X1Y108_IPAD,
  input RIOB33_X105Y109_IOB_X1Y109_IPAD,
  input RIOB33_X105Y109_IOB_X1Y110_IPAD,
  input RIOB33_X105Y111_IOB_X1Y111_IPAD,
  input RIOB33_X105Y111_IOB_X1Y112_IPAD,
  input RIOB33_X105Y113_IOB_X1Y113_IPAD,
  input RIOB33_X105Y113_IOB_X1Y114_IPAD,
  input RIOB33_X105Y115_IOB_X1Y115_IPAD,
  input RIOB33_X105Y115_IOB_X1Y116_IPAD,
  input RIOB33_X105Y117_IOB_X1Y117_IPAD,
  input RIOB33_X105Y117_IOB_X1Y118_IPAD,
  input RIOB33_X105Y119_IOB_X1Y119_IPAD,
  input RIOB33_X105Y119_IOB_X1Y120_IPAD,
  input RIOB33_X105Y121_IOB_X1Y121_IPAD,
  input RIOB33_X105Y121_IOB_X1Y122_IPAD,
  input RIOB33_X105Y123_IOB_X1Y123_IPAD,
  input RIOB33_X105Y123_IOB_X1Y124_IPAD,
  input RIOB33_X105Y125_IOB_X1Y125_IPAD,
  input RIOB33_X105Y125_IOB_X1Y126_IPAD,
  input RIOB33_X105Y127_IOB_X1Y127_IPAD,
  input RIOB33_X105Y127_IOB_X1Y128_IPAD,
  input RIOB33_X105Y129_IOB_X1Y129_IPAD,
  input RIOB33_X105Y129_IOB_X1Y130_IPAD,
  input RIOB33_X105Y131_IOB_X1Y131_IPAD,
  input RIOB33_X105Y131_IOB_X1Y132_IPAD,
  input RIOB33_X105Y133_IOB_X1Y133_IPAD,
  input RIOB33_X105Y133_IOB_X1Y134_IPAD,
  input RIOB33_X105Y135_IOB_X1Y135_IPAD,
  input RIOB33_X105Y135_IOB_X1Y136_IPAD,
  input RIOB33_X105Y137_IOB_X1Y137_IPAD,
  input RIOB33_X105Y137_IOB_X1Y138_IPAD,
  input RIOB33_X105Y139_IOB_X1Y139_IPAD,
  input RIOB33_X105Y139_IOB_X1Y140_IPAD,
  input RIOB33_X105Y141_IOB_X1Y141_IPAD,
  input RIOB33_X105Y141_IOB_X1Y142_IPAD,
  input RIOB33_X105Y143_IOB_X1Y143_IPAD,
  input RIOB33_X105Y143_IOB_X1Y144_IPAD,
  input RIOB33_X105Y145_IOB_X1Y145_IPAD,
  input RIOB33_X105Y145_IOB_X1Y146_IPAD,
  input RIOB33_X105Y147_IOB_X1Y147_IPAD,
  input RIOB33_X105Y147_IOB_X1Y148_IPAD,
  output LIOB33_SING_X0Y100_IOB_X0Y100_OPAD,
  output LIOB33_SING_X0Y149_IOB_X0Y149_OPAD,
  output LIOB33_SING_X0Y150_IOB_X0Y150_OPAD,
  output LIOB33_SING_X0Y199_IOB_X0Y199_OPAD,
  output LIOB33_X0Y101_IOB_X0Y101_OPAD,
  output LIOB33_X0Y101_IOB_X0Y102_OPAD,
  output LIOB33_X0Y103_IOB_X0Y103_OPAD,
  output LIOB33_X0Y103_IOB_X0Y104_OPAD,
  output LIOB33_X0Y105_IOB_X0Y105_OPAD,
  output LIOB33_X0Y105_IOB_X0Y106_OPAD,
  output LIOB33_X0Y107_IOB_X0Y107_OPAD,
  output LIOB33_X0Y107_IOB_X0Y108_OPAD,
  output LIOB33_X0Y109_IOB_X0Y109_OPAD,
  output LIOB33_X0Y109_IOB_X0Y110_OPAD,
  output LIOB33_X0Y111_IOB_X0Y111_OPAD,
  output LIOB33_X0Y111_IOB_X0Y112_OPAD,
  output LIOB33_X0Y113_IOB_X0Y113_OPAD,
  output LIOB33_X0Y113_IOB_X0Y114_OPAD,
  output LIOB33_X0Y115_IOB_X0Y115_OPAD,
  output LIOB33_X0Y115_IOB_X0Y116_OPAD,
  output LIOB33_X0Y117_IOB_X0Y117_OPAD,
  output LIOB33_X0Y117_IOB_X0Y118_OPAD,
  output LIOB33_X0Y119_IOB_X0Y119_OPAD,
  output LIOB33_X0Y119_IOB_X0Y120_OPAD,
  output LIOB33_X0Y121_IOB_X0Y121_OPAD,
  output LIOB33_X0Y121_IOB_X0Y122_OPAD,
  output LIOB33_X0Y123_IOB_X0Y123_OPAD,
  output LIOB33_X0Y123_IOB_X0Y124_OPAD,
  output LIOB33_X0Y125_IOB_X0Y125_OPAD,
  output LIOB33_X0Y125_IOB_X0Y126_OPAD,
  output LIOB33_X0Y127_IOB_X0Y127_OPAD,
  output LIOB33_X0Y127_IOB_X0Y128_OPAD,
  output LIOB33_X0Y129_IOB_X0Y129_OPAD,
  output LIOB33_X0Y129_IOB_X0Y130_OPAD,
  output LIOB33_X0Y131_IOB_X0Y131_OPAD,
  output LIOB33_X0Y131_IOB_X0Y132_OPAD,
  output LIOB33_X0Y133_IOB_X0Y133_OPAD,
  output LIOB33_X0Y133_IOB_X0Y134_OPAD,
  output LIOB33_X0Y135_IOB_X0Y135_OPAD,
  output LIOB33_X0Y135_IOB_X0Y136_OPAD,
  output LIOB33_X0Y137_IOB_X0Y137_OPAD,
  output LIOB33_X0Y137_IOB_X0Y138_OPAD,
  output LIOB33_X0Y139_IOB_X0Y139_OPAD,
  output LIOB33_X0Y139_IOB_X0Y140_OPAD,
  output LIOB33_X0Y141_IOB_X0Y141_OPAD,
  output LIOB33_X0Y141_IOB_X0Y142_OPAD,
  output LIOB33_X0Y143_IOB_X0Y143_OPAD,
  output LIOB33_X0Y145_IOB_X0Y145_OPAD,
  output LIOB33_X0Y145_IOB_X0Y146_OPAD,
  output LIOB33_X0Y147_IOB_X0Y147_OPAD,
  output LIOB33_X0Y147_IOB_X0Y148_OPAD,
  output LIOB33_X0Y151_IOB_X0Y151_OPAD,
  output LIOB33_X0Y151_IOB_X0Y152_OPAD,
  output LIOB33_X0Y153_IOB_X0Y153_OPAD,
  output LIOB33_X0Y153_IOB_X0Y154_OPAD,
  output LIOB33_X0Y155_IOB_X0Y155_OPAD,
  output LIOB33_X0Y155_IOB_X0Y156_OPAD,
  output LIOB33_X0Y157_IOB_X0Y157_OPAD,
  output LIOB33_X0Y157_IOB_X0Y158_OPAD,
  output LIOB33_X0Y159_IOB_X0Y159_OPAD,
  output LIOB33_X0Y159_IOB_X0Y160_OPAD,
  output LIOB33_X0Y161_IOB_X0Y161_OPAD,
  output LIOB33_X0Y161_IOB_X0Y162_OPAD,
  output LIOB33_X0Y163_IOB_X0Y163_OPAD,
  output LIOB33_X0Y163_IOB_X0Y164_OPAD,
  output LIOB33_X0Y165_IOB_X0Y165_OPAD,
  output LIOB33_X0Y165_IOB_X0Y166_OPAD,
  output LIOB33_X0Y167_IOB_X0Y167_OPAD,
  output LIOB33_X0Y167_IOB_X0Y168_OPAD,
  output LIOB33_X0Y169_IOB_X0Y169_OPAD,
  output LIOB33_X0Y169_IOB_X0Y170_OPAD,
  output LIOB33_X0Y171_IOB_X0Y171_OPAD,
  output LIOB33_X0Y171_IOB_X0Y172_OPAD,
  output LIOB33_X0Y173_IOB_X0Y173_OPAD,
  output LIOB33_X0Y173_IOB_X0Y174_OPAD,
  output LIOB33_X0Y175_IOB_X0Y175_OPAD,
  output LIOB33_X0Y175_IOB_X0Y176_OPAD,
  output LIOB33_X0Y177_IOB_X0Y177_OPAD,
  output LIOB33_X0Y177_IOB_X0Y178_OPAD,
  output LIOB33_X0Y179_IOB_X0Y179_OPAD,
  output LIOB33_X0Y179_IOB_X0Y180_OPAD,
  output LIOB33_X0Y181_IOB_X0Y181_OPAD,
  output LIOB33_X0Y181_IOB_X0Y182_OPAD,
  output LIOB33_X0Y183_IOB_X0Y183_OPAD,
  output LIOB33_X0Y183_IOB_X0Y184_OPAD,
  output LIOB33_X0Y185_IOB_X0Y185_OPAD,
  output LIOB33_X0Y185_IOB_X0Y186_OPAD,
  output LIOB33_X0Y187_IOB_X0Y187_OPAD,
  output LIOB33_X0Y187_IOB_X0Y188_OPAD,
  output LIOB33_X0Y189_IOB_X0Y189_OPAD,
  output LIOB33_X0Y189_IOB_X0Y190_OPAD,
  output LIOB33_X0Y191_IOB_X0Y191_OPAD,
  output LIOB33_X0Y191_IOB_X0Y192_OPAD,
  output LIOB33_X0Y193_IOB_X0Y193_OPAD,
  output LIOB33_X0Y193_IOB_X0Y194_OPAD,
  output LIOB33_X0Y195_IOB_X0Y195_OPAD,
  output LIOB33_X0Y195_IOB_X0Y196_OPAD,
  output LIOB33_X0Y197_IOB_X0Y197_OPAD,
  output LIOB33_X0Y197_IOB_X0Y198_OPAD,
  output LIOB33_X0Y63_IOB_X0Y64_OPAD,
  output LIOB33_X0Y65_IOB_X0Y65_OPAD,
  output LIOB33_X0Y65_IOB_X0Y66_OPAD,
  output RIOB33_SING_X105Y150_IOB_X1Y150_OPAD,
  output RIOB33_SING_X105Y199_IOB_X1Y199_OPAD,
  output RIOB33_X105Y151_IOB_X1Y151_OPAD,
  output RIOB33_X105Y151_IOB_X1Y152_OPAD,
  output RIOB33_X105Y153_IOB_X1Y153_OPAD,
  output RIOB33_X105Y153_IOB_X1Y154_OPAD,
  output RIOB33_X105Y155_IOB_X1Y155_OPAD,
  output RIOB33_X105Y155_IOB_X1Y156_OPAD,
  output RIOB33_X105Y157_IOB_X1Y157_OPAD,
  output RIOB33_X105Y157_IOB_X1Y158_OPAD,
  output RIOB33_X105Y159_IOB_X1Y159_OPAD,
  output RIOB33_X105Y159_IOB_X1Y160_OPAD,
  output RIOB33_X105Y161_IOB_X1Y161_OPAD,
  output RIOB33_X105Y161_IOB_X1Y162_OPAD,
  output RIOB33_X105Y163_IOB_X1Y163_OPAD,
  output RIOB33_X105Y163_IOB_X1Y164_OPAD,
  output RIOB33_X105Y165_IOB_X1Y165_OPAD,
  output RIOB33_X105Y165_IOB_X1Y166_OPAD,
  output RIOB33_X105Y167_IOB_X1Y167_OPAD,
  output RIOB33_X105Y167_IOB_X1Y168_OPAD,
  output RIOB33_X105Y169_IOB_X1Y169_OPAD,
  output RIOB33_X105Y169_IOB_X1Y170_OPAD,
  output RIOB33_X105Y171_IOB_X1Y171_OPAD,
  output RIOB33_X105Y171_IOB_X1Y172_OPAD,
  output RIOB33_X105Y173_IOB_X1Y173_OPAD,
  output RIOB33_X105Y173_IOB_X1Y174_OPAD,
  output RIOB33_X105Y175_IOB_X1Y175_OPAD,
  output RIOB33_X105Y175_IOB_X1Y176_OPAD,
  output RIOB33_X105Y177_IOB_X1Y177_OPAD,
  output RIOB33_X105Y177_IOB_X1Y178_OPAD,
  output RIOB33_X105Y179_IOB_X1Y179_OPAD,
  output RIOB33_X105Y179_IOB_X1Y180_OPAD,
  output RIOB33_X105Y181_IOB_X1Y181_OPAD,
  output RIOB33_X105Y181_IOB_X1Y182_OPAD,
  output RIOB33_X105Y183_IOB_X1Y183_OPAD,
  output RIOB33_X105Y183_IOB_X1Y184_OPAD,
  output RIOB33_X105Y185_IOB_X1Y185_OPAD,
  output RIOB33_X105Y185_IOB_X1Y186_OPAD,
  output RIOB33_X105Y187_IOB_X1Y187_OPAD,
  output RIOB33_X105Y187_IOB_X1Y188_OPAD,
  output RIOB33_X105Y189_IOB_X1Y189_OPAD,
  output RIOB33_X105Y189_IOB_X1Y190_OPAD,
  output RIOB33_X105Y191_IOB_X1Y191_OPAD,
  output RIOB33_X105Y191_IOB_X1Y192_OPAD,
  output RIOB33_X105Y193_IOB_X1Y193_OPAD,
  output RIOB33_X105Y193_IOB_X1Y194_OPAD,
  output RIOB33_X105Y195_IOB_X1Y195_OPAD,
  output RIOB33_X105Y195_IOB_X1Y196_OPAD,
  output RIOB33_X105Y197_IOB_X1Y197_OPAD,
  output RIOB33_X105Y197_IOB_X1Y198_OPAD
  );
  wire [0:0] CLBLL_L_X2Y144_SLICE_X0Y144_A;
  wire [0:0] CLBLL_L_X2Y144_SLICE_X0Y144_A1;
  wire [0:0] CLBLL_L_X2Y144_SLICE_X0Y144_A2;
  wire [0:0] CLBLL_L_X2Y144_SLICE_X0Y144_A3;
  wire [0:0] CLBLL_L_X2Y144_SLICE_X0Y144_A4;
  wire [0:0] CLBLL_L_X2Y144_SLICE_X0Y144_A5;
  wire [0:0] CLBLL_L_X2Y144_SLICE_X0Y144_A6;
  wire [0:0] CLBLL_L_X2Y144_SLICE_X0Y144_AO5;
  wire [0:0] CLBLL_L_X2Y144_SLICE_X0Y144_AO6;
  wire [0:0] CLBLL_L_X2Y144_SLICE_X0Y144_A_CY;
  wire [0:0] CLBLL_L_X2Y144_SLICE_X0Y144_A_XOR;
  wire [0:0] CLBLL_L_X2Y144_SLICE_X0Y144_B;
  wire [0:0] CLBLL_L_X2Y144_SLICE_X0Y144_B1;
  wire [0:0] CLBLL_L_X2Y144_SLICE_X0Y144_B2;
  wire [0:0] CLBLL_L_X2Y144_SLICE_X0Y144_B3;
  wire [0:0] CLBLL_L_X2Y144_SLICE_X0Y144_B4;
  wire [0:0] CLBLL_L_X2Y144_SLICE_X0Y144_B5;
  wire [0:0] CLBLL_L_X2Y144_SLICE_X0Y144_B6;
  wire [0:0] CLBLL_L_X2Y144_SLICE_X0Y144_BO5;
  wire [0:0] CLBLL_L_X2Y144_SLICE_X0Y144_BO6;
  wire [0:0] CLBLL_L_X2Y144_SLICE_X0Y144_B_CY;
  wire [0:0] CLBLL_L_X2Y144_SLICE_X0Y144_B_XOR;
  wire [0:0] CLBLL_L_X2Y144_SLICE_X0Y144_C;
  wire [0:0] CLBLL_L_X2Y144_SLICE_X0Y144_C1;
  wire [0:0] CLBLL_L_X2Y144_SLICE_X0Y144_C2;
  wire [0:0] CLBLL_L_X2Y144_SLICE_X0Y144_C3;
  wire [0:0] CLBLL_L_X2Y144_SLICE_X0Y144_C4;
  wire [0:0] CLBLL_L_X2Y144_SLICE_X0Y144_C5;
  wire [0:0] CLBLL_L_X2Y144_SLICE_X0Y144_C6;
  wire [0:0] CLBLL_L_X2Y144_SLICE_X0Y144_CO5;
  wire [0:0] CLBLL_L_X2Y144_SLICE_X0Y144_CO6;
  wire [0:0] CLBLL_L_X2Y144_SLICE_X0Y144_C_CY;
  wire [0:0] CLBLL_L_X2Y144_SLICE_X0Y144_C_XOR;
  wire [0:0] CLBLL_L_X2Y144_SLICE_X0Y144_D;
  wire [0:0] CLBLL_L_X2Y144_SLICE_X0Y144_D1;
  wire [0:0] CLBLL_L_X2Y144_SLICE_X0Y144_D2;
  wire [0:0] CLBLL_L_X2Y144_SLICE_X0Y144_D3;
  wire [0:0] CLBLL_L_X2Y144_SLICE_X0Y144_D4;
  wire [0:0] CLBLL_L_X2Y144_SLICE_X0Y144_D5;
  wire [0:0] CLBLL_L_X2Y144_SLICE_X0Y144_D6;
  wire [0:0] CLBLL_L_X2Y144_SLICE_X0Y144_DO5;
  wire [0:0] CLBLL_L_X2Y144_SLICE_X0Y144_DO6;
  wire [0:0] CLBLL_L_X2Y144_SLICE_X0Y144_D_CY;
  wire [0:0] CLBLL_L_X2Y144_SLICE_X0Y144_D_XOR;
  wire [0:0] CLBLL_L_X2Y144_SLICE_X1Y144_A;
  wire [0:0] CLBLL_L_X2Y144_SLICE_X1Y144_A1;
  wire [0:0] CLBLL_L_X2Y144_SLICE_X1Y144_A2;
  wire [0:0] CLBLL_L_X2Y144_SLICE_X1Y144_A3;
  wire [0:0] CLBLL_L_X2Y144_SLICE_X1Y144_A4;
  wire [0:0] CLBLL_L_X2Y144_SLICE_X1Y144_A5;
  wire [0:0] CLBLL_L_X2Y144_SLICE_X1Y144_A6;
  wire [0:0] CLBLL_L_X2Y144_SLICE_X1Y144_AO5;
  wire [0:0] CLBLL_L_X2Y144_SLICE_X1Y144_AO6;
  wire [0:0] CLBLL_L_X2Y144_SLICE_X1Y144_A_CY;
  wire [0:0] CLBLL_L_X2Y144_SLICE_X1Y144_A_XOR;
  wire [0:0] CLBLL_L_X2Y144_SLICE_X1Y144_B;
  wire [0:0] CLBLL_L_X2Y144_SLICE_X1Y144_B1;
  wire [0:0] CLBLL_L_X2Y144_SLICE_X1Y144_B2;
  wire [0:0] CLBLL_L_X2Y144_SLICE_X1Y144_B3;
  wire [0:0] CLBLL_L_X2Y144_SLICE_X1Y144_B4;
  wire [0:0] CLBLL_L_X2Y144_SLICE_X1Y144_B5;
  wire [0:0] CLBLL_L_X2Y144_SLICE_X1Y144_B6;
  wire [0:0] CLBLL_L_X2Y144_SLICE_X1Y144_BO5;
  wire [0:0] CLBLL_L_X2Y144_SLICE_X1Y144_BO6;
  wire [0:0] CLBLL_L_X2Y144_SLICE_X1Y144_B_CY;
  wire [0:0] CLBLL_L_X2Y144_SLICE_X1Y144_B_XOR;
  wire [0:0] CLBLL_L_X2Y144_SLICE_X1Y144_C;
  wire [0:0] CLBLL_L_X2Y144_SLICE_X1Y144_C1;
  wire [0:0] CLBLL_L_X2Y144_SLICE_X1Y144_C2;
  wire [0:0] CLBLL_L_X2Y144_SLICE_X1Y144_C3;
  wire [0:0] CLBLL_L_X2Y144_SLICE_X1Y144_C4;
  wire [0:0] CLBLL_L_X2Y144_SLICE_X1Y144_C5;
  wire [0:0] CLBLL_L_X2Y144_SLICE_X1Y144_C6;
  wire [0:0] CLBLL_L_X2Y144_SLICE_X1Y144_CO5;
  wire [0:0] CLBLL_L_X2Y144_SLICE_X1Y144_CO6;
  wire [0:0] CLBLL_L_X2Y144_SLICE_X1Y144_C_CY;
  wire [0:0] CLBLL_L_X2Y144_SLICE_X1Y144_C_XOR;
  wire [0:0] CLBLL_L_X2Y144_SLICE_X1Y144_D;
  wire [0:0] CLBLL_L_X2Y144_SLICE_X1Y144_D1;
  wire [0:0] CLBLL_L_X2Y144_SLICE_X1Y144_D2;
  wire [0:0] CLBLL_L_X2Y144_SLICE_X1Y144_D3;
  wire [0:0] CLBLL_L_X2Y144_SLICE_X1Y144_D4;
  wire [0:0] CLBLL_L_X2Y144_SLICE_X1Y144_D5;
  wire [0:0] CLBLL_L_X2Y144_SLICE_X1Y144_D6;
  wire [0:0] CLBLL_L_X2Y144_SLICE_X1Y144_DO5;
  wire [0:0] CLBLL_L_X2Y144_SLICE_X1Y144_DO6;
  wire [0:0] CLBLL_L_X2Y144_SLICE_X1Y144_D_CY;
  wire [0:0] CLBLL_L_X2Y144_SLICE_X1Y144_D_XOR;
  wire [0:0] CLBLL_L_X2Y145_SLICE_X0Y145_A;
  wire [0:0] CLBLL_L_X2Y145_SLICE_X0Y145_A1;
  wire [0:0] CLBLL_L_X2Y145_SLICE_X0Y145_A2;
  wire [0:0] CLBLL_L_X2Y145_SLICE_X0Y145_A3;
  wire [0:0] CLBLL_L_X2Y145_SLICE_X0Y145_A4;
  wire [0:0] CLBLL_L_X2Y145_SLICE_X0Y145_A5;
  wire [0:0] CLBLL_L_X2Y145_SLICE_X0Y145_A6;
  wire [0:0] CLBLL_L_X2Y145_SLICE_X0Y145_AO5;
  wire [0:0] CLBLL_L_X2Y145_SLICE_X0Y145_AO6;
  wire [0:0] CLBLL_L_X2Y145_SLICE_X0Y145_AQ;
  wire [0:0] CLBLL_L_X2Y145_SLICE_X0Y145_A_CY;
  wire [0:0] CLBLL_L_X2Y145_SLICE_X0Y145_A_XOR;
  wire [0:0] CLBLL_L_X2Y145_SLICE_X0Y145_B;
  wire [0:0] CLBLL_L_X2Y145_SLICE_X0Y145_B1;
  wire [0:0] CLBLL_L_X2Y145_SLICE_X0Y145_B2;
  wire [0:0] CLBLL_L_X2Y145_SLICE_X0Y145_B3;
  wire [0:0] CLBLL_L_X2Y145_SLICE_X0Y145_B4;
  wire [0:0] CLBLL_L_X2Y145_SLICE_X0Y145_B5;
  wire [0:0] CLBLL_L_X2Y145_SLICE_X0Y145_B6;
  wire [0:0] CLBLL_L_X2Y145_SLICE_X0Y145_BO5;
  wire [0:0] CLBLL_L_X2Y145_SLICE_X0Y145_BO6;
  wire [0:0] CLBLL_L_X2Y145_SLICE_X0Y145_BQ;
  wire [0:0] CLBLL_L_X2Y145_SLICE_X0Y145_B_CY;
  wire [0:0] CLBLL_L_X2Y145_SLICE_X0Y145_B_XOR;
  wire [0:0] CLBLL_L_X2Y145_SLICE_X0Y145_C;
  wire [0:0] CLBLL_L_X2Y145_SLICE_X0Y145_C1;
  wire [0:0] CLBLL_L_X2Y145_SLICE_X0Y145_C2;
  wire [0:0] CLBLL_L_X2Y145_SLICE_X0Y145_C3;
  wire [0:0] CLBLL_L_X2Y145_SLICE_X0Y145_C4;
  wire [0:0] CLBLL_L_X2Y145_SLICE_X0Y145_C5;
  wire [0:0] CLBLL_L_X2Y145_SLICE_X0Y145_C6;
  wire [0:0] CLBLL_L_X2Y145_SLICE_X0Y145_CLK;
  wire [0:0] CLBLL_L_X2Y145_SLICE_X0Y145_CO5;
  wire [0:0] CLBLL_L_X2Y145_SLICE_X0Y145_CO6;
  wire [0:0] CLBLL_L_X2Y145_SLICE_X0Y145_C_CY;
  wire [0:0] CLBLL_L_X2Y145_SLICE_X0Y145_C_XOR;
  wire [0:0] CLBLL_L_X2Y145_SLICE_X0Y145_D;
  wire [0:0] CLBLL_L_X2Y145_SLICE_X0Y145_D1;
  wire [0:0] CLBLL_L_X2Y145_SLICE_X0Y145_D2;
  wire [0:0] CLBLL_L_X2Y145_SLICE_X0Y145_D3;
  wire [0:0] CLBLL_L_X2Y145_SLICE_X0Y145_D4;
  wire [0:0] CLBLL_L_X2Y145_SLICE_X0Y145_D5;
  wire [0:0] CLBLL_L_X2Y145_SLICE_X0Y145_D6;
  wire [0:0] CLBLL_L_X2Y145_SLICE_X0Y145_DO5;
  wire [0:0] CLBLL_L_X2Y145_SLICE_X0Y145_DO6;
  wire [0:0] CLBLL_L_X2Y145_SLICE_X0Y145_D_CY;
  wire [0:0] CLBLL_L_X2Y145_SLICE_X0Y145_D_XOR;
  wire [0:0] CLBLL_L_X2Y145_SLICE_X1Y145_A;
  wire [0:0] CLBLL_L_X2Y145_SLICE_X1Y145_A1;
  wire [0:0] CLBLL_L_X2Y145_SLICE_X1Y145_A2;
  wire [0:0] CLBLL_L_X2Y145_SLICE_X1Y145_A3;
  wire [0:0] CLBLL_L_X2Y145_SLICE_X1Y145_A4;
  wire [0:0] CLBLL_L_X2Y145_SLICE_X1Y145_A5;
  wire [0:0] CLBLL_L_X2Y145_SLICE_X1Y145_A6;
  wire [0:0] CLBLL_L_X2Y145_SLICE_X1Y145_AO5;
  wire [0:0] CLBLL_L_X2Y145_SLICE_X1Y145_AO6;
  wire [0:0] CLBLL_L_X2Y145_SLICE_X1Y145_AQ;
  wire [0:0] CLBLL_L_X2Y145_SLICE_X1Y145_A_CY;
  wire [0:0] CLBLL_L_X2Y145_SLICE_X1Y145_A_XOR;
  wire [0:0] CLBLL_L_X2Y145_SLICE_X1Y145_B;
  wire [0:0] CLBLL_L_X2Y145_SLICE_X1Y145_B1;
  wire [0:0] CLBLL_L_X2Y145_SLICE_X1Y145_B2;
  wire [0:0] CLBLL_L_X2Y145_SLICE_X1Y145_B3;
  wire [0:0] CLBLL_L_X2Y145_SLICE_X1Y145_B4;
  wire [0:0] CLBLL_L_X2Y145_SLICE_X1Y145_B5;
  wire [0:0] CLBLL_L_X2Y145_SLICE_X1Y145_B6;
  wire [0:0] CLBLL_L_X2Y145_SLICE_X1Y145_BO5;
  wire [0:0] CLBLL_L_X2Y145_SLICE_X1Y145_BO6;
  wire [0:0] CLBLL_L_X2Y145_SLICE_X1Y145_BQ;
  wire [0:0] CLBLL_L_X2Y145_SLICE_X1Y145_B_CY;
  wire [0:0] CLBLL_L_X2Y145_SLICE_X1Y145_B_XOR;
  wire [0:0] CLBLL_L_X2Y145_SLICE_X1Y145_C;
  wire [0:0] CLBLL_L_X2Y145_SLICE_X1Y145_C1;
  wire [0:0] CLBLL_L_X2Y145_SLICE_X1Y145_C2;
  wire [0:0] CLBLL_L_X2Y145_SLICE_X1Y145_C3;
  wire [0:0] CLBLL_L_X2Y145_SLICE_X1Y145_C4;
  wire [0:0] CLBLL_L_X2Y145_SLICE_X1Y145_C5;
  wire [0:0] CLBLL_L_X2Y145_SLICE_X1Y145_C6;
  wire [0:0] CLBLL_L_X2Y145_SLICE_X1Y145_CLK;
  wire [0:0] CLBLL_L_X2Y145_SLICE_X1Y145_CO5;
  wire [0:0] CLBLL_L_X2Y145_SLICE_X1Y145_CO6;
  wire [0:0] CLBLL_L_X2Y145_SLICE_X1Y145_CQ;
  wire [0:0] CLBLL_L_X2Y145_SLICE_X1Y145_C_CY;
  wire [0:0] CLBLL_L_X2Y145_SLICE_X1Y145_C_XOR;
  wire [0:0] CLBLL_L_X2Y145_SLICE_X1Y145_D;
  wire [0:0] CLBLL_L_X2Y145_SLICE_X1Y145_D1;
  wire [0:0] CLBLL_L_X2Y145_SLICE_X1Y145_D2;
  wire [0:0] CLBLL_L_X2Y145_SLICE_X1Y145_D3;
  wire [0:0] CLBLL_L_X2Y145_SLICE_X1Y145_D4;
  wire [0:0] CLBLL_L_X2Y145_SLICE_X1Y145_D5;
  wire [0:0] CLBLL_L_X2Y145_SLICE_X1Y145_D6;
  wire [0:0] CLBLL_L_X2Y145_SLICE_X1Y145_DMUX;
  wire [0:0] CLBLL_L_X2Y145_SLICE_X1Y145_DO5;
  wire [0:0] CLBLL_L_X2Y145_SLICE_X1Y145_DO6;
  wire [0:0] CLBLL_L_X2Y145_SLICE_X1Y145_D_CY;
  wire [0:0] CLBLL_L_X2Y145_SLICE_X1Y145_D_XOR;
  wire [0:0] CLBLL_L_X2Y146_SLICE_X0Y146_A;
  wire [0:0] CLBLL_L_X2Y146_SLICE_X0Y146_A1;
  wire [0:0] CLBLL_L_X2Y146_SLICE_X0Y146_A2;
  wire [0:0] CLBLL_L_X2Y146_SLICE_X0Y146_A3;
  wire [0:0] CLBLL_L_X2Y146_SLICE_X0Y146_A4;
  wire [0:0] CLBLL_L_X2Y146_SLICE_X0Y146_A5;
  wire [0:0] CLBLL_L_X2Y146_SLICE_X0Y146_A6;
  wire [0:0] CLBLL_L_X2Y146_SLICE_X0Y146_AO5;
  wire [0:0] CLBLL_L_X2Y146_SLICE_X0Y146_AO6;
  wire [0:0] CLBLL_L_X2Y146_SLICE_X0Y146_AQ;
  wire [0:0] CLBLL_L_X2Y146_SLICE_X0Y146_A_CY;
  wire [0:0] CLBLL_L_X2Y146_SLICE_X0Y146_A_XOR;
  wire [0:0] CLBLL_L_X2Y146_SLICE_X0Y146_B;
  wire [0:0] CLBLL_L_X2Y146_SLICE_X0Y146_B1;
  wire [0:0] CLBLL_L_X2Y146_SLICE_X0Y146_B2;
  wire [0:0] CLBLL_L_X2Y146_SLICE_X0Y146_B3;
  wire [0:0] CLBLL_L_X2Y146_SLICE_X0Y146_B4;
  wire [0:0] CLBLL_L_X2Y146_SLICE_X0Y146_B5;
  wire [0:0] CLBLL_L_X2Y146_SLICE_X0Y146_B6;
  wire [0:0] CLBLL_L_X2Y146_SLICE_X0Y146_BO5;
  wire [0:0] CLBLL_L_X2Y146_SLICE_X0Y146_BO6;
  wire [0:0] CLBLL_L_X2Y146_SLICE_X0Y146_BQ;
  wire [0:0] CLBLL_L_X2Y146_SLICE_X0Y146_B_CY;
  wire [0:0] CLBLL_L_X2Y146_SLICE_X0Y146_B_XOR;
  wire [0:0] CLBLL_L_X2Y146_SLICE_X0Y146_C;
  wire [0:0] CLBLL_L_X2Y146_SLICE_X0Y146_C1;
  wire [0:0] CLBLL_L_X2Y146_SLICE_X0Y146_C2;
  wire [0:0] CLBLL_L_X2Y146_SLICE_X0Y146_C3;
  wire [0:0] CLBLL_L_X2Y146_SLICE_X0Y146_C4;
  wire [0:0] CLBLL_L_X2Y146_SLICE_X0Y146_C5;
  wire [0:0] CLBLL_L_X2Y146_SLICE_X0Y146_C6;
  wire [0:0] CLBLL_L_X2Y146_SLICE_X0Y146_CLK;
  wire [0:0] CLBLL_L_X2Y146_SLICE_X0Y146_CO5;
  wire [0:0] CLBLL_L_X2Y146_SLICE_X0Y146_CO6;
  wire [0:0] CLBLL_L_X2Y146_SLICE_X0Y146_CQ;
  wire [0:0] CLBLL_L_X2Y146_SLICE_X0Y146_C_CY;
  wire [0:0] CLBLL_L_X2Y146_SLICE_X0Y146_C_XOR;
  wire [0:0] CLBLL_L_X2Y146_SLICE_X0Y146_D;
  wire [0:0] CLBLL_L_X2Y146_SLICE_X0Y146_D1;
  wire [0:0] CLBLL_L_X2Y146_SLICE_X0Y146_D2;
  wire [0:0] CLBLL_L_X2Y146_SLICE_X0Y146_D3;
  wire [0:0] CLBLL_L_X2Y146_SLICE_X0Y146_D4;
  wire [0:0] CLBLL_L_X2Y146_SLICE_X0Y146_D5;
  wire [0:0] CLBLL_L_X2Y146_SLICE_X0Y146_D6;
  wire [0:0] CLBLL_L_X2Y146_SLICE_X0Y146_DO5;
  wire [0:0] CLBLL_L_X2Y146_SLICE_X0Y146_DO6;
  wire [0:0] CLBLL_L_X2Y146_SLICE_X0Y146_DQ;
  wire [0:0] CLBLL_L_X2Y146_SLICE_X0Y146_D_CY;
  wire [0:0] CLBLL_L_X2Y146_SLICE_X0Y146_D_XOR;
  wire [0:0] CLBLL_L_X2Y146_SLICE_X1Y146_A;
  wire [0:0] CLBLL_L_X2Y146_SLICE_X1Y146_A1;
  wire [0:0] CLBLL_L_X2Y146_SLICE_X1Y146_A2;
  wire [0:0] CLBLL_L_X2Y146_SLICE_X1Y146_A3;
  wire [0:0] CLBLL_L_X2Y146_SLICE_X1Y146_A4;
  wire [0:0] CLBLL_L_X2Y146_SLICE_X1Y146_A5;
  wire [0:0] CLBLL_L_X2Y146_SLICE_X1Y146_A6;
  wire [0:0] CLBLL_L_X2Y146_SLICE_X1Y146_AO5;
  wire [0:0] CLBLL_L_X2Y146_SLICE_X1Y146_AO6;
  wire [0:0] CLBLL_L_X2Y146_SLICE_X1Y146_AQ;
  wire [0:0] CLBLL_L_X2Y146_SLICE_X1Y146_A_CY;
  wire [0:0] CLBLL_L_X2Y146_SLICE_X1Y146_A_XOR;
  wire [0:0] CLBLL_L_X2Y146_SLICE_X1Y146_B;
  wire [0:0] CLBLL_L_X2Y146_SLICE_X1Y146_B1;
  wire [0:0] CLBLL_L_X2Y146_SLICE_X1Y146_B2;
  wire [0:0] CLBLL_L_X2Y146_SLICE_X1Y146_B3;
  wire [0:0] CLBLL_L_X2Y146_SLICE_X1Y146_B4;
  wire [0:0] CLBLL_L_X2Y146_SLICE_X1Y146_B5;
  wire [0:0] CLBLL_L_X2Y146_SLICE_X1Y146_B5Q;
  wire [0:0] CLBLL_L_X2Y146_SLICE_X1Y146_B6;
  wire [0:0] CLBLL_L_X2Y146_SLICE_X1Y146_BMUX;
  wire [0:0] CLBLL_L_X2Y146_SLICE_X1Y146_BO5;
  wire [0:0] CLBLL_L_X2Y146_SLICE_X1Y146_BO6;
  wire [0:0] CLBLL_L_X2Y146_SLICE_X1Y146_BQ;
  wire [0:0] CLBLL_L_X2Y146_SLICE_X1Y146_B_CY;
  wire [0:0] CLBLL_L_X2Y146_SLICE_X1Y146_B_XOR;
  wire [0:0] CLBLL_L_X2Y146_SLICE_X1Y146_C;
  wire [0:0] CLBLL_L_X2Y146_SLICE_X1Y146_C1;
  wire [0:0] CLBLL_L_X2Y146_SLICE_X1Y146_C2;
  wire [0:0] CLBLL_L_X2Y146_SLICE_X1Y146_C3;
  wire [0:0] CLBLL_L_X2Y146_SLICE_X1Y146_C4;
  wire [0:0] CLBLL_L_X2Y146_SLICE_X1Y146_C5;
  wire [0:0] CLBLL_L_X2Y146_SLICE_X1Y146_C6;
  wire [0:0] CLBLL_L_X2Y146_SLICE_X1Y146_CLK;
  wire [0:0] CLBLL_L_X2Y146_SLICE_X1Y146_CMUX;
  wire [0:0] CLBLL_L_X2Y146_SLICE_X1Y146_CO5;
  wire [0:0] CLBLL_L_X2Y146_SLICE_X1Y146_CO6;
  wire [0:0] CLBLL_L_X2Y146_SLICE_X1Y146_C_CY;
  wire [0:0] CLBLL_L_X2Y146_SLICE_X1Y146_C_XOR;
  wire [0:0] CLBLL_L_X2Y146_SLICE_X1Y146_D;
  wire [0:0] CLBLL_L_X2Y146_SLICE_X1Y146_D1;
  wire [0:0] CLBLL_L_X2Y146_SLICE_X1Y146_D2;
  wire [0:0] CLBLL_L_X2Y146_SLICE_X1Y146_D3;
  wire [0:0] CLBLL_L_X2Y146_SLICE_X1Y146_D4;
  wire [0:0] CLBLL_L_X2Y146_SLICE_X1Y146_D5;
  wire [0:0] CLBLL_L_X2Y146_SLICE_X1Y146_D6;
  wire [0:0] CLBLL_L_X2Y146_SLICE_X1Y146_DO5;
  wire [0:0] CLBLL_L_X2Y146_SLICE_X1Y146_DO6;
  wire [0:0] CLBLL_L_X2Y146_SLICE_X1Y146_D_CY;
  wire [0:0] CLBLL_L_X2Y146_SLICE_X1Y146_D_XOR;
  wire [0:0] CLBLL_L_X2Y147_SLICE_X0Y147_A;
  wire [0:0] CLBLL_L_X2Y147_SLICE_X0Y147_A1;
  wire [0:0] CLBLL_L_X2Y147_SLICE_X0Y147_A2;
  wire [0:0] CLBLL_L_X2Y147_SLICE_X0Y147_A3;
  wire [0:0] CLBLL_L_X2Y147_SLICE_X0Y147_A4;
  wire [0:0] CLBLL_L_X2Y147_SLICE_X0Y147_A5;
  wire [0:0] CLBLL_L_X2Y147_SLICE_X0Y147_A6;
  wire [0:0] CLBLL_L_X2Y147_SLICE_X0Y147_AO5;
  wire [0:0] CLBLL_L_X2Y147_SLICE_X0Y147_AO6;
  wire [0:0] CLBLL_L_X2Y147_SLICE_X0Y147_A_CY;
  wire [0:0] CLBLL_L_X2Y147_SLICE_X0Y147_A_XOR;
  wire [0:0] CLBLL_L_X2Y147_SLICE_X0Y147_B;
  wire [0:0] CLBLL_L_X2Y147_SLICE_X0Y147_B1;
  wire [0:0] CLBLL_L_X2Y147_SLICE_X0Y147_B2;
  wire [0:0] CLBLL_L_X2Y147_SLICE_X0Y147_B3;
  wire [0:0] CLBLL_L_X2Y147_SLICE_X0Y147_B4;
  wire [0:0] CLBLL_L_X2Y147_SLICE_X0Y147_B5;
  wire [0:0] CLBLL_L_X2Y147_SLICE_X0Y147_B6;
  wire [0:0] CLBLL_L_X2Y147_SLICE_X0Y147_BO5;
  wire [0:0] CLBLL_L_X2Y147_SLICE_X0Y147_BO6;
  wire [0:0] CLBLL_L_X2Y147_SLICE_X0Y147_B_CY;
  wire [0:0] CLBLL_L_X2Y147_SLICE_X0Y147_B_XOR;
  wire [0:0] CLBLL_L_X2Y147_SLICE_X0Y147_C;
  wire [0:0] CLBLL_L_X2Y147_SLICE_X0Y147_C1;
  wire [0:0] CLBLL_L_X2Y147_SLICE_X0Y147_C2;
  wire [0:0] CLBLL_L_X2Y147_SLICE_X0Y147_C3;
  wire [0:0] CLBLL_L_X2Y147_SLICE_X0Y147_C4;
  wire [0:0] CLBLL_L_X2Y147_SLICE_X0Y147_C5;
  wire [0:0] CLBLL_L_X2Y147_SLICE_X0Y147_C6;
  wire [0:0] CLBLL_L_X2Y147_SLICE_X0Y147_CO5;
  wire [0:0] CLBLL_L_X2Y147_SLICE_X0Y147_CO6;
  wire [0:0] CLBLL_L_X2Y147_SLICE_X0Y147_C_CY;
  wire [0:0] CLBLL_L_X2Y147_SLICE_X0Y147_C_XOR;
  wire [0:0] CLBLL_L_X2Y147_SLICE_X0Y147_D;
  wire [0:0] CLBLL_L_X2Y147_SLICE_X0Y147_D1;
  wire [0:0] CLBLL_L_X2Y147_SLICE_X0Y147_D2;
  wire [0:0] CLBLL_L_X2Y147_SLICE_X0Y147_D3;
  wire [0:0] CLBLL_L_X2Y147_SLICE_X0Y147_D4;
  wire [0:0] CLBLL_L_X2Y147_SLICE_X0Y147_D5;
  wire [0:0] CLBLL_L_X2Y147_SLICE_X0Y147_D6;
  wire [0:0] CLBLL_L_X2Y147_SLICE_X0Y147_DO5;
  wire [0:0] CLBLL_L_X2Y147_SLICE_X0Y147_DO6;
  wire [0:0] CLBLL_L_X2Y147_SLICE_X0Y147_D_CY;
  wire [0:0] CLBLL_L_X2Y147_SLICE_X0Y147_D_XOR;
  wire [0:0] CLBLL_L_X2Y147_SLICE_X1Y147_A;
  wire [0:0] CLBLL_L_X2Y147_SLICE_X1Y147_A1;
  wire [0:0] CLBLL_L_X2Y147_SLICE_X1Y147_A2;
  wire [0:0] CLBLL_L_X2Y147_SLICE_X1Y147_A3;
  wire [0:0] CLBLL_L_X2Y147_SLICE_X1Y147_A4;
  wire [0:0] CLBLL_L_X2Y147_SLICE_X1Y147_A5;
  wire [0:0] CLBLL_L_X2Y147_SLICE_X1Y147_A6;
  wire [0:0] CLBLL_L_X2Y147_SLICE_X1Y147_AO5;
  wire [0:0] CLBLL_L_X2Y147_SLICE_X1Y147_AO6;
  wire [0:0] CLBLL_L_X2Y147_SLICE_X1Y147_A_CY;
  wire [0:0] CLBLL_L_X2Y147_SLICE_X1Y147_A_XOR;
  wire [0:0] CLBLL_L_X2Y147_SLICE_X1Y147_B;
  wire [0:0] CLBLL_L_X2Y147_SLICE_X1Y147_B1;
  wire [0:0] CLBLL_L_X2Y147_SLICE_X1Y147_B2;
  wire [0:0] CLBLL_L_X2Y147_SLICE_X1Y147_B3;
  wire [0:0] CLBLL_L_X2Y147_SLICE_X1Y147_B4;
  wire [0:0] CLBLL_L_X2Y147_SLICE_X1Y147_B5;
  wire [0:0] CLBLL_L_X2Y147_SLICE_X1Y147_B6;
  wire [0:0] CLBLL_L_X2Y147_SLICE_X1Y147_BO5;
  wire [0:0] CLBLL_L_X2Y147_SLICE_X1Y147_BO6;
  wire [0:0] CLBLL_L_X2Y147_SLICE_X1Y147_B_CY;
  wire [0:0] CLBLL_L_X2Y147_SLICE_X1Y147_B_XOR;
  wire [0:0] CLBLL_L_X2Y147_SLICE_X1Y147_C;
  wire [0:0] CLBLL_L_X2Y147_SLICE_X1Y147_C1;
  wire [0:0] CLBLL_L_X2Y147_SLICE_X1Y147_C2;
  wire [0:0] CLBLL_L_X2Y147_SLICE_X1Y147_C3;
  wire [0:0] CLBLL_L_X2Y147_SLICE_X1Y147_C4;
  wire [0:0] CLBLL_L_X2Y147_SLICE_X1Y147_C5;
  wire [0:0] CLBLL_L_X2Y147_SLICE_X1Y147_C6;
  wire [0:0] CLBLL_L_X2Y147_SLICE_X1Y147_CO5;
  wire [0:0] CLBLL_L_X2Y147_SLICE_X1Y147_CO6;
  wire [0:0] CLBLL_L_X2Y147_SLICE_X1Y147_C_CY;
  wire [0:0] CLBLL_L_X2Y147_SLICE_X1Y147_C_XOR;
  wire [0:0] CLBLL_L_X2Y147_SLICE_X1Y147_D;
  wire [0:0] CLBLL_L_X2Y147_SLICE_X1Y147_D1;
  wire [0:0] CLBLL_L_X2Y147_SLICE_X1Y147_D2;
  wire [0:0] CLBLL_L_X2Y147_SLICE_X1Y147_D3;
  wire [0:0] CLBLL_L_X2Y147_SLICE_X1Y147_D4;
  wire [0:0] CLBLL_L_X2Y147_SLICE_X1Y147_D5;
  wire [0:0] CLBLL_L_X2Y147_SLICE_X1Y147_D6;
  wire [0:0] CLBLL_L_X2Y147_SLICE_X1Y147_DO5;
  wire [0:0] CLBLL_L_X2Y147_SLICE_X1Y147_DO6;
  wire [0:0] CLBLL_L_X2Y147_SLICE_X1Y147_D_CY;
  wire [0:0] CLBLL_L_X2Y147_SLICE_X1Y147_D_XOR;
  wire [0:0] CLBLL_L_X2Y148_SLICE_X0Y148_A;
  wire [0:0] CLBLL_L_X2Y148_SLICE_X0Y148_A1;
  wire [0:0] CLBLL_L_X2Y148_SLICE_X0Y148_A2;
  wire [0:0] CLBLL_L_X2Y148_SLICE_X0Y148_A3;
  wire [0:0] CLBLL_L_X2Y148_SLICE_X0Y148_A4;
  wire [0:0] CLBLL_L_X2Y148_SLICE_X0Y148_A5;
  wire [0:0] CLBLL_L_X2Y148_SLICE_X0Y148_A6;
  wire [0:0] CLBLL_L_X2Y148_SLICE_X0Y148_AO5;
  wire [0:0] CLBLL_L_X2Y148_SLICE_X0Y148_AO6;
  wire [0:0] CLBLL_L_X2Y148_SLICE_X0Y148_AQ;
  wire [0:0] CLBLL_L_X2Y148_SLICE_X0Y148_AX;
  wire [0:0] CLBLL_L_X2Y148_SLICE_X0Y148_A_CY;
  wire [0:0] CLBLL_L_X2Y148_SLICE_X0Y148_A_XOR;
  wire [0:0] CLBLL_L_X2Y148_SLICE_X0Y148_B;
  wire [0:0] CLBLL_L_X2Y148_SLICE_X0Y148_B1;
  wire [0:0] CLBLL_L_X2Y148_SLICE_X0Y148_B2;
  wire [0:0] CLBLL_L_X2Y148_SLICE_X0Y148_B3;
  wire [0:0] CLBLL_L_X2Y148_SLICE_X0Y148_B4;
  wire [0:0] CLBLL_L_X2Y148_SLICE_X0Y148_B5;
  wire [0:0] CLBLL_L_X2Y148_SLICE_X0Y148_B6;
  wire [0:0] CLBLL_L_X2Y148_SLICE_X0Y148_BO5;
  wire [0:0] CLBLL_L_X2Y148_SLICE_X0Y148_BO6;
  wire [0:0] CLBLL_L_X2Y148_SLICE_X0Y148_B_CY;
  wire [0:0] CLBLL_L_X2Y148_SLICE_X0Y148_B_XOR;
  wire [0:0] CLBLL_L_X2Y148_SLICE_X0Y148_C;
  wire [0:0] CLBLL_L_X2Y148_SLICE_X0Y148_C1;
  wire [0:0] CLBLL_L_X2Y148_SLICE_X0Y148_C2;
  wire [0:0] CLBLL_L_X2Y148_SLICE_X0Y148_C3;
  wire [0:0] CLBLL_L_X2Y148_SLICE_X0Y148_C4;
  wire [0:0] CLBLL_L_X2Y148_SLICE_X0Y148_C5;
  wire [0:0] CLBLL_L_X2Y148_SLICE_X0Y148_C6;
  wire [0:0] CLBLL_L_X2Y148_SLICE_X0Y148_CE;
  wire [0:0] CLBLL_L_X2Y148_SLICE_X0Y148_CLK;
  wire [0:0] CLBLL_L_X2Y148_SLICE_X0Y148_CO5;
  wire [0:0] CLBLL_L_X2Y148_SLICE_X0Y148_CO6;
  wire [0:0] CLBLL_L_X2Y148_SLICE_X0Y148_C_CY;
  wire [0:0] CLBLL_L_X2Y148_SLICE_X0Y148_C_XOR;
  wire [0:0] CLBLL_L_X2Y148_SLICE_X0Y148_D;
  wire [0:0] CLBLL_L_X2Y148_SLICE_X0Y148_D1;
  wire [0:0] CLBLL_L_X2Y148_SLICE_X0Y148_D2;
  wire [0:0] CLBLL_L_X2Y148_SLICE_X0Y148_D3;
  wire [0:0] CLBLL_L_X2Y148_SLICE_X0Y148_D4;
  wire [0:0] CLBLL_L_X2Y148_SLICE_X0Y148_D5;
  wire [0:0] CLBLL_L_X2Y148_SLICE_X0Y148_D6;
  wire [0:0] CLBLL_L_X2Y148_SLICE_X0Y148_DO5;
  wire [0:0] CLBLL_L_X2Y148_SLICE_X0Y148_DO6;
  wire [0:0] CLBLL_L_X2Y148_SLICE_X0Y148_D_CY;
  wire [0:0] CLBLL_L_X2Y148_SLICE_X0Y148_D_XOR;
  wire [0:0] CLBLL_L_X2Y148_SLICE_X1Y148_A;
  wire [0:0] CLBLL_L_X2Y148_SLICE_X1Y148_A1;
  wire [0:0] CLBLL_L_X2Y148_SLICE_X1Y148_A2;
  wire [0:0] CLBLL_L_X2Y148_SLICE_X1Y148_A3;
  wire [0:0] CLBLL_L_X2Y148_SLICE_X1Y148_A4;
  wire [0:0] CLBLL_L_X2Y148_SLICE_X1Y148_A5;
  wire [0:0] CLBLL_L_X2Y148_SLICE_X1Y148_A6;
  wire [0:0] CLBLL_L_X2Y148_SLICE_X1Y148_AO5;
  wire [0:0] CLBLL_L_X2Y148_SLICE_X1Y148_AO6;
  wire [0:0] CLBLL_L_X2Y148_SLICE_X1Y148_A_CY;
  wire [0:0] CLBLL_L_X2Y148_SLICE_X1Y148_A_XOR;
  wire [0:0] CLBLL_L_X2Y148_SLICE_X1Y148_B;
  wire [0:0] CLBLL_L_X2Y148_SLICE_X1Y148_B1;
  wire [0:0] CLBLL_L_X2Y148_SLICE_X1Y148_B2;
  wire [0:0] CLBLL_L_X2Y148_SLICE_X1Y148_B3;
  wire [0:0] CLBLL_L_X2Y148_SLICE_X1Y148_B4;
  wire [0:0] CLBLL_L_X2Y148_SLICE_X1Y148_B5;
  wire [0:0] CLBLL_L_X2Y148_SLICE_X1Y148_B6;
  wire [0:0] CLBLL_L_X2Y148_SLICE_X1Y148_BO5;
  wire [0:0] CLBLL_L_X2Y148_SLICE_X1Y148_BO6;
  wire [0:0] CLBLL_L_X2Y148_SLICE_X1Y148_B_CY;
  wire [0:0] CLBLL_L_X2Y148_SLICE_X1Y148_B_XOR;
  wire [0:0] CLBLL_L_X2Y148_SLICE_X1Y148_C;
  wire [0:0] CLBLL_L_X2Y148_SLICE_X1Y148_C1;
  wire [0:0] CLBLL_L_X2Y148_SLICE_X1Y148_C2;
  wire [0:0] CLBLL_L_X2Y148_SLICE_X1Y148_C3;
  wire [0:0] CLBLL_L_X2Y148_SLICE_X1Y148_C4;
  wire [0:0] CLBLL_L_X2Y148_SLICE_X1Y148_C5;
  wire [0:0] CLBLL_L_X2Y148_SLICE_X1Y148_C6;
  wire [0:0] CLBLL_L_X2Y148_SLICE_X1Y148_CO5;
  wire [0:0] CLBLL_L_X2Y148_SLICE_X1Y148_CO6;
  wire [0:0] CLBLL_L_X2Y148_SLICE_X1Y148_C_CY;
  wire [0:0] CLBLL_L_X2Y148_SLICE_X1Y148_C_XOR;
  wire [0:0] CLBLL_L_X2Y148_SLICE_X1Y148_D;
  wire [0:0] CLBLL_L_X2Y148_SLICE_X1Y148_D1;
  wire [0:0] CLBLL_L_X2Y148_SLICE_X1Y148_D2;
  wire [0:0] CLBLL_L_X2Y148_SLICE_X1Y148_D3;
  wire [0:0] CLBLL_L_X2Y148_SLICE_X1Y148_D4;
  wire [0:0] CLBLL_L_X2Y148_SLICE_X1Y148_D5;
  wire [0:0] CLBLL_L_X2Y148_SLICE_X1Y148_D6;
  wire [0:0] CLBLL_L_X2Y148_SLICE_X1Y148_DO5;
  wire [0:0] CLBLL_L_X2Y148_SLICE_X1Y148_DO6;
  wire [0:0] CLBLL_L_X2Y148_SLICE_X1Y148_D_CY;
  wire [0:0] CLBLL_L_X2Y148_SLICE_X1Y148_D_XOR;
  wire [0:0] CLBLL_L_X2Y150_SLICE_X0Y150_A;
  wire [0:0] CLBLL_L_X2Y150_SLICE_X0Y150_A1;
  wire [0:0] CLBLL_L_X2Y150_SLICE_X0Y150_A2;
  wire [0:0] CLBLL_L_X2Y150_SLICE_X0Y150_A3;
  wire [0:0] CLBLL_L_X2Y150_SLICE_X0Y150_A4;
  wire [0:0] CLBLL_L_X2Y150_SLICE_X0Y150_A5;
  wire [0:0] CLBLL_L_X2Y150_SLICE_X0Y150_A6;
  wire [0:0] CLBLL_L_X2Y150_SLICE_X0Y150_AO5;
  wire [0:0] CLBLL_L_X2Y150_SLICE_X0Y150_AO6;
  wire [0:0] CLBLL_L_X2Y150_SLICE_X0Y150_A_CY;
  wire [0:0] CLBLL_L_X2Y150_SLICE_X0Y150_A_XOR;
  wire [0:0] CLBLL_L_X2Y150_SLICE_X0Y150_B;
  wire [0:0] CLBLL_L_X2Y150_SLICE_X0Y150_B1;
  wire [0:0] CLBLL_L_X2Y150_SLICE_X0Y150_B2;
  wire [0:0] CLBLL_L_X2Y150_SLICE_X0Y150_B3;
  wire [0:0] CLBLL_L_X2Y150_SLICE_X0Y150_B4;
  wire [0:0] CLBLL_L_X2Y150_SLICE_X0Y150_B5;
  wire [0:0] CLBLL_L_X2Y150_SLICE_X0Y150_B6;
  wire [0:0] CLBLL_L_X2Y150_SLICE_X0Y150_BO5;
  wire [0:0] CLBLL_L_X2Y150_SLICE_X0Y150_BO6;
  wire [0:0] CLBLL_L_X2Y150_SLICE_X0Y150_B_CY;
  wire [0:0] CLBLL_L_X2Y150_SLICE_X0Y150_B_XOR;
  wire [0:0] CLBLL_L_X2Y150_SLICE_X0Y150_C;
  wire [0:0] CLBLL_L_X2Y150_SLICE_X0Y150_C1;
  wire [0:0] CLBLL_L_X2Y150_SLICE_X0Y150_C2;
  wire [0:0] CLBLL_L_X2Y150_SLICE_X0Y150_C3;
  wire [0:0] CLBLL_L_X2Y150_SLICE_X0Y150_C4;
  wire [0:0] CLBLL_L_X2Y150_SLICE_X0Y150_C5;
  wire [0:0] CLBLL_L_X2Y150_SLICE_X0Y150_C6;
  wire [0:0] CLBLL_L_X2Y150_SLICE_X0Y150_CO5;
  wire [0:0] CLBLL_L_X2Y150_SLICE_X0Y150_CO6;
  wire [0:0] CLBLL_L_X2Y150_SLICE_X0Y150_C_CY;
  wire [0:0] CLBLL_L_X2Y150_SLICE_X0Y150_C_XOR;
  wire [0:0] CLBLL_L_X2Y150_SLICE_X0Y150_D;
  wire [0:0] CLBLL_L_X2Y150_SLICE_X0Y150_D1;
  wire [0:0] CLBLL_L_X2Y150_SLICE_X0Y150_D2;
  wire [0:0] CLBLL_L_X2Y150_SLICE_X0Y150_D3;
  wire [0:0] CLBLL_L_X2Y150_SLICE_X0Y150_D4;
  wire [0:0] CLBLL_L_X2Y150_SLICE_X0Y150_D5;
  wire [0:0] CLBLL_L_X2Y150_SLICE_X0Y150_D6;
  wire [0:0] CLBLL_L_X2Y150_SLICE_X0Y150_DO5;
  wire [0:0] CLBLL_L_X2Y150_SLICE_X0Y150_DO6;
  wire [0:0] CLBLL_L_X2Y150_SLICE_X0Y150_D_CY;
  wire [0:0] CLBLL_L_X2Y150_SLICE_X0Y150_D_XOR;
  wire [0:0] CLBLL_L_X2Y150_SLICE_X1Y150_A;
  wire [0:0] CLBLL_L_X2Y150_SLICE_X1Y150_A1;
  wire [0:0] CLBLL_L_X2Y150_SLICE_X1Y150_A2;
  wire [0:0] CLBLL_L_X2Y150_SLICE_X1Y150_A3;
  wire [0:0] CLBLL_L_X2Y150_SLICE_X1Y150_A4;
  wire [0:0] CLBLL_L_X2Y150_SLICE_X1Y150_A5;
  wire [0:0] CLBLL_L_X2Y150_SLICE_X1Y150_A6;
  wire [0:0] CLBLL_L_X2Y150_SLICE_X1Y150_AO5;
  wire [0:0] CLBLL_L_X2Y150_SLICE_X1Y150_AO6;
  wire [0:0] CLBLL_L_X2Y150_SLICE_X1Y150_AQ;
  wire [0:0] CLBLL_L_X2Y150_SLICE_X1Y150_A_CY;
  wire [0:0] CLBLL_L_X2Y150_SLICE_X1Y150_A_XOR;
  wire [0:0] CLBLL_L_X2Y150_SLICE_X1Y150_B;
  wire [0:0] CLBLL_L_X2Y150_SLICE_X1Y150_B1;
  wire [0:0] CLBLL_L_X2Y150_SLICE_X1Y150_B2;
  wire [0:0] CLBLL_L_X2Y150_SLICE_X1Y150_B3;
  wire [0:0] CLBLL_L_X2Y150_SLICE_X1Y150_B4;
  wire [0:0] CLBLL_L_X2Y150_SLICE_X1Y150_B5;
  wire [0:0] CLBLL_L_X2Y150_SLICE_X1Y150_B6;
  wire [0:0] CLBLL_L_X2Y150_SLICE_X1Y150_BO5;
  wire [0:0] CLBLL_L_X2Y150_SLICE_X1Y150_BO6;
  wire [0:0] CLBLL_L_X2Y150_SLICE_X1Y150_B_CY;
  wire [0:0] CLBLL_L_X2Y150_SLICE_X1Y150_B_XOR;
  wire [0:0] CLBLL_L_X2Y150_SLICE_X1Y150_C;
  wire [0:0] CLBLL_L_X2Y150_SLICE_X1Y150_C1;
  wire [0:0] CLBLL_L_X2Y150_SLICE_X1Y150_C2;
  wire [0:0] CLBLL_L_X2Y150_SLICE_X1Y150_C3;
  wire [0:0] CLBLL_L_X2Y150_SLICE_X1Y150_C4;
  wire [0:0] CLBLL_L_X2Y150_SLICE_X1Y150_C5;
  wire [0:0] CLBLL_L_X2Y150_SLICE_X1Y150_C6;
  wire [0:0] CLBLL_L_X2Y150_SLICE_X1Y150_CLK;
  wire [0:0] CLBLL_L_X2Y150_SLICE_X1Y150_CO5;
  wire [0:0] CLBLL_L_X2Y150_SLICE_X1Y150_CO6;
  wire [0:0] CLBLL_L_X2Y150_SLICE_X1Y150_C_CY;
  wire [0:0] CLBLL_L_X2Y150_SLICE_X1Y150_C_XOR;
  wire [0:0] CLBLL_L_X2Y150_SLICE_X1Y150_D;
  wire [0:0] CLBLL_L_X2Y150_SLICE_X1Y150_D1;
  wire [0:0] CLBLL_L_X2Y150_SLICE_X1Y150_D2;
  wire [0:0] CLBLL_L_X2Y150_SLICE_X1Y150_D3;
  wire [0:0] CLBLL_L_X2Y150_SLICE_X1Y150_D4;
  wire [0:0] CLBLL_L_X2Y150_SLICE_X1Y150_D5;
  wire [0:0] CLBLL_L_X2Y150_SLICE_X1Y150_D6;
  wire [0:0] CLBLL_L_X2Y150_SLICE_X1Y150_DO5;
  wire [0:0] CLBLL_L_X2Y150_SLICE_X1Y150_DO6;
  wire [0:0] CLBLL_L_X2Y150_SLICE_X1Y150_D_CY;
  wire [0:0] CLBLL_L_X2Y150_SLICE_X1Y150_D_XOR;
  wire [0:0] CLBLL_L_X2Y166_SLICE_X0Y166_A;
  wire [0:0] CLBLL_L_X2Y166_SLICE_X0Y166_A1;
  wire [0:0] CLBLL_L_X2Y166_SLICE_X0Y166_A2;
  wire [0:0] CLBLL_L_X2Y166_SLICE_X0Y166_A3;
  wire [0:0] CLBLL_L_X2Y166_SLICE_X0Y166_A4;
  wire [0:0] CLBLL_L_X2Y166_SLICE_X0Y166_A5;
  wire [0:0] CLBLL_L_X2Y166_SLICE_X0Y166_A6;
  wire [0:0] CLBLL_L_X2Y166_SLICE_X0Y166_AO5;
  wire [0:0] CLBLL_L_X2Y166_SLICE_X0Y166_AO6;
  wire [0:0] CLBLL_L_X2Y166_SLICE_X0Y166_A_CY;
  wire [0:0] CLBLL_L_X2Y166_SLICE_X0Y166_A_XOR;
  wire [0:0] CLBLL_L_X2Y166_SLICE_X0Y166_B;
  wire [0:0] CLBLL_L_X2Y166_SLICE_X0Y166_B1;
  wire [0:0] CLBLL_L_X2Y166_SLICE_X0Y166_B2;
  wire [0:0] CLBLL_L_X2Y166_SLICE_X0Y166_B3;
  wire [0:0] CLBLL_L_X2Y166_SLICE_X0Y166_B4;
  wire [0:0] CLBLL_L_X2Y166_SLICE_X0Y166_B5;
  wire [0:0] CLBLL_L_X2Y166_SLICE_X0Y166_B6;
  wire [0:0] CLBLL_L_X2Y166_SLICE_X0Y166_BO5;
  wire [0:0] CLBLL_L_X2Y166_SLICE_X0Y166_BO6;
  wire [0:0] CLBLL_L_X2Y166_SLICE_X0Y166_B_CY;
  wire [0:0] CLBLL_L_X2Y166_SLICE_X0Y166_B_XOR;
  wire [0:0] CLBLL_L_X2Y166_SLICE_X0Y166_C;
  wire [0:0] CLBLL_L_X2Y166_SLICE_X0Y166_C1;
  wire [0:0] CLBLL_L_X2Y166_SLICE_X0Y166_C2;
  wire [0:0] CLBLL_L_X2Y166_SLICE_X0Y166_C3;
  wire [0:0] CLBLL_L_X2Y166_SLICE_X0Y166_C4;
  wire [0:0] CLBLL_L_X2Y166_SLICE_X0Y166_C5;
  wire [0:0] CLBLL_L_X2Y166_SLICE_X0Y166_C6;
  wire [0:0] CLBLL_L_X2Y166_SLICE_X0Y166_CO5;
  wire [0:0] CLBLL_L_X2Y166_SLICE_X0Y166_CO6;
  wire [0:0] CLBLL_L_X2Y166_SLICE_X0Y166_C_CY;
  wire [0:0] CLBLL_L_X2Y166_SLICE_X0Y166_C_XOR;
  wire [0:0] CLBLL_L_X2Y166_SLICE_X0Y166_D;
  wire [0:0] CLBLL_L_X2Y166_SLICE_X0Y166_D1;
  wire [0:0] CLBLL_L_X2Y166_SLICE_X0Y166_D2;
  wire [0:0] CLBLL_L_X2Y166_SLICE_X0Y166_D3;
  wire [0:0] CLBLL_L_X2Y166_SLICE_X0Y166_D4;
  wire [0:0] CLBLL_L_X2Y166_SLICE_X0Y166_D5;
  wire [0:0] CLBLL_L_X2Y166_SLICE_X0Y166_D6;
  wire [0:0] CLBLL_L_X2Y166_SLICE_X0Y166_DO5;
  wire [0:0] CLBLL_L_X2Y166_SLICE_X0Y166_DO6;
  wire [0:0] CLBLL_L_X2Y166_SLICE_X0Y166_D_CY;
  wire [0:0] CLBLL_L_X2Y166_SLICE_X0Y166_D_XOR;
  wire [0:0] CLBLL_L_X2Y166_SLICE_X1Y166_A;
  wire [0:0] CLBLL_L_X2Y166_SLICE_X1Y166_A1;
  wire [0:0] CLBLL_L_X2Y166_SLICE_X1Y166_A2;
  wire [0:0] CLBLL_L_X2Y166_SLICE_X1Y166_A3;
  wire [0:0] CLBLL_L_X2Y166_SLICE_X1Y166_A4;
  wire [0:0] CLBLL_L_X2Y166_SLICE_X1Y166_A5;
  wire [0:0] CLBLL_L_X2Y166_SLICE_X1Y166_A6;
  wire [0:0] CLBLL_L_X2Y166_SLICE_X1Y166_AO5;
  wire [0:0] CLBLL_L_X2Y166_SLICE_X1Y166_AO6;
  wire [0:0] CLBLL_L_X2Y166_SLICE_X1Y166_A_CY;
  wire [0:0] CLBLL_L_X2Y166_SLICE_X1Y166_A_XOR;
  wire [0:0] CLBLL_L_X2Y166_SLICE_X1Y166_B;
  wire [0:0] CLBLL_L_X2Y166_SLICE_X1Y166_B1;
  wire [0:0] CLBLL_L_X2Y166_SLICE_X1Y166_B2;
  wire [0:0] CLBLL_L_X2Y166_SLICE_X1Y166_B3;
  wire [0:0] CLBLL_L_X2Y166_SLICE_X1Y166_B4;
  wire [0:0] CLBLL_L_X2Y166_SLICE_X1Y166_B5;
  wire [0:0] CLBLL_L_X2Y166_SLICE_X1Y166_B6;
  wire [0:0] CLBLL_L_X2Y166_SLICE_X1Y166_BO5;
  wire [0:0] CLBLL_L_X2Y166_SLICE_X1Y166_BO6;
  wire [0:0] CLBLL_L_X2Y166_SLICE_X1Y166_B_CY;
  wire [0:0] CLBLL_L_X2Y166_SLICE_X1Y166_B_XOR;
  wire [0:0] CLBLL_L_X2Y166_SLICE_X1Y166_C;
  wire [0:0] CLBLL_L_X2Y166_SLICE_X1Y166_C1;
  wire [0:0] CLBLL_L_X2Y166_SLICE_X1Y166_C2;
  wire [0:0] CLBLL_L_X2Y166_SLICE_X1Y166_C3;
  wire [0:0] CLBLL_L_X2Y166_SLICE_X1Y166_C4;
  wire [0:0] CLBLL_L_X2Y166_SLICE_X1Y166_C5;
  wire [0:0] CLBLL_L_X2Y166_SLICE_X1Y166_C6;
  wire [0:0] CLBLL_L_X2Y166_SLICE_X1Y166_CO5;
  wire [0:0] CLBLL_L_X2Y166_SLICE_X1Y166_CO6;
  wire [0:0] CLBLL_L_X2Y166_SLICE_X1Y166_C_CY;
  wire [0:0] CLBLL_L_X2Y166_SLICE_X1Y166_C_XOR;
  wire [0:0] CLBLL_L_X2Y166_SLICE_X1Y166_D;
  wire [0:0] CLBLL_L_X2Y166_SLICE_X1Y166_D1;
  wire [0:0] CLBLL_L_X2Y166_SLICE_X1Y166_D2;
  wire [0:0] CLBLL_L_X2Y166_SLICE_X1Y166_D3;
  wire [0:0] CLBLL_L_X2Y166_SLICE_X1Y166_D4;
  wire [0:0] CLBLL_L_X2Y166_SLICE_X1Y166_D5;
  wire [0:0] CLBLL_L_X2Y166_SLICE_X1Y166_D6;
  wire [0:0] CLBLL_L_X2Y166_SLICE_X1Y166_DO5;
  wire [0:0] CLBLL_L_X2Y166_SLICE_X1Y166_DO6;
  wire [0:0] CLBLL_L_X2Y166_SLICE_X1Y166_D_CY;
  wire [0:0] CLBLL_L_X2Y166_SLICE_X1Y166_D_XOR;
  wire [0:0] CLBLL_L_X2Y75_SLICE_X0Y75_A;
  wire [0:0] CLBLL_L_X2Y75_SLICE_X0Y75_A1;
  wire [0:0] CLBLL_L_X2Y75_SLICE_X0Y75_A2;
  wire [0:0] CLBLL_L_X2Y75_SLICE_X0Y75_A3;
  wire [0:0] CLBLL_L_X2Y75_SLICE_X0Y75_A4;
  wire [0:0] CLBLL_L_X2Y75_SLICE_X0Y75_A5;
  wire [0:0] CLBLL_L_X2Y75_SLICE_X0Y75_A6;
  wire [0:0] CLBLL_L_X2Y75_SLICE_X0Y75_AO5;
  wire [0:0] CLBLL_L_X2Y75_SLICE_X0Y75_AO6;
  wire [0:0] CLBLL_L_X2Y75_SLICE_X0Y75_A_CY;
  wire [0:0] CLBLL_L_X2Y75_SLICE_X0Y75_A_XOR;
  wire [0:0] CLBLL_L_X2Y75_SLICE_X0Y75_B;
  wire [0:0] CLBLL_L_X2Y75_SLICE_X0Y75_B1;
  wire [0:0] CLBLL_L_X2Y75_SLICE_X0Y75_B2;
  wire [0:0] CLBLL_L_X2Y75_SLICE_X0Y75_B3;
  wire [0:0] CLBLL_L_X2Y75_SLICE_X0Y75_B4;
  wire [0:0] CLBLL_L_X2Y75_SLICE_X0Y75_B5;
  wire [0:0] CLBLL_L_X2Y75_SLICE_X0Y75_B6;
  wire [0:0] CLBLL_L_X2Y75_SLICE_X0Y75_BO5;
  wire [0:0] CLBLL_L_X2Y75_SLICE_X0Y75_BO6;
  wire [0:0] CLBLL_L_X2Y75_SLICE_X0Y75_B_CY;
  wire [0:0] CLBLL_L_X2Y75_SLICE_X0Y75_B_XOR;
  wire [0:0] CLBLL_L_X2Y75_SLICE_X0Y75_C;
  wire [0:0] CLBLL_L_X2Y75_SLICE_X0Y75_C1;
  wire [0:0] CLBLL_L_X2Y75_SLICE_X0Y75_C2;
  wire [0:0] CLBLL_L_X2Y75_SLICE_X0Y75_C3;
  wire [0:0] CLBLL_L_X2Y75_SLICE_X0Y75_C4;
  wire [0:0] CLBLL_L_X2Y75_SLICE_X0Y75_C5;
  wire [0:0] CLBLL_L_X2Y75_SLICE_X0Y75_C6;
  wire [0:0] CLBLL_L_X2Y75_SLICE_X0Y75_CO5;
  wire [0:0] CLBLL_L_X2Y75_SLICE_X0Y75_CO6;
  wire [0:0] CLBLL_L_X2Y75_SLICE_X0Y75_C_CY;
  wire [0:0] CLBLL_L_X2Y75_SLICE_X0Y75_C_XOR;
  wire [0:0] CLBLL_L_X2Y75_SLICE_X0Y75_D;
  wire [0:0] CLBLL_L_X2Y75_SLICE_X0Y75_D1;
  wire [0:0] CLBLL_L_X2Y75_SLICE_X0Y75_D2;
  wire [0:0] CLBLL_L_X2Y75_SLICE_X0Y75_D3;
  wire [0:0] CLBLL_L_X2Y75_SLICE_X0Y75_D4;
  wire [0:0] CLBLL_L_X2Y75_SLICE_X0Y75_D5;
  wire [0:0] CLBLL_L_X2Y75_SLICE_X0Y75_D6;
  wire [0:0] CLBLL_L_X2Y75_SLICE_X0Y75_DO5;
  wire [0:0] CLBLL_L_X2Y75_SLICE_X0Y75_DO6;
  wire [0:0] CLBLL_L_X2Y75_SLICE_X0Y75_D_CY;
  wire [0:0] CLBLL_L_X2Y75_SLICE_X0Y75_D_XOR;
  wire [0:0] CLBLL_L_X2Y75_SLICE_X1Y75_A;
  wire [0:0] CLBLL_L_X2Y75_SLICE_X1Y75_A1;
  wire [0:0] CLBLL_L_X2Y75_SLICE_X1Y75_A2;
  wire [0:0] CLBLL_L_X2Y75_SLICE_X1Y75_A3;
  wire [0:0] CLBLL_L_X2Y75_SLICE_X1Y75_A4;
  wire [0:0] CLBLL_L_X2Y75_SLICE_X1Y75_A5;
  wire [0:0] CLBLL_L_X2Y75_SLICE_X1Y75_A6;
  wire [0:0] CLBLL_L_X2Y75_SLICE_X1Y75_AO5;
  wire [0:0] CLBLL_L_X2Y75_SLICE_X1Y75_AO6;
  wire [0:0] CLBLL_L_X2Y75_SLICE_X1Y75_A_CY;
  wire [0:0] CLBLL_L_X2Y75_SLICE_X1Y75_A_XOR;
  wire [0:0] CLBLL_L_X2Y75_SLICE_X1Y75_B;
  wire [0:0] CLBLL_L_X2Y75_SLICE_X1Y75_B1;
  wire [0:0] CLBLL_L_X2Y75_SLICE_X1Y75_B2;
  wire [0:0] CLBLL_L_X2Y75_SLICE_X1Y75_B3;
  wire [0:0] CLBLL_L_X2Y75_SLICE_X1Y75_B4;
  wire [0:0] CLBLL_L_X2Y75_SLICE_X1Y75_B5;
  wire [0:0] CLBLL_L_X2Y75_SLICE_X1Y75_B6;
  wire [0:0] CLBLL_L_X2Y75_SLICE_X1Y75_BO5;
  wire [0:0] CLBLL_L_X2Y75_SLICE_X1Y75_BO6;
  wire [0:0] CLBLL_L_X2Y75_SLICE_X1Y75_B_CY;
  wire [0:0] CLBLL_L_X2Y75_SLICE_X1Y75_B_XOR;
  wire [0:0] CLBLL_L_X2Y75_SLICE_X1Y75_C;
  wire [0:0] CLBLL_L_X2Y75_SLICE_X1Y75_C1;
  wire [0:0] CLBLL_L_X2Y75_SLICE_X1Y75_C2;
  wire [0:0] CLBLL_L_X2Y75_SLICE_X1Y75_C3;
  wire [0:0] CLBLL_L_X2Y75_SLICE_X1Y75_C4;
  wire [0:0] CLBLL_L_X2Y75_SLICE_X1Y75_C5;
  wire [0:0] CLBLL_L_X2Y75_SLICE_X1Y75_C6;
  wire [0:0] CLBLL_L_X2Y75_SLICE_X1Y75_CO5;
  wire [0:0] CLBLL_L_X2Y75_SLICE_X1Y75_CO6;
  wire [0:0] CLBLL_L_X2Y75_SLICE_X1Y75_C_CY;
  wire [0:0] CLBLL_L_X2Y75_SLICE_X1Y75_C_XOR;
  wire [0:0] CLBLL_L_X2Y75_SLICE_X1Y75_D;
  wire [0:0] CLBLL_L_X2Y75_SLICE_X1Y75_D1;
  wire [0:0] CLBLL_L_X2Y75_SLICE_X1Y75_D2;
  wire [0:0] CLBLL_L_X2Y75_SLICE_X1Y75_D3;
  wire [0:0] CLBLL_L_X2Y75_SLICE_X1Y75_D4;
  wire [0:0] CLBLL_L_X2Y75_SLICE_X1Y75_D5;
  wire [0:0] CLBLL_L_X2Y75_SLICE_X1Y75_D6;
  wire [0:0] CLBLL_L_X2Y75_SLICE_X1Y75_DO5;
  wire [0:0] CLBLL_L_X2Y75_SLICE_X1Y75_DO6;
  wire [0:0] CLBLL_L_X2Y75_SLICE_X1Y75_D_CY;
  wire [0:0] CLBLL_L_X2Y75_SLICE_X1Y75_D_XOR;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X4Y140_A;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X4Y140_A1;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X4Y140_A2;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X4Y140_A3;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X4Y140_A4;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X4Y140_A5;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X4Y140_A5Q;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X4Y140_A6;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X4Y140_AMUX;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X4Y140_AO5;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X4Y140_AO6;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X4Y140_AQ;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X4Y140_AX;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X4Y140_A_CY;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X4Y140_A_XOR;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X4Y140_B;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X4Y140_B1;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X4Y140_B2;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X4Y140_B3;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X4Y140_B4;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X4Y140_B5;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X4Y140_B6;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X4Y140_BMUX;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X4Y140_BO5;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X4Y140_BO6;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X4Y140_B_CY;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X4Y140_B_XOR;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X4Y140_C;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X4Y140_C1;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X4Y140_C2;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X4Y140_C3;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X4Y140_C4;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X4Y140_C5;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X4Y140_C6;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X4Y140_CLK;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X4Y140_CO5;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X4Y140_CO6;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X4Y140_C_CY;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X4Y140_C_XOR;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X4Y140_D;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X4Y140_D1;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X4Y140_D2;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X4Y140_D3;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X4Y140_D4;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X4Y140_D5;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X4Y140_D6;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X4Y140_DO5;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X4Y140_DO6;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X4Y140_D_CY;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X4Y140_D_XOR;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X5Y140_A;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X5Y140_A1;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X5Y140_A2;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X5Y140_A3;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X5Y140_A4;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X5Y140_A5;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X5Y140_A6;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X5Y140_AO5;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X5Y140_AO6;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X5Y140_AQ;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X5Y140_A_CY;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X5Y140_A_XOR;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X5Y140_B;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X5Y140_B1;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X5Y140_B2;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X5Y140_B3;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X5Y140_B4;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X5Y140_B5;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X5Y140_B6;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X5Y140_BO5;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X5Y140_BO6;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X5Y140_BQ;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X5Y140_B_CY;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X5Y140_B_XOR;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X5Y140_C;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X5Y140_C1;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X5Y140_C2;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X5Y140_C3;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X5Y140_C4;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X5Y140_C5;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X5Y140_C6;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X5Y140_CLK;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X5Y140_CMUX;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X5Y140_CO5;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X5Y140_CO6;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X5Y140_C_CY;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X5Y140_C_XOR;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X5Y140_D;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X5Y140_D1;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X5Y140_D2;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X5Y140_D3;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X5Y140_D4;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X5Y140_D5;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X5Y140_D6;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X5Y140_DO5;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X5Y140_DO6;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X5Y140_D_CY;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X5Y140_D_XOR;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X4Y142_A;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X4Y142_A1;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X4Y142_A2;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X4Y142_A3;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X4Y142_A4;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X4Y142_A5;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X4Y142_A5Q;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X4Y142_A6;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X4Y142_AMUX;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X4Y142_AO5;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X4Y142_AO6;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X4Y142_AQ;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X4Y142_AX;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X4Y142_A_CY;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X4Y142_A_XOR;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X4Y142_B;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X4Y142_B1;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X4Y142_B2;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X4Y142_B3;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X4Y142_B4;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X4Y142_B5;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X4Y142_B6;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X4Y142_BO5;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X4Y142_BO6;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X4Y142_BQ;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X4Y142_B_CY;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X4Y142_B_XOR;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X4Y142_C;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X4Y142_C1;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X4Y142_C2;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X4Y142_C3;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X4Y142_C4;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X4Y142_C5;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X4Y142_C6;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X4Y142_CLK;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X4Y142_CO5;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X4Y142_CO6;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X4Y142_CQ;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X4Y142_C_CY;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X4Y142_C_XOR;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X4Y142_D;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X4Y142_D1;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X4Y142_D2;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X4Y142_D3;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X4Y142_D4;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X4Y142_D5;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X4Y142_D6;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X4Y142_DO5;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X4Y142_DO6;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X4Y142_D_CY;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X4Y142_D_XOR;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X5Y142_A;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X5Y142_A1;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X5Y142_A2;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X5Y142_A3;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X5Y142_A4;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X5Y142_A5;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X5Y142_A6;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X5Y142_AO5;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X5Y142_AO6;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X5Y142_AQ;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X5Y142_A_CY;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X5Y142_A_XOR;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X5Y142_B;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X5Y142_B1;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X5Y142_B2;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X5Y142_B3;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X5Y142_B4;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X5Y142_B5;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X5Y142_B6;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X5Y142_BO5;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X5Y142_BO6;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X5Y142_BQ;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X5Y142_B_CY;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X5Y142_B_XOR;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X5Y142_C;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X5Y142_C1;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X5Y142_C2;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X5Y142_C3;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X5Y142_C4;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X5Y142_C5;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X5Y142_C5Q;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X5Y142_C6;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X5Y142_CLK;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X5Y142_CMUX;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X5Y142_CO5;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X5Y142_CO6;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X5Y142_CQ;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X5Y142_C_CY;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X5Y142_C_XOR;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X5Y142_D;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X5Y142_D1;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X5Y142_D2;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X5Y142_D3;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X5Y142_D4;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X5Y142_D5;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X5Y142_D5Q;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X5Y142_D6;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X5Y142_DMUX;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X5Y142_DO5;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X5Y142_DO6;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X5Y142_DQ;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X5Y142_D_CY;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X5Y142_D_XOR;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X4Y143_A;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X4Y143_A1;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X4Y143_A2;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X4Y143_A3;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X4Y143_A4;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X4Y143_A5;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X4Y143_A5Q;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X4Y143_A6;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X4Y143_AMUX;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X4Y143_AO5;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X4Y143_AO6;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X4Y143_AQ;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X4Y143_AX;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X4Y143_A_CY;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X4Y143_A_XOR;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X4Y143_B;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X4Y143_B1;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X4Y143_B2;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X4Y143_B3;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X4Y143_B4;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X4Y143_B5;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X4Y143_B6;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X4Y143_BMUX;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X4Y143_BO5;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X4Y143_BO6;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X4Y143_BQ;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X4Y143_B_CY;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X4Y143_B_XOR;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X4Y143_C;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X4Y143_C1;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X4Y143_C2;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X4Y143_C3;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X4Y143_C4;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X4Y143_C5;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X4Y143_C5Q;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X4Y143_C6;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X4Y143_CLK;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X4Y143_CMUX;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X4Y143_CO5;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X4Y143_CO6;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X4Y143_CQ;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X4Y143_C_CY;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X4Y143_C_XOR;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X4Y143_D;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X4Y143_D1;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X4Y143_D2;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X4Y143_D3;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X4Y143_D4;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X4Y143_D5;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X4Y143_D5Q;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X4Y143_D6;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X4Y143_DMUX;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X4Y143_DO5;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X4Y143_DO6;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X4Y143_DQ;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X4Y143_D_CY;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X4Y143_D_XOR;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X5Y143_A;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X5Y143_A1;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X5Y143_A2;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X5Y143_A3;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X5Y143_A4;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X5Y143_A5;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X5Y143_A6;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X5Y143_AO5;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X5Y143_AO6;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X5Y143_AQ;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X5Y143_A_CY;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X5Y143_A_XOR;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X5Y143_B;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X5Y143_B1;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X5Y143_B2;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X5Y143_B3;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X5Y143_B4;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X5Y143_B5;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X5Y143_B5Q;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X5Y143_B6;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X5Y143_BMUX;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X5Y143_BO5;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X5Y143_BO6;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X5Y143_BQ;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X5Y143_B_CY;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X5Y143_B_XOR;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X5Y143_C;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X5Y143_C1;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X5Y143_C2;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X5Y143_C3;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X5Y143_C4;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X5Y143_C5;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X5Y143_C6;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X5Y143_CLK;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X5Y143_CMUX;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X5Y143_CO5;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X5Y143_CO6;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X5Y143_C_CY;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X5Y143_C_XOR;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X5Y143_D;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X5Y143_D1;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X5Y143_D2;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X5Y143_D3;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X5Y143_D4;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X5Y143_D5;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X5Y143_D5Q;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X5Y143_D6;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X5Y143_DMUX;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X5Y143_DO5;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X5Y143_DO6;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X5Y143_DQ;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X5Y143_D_CY;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X5Y143_D_XOR;
  wire [0:0] CLBLL_L_X4Y144_SLICE_X4Y144_A;
  wire [0:0] CLBLL_L_X4Y144_SLICE_X4Y144_A1;
  wire [0:0] CLBLL_L_X4Y144_SLICE_X4Y144_A2;
  wire [0:0] CLBLL_L_X4Y144_SLICE_X4Y144_A3;
  wire [0:0] CLBLL_L_X4Y144_SLICE_X4Y144_A4;
  wire [0:0] CLBLL_L_X4Y144_SLICE_X4Y144_A5;
  wire [0:0] CLBLL_L_X4Y144_SLICE_X4Y144_A6;
  wire [0:0] CLBLL_L_X4Y144_SLICE_X4Y144_AO5;
  wire [0:0] CLBLL_L_X4Y144_SLICE_X4Y144_AO6;
  wire [0:0] CLBLL_L_X4Y144_SLICE_X4Y144_AQ;
  wire [0:0] CLBLL_L_X4Y144_SLICE_X4Y144_A_CY;
  wire [0:0] CLBLL_L_X4Y144_SLICE_X4Y144_A_XOR;
  wire [0:0] CLBLL_L_X4Y144_SLICE_X4Y144_B;
  wire [0:0] CLBLL_L_X4Y144_SLICE_X4Y144_B1;
  wire [0:0] CLBLL_L_X4Y144_SLICE_X4Y144_B2;
  wire [0:0] CLBLL_L_X4Y144_SLICE_X4Y144_B3;
  wire [0:0] CLBLL_L_X4Y144_SLICE_X4Y144_B4;
  wire [0:0] CLBLL_L_X4Y144_SLICE_X4Y144_B5;
  wire [0:0] CLBLL_L_X4Y144_SLICE_X4Y144_B5Q;
  wire [0:0] CLBLL_L_X4Y144_SLICE_X4Y144_B6;
  wire [0:0] CLBLL_L_X4Y144_SLICE_X4Y144_BMUX;
  wire [0:0] CLBLL_L_X4Y144_SLICE_X4Y144_BO5;
  wire [0:0] CLBLL_L_X4Y144_SLICE_X4Y144_BO6;
  wire [0:0] CLBLL_L_X4Y144_SLICE_X4Y144_BQ;
  wire [0:0] CLBLL_L_X4Y144_SLICE_X4Y144_B_CY;
  wire [0:0] CLBLL_L_X4Y144_SLICE_X4Y144_B_XOR;
  wire [0:0] CLBLL_L_X4Y144_SLICE_X4Y144_C;
  wire [0:0] CLBLL_L_X4Y144_SLICE_X4Y144_C1;
  wire [0:0] CLBLL_L_X4Y144_SLICE_X4Y144_C2;
  wire [0:0] CLBLL_L_X4Y144_SLICE_X4Y144_C3;
  wire [0:0] CLBLL_L_X4Y144_SLICE_X4Y144_C4;
  wire [0:0] CLBLL_L_X4Y144_SLICE_X4Y144_C5;
  wire [0:0] CLBLL_L_X4Y144_SLICE_X4Y144_C5Q;
  wire [0:0] CLBLL_L_X4Y144_SLICE_X4Y144_C6;
  wire [0:0] CLBLL_L_X4Y144_SLICE_X4Y144_CLK;
  wire [0:0] CLBLL_L_X4Y144_SLICE_X4Y144_CMUX;
  wire [0:0] CLBLL_L_X4Y144_SLICE_X4Y144_CO5;
  wire [0:0] CLBLL_L_X4Y144_SLICE_X4Y144_CO6;
  wire [0:0] CLBLL_L_X4Y144_SLICE_X4Y144_CQ;
  wire [0:0] CLBLL_L_X4Y144_SLICE_X4Y144_C_CY;
  wire [0:0] CLBLL_L_X4Y144_SLICE_X4Y144_C_XOR;
  wire [0:0] CLBLL_L_X4Y144_SLICE_X4Y144_D;
  wire [0:0] CLBLL_L_X4Y144_SLICE_X4Y144_D1;
  wire [0:0] CLBLL_L_X4Y144_SLICE_X4Y144_D2;
  wire [0:0] CLBLL_L_X4Y144_SLICE_X4Y144_D3;
  wire [0:0] CLBLL_L_X4Y144_SLICE_X4Y144_D4;
  wire [0:0] CLBLL_L_X4Y144_SLICE_X4Y144_D5;
  wire [0:0] CLBLL_L_X4Y144_SLICE_X4Y144_D5Q;
  wire [0:0] CLBLL_L_X4Y144_SLICE_X4Y144_D6;
  wire [0:0] CLBLL_L_X4Y144_SLICE_X4Y144_DMUX;
  wire [0:0] CLBLL_L_X4Y144_SLICE_X4Y144_DO5;
  wire [0:0] CLBLL_L_X4Y144_SLICE_X4Y144_DO6;
  wire [0:0] CLBLL_L_X4Y144_SLICE_X4Y144_DQ;
  wire [0:0] CLBLL_L_X4Y144_SLICE_X4Y144_D_CY;
  wire [0:0] CLBLL_L_X4Y144_SLICE_X4Y144_D_XOR;
  wire [0:0] CLBLL_L_X4Y144_SLICE_X5Y144_A;
  wire [0:0] CLBLL_L_X4Y144_SLICE_X5Y144_A1;
  wire [0:0] CLBLL_L_X4Y144_SLICE_X5Y144_A2;
  wire [0:0] CLBLL_L_X4Y144_SLICE_X5Y144_A3;
  wire [0:0] CLBLL_L_X4Y144_SLICE_X5Y144_A4;
  wire [0:0] CLBLL_L_X4Y144_SLICE_X5Y144_A5;
  wire [0:0] CLBLL_L_X4Y144_SLICE_X5Y144_A6;
  wire [0:0] CLBLL_L_X4Y144_SLICE_X5Y144_AO5;
  wire [0:0] CLBLL_L_X4Y144_SLICE_X5Y144_AO6;
  wire [0:0] CLBLL_L_X4Y144_SLICE_X5Y144_AQ;
  wire [0:0] CLBLL_L_X4Y144_SLICE_X5Y144_A_CY;
  wire [0:0] CLBLL_L_X4Y144_SLICE_X5Y144_A_XOR;
  wire [0:0] CLBLL_L_X4Y144_SLICE_X5Y144_B;
  wire [0:0] CLBLL_L_X4Y144_SLICE_X5Y144_B1;
  wire [0:0] CLBLL_L_X4Y144_SLICE_X5Y144_B2;
  wire [0:0] CLBLL_L_X4Y144_SLICE_X5Y144_B3;
  wire [0:0] CLBLL_L_X4Y144_SLICE_X5Y144_B4;
  wire [0:0] CLBLL_L_X4Y144_SLICE_X5Y144_B5;
  wire [0:0] CLBLL_L_X4Y144_SLICE_X5Y144_B6;
  wire [0:0] CLBLL_L_X4Y144_SLICE_X5Y144_BO5;
  wire [0:0] CLBLL_L_X4Y144_SLICE_X5Y144_BO6;
  wire [0:0] CLBLL_L_X4Y144_SLICE_X5Y144_BQ;
  wire [0:0] CLBLL_L_X4Y144_SLICE_X5Y144_B_CY;
  wire [0:0] CLBLL_L_X4Y144_SLICE_X5Y144_B_XOR;
  wire [0:0] CLBLL_L_X4Y144_SLICE_X5Y144_C;
  wire [0:0] CLBLL_L_X4Y144_SLICE_X5Y144_C1;
  wire [0:0] CLBLL_L_X4Y144_SLICE_X5Y144_C2;
  wire [0:0] CLBLL_L_X4Y144_SLICE_X5Y144_C3;
  wire [0:0] CLBLL_L_X4Y144_SLICE_X5Y144_C4;
  wire [0:0] CLBLL_L_X4Y144_SLICE_X5Y144_C5;
  wire [0:0] CLBLL_L_X4Y144_SLICE_X5Y144_C6;
  wire [0:0] CLBLL_L_X4Y144_SLICE_X5Y144_CLK;
  wire [0:0] CLBLL_L_X4Y144_SLICE_X5Y144_CO5;
  wire [0:0] CLBLL_L_X4Y144_SLICE_X5Y144_CO6;
  wire [0:0] CLBLL_L_X4Y144_SLICE_X5Y144_CQ;
  wire [0:0] CLBLL_L_X4Y144_SLICE_X5Y144_C_CY;
  wire [0:0] CLBLL_L_X4Y144_SLICE_X5Y144_C_XOR;
  wire [0:0] CLBLL_L_X4Y144_SLICE_X5Y144_D;
  wire [0:0] CLBLL_L_X4Y144_SLICE_X5Y144_D1;
  wire [0:0] CLBLL_L_X4Y144_SLICE_X5Y144_D2;
  wire [0:0] CLBLL_L_X4Y144_SLICE_X5Y144_D3;
  wire [0:0] CLBLL_L_X4Y144_SLICE_X5Y144_D4;
  wire [0:0] CLBLL_L_X4Y144_SLICE_X5Y144_D5;
  wire [0:0] CLBLL_L_X4Y144_SLICE_X5Y144_D5Q;
  wire [0:0] CLBLL_L_X4Y144_SLICE_X5Y144_D6;
  wire [0:0] CLBLL_L_X4Y144_SLICE_X5Y144_DMUX;
  wire [0:0] CLBLL_L_X4Y144_SLICE_X5Y144_DO5;
  wire [0:0] CLBLL_L_X4Y144_SLICE_X5Y144_DO6;
  wire [0:0] CLBLL_L_X4Y144_SLICE_X5Y144_DQ;
  wire [0:0] CLBLL_L_X4Y144_SLICE_X5Y144_D_CY;
  wire [0:0] CLBLL_L_X4Y144_SLICE_X5Y144_D_XOR;
  wire [0:0] CLBLL_L_X4Y145_SLICE_X4Y145_A;
  wire [0:0] CLBLL_L_X4Y145_SLICE_X4Y145_A1;
  wire [0:0] CLBLL_L_X4Y145_SLICE_X4Y145_A2;
  wire [0:0] CLBLL_L_X4Y145_SLICE_X4Y145_A3;
  wire [0:0] CLBLL_L_X4Y145_SLICE_X4Y145_A4;
  wire [0:0] CLBLL_L_X4Y145_SLICE_X4Y145_A5;
  wire [0:0] CLBLL_L_X4Y145_SLICE_X4Y145_A6;
  wire [0:0] CLBLL_L_X4Y145_SLICE_X4Y145_AO5;
  wire [0:0] CLBLL_L_X4Y145_SLICE_X4Y145_AO6;
  wire [0:0] CLBLL_L_X4Y145_SLICE_X4Y145_AQ;
  wire [0:0] CLBLL_L_X4Y145_SLICE_X4Y145_A_CY;
  wire [0:0] CLBLL_L_X4Y145_SLICE_X4Y145_A_XOR;
  wire [0:0] CLBLL_L_X4Y145_SLICE_X4Y145_B;
  wire [0:0] CLBLL_L_X4Y145_SLICE_X4Y145_B1;
  wire [0:0] CLBLL_L_X4Y145_SLICE_X4Y145_B2;
  wire [0:0] CLBLL_L_X4Y145_SLICE_X4Y145_B3;
  wire [0:0] CLBLL_L_X4Y145_SLICE_X4Y145_B4;
  wire [0:0] CLBLL_L_X4Y145_SLICE_X4Y145_B5;
  wire [0:0] CLBLL_L_X4Y145_SLICE_X4Y145_B5Q;
  wire [0:0] CLBLL_L_X4Y145_SLICE_X4Y145_B6;
  wire [0:0] CLBLL_L_X4Y145_SLICE_X4Y145_BMUX;
  wire [0:0] CLBLL_L_X4Y145_SLICE_X4Y145_BO5;
  wire [0:0] CLBLL_L_X4Y145_SLICE_X4Y145_BO6;
  wire [0:0] CLBLL_L_X4Y145_SLICE_X4Y145_BQ;
  wire [0:0] CLBLL_L_X4Y145_SLICE_X4Y145_B_CY;
  wire [0:0] CLBLL_L_X4Y145_SLICE_X4Y145_B_XOR;
  wire [0:0] CLBLL_L_X4Y145_SLICE_X4Y145_C;
  wire [0:0] CLBLL_L_X4Y145_SLICE_X4Y145_C1;
  wire [0:0] CLBLL_L_X4Y145_SLICE_X4Y145_C2;
  wire [0:0] CLBLL_L_X4Y145_SLICE_X4Y145_C3;
  wire [0:0] CLBLL_L_X4Y145_SLICE_X4Y145_C4;
  wire [0:0] CLBLL_L_X4Y145_SLICE_X4Y145_C5;
  wire [0:0] CLBLL_L_X4Y145_SLICE_X4Y145_C5Q;
  wire [0:0] CLBLL_L_X4Y145_SLICE_X4Y145_C6;
  wire [0:0] CLBLL_L_X4Y145_SLICE_X4Y145_CLK;
  wire [0:0] CLBLL_L_X4Y145_SLICE_X4Y145_CMUX;
  wire [0:0] CLBLL_L_X4Y145_SLICE_X4Y145_CO5;
  wire [0:0] CLBLL_L_X4Y145_SLICE_X4Y145_CO6;
  wire [0:0] CLBLL_L_X4Y145_SLICE_X4Y145_CQ;
  wire [0:0] CLBLL_L_X4Y145_SLICE_X4Y145_C_CY;
  wire [0:0] CLBLL_L_X4Y145_SLICE_X4Y145_C_XOR;
  wire [0:0] CLBLL_L_X4Y145_SLICE_X4Y145_D;
  wire [0:0] CLBLL_L_X4Y145_SLICE_X4Y145_D1;
  wire [0:0] CLBLL_L_X4Y145_SLICE_X4Y145_D2;
  wire [0:0] CLBLL_L_X4Y145_SLICE_X4Y145_D3;
  wire [0:0] CLBLL_L_X4Y145_SLICE_X4Y145_D4;
  wire [0:0] CLBLL_L_X4Y145_SLICE_X4Y145_D5;
  wire [0:0] CLBLL_L_X4Y145_SLICE_X4Y145_D6;
  wire [0:0] CLBLL_L_X4Y145_SLICE_X4Y145_DMUX;
  wire [0:0] CLBLL_L_X4Y145_SLICE_X4Y145_DO5;
  wire [0:0] CLBLL_L_X4Y145_SLICE_X4Y145_DO6;
  wire [0:0] CLBLL_L_X4Y145_SLICE_X4Y145_D_CY;
  wire [0:0] CLBLL_L_X4Y145_SLICE_X4Y145_D_XOR;
  wire [0:0] CLBLL_L_X4Y145_SLICE_X5Y145_A;
  wire [0:0] CLBLL_L_X4Y145_SLICE_X5Y145_A1;
  wire [0:0] CLBLL_L_X4Y145_SLICE_X5Y145_A2;
  wire [0:0] CLBLL_L_X4Y145_SLICE_X5Y145_A3;
  wire [0:0] CLBLL_L_X4Y145_SLICE_X5Y145_A4;
  wire [0:0] CLBLL_L_X4Y145_SLICE_X5Y145_A5;
  wire [0:0] CLBLL_L_X4Y145_SLICE_X5Y145_A6;
  wire [0:0] CLBLL_L_X4Y145_SLICE_X5Y145_AO5;
  wire [0:0] CLBLL_L_X4Y145_SLICE_X5Y145_AO6;
  wire [0:0] CLBLL_L_X4Y145_SLICE_X5Y145_AQ;
  wire [0:0] CLBLL_L_X4Y145_SLICE_X5Y145_A_CY;
  wire [0:0] CLBLL_L_X4Y145_SLICE_X5Y145_A_XOR;
  wire [0:0] CLBLL_L_X4Y145_SLICE_X5Y145_B;
  wire [0:0] CLBLL_L_X4Y145_SLICE_X5Y145_B1;
  wire [0:0] CLBLL_L_X4Y145_SLICE_X5Y145_B2;
  wire [0:0] CLBLL_L_X4Y145_SLICE_X5Y145_B3;
  wire [0:0] CLBLL_L_X4Y145_SLICE_X5Y145_B4;
  wire [0:0] CLBLL_L_X4Y145_SLICE_X5Y145_B5;
  wire [0:0] CLBLL_L_X4Y145_SLICE_X5Y145_B6;
  wire [0:0] CLBLL_L_X4Y145_SLICE_X5Y145_BO5;
  wire [0:0] CLBLL_L_X4Y145_SLICE_X5Y145_BO6;
  wire [0:0] CLBLL_L_X4Y145_SLICE_X5Y145_BQ;
  wire [0:0] CLBLL_L_X4Y145_SLICE_X5Y145_B_CY;
  wire [0:0] CLBLL_L_X4Y145_SLICE_X5Y145_B_XOR;
  wire [0:0] CLBLL_L_X4Y145_SLICE_X5Y145_C;
  wire [0:0] CLBLL_L_X4Y145_SLICE_X5Y145_C1;
  wire [0:0] CLBLL_L_X4Y145_SLICE_X5Y145_C2;
  wire [0:0] CLBLL_L_X4Y145_SLICE_X5Y145_C3;
  wire [0:0] CLBLL_L_X4Y145_SLICE_X5Y145_C4;
  wire [0:0] CLBLL_L_X4Y145_SLICE_X5Y145_C5;
  wire [0:0] CLBLL_L_X4Y145_SLICE_X5Y145_C5Q;
  wire [0:0] CLBLL_L_X4Y145_SLICE_X5Y145_C6;
  wire [0:0] CLBLL_L_X4Y145_SLICE_X5Y145_CLK;
  wire [0:0] CLBLL_L_X4Y145_SLICE_X5Y145_CMUX;
  wire [0:0] CLBLL_L_X4Y145_SLICE_X5Y145_CO5;
  wire [0:0] CLBLL_L_X4Y145_SLICE_X5Y145_CO6;
  wire [0:0] CLBLL_L_X4Y145_SLICE_X5Y145_CQ;
  wire [0:0] CLBLL_L_X4Y145_SLICE_X5Y145_C_CY;
  wire [0:0] CLBLL_L_X4Y145_SLICE_X5Y145_C_XOR;
  wire [0:0] CLBLL_L_X4Y145_SLICE_X5Y145_D;
  wire [0:0] CLBLL_L_X4Y145_SLICE_X5Y145_D1;
  wire [0:0] CLBLL_L_X4Y145_SLICE_X5Y145_D2;
  wire [0:0] CLBLL_L_X4Y145_SLICE_X5Y145_D3;
  wire [0:0] CLBLL_L_X4Y145_SLICE_X5Y145_D4;
  wire [0:0] CLBLL_L_X4Y145_SLICE_X5Y145_D5;
  wire [0:0] CLBLL_L_X4Y145_SLICE_X5Y145_D6;
  wire [0:0] CLBLL_L_X4Y145_SLICE_X5Y145_DO5;
  wire [0:0] CLBLL_L_X4Y145_SLICE_X5Y145_DO6;
  wire [0:0] CLBLL_L_X4Y145_SLICE_X5Y145_D_CY;
  wire [0:0] CLBLL_L_X4Y145_SLICE_X5Y145_D_XOR;
  wire [0:0] CLBLL_L_X4Y146_SLICE_X4Y146_A;
  wire [0:0] CLBLL_L_X4Y146_SLICE_X4Y146_A1;
  wire [0:0] CLBLL_L_X4Y146_SLICE_X4Y146_A2;
  wire [0:0] CLBLL_L_X4Y146_SLICE_X4Y146_A3;
  wire [0:0] CLBLL_L_X4Y146_SLICE_X4Y146_A4;
  wire [0:0] CLBLL_L_X4Y146_SLICE_X4Y146_A5;
  wire [0:0] CLBLL_L_X4Y146_SLICE_X4Y146_A6;
  wire [0:0] CLBLL_L_X4Y146_SLICE_X4Y146_AO5;
  wire [0:0] CLBLL_L_X4Y146_SLICE_X4Y146_AO6;
  wire [0:0] CLBLL_L_X4Y146_SLICE_X4Y146_AQ;
  wire [0:0] CLBLL_L_X4Y146_SLICE_X4Y146_A_CY;
  wire [0:0] CLBLL_L_X4Y146_SLICE_X4Y146_A_XOR;
  wire [0:0] CLBLL_L_X4Y146_SLICE_X4Y146_B;
  wire [0:0] CLBLL_L_X4Y146_SLICE_X4Y146_B1;
  wire [0:0] CLBLL_L_X4Y146_SLICE_X4Y146_B2;
  wire [0:0] CLBLL_L_X4Y146_SLICE_X4Y146_B3;
  wire [0:0] CLBLL_L_X4Y146_SLICE_X4Y146_B4;
  wire [0:0] CLBLL_L_X4Y146_SLICE_X4Y146_B5;
  wire [0:0] CLBLL_L_X4Y146_SLICE_X4Y146_B5Q;
  wire [0:0] CLBLL_L_X4Y146_SLICE_X4Y146_B6;
  wire [0:0] CLBLL_L_X4Y146_SLICE_X4Y146_BMUX;
  wire [0:0] CLBLL_L_X4Y146_SLICE_X4Y146_BO5;
  wire [0:0] CLBLL_L_X4Y146_SLICE_X4Y146_BO6;
  wire [0:0] CLBLL_L_X4Y146_SLICE_X4Y146_BQ;
  wire [0:0] CLBLL_L_X4Y146_SLICE_X4Y146_B_CY;
  wire [0:0] CLBLL_L_X4Y146_SLICE_X4Y146_B_XOR;
  wire [0:0] CLBLL_L_X4Y146_SLICE_X4Y146_C;
  wire [0:0] CLBLL_L_X4Y146_SLICE_X4Y146_C1;
  wire [0:0] CLBLL_L_X4Y146_SLICE_X4Y146_C2;
  wire [0:0] CLBLL_L_X4Y146_SLICE_X4Y146_C3;
  wire [0:0] CLBLL_L_X4Y146_SLICE_X4Y146_C4;
  wire [0:0] CLBLL_L_X4Y146_SLICE_X4Y146_C5;
  wire [0:0] CLBLL_L_X4Y146_SLICE_X4Y146_C5Q;
  wire [0:0] CLBLL_L_X4Y146_SLICE_X4Y146_C6;
  wire [0:0] CLBLL_L_X4Y146_SLICE_X4Y146_CLK;
  wire [0:0] CLBLL_L_X4Y146_SLICE_X4Y146_CMUX;
  wire [0:0] CLBLL_L_X4Y146_SLICE_X4Y146_CO5;
  wire [0:0] CLBLL_L_X4Y146_SLICE_X4Y146_CO6;
  wire [0:0] CLBLL_L_X4Y146_SLICE_X4Y146_CQ;
  wire [0:0] CLBLL_L_X4Y146_SLICE_X4Y146_C_CY;
  wire [0:0] CLBLL_L_X4Y146_SLICE_X4Y146_C_XOR;
  wire [0:0] CLBLL_L_X4Y146_SLICE_X4Y146_D;
  wire [0:0] CLBLL_L_X4Y146_SLICE_X4Y146_D1;
  wire [0:0] CLBLL_L_X4Y146_SLICE_X4Y146_D2;
  wire [0:0] CLBLL_L_X4Y146_SLICE_X4Y146_D3;
  wire [0:0] CLBLL_L_X4Y146_SLICE_X4Y146_D4;
  wire [0:0] CLBLL_L_X4Y146_SLICE_X4Y146_D5;
  wire [0:0] CLBLL_L_X4Y146_SLICE_X4Y146_D6;
  wire [0:0] CLBLL_L_X4Y146_SLICE_X4Y146_DMUX;
  wire [0:0] CLBLL_L_X4Y146_SLICE_X4Y146_DO5;
  wire [0:0] CLBLL_L_X4Y146_SLICE_X4Y146_DO6;
  wire [0:0] CLBLL_L_X4Y146_SLICE_X4Y146_D_CY;
  wire [0:0] CLBLL_L_X4Y146_SLICE_X4Y146_D_XOR;
  wire [0:0] CLBLL_L_X4Y146_SLICE_X5Y146_A;
  wire [0:0] CLBLL_L_X4Y146_SLICE_X5Y146_A1;
  wire [0:0] CLBLL_L_X4Y146_SLICE_X5Y146_A2;
  wire [0:0] CLBLL_L_X4Y146_SLICE_X5Y146_A3;
  wire [0:0] CLBLL_L_X4Y146_SLICE_X5Y146_A4;
  wire [0:0] CLBLL_L_X4Y146_SLICE_X5Y146_A5;
  wire [0:0] CLBLL_L_X4Y146_SLICE_X5Y146_A6;
  wire [0:0] CLBLL_L_X4Y146_SLICE_X5Y146_AMUX;
  wire [0:0] CLBLL_L_X4Y146_SLICE_X5Y146_AO5;
  wire [0:0] CLBLL_L_X4Y146_SLICE_X5Y146_AO6;
  wire [0:0] CLBLL_L_X4Y146_SLICE_X5Y146_AQ;
  wire [0:0] CLBLL_L_X4Y146_SLICE_X5Y146_A_CY;
  wire [0:0] CLBLL_L_X4Y146_SLICE_X5Y146_A_XOR;
  wire [0:0] CLBLL_L_X4Y146_SLICE_X5Y146_B;
  wire [0:0] CLBLL_L_X4Y146_SLICE_X5Y146_B1;
  wire [0:0] CLBLL_L_X4Y146_SLICE_X5Y146_B2;
  wire [0:0] CLBLL_L_X4Y146_SLICE_X5Y146_B3;
  wire [0:0] CLBLL_L_X4Y146_SLICE_X5Y146_B4;
  wire [0:0] CLBLL_L_X4Y146_SLICE_X5Y146_B5;
  wire [0:0] CLBLL_L_X4Y146_SLICE_X5Y146_B6;
  wire [0:0] CLBLL_L_X4Y146_SLICE_X5Y146_BO5;
  wire [0:0] CLBLL_L_X4Y146_SLICE_X5Y146_BO6;
  wire [0:0] CLBLL_L_X4Y146_SLICE_X5Y146_BQ;
  wire [0:0] CLBLL_L_X4Y146_SLICE_X5Y146_B_CY;
  wire [0:0] CLBLL_L_X4Y146_SLICE_X5Y146_B_XOR;
  wire [0:0] CLBLL_L_X4Y146_SLICE_X5Y146_C;
  wire [0:0] CLBLL_L_X4Y146_SLICE_X5Y146_C1;
  wire [0:0] CLBLL_L_X4Y146_SLICE_X5Y146_C2;
  wire [0:0] CLBLL_L_X4Y146_SLICE_X5Y146_C3;
  wire [0:0] CLBLL_L_X4Y146_SLICE_X5Y146_C4;
  wire [0:0] CLBLL_L_X4Y146_SLICE_X5Y146_C5;
  wire [0:0] CLBLL_L_X4Y146_SLICE_X5Y146_C6;
  wire [0:0] CLBLL_L_X4Y146_SLICE_X5Y146_CLK;
  wire [0:0] CLBLL_L_X4Y146_SLICE_X5Y146_CO5;
  wire [0:0] CLBLL_L_X4Y146_SLICE_X5Y146_CO6;
  wire [0:0] CLBLL_L_X4Y146_SLICE_X5Y146_CQ;
  wire [0:0] CLBLL_L_X4Y146_SLICE_X5Y146_C_CY;
  wire [0:0] CLBLL_L_X4Y146_SLICE_X5Y146_C_XOR;
  wire [0:0] CLBLL_L_X4Y146_SLICE_X5Y146_D;
  wire [0:0] CLBLL_L_X4Y146_SLICE_X5Y146_D1;
  wire [0:0] CLBLL_L_X4Y146_SLICE_X5Y146_D2;
  wire [0:0] CLBLL_L_X4Y146_SLICE_X5Y146_D3;
  wire [0:0] CLBLL_L_X4Y146_SLICE_X5Y146_D4;
  wire [0:0] CLBLL_L_X4Y146_SLICE_X5Y146_D5;
  wire [0:0] CLBLL_L_X4Y146_SLICE_X5Y146_D6;
  wire [0:0] CLBLL_L_X4Y146_SLICE_X5Y146_DO5;
  wire [0:0] CLBLL_L_X4Y146_SLICE_X5Y146_DO6;
  wire [0:0] CLBLL_L_X4Y146_SLICE_X5Y146_DQ;
  wire [0:0] CLBLL_L_X4Y146_SLICE_X5Y146_D_CY;
  wire [0:0] CLBLL_L_X4Y146_SLICE_X5Y146_D_XOR;
  wire [0:0] CLBLL_L_X4Y147_SLICE_X4Y147_A;
  wire [0:0] CLBLL_L_X4Y147_SLICE_X4Y147_A1;
  wire [0:0] CLBLL_L_X4Y147_SLICE_X4Y147_A2;
  wire [0:0] CLBLL_L_X4Y147_SLICE_X4Y147_A3;
  wire [0:0] CLBLL_L_X4Y147_SLICE_X4Y147_A4;
  wire [0:0] CLBLL_L_X4Y147_SLICE_X4Y147_A5;
  wire [0:0] CLBLL_L_X4Y147_SLICE_X4Y147_A6;
  wire [0:0] CLBLL_L_X4Y147_SLICE_X4Y147_AO5;
  wire [0:0] CLBLL_L_X4Y147_SLICE_X4Y147_AO6;
  wire [0:0] CLBLL_L_X4Y147_SLICE_X4Y147_AQ;
  wire [0:0] CLBLL_L_X4Y147_SLICE_X4Y147_A_CY;
  wire [0:0] CLBLL_L_X4Y147_SLICE_X4Y147_A_XOR;
  wire [0:0] CLBLL_L_X4Y147_SLICE_X4Y147_B;
  wire [0:0] CLBLL_L_X4Y147_SLICE_X4Y147_B1;
  wire [0:0] CLBLL_L_X4Y147_SLICE_X4Y147_B2;
  wire [0:0] CLBLL_L_X4Y147_SLICE_X4Y147_B3;
  wire [0:0] CLBLL_L_X4Y147_SLICE_X4Y147_B4;
  wire [0:0] CLBLL_L_X4Y147_SLICE_X4Y147_B5;
  wire [0:0] CLBLL_L_X4Y147_SLICE_X4Y147_B5Q;
  wire [0:0] CLBLL_L_X4Y147_SLICE_X4Y147_B6;
  wire [0:0] CLBLL_L_X4Y147_SLICE_X4Y147_BMUX;
  wire [0:0] CLBLL_L_X4Y147_SLICE_X4Y147_BO5;
  wire [0:0] CLBLL_L_X4Y147_SLICE_X4Y147_BO6;
  wire [0:0] CLBLL_L_X4Y147_SLICE_X4Y147_BQ;
  wire [0:0] CLBLL_L_X4Y147_SLICE_X4Y147_B_CY;
  wire [0:0] CLBLL_L_X4Y147_SLICE_X4Y147_B_XOR;
  wire [0:0] CLBLL_L_X4Y147_SLICE_X4Y147_C;
  wire [0:0] CLBLL_L_X4Y147_SLICE_X4Y147_C1;
  wire [0:0] CLBLL_L_X4Y147_SLICE_X4Y147_C2;
  wire [0:0] CLBLL_L_X4Y147_SLICE_X4Y147_C3;
  wire [0:0] CLBLL_L_X4Y147_SLICE_X4Y147_C4;
  wire [0:0] CLBLL_L_X4Y147_SLICE_X4Y147_C5;
  wire [0:0] CLBLL_L_X4Y147_SLICE_X4Y147_C5Q;
  wire [0:0] CLBLL_L_X4Y147_SLICE_X4Y147_C6;
  wire [0:0] CLBLL_L_X4Y147_SLICE_X4Y147_CLK;
  wire [0:0] CLBLL_L_X4Y147_SLICE_X4Y147_CMUX;
  wire [0:0] CLBLL_L_X4Y147_SLICE_X4Y147_CO5;
  wire [0:0] CLBLL_L_X4Y147_SLICE_X4Y147_CO6;
  wire [0:0] CLBLL_L_X4Y147_SLICE_X4Y147_CQ;
  wire [0:0] CLBLL_L_X4Y147_SLICE_X4Y147_C_CY;
  wire [0:0] CLBLL_L_X4Y147_SLICE_X4Y147_C_XOR;
  wire [0:0] CLBLL_L_X4Y147_SLICE_X4Y147_D;
  wire [0:0] CLBLL_L_X4Y147_SLICE_X4Y147_D1;
  wire [0:0] CLBLL_L_X4Y147_SLICE_X4Y147_D2;
  wire [0:0] CLBLL_L_X4Y147_SLICE_X4Y147_D3;
  wire [0:0] CLBLL_L_X4Y147_SLICE_X4Y147_D4;
  wire [0:0] CLBLL_L_X4Y147_SLICE_X4Y147_D5;
  wire [0:0] CLBLL_L_X4Y147_SLICE_X4Y147_D5Q;
  wire [0:0] CLBLL_L_X4Y147_SLICE_X4Y147_D6;
  wire [0:0] CLBLL_L_X4Y147_SLICE_X4Y147_DMUX;
  wire [0:0] CLBLL_L_X4Y147_SLICE_X4Y147_DO5;
  wire [0:0] CLBLL_L_X4Y147_SLICE_X4Y147_DO6;
  wire [0:0] CLBLL_L_X4Y147_SLICE_X4Y147_DQ;
  wire [0:0] CLBLL_L_X4Y147_SLICE_X4Y147_D_CY;
  wire [0:0] CLBLL_L_X4Y147_SLICE_X4Y147_D_XOR;
  wire [0:0] CLBLL_L_X4Y147_SLICE_X5Y147_A;
  wire [0:0] CLBLL_L_X4Y147_SLICE_X5Y147_A1;
  wire [0:0] CLBLL_L_X4Y147_SLICE_X5Y147_A2;
  wire [0:0] CLBLL_L_X4Y147_SLICE_X5Y147_A3;
  wire [0:0] CLBLL_L_X4Y147_SLICE_X5Y147_A4;
  wire [0:0] CLBLL_L_X4Y147_SLICE_X5Y147_A5;
  wire [0:0] CLBLL_L_X4Y147_SLICE_X5Y147_A6;
  wire [0:0] CLBLL_L_X4Y147_SLICE_X5Y147_AO5;
  wire [0:0] CLBLL_L_X4Y147_SLICE_X5Y147_AO6;
  wire [0:0] CLBLL_L_X4Y147_SLICE_X5Y147_AQ;
  wire [0:0] CLBLL_L_X4Y147_SLICE_X5Y147_A_CY;
  wire [0:0] CLBLL_L_X4Y147_SLICE_X5Y147_A_XOR;
  wire [0:0] CLBLL_L_X4Y147_SLICE_X5Y147_B;
  wire [0:0] CLBLL_L_X4Y147_SLICE_X5Y147_B1;
  wire [0:0] CLBLL_L_X4Y147_SLICE_X5Y147_B2;
  wire [0:0] CLBLL_L_X4Y147_SLICE_X5Y147_B3;
  wire [0:0] CLBLL_L_X4Y147_SLICE_X5Y147_B4;
  wire [0:0] CLBLL_L_X4Y147_SLICE_X5Y147_B5;
  wire [0:0] CLBLL_L_X4Y147_SLICE_X5Y147_B5Q;
  wire [0:0] CLBLL_L_X4Y147_SLICE_X5Y147_B6;
  wire [0:0] CLBLL_L_X4Y147_SLICE_X5Y147_BMUX;
  wire [0:0] CLBLL_L_X4Y147_SLICE_X5Y147_BO5;
  wire [0:0] CLBLL_L_X4Y147_SLICE_X5Y147_BO6;
  wire [0:0] CLBLL_L_X4Y147_SLICE_X5Y147_BQ;
  wire [0:0] CLBLL_L_X4Y147_SLICE_X5Y147_B_CY;
  wire [0:0] CLBLL_L_X4Y147_SLICE_X5Y147_B_XOR;
  wire [0:0] CLBLL_L_X4Y147_SLICE_X5Y147_C;
  wire [0:0] CLBLL_L_X4Y147_SLICE_X5Y147_C1;
  wire [0:0] CLBLL_L_X4Y147_SLICE_X5Y147_C2;
  wire [0:0] CLBLL_L_X4Y147_SLICE_X5Y147_C3;
  wire [0:0] CLBLL_L_X4Y147_SLICE_X5Y147_C4;
  wire [0:0] CLBLL_L_X4Y147_SLICE_X5Y147_C5;
  wire [0:0] CLBLL_L_X4Y147_SLICE_X5Y147_C5Q;
  wire [0:0] CLBLL_L_X4Y147_SLICE_X5Y147_C6;
  wire [0:0] CLBLL_L_X4Y147_SLICE_X5Y147_CLK;
  wire [0:0] CLBLL_L_X4Y147_SLICE_X5Y147_CMUX;
  wire [0:0] CLBLL_L_X4Y147_SLICE_X5Y147_CO5;
  wire [0:0] CLBLL_L_X4Y147_SLICE_X5Y147_CO6;
  wire [0:0] CLBLL_L_X4Y147_SLICE_X5Y147_CQ;
  wire [0:0] CLBLL_L_X4Y147_SLICE_X5Y147_C_CY;
  wire [0:0] CLBLL_L_X4Y147_SLICE_X5Y147_C_XOR;
  wire [0:0] CLBLL_L_X4Y147_SLICE_X5Y147_D;
  wire [0:0] CLBLL_L_X4Y147_SLICE_X5Y147_D1;
  wire [0:0] CLBLL_L_X4Y147_SLICE_X5Y147_D2;
  wire [0:0] CLBLL_L_X4Y147_SLICE_X5Y147_D3;
  wire [0:0] CLBLL_L_X4Y147_SLICE_X5Y147_D4;
  wire [0:0] CLBLL_L_X4Y147_SLICE_X5Y147_D5;
  wire [0:0] CLBLL_L_X4Y147_SLICE_X5Y147_D6;
  wire [0:0] CLBLL_L_X4Y147_SLICE_X5Y147_DMUX;
  wire [0:0] CLBLL_L_X4Y147_SLICE_X5Y147_DO5;
  wire [0:0] CLBLL_L_X4Y147_SLICE_X5Y147_DO6;
  wire [0:0] CLBLL_L_X4Y147_SLICE_X5Y147_D_CY;
  wire [0:0] CLBLL_L_X4Y147_SLICE_X5Y147_D_XOR;
  wire [0:0] CLBLL_L_X4Y148_SLICE_X4Y148_A;
  wire [0:0] CLBLL_L_X4Y148_SLICE_X4Y148_A1;
  wire [0:0] CLBLL_L_X4Y148_SLICE_X4Y148_A2;
  wire [0:0] CLBLL_L_X4Y148_SLICE_X4Y148_A3;
  wire [0:0] CLBLL_L_X4Y148_SLICE_X4Y148_A4;
  wire [0:0] CLBLL_L_X4Y148_SLICE_X4Y148_A5;
  wire [0:0] CLBLL_L_X4Y148_SLICE_X4Y148_A6;
  wire [0:0] CLBLL_L_X4Y148_SLICE_X4Y148_AO5;
  wire [0:0] CLBLL_L_X4Y148_SLICE_X4Y148_AO6;
  wire [0:0] CLBLL_L_X4Y148_SLICE_X4Y148_AQ;
  wire [0:0] CLBLL_L_X4Y148_SLICE_X4Y148_A_CY;
  wire [0:0] CLBLL_L_X4Y148_SLICE_X4Y148_A_XOR;
  wire [0:0] CLBLL_L_X4Y148_SLICE_X4Y148_B;
  wire [0:0] CLBLL_L_X4Y148_SLICE_X4Y148_B1;
  wire [0:0] CLBLL_L_X4Y148_SLICE_X4Y148_B2;
  wire [0:0] CLBLL_L_X4Y148_SLICE_X4Y148_B3;
  wire [0:0] CLBLL_L_X4Y148_SLICE_X4Y148_B4;
  wire [0:0] CLBLL_L_X4Y148_SLICE_X4Y148_B5;
  wire [0:0] CLBLL_L_X4Y148_SLICE_X4Y148_B6;
  wire [0:0] CLBLL_L_X4Y148_SLICE_X4Y148_BO5;
  wire [0:0] CLBLL_L_X4Y148_SLICE_X4Y148_BO6;
  wire [0:0] CLBLL_L_X4Y148_SLICE_X4Y148_BQ;
  wire [0:0] CLBLL_L_X4Y148_SLICE_X4Y148_B_CY;
  wire [0:0] CLBLL_L_X4Y148_SLICE_X4Y148_B_XOR;
  wire [0:0] CLBLL_L_X4Y148_SLICE_X4Y148_C;
  wire [0:0] CLBLL_L_X4Y148_SLICE_X4Y148_C1;
  wire [0:0] CLBLL_L_X4Y148_SLICE_X4Y148_C2;
  wire [0:0] CLBLL_L_X4Y148_SLICE_X4Y148_C3;
  wire [0:0] CLBLL_L_X4Y148_SLICE_X4Y148_C4;
  wire [0:0] CLBLL_L_X4Y148_SLICE_X4Y148_C5;
  wire [0:0] CLBLL_L_X4Y148_SLICE_X4Y148_C5Q;
  wire [0:0] CLBLL_L_X4Y148_SLICE_X4Y148_C6;
  wire [0:0] CLBLL_L_X4Y148_SLICE_X4Y148_CLK;
  wire [0:0] CLBLL_L_X4Y148_SLICE_X4Y148_CMUX;
  wire [0:0] CLBLL_L_X4Y148_SLICE_X4Y148_CO5;
  wire [0:0] CLBLL_L_X4Y148_SLICE_X4Y148_CO6;
  wire [0:0] CLBLL_L_X4Y148_SLICE_X4Y148_CQ;
  wire [0:0] CLBLL_L_X4Y148_SLICE_X4Y148_C_CY;
  wire [0:0] CLBLL_L_X4Y148_SLICE_X4Y148_C_XOR;
  wire [0:0] CLBLL_L_X4Y148_SLICE_X4Y148_D;
  wire [0:0] CLBLL_L_X4Y148_SLICE_X4Y148_D1;
  wire [0:0] CLBLL_L_X4Y148_SLICE_X4Y148_D2;
  wire [0:0] CLBLL_L_X4Y148_SLICE_X4Y148_D3;
  wire [0:0] CLBLL_L_X4Y148_SLICE_X4Y148_D4;
  wire [0:0] CLBLL_L_X4Y148_SLICE_X4Y148_D5;
  wire [0:0] CLBLL_L_X4Y148_SLICE_X4Y148_D6;
  wire [0:0] CLBLL_L_X4Y148_SLICE_X4Y148_DO5;
  wire [0:0] CLBLL_L_X4Y148_SLICE_X4Y148_DO6;
  wire [0:0] CLBLL_L_X4Y148_SLICE_X4Y148_D_CY;
  wire [0:0] CLBLL_L_X4Y148_SLICE_X4Y148_D_XOR;
  wire [0:0] CLBLL_L_X4Y148_SLICE_X5Y148_A;
  wire [0:0] CLBLL_L_X4Y148_SLICE_X5Y148_A1;
  wire [0:0] CLBLL_L_X4Y148_SLICE_X5Y148_A2;
  wire [0:0] CLBLL_L_X4Y148_SLICE_X5Y148_A3;
  wire [0:0] CLBLL_L_X4Y148_SLICE_X5Y148_A4;
  wire [0:0] CLBLL_L_X4Y148_SLICE_X5Y148_A5;
  wire [0:0] CLBLL_L_X4Y148_SLICE_X5Y148_A5Q;
  wire [0:0] CLBLL_L_X4Y148_SLICE_X5Y148_A6;
  wire [0:0] CLBLL_L_X4Y148_SLICE_X5Y148_AMUX;
  wire [0:0] CLBLL_L_X4Y148_SLICE_X5Y148_AO5;
  wire [0:0] CLBLL_L_X4Y148_SLICE_X5Y148_AO6;
  wire [0:0] CLBLL_L_X4Y148_SLICE_X5Y148_AQ;
  wire [0:0] CLBLL_L_X4Y148_SLICE_X5Y148_A_CY;
  wire [0:0] CLBLL_L_X4Y148_SLICE_X5Y148_A_XOR;
  wire [0:0] CLBLL_L_X4Y148_SLICE_X5Y148_B;
  wire [0:0] CLBLL_L_X4Y148_SLICE_X5Y148_B1;
  wire [0:0] CLBLL_L_X4Y148_SLICE_X5Y148_B2;
  wire [0:0] CLBLL_L_X4Y148_SLICE_X5Y148_B3;
  wire [0:0] CLBLL_L_X4Y148_SLICE_X5Y148_B4;
  wire [0:0] CLBLL_L_X4Y148_SLICE_X5Y148_B5;
  wire [0:0] CLBLL_L_X4Y148_SLICE_X5Y148_B5Q;
  wire [0:0] CLBLL_L_X4Y148_SLICE_X5Y148_B6;
  wire [0:0] CLBLL_L_X4Y148_SLICE_X5Y148_BMUX;
  wire [0:0] CLBLL_L_X4Y148_SLICE_X5Y148_BO5;
  wire [0:0] CLBLL_L_X4Y148_SLICE_X5Y148_BO6;
  wire [0:0] CLBLL_L_X4Y148_SLICE_X5Y148_BQ;
  wire [0:0] CLBLL_L_X4Y148_SLICE_X5Y148_B_CY;
  wire [0:0] CLBLL_L_X4Y148_SLICE_X5Y148_B_XOR;
  wire [0:0] CLBLL_L_X4Y148_SLICE_X5Y148_C;
  wire [0:0] CLBLL_L_X4Y148_SLICE_X5Y148_C1;
  wire [0:0] CLBLL_L_X4Y148_SLICE_X5Y148_C2;
  wire [0:0] CLBLL_L_X4Y148_SLICE_X5Y148_C3;
  wire [0:0] CLBLL_L_X4Y148_SLICE_X5Y148_C4;
  wire [0:0] CLBLL_L_X4Y148_SLICE_X5Y148_C5;
  wire [0:0] CLBLL_L_X4Y148_SLICE_X5Y148_C6;
  wire [0:0] CLBLL_L_X4Y148_SLICE_X5Y148_CLK;
  wire [0:0] CLBLL_L_X4Y148_SLICE_X5Y148_CO5;
  wire [0:0] CLBLL_L_X4Y148_SLICE_X5Y148_CO6;
  wire [0:0] CLBLL_L_X4Y148_SLICE_X5Y148_CQ;
  wire [0:0] CLBLL_L_X4Y148_SLICE_X5Y148_C_CY;
  wire [0:0] CLBLL_L_X4Y148_SLICE_X5Y148_C_XOR;
  wire [0:0] CLBLL_L_X4Y148_SLICE_X5Y148_D;
  wire [0:0] CLBLL_L_X4Y148_SLICE_X5Y148_D1;
  wire [0:0] CLBLL_L_X4Y148_SLICE_X5Y148_D2;
  wire [0:0] CLBLL_L_X4Y148_SLICE_X5Y148_D3;
  wire [0:0] CLBLL_L_X4Y148_SLICE_X5Y148_D4;
  wire [0:0] CLBLL_L_X4Y148_SLICE_X5Y148_D5;
  wire [0:0] CLBLL_L_X4Y148_SLICE_X5Y148_D5Q;
  wire [0:0] CLBLL_L_X4Y148_SLICE_X5Y148_D6;
  wire [0:0] CLBLL_L_X4Y148_SLICE_X5Y148_DMUX;
  wire [0:0] CLBLL_L_X4Y148_SLICE_X5Y148_DO5;
  wire [0:0] CLBLL_L_X4Y148_SLICE_X5Y148_DO6;
  wire [0:0] CLBLL_L_X4Y148_SLICE_X5Y148_DQ;
  wire [0:0] CLBLL_L_X4Y148_SLICE_X5Y148_D_CY;
  wire [0:0] CLBLL_L_X4Y148_SLICE_X5Y148_D_XOR;
  wire [0:0] CLBLL_L_X4Y149_SLICE_X4Y149_A;
  wire [0:0] CLBLL_L_X4Y149_SLICE_X4Y149_A1;
  wire [0:0] CLBLL_L_X4Y149_SLICE_X4Y149_A2;
  wire [0:0] CLBLL_L_X4Y149_SLICE_X4Y149_A3;
  wire [0:0] CLBLL_L_X4Y149_SLICE_X4Y149_A4;
  wire [0:0] CLBLL_L_X4Y149_SLICE_X4Y149_A5;
  wire [0:0] CLBLL_L_X4Y149_SLICE_X4Y149_A6;
  wire [0:0] CLBLL_L_X4Y149_SLICE_X4Y149_AO5;
  wire [0:0] CLBLL_L_X4Y149_SLICE_X4Y149_AO6;
  wire [0:0] CLBLL_L_X4Y149_SLICE_X4Y149_AQ;
  wire [0:0] CLBLL_L_X4Y149_SLICE_X4Y149_A_CY;
  wire [0:0] CLBLL_L_X4Y149_SLICE_X4Y149_A_XOR;
  wire [0:0] CLBLL_L_X4Y149_SLICE_X4Y149_B;
  wire [0:0] CLBLL_L_X4Y149_SLICE_X4Y149_B1;
  wire [0:0] CLBLL_L_X4Y149_SLICE_X4Y149_B2;
  wire [0:0] CLBLL_L_X4Y149_SLICE_X4Y149_B3;
  wire [0:0] CLBLL_L_X4Y149_SLICE_X4Y149_B4;
  wire [0:0] CLBLL_L_X4Y149_SLICE_X4Y149_B5;
  wire [0:0] CLBLL_L_X4Y149_SLICE_X4Y149_B5Q;
  wire [0:0] CLBLL_L_X4Y149_SLICE_X4Y149_B6;
  wire [0:0] CLBLL_L_X4Y149_SLICE_X4Y149_BMUX;
  wire [0:0] CLBLL_L_X4Y149_SLICE_X4Y149_BO5;
  wire [0:0] CLBLL_L_X4Y149_SLICE_X4Y149_BO6;
  wire [0:0] CLBLL_L_X4Y149_SLICE_X4Y149_BQ;
  wire [0:0] CLBLL_L_X4Y149_SLICE_X4Y149_B_CY;
  wire [0:0] CLBLL_L_X4Y149_SLICE_X4Y149_B_XOR;
  wire [0:0] CLBLL_L_X4Y149_SLICE_X4Y149_C;
  wire [0:0] CLBLL_L_X4Y149_SLICE_X4Y149_C1;
  wire [0:0] CLBLL_L_X4Y149_SLICE_X4Y149_C2;
  wire [0:0] CLBLL_L_X4Y149_SLICE_X4Y149_C3;
  wire [0:0] CLBLL_L_X4Y149_SLICE_X4Y149_C4;
  wire [0:0] CLBLL_L_X4Y149_SLICE_X4Y149_C5;
  wire [0:0] CLBLL_L_X4Y149_SLICE_X4Y149_C6;
  wire [0:0] CLBLL_L_X4Y149_SLICE_X4Y149_CLK;
  wire [0:0] CLBLL_L_X4Y149_SLICE_X4Y149_CO5;
  wire [0:0] CLBLL_L_X4Y149_SLICE_X4Y149_CO6;
  wire [0:0] CLBLL_L_X4Y149_SLICE_X4Y149_CQ;
  wire [0:0] CLBLL_L_X4Y149_SLICE_X4Y149_C_CY;
  wire [0:0] CLBLL_L_X4Y149_SLICE_X4Y149_C_XOR;
  wire [0:0] CLBLL_L_X4Y149_SLICE_X4Y149_D;
  wire [0:0] CLBLL_L_X4Y149_SLICE_X4Y149_D1;
  wire [0:0] CLBLL_L_X4Y149_SLICE_X4Y149_D2;
  wire [0:0] CLBLL_L_X4Y149_SLICE_X4Y149_D3;
  wire [0:0] CLBLL_L_X4Y149_SLICE_X4Y149_D4;
  wire [0:0] CLBLL_L_X4Y149_SLICE_X4Y149_D5;
  wire [0:0] CLBLL_L_X4Y149_SLICE_X4Y149_D5Q;
  wire [0:0] CLBLL_L_X4Y149_SLICE_X4Y149_D6;
  wire [0:0] CLBLL_L_X4Y149_SLICE_X4Y149_DMUX;
  wire [0:0] CLBLL_L_X4Y149_SLICE_X4Y149_DO5;
  wire [0:0] CLBLL_L_X4Y149_SLICE_X4Y149_DO6;
  wire [0:0] CLBLL_L_X4Y149_SLICE_X4Y149_DQ;
  wire [0:0] CLBLL_L_X4Y149_SLICE_X4Y149_D_CY;
  wire [0:0] CLBLL_L_X4Y149_SLICE_X4Y149_D_XOR;
  wire [0:0] CLBLL_L_X4Y149_SLICE_X5Y149_A;
  wire [0:0] CLBLL_L_X4Y149_SLICE_X5Y149_A1;
  wire [0:0] CLBLL_L_X4Y149_SLICE_X5Y149_A2;
  wire [0:0] CLBLL_L_X4Y149_SLICE_X5Y149_A3;
  wire [0:0] CLBLL_L_X4Y149_SLICE_X5Y149_A4;
  wire [0:0] CLBLL_L_X4Y149_SLICE_X5Y149_A5;
  wire [0:0] CLBLL_L_X4Y149_SLICE_X5Y149_A6;
  wire [0:0] CLBLL_L_X4Y149_SLICE_X5Y149_AO5;
  wire [0:0] CLBLL_L_X4Y149_SLICE_X5Y149_AO6;
  wire [0:0] CLBLL_L_X4Y149_SLICE_X5Y149_AQ;
  wire [0:0] CLBLL_L_X4Y149_SLICE_X5Y149_A_CY;
  wire [0:0] CLBLL_L_X4Y149_SLICE_X5Y149_A_XOR;
  wire [0:0] CLBLL_L_X4Y149_SLICE_X5Y149_B;
  wire [0:0] CLBLL_L_X4Y149_SLICE_X5Y149_B1;
  wire [0:0] CLBLL_L_X4Y149_SLICE_X5Y149_B2;
  wire [0:0] CLBLL_L_X4Y149_SLICE_X5Y149_B3;
  wire [0:0] CLBLL_L_X4Y149_SLICE_X5Y149_B4;
  wire [0:0] CLBLL_L_X4Y149_SLICE_X5Y149_B5;
  wire [0:0] CLBLL_L_X4Y149_SLICE_X5Y149_B6;
  wire [0:0] CLBLL_L_X4Y149_SLICE_X5Y149_BO5;
  wire [0:0] CLBLL_L_X4Y149_SLICE_X5Y149_BO6;
  wire [0:0] CLBLL_L_X4Y149_SLICE_X5Y149_BQ;
  wire [0:0] CLBLL_L_X4Y149_SLICE_X5Y149_B_CY;
  wire [0:0] CLBLL_L_X4Y149_SLICE_X5Y149_B_XOR;
  wire [0:0] CLBLL_L_X4Y149_SLICE_X5Y149_C;
  wire [0:0] CLBLL_L_X4Y149_SLICE_X5Y149_C1;
  wire [0:0] CLBLL_L_X4Y149_SLICE_X5Y149_C2;
  wire [0:0] CLBLL_L_X4Y149_SLICE_X5Y149_C3;
  wire [0:0] CLBLL_L_X4Y149_SLICE_X5Y149_C4;
  wire [0:0] CLBLL_L_X4Y149_SLICE_X5Y149_C5;
  wire [0:0] CLBLL_L_X4Y149_SLICE_X5Y149_C5Q;
  wire [0:0] CLBLL_L_X4Y149_SLICE_X5Y149_C6;
  wire [0:0] CLBLL_L_X4Y149_SLICE_X5Y149_CLK;
  wire [0:0] CLBLL_L_X4Y149_SLICE_X5Y149_CMUX;
  wire [0:0] CLBLL_L_X4Y149_SLICE_X5Y149_CO5;
  wire [0:0] CLBLL_L_X4Y149_SLICE_X5Y149_CO6;
  wire [0:0] CLBLL_L_X4Y149_SLICE_X5Y149_CQ;
  wire [0:0] CLBLL_L_X4Y149_SLICE_X5Y149_C_CY;
  wire [0:0] CLBLL_L_X4Y149_SLICE_X5Y149_C_XOR;
  wire [0:0] CLBLL_L_X4Y149_SLICE_X5Y149_D;
  wire [0:0] CLBLL_L_X4Y149_SLICE_X5Y149_D1;
  wire [0:0] CLBLL_L_X4Y149_SLICE_X5Y149_D2;
  wire [0:0] CLBLL_L_X4Y149_SLICE_X5Y149_D3;
  wire [0:0] CLBLL_L_X4Y149_SLICE_X5Y149_D4;
  wire [0:0] CLBLL_L_X4Y149_SLICE_X5Y149_D5;
  wire [0:0] CLBLL_L_X4Y149_SLICE_X5Y149_D6;
  wire [0:0] CLBLL_L_X4Y149_SLICE_X5Y149_DO5;
  wire [0:0] CLBLL_L_X4Y149_SLICE_X5Y149_DO6;
  wire [0:0] CLBLL_L_X4Y149_SLICE_X5Y149_DQ;
  wire [0:0] CLBLL_L_X4Y149_SLICE_X5Y149_D_CY;
  wire [0:0] CLBLL_L_X4Y149_SLICE_X5Y149_D_XOR;
  wire [0:0] CLBLL_L_X4Y150_SLICE_X4Y150_A;
  wire [0:0] CLBLL_L_X4Y150_SLICE_X4Y150_A1;
  wire [0:0] CLBLL_L_X4Y150_SLICE_X4Y150_A2;
  wire [0:0] CLBLL_L_X4Y150_SLICE_X4Y150_A3;
  wire [0:0] CLBLL_L_X4Y150_SLICE_X4Y150_A4;
  wire [0:0] CLBLL_L_X4Y150_SLICE_X4Y150_A5;
  wire [0:0] CLBLL_L_X4Y150_SLICE_X4Y150_A5Q;
  wire [0:0] CLBLL_L_X4Y150_SLICE_X4Y150_A6;
  wire [0:0] CLBLL_L_X4Y150_SLICE_X4Y150_AMUX;
  wire [0:0] CLBLL_L_X4Y150_SLICE_X4Y150_AO5;
  wire [0:0] CLBLL_L_X4Y150_SLICE_X4Y150_AO6;
  wire [0:0] CLBLL_L_X4Y150_SLICE_X4Y150_AQ;
  wire [0:0] CLBLL_L_X4Y150_SLICE_X4Y150_A_CY;
  wire [0:0] CLBLL_L_X4Y150_SLICE_X4Y150_A_XOR;
  wire [0:0] CLBLL_L_X4Y150_SLICE_X4Y150_B;
  wire [0:0] CLBLL_L_X4Y150_SLICE_X4Y150_B1;
  wire [0:0] CLBLL_L_X4Y150_SLICE_X4Y150_B2;
  wire [0:0] CLBLL_L_X4Y150_SLICE_X4Y150_B3;
  wire [0:0] CLBLL_L_X4Y150_SLICE_X4Y150_B4;
  wire [0:0] CLBLL_L_X4Y150_SLICE_X4Y150_B5;
  wire [0:0] CLBLL_L_X4Y150_SLICE_X4Y150_B5Q;
  wire [0:0] CLBLL_L_X4Y150_SLICE_X4Y150_B6;
  wire [0:0] CLBLL_L_X4Y150_SLICE_X4Y150_BMUX;
  wire [0:0] CLBLL_L_X4Y150_SLICE_X4Y150_BO5;
  wire [0:0] CLBLL_L_X4Y150_SLICE_X4Y150_BO6;
  wire [0:0] CLBLL_L_X4Y150_SLICE_X4Y150_BQ;
  wire [0:0] CLBLL_L_X4Y150_SLICE_X4Y150_B_CY;
  wire [0:0] CLBLL_L_X4Y150_SLICE_X4Y150_B_XOR;
  wire [0:0] CLBLL_L_X4Y150_SLICE_X4Y150_C;
  wire [0:0] CLBLL_L_X4Y150_SLICE_X4Y150_C1;
  wire [0:0] CLBLL_L_X4Y150_SLICE_X4Y150_C2;
  wire [0:0] CLBLL_L_X4Y150_SLICE_X4Y150_C3;
  wire [0:0] CLBLL_L_X4Y150_SLICE_X4Y150_C4;
  wire [0:0] CLBLL_L_X4Y150_SLICE_X4Y150_C5;
  wire [0:0] CLBLL_L_X4Y150_SLICE_X4Y150_C5Q;
  wire [0:0] CLBLL_L_X4Y150_SLICE_X4Y150_C6;
  wire [0:0] CLBLL_L_X4Y150_SLICE_X4Y150_CLK;
  wire [0:0] CLBLL_L_X4Y150_SLICE_X4Y150_CMUX;
  wire [0:0] CLBLL_L_X4Y150_SLICE_X4Y150_CO5;
  wire [0:0] CLBLL_L_X4Y150_SLICE_X4Y150_CO6;
  wire [0:0] CLBLL_L_X4Y150_SLICE_X4Y150_CQ;
  wire [0:0] CLBLL_L_X4Y150_SLICE_X4Y150_C_CY;
  wire [0:0] CLBLL_L_X4Y150_SLICE_X4Y150_C_XOR;
  wire [0:0] CLBLL_L_X4Y150_SLICE_X4Y150_D;
  wire [0:0] CLBLL_L_X4Y150_SLICE_X4Y150_D1;
  wire [0:0] CLBLL_L_X4Y150_SLICE_X4Y150_D2;
  wire [0:0] CLBLL_L_X4Y150_SLICE_X4Y150_D3;
  wire [0:0] CLBLL_L_X4Y150_SLICE_X4Y150_D4;
  wire [0:0] CLBLL_L_X4Y150_SLICE_X4Y150_D5;
  wire [0:0] CLBLL_L_X4Y150_SLICE_X4Y150_D6;
  wire [0:0] CLBLL_L_X4Y150_SLICE_X4Y150_DO5;
  wire [0:0] CLBLL_L_X4Y150_SLICE_X4Y150_DO6;
  wire [0:0] CLBLL_L_X4Y150_SLICE_X4Y150_D_CY;
  wire [0:0] CLBLL_L_X4Y150_SLICE_X4Y150_D_XOR;
  wire [0:0] CLBLL_L_X4Y150_SLICE_X5Y150_A;
  wire [0:0] CLBLL_L_X4Y150_SLICE_X5Y150_A1;
  wire [0:0] CLBLL_L_X4Y150_SLICE_X5Y150_A2;
  wire [0:0] CLBLL_L_X4Y150_SLICE_X5Y150_A3;
  wire [0:0] CLBLL_L_X4Y150_SLICE_X5Y150_A4;
  wire [0:0] CLBLL_L_X4Y150_SLICE_X5Y150_A5;
  wire [0:0] CLBLL_L_X4Y150_SLICE_X5Y150_A5Q;
  wire [0:0] CLBLL_L_X4Y150_SLICE_X5Y150_A6;
  wire [0:0] CLBLL_L_X4Y150_SLICE_X5Y150_AMUX;
  wire [0:0] CLBLL_L_X4Y150_SLICE_X5Y150_AO5;
  wire [0:0] CLBLL_L_X4Y150_SLICE_X5Y150_AO6;
  wire [0:0] CLBLL_L_X4Y150_SLICE_X5Y150_AQ;
  wire [0:0] CLBLL_L_X4Y150_SLICE_X5Y150_AX;
  wire [0:0] CLBLL_L_X4Y150_SLICE_X5Y150_A_CY;
  wire [0:0] CLBLL_L_X4Y150_SLICE_X5Y150_A_XOR;
  wire [0:0] CLBLL_L_X4Y150_SLICE_X5Y150_B;
  wire [0:0] CLBLL_L_X4Y150_SLICE_X5Y150_B1;
  wire [0:0] CLBLL_L_X4Y150_SLICE_X5Y150_B2;
  wire [0:0] CLBLL_L_X4Y150_SLICE_X5Y150_B3;
  wire [0:0] CLBLL_L_X4Y150_SLICE_X5Y150_B4;
  wire [0:0] CLBLL_L_X4Y150_SLICE_X5Y150_B5;
  wire [0:0] CLBLL_L_X4Y150_SLICE_X5Y150_B6;
  wire [0:0] CLBLL_L_X4Y150_SLICE_X5Y150_BO5;
  wire [0:0] CLBLL_L_X4Y150_SLICE_X5Y150_BO6;
  wire [0:0] CLBLL_L_X4Y150_SLICE_X5Y150_BQ;
  wire [0:0] CLBLL_L_X4Y150_SLICE_X5Y150_B_CY;
  wire [0:0] CLBLL_L_X4Y150_SLICE_X5Y150_B_XOR;
  wire [0:0] CLBLL_L_X4Y150_SLICE_X5Y150_C;
  wire [0:0] CLBLL_L_X4Y150_SLICE_X5Y150_C1;
  wire [0:0] CLBLL_L_X4Y150_SLICE_X5Y150_C2;
  wire [0:0] CLBLL_L_X4Y150_SLICE_X5Y150_C3;
  wire [0:0] CLBLL_L_X4Y150_SLICE_X5Y150_C4;
  wire [0:0] CLBLL_L_X4Y150_SLICE_X5Y150_C5;
  wire [0:0] CLBLL_L_X4Y150_SLICE_X5Y150_C6;
  wire [0:0] CLBLL_L_X4Y150_SLICE_X5Y150_CLK;
  wire [0:0] CLBLL_L_X4Y150_SLICE_X5Y150_CMUX;
  wire [0:0] CLBLL_L_X4Y150_SLICE_X5Y150_CO5;
  wire [0:0] CLBLL_L_X4Y150_SLICE_X5Y150_CO6;
  wire [0:0] CLBLL_L_X4Y150_SLICE_X5Y150_C_CY;
  wire [0:0] CLBLL_L_X4Y150_SLICE_X5Y150_C_XOR;
  wire [0:0] CLBLL_L_X4Y150_SLICE_X5Y150_D;
  wire [0:0] CLBLL_L_X4Y150_SLICE_X5Y150_D1;
  wire [0:0] CLBLL_L_X4Y150_SLICE_X5Y150_D2;
  wire [0:0] CLBLL_L_X4Y150_SLICE_X5Y150_D3;
  wire [0:0] CLBLL_L_X4Y150_SLICE_X5Y150_D4;
  wire [0:0] CLBLL_L_X4Y150_SLICE_X5Y150_D5;
  wire [0:0] CLBLL_L_X4Y150_SLICE_X5Y150_D6;
  wire [0:0] CLBLL_L_X4Y150_SLICE_X5Y150_DO5;
  wire [0:0] CLBLL_L_X4Y150_SLICE_X5Y150_DO6;
  wire [0:0] CLBLL_L_X4Y150_SLICE_X5Y150_D_CY;
  wire [0:0] CLBLL_L_X4Y150_SLICE_X5Y150_D_XOR;
  wire [0:0] CLBLL_L_X4Y151_SLICE_X4Y151_A;
  wire [0:0] CLBLL_L_X4Y151_SLICE_X4Y151_A1;
  wire [0:0] CLBLL_L_X4Y151_SLICE_X4Y151_A2;
  wire [0:0] CLBLL_L_X4Y151_SLICE_X4Y151_A3;
  wire [0:0] CLBLL_L_X4Y151_SLICE_X4Y151_A4;
  wire [0:0] CLBLL_L_X4Y151_SLICE_X4Y151_A5;
  wire [0:0] CLBLL_L_X4Y151_SLICE_X4Y151_A5Q;
  wire [0:0] CLBLL_L_X4Y151_SLICE_X4Y151_A6;
  wire [0:0] CLBLL_L_X4Y151_SLICE_X4Y151_AMUX;
  wire [0:0] CLBLL_L_X4Y151_SLICE_X4Y151_AO5;
  wire [0:0] CLBLL_L_X4Y151_SLICE_X4Y151_AO6;
  wire [0:0] CLBLL_L_X4Y151_SLICE_X4Y151_AQ;
  wire [0:0] CLBLL_L_X4Y151_SLICE_X4Y151_AX;
  wire [0:0] CLBLL_L_X4Y151_SLICE_X4Y151_A_CY;
  wire [0:0] CLBLL_L_X4Y151_SLICE_X4Y151_A_XOR;
  wire [0:0] CLBLL_L_X4Y151_SLICE_X4Y151_B;
  wire [0:0] CLBLL_L_X4Y151_SLICE_X4Y151_B1;
  wire [0:0] CLBLL_L_X4Y151_SLICE_X4Y151_B2;
  wire [0:0] CLBLL_L_X4Y151_SLICE_X4Y151_B3;
  wire [0:0] CLBLL_L_X4Y151_SLICE_X4Y151_B4;
  wire [0:0] CLBLL_L_X4Y151_SLICE_X4Y151_B5;
  wire [0:0] CLBLL_L_X4Y151_SLICE_X4Y151_B5Q;
  wire [0:0] CLBLL_L_X4Y151_SLICE_X4Y151_B6;
  wire [0:0] CLBLL_L_X4Y151_SLICE_X4Y151_BMUX;
  wire [0:0] CLBLL_L_X4Y151_SLICE_X4Y151_BO5;
  wire [0:0] CLBLL_L_X4Y151_SLICE_X4Y151_BO6;
  wire [0:0] CLBLL_L_X4Y151_SLICE_X4Y151_BQ;
  wire [0:0] CLBLL_L_X4Y151_SLICE_X4Y151_B_CY;
  wire [0:0] CLBLL_L_X4Y151_SLICE_X4Y151_B_XOR;
  wire [0:0] CLBLL_L_X4Y151_SLICE_X4Y151_C;
  wire [0:0] CLBLL_L_X4Y151_SLICE_X4Y151_C1;
  wire [0:0] CLBLL_L_X4Y151_SLICE_X4Y151_C2;
  wire [0:0] CLBLL_L_X4Y151_SLICE_X4Y151_C3;
  wire [0:0] CLBLL_L_X4Y151_SLICE_X4Y151_C4;
  wire [0:0] CLBLL_L_X4Y151_SLICE_X4Y151_C5;
  wire [0:0] CLBLL_L_X4Y151_SLICE_X4Y151_C5Q;
  wire [0:0] CLBLL_L_X4Y151_SLICE_X4Y151_C6;
  wire [0:0] CLBLL_L_X4Y151_SLICE_X4Y151_CLK;
  wire [0:0] CLBLL_L_X4Y151_SLICE_X4Y151_CMUX;
  wire [0:0] CLBLL_L_X4Y151_SLICE_X4Y151_CO5;
  wire [0:0] CLBLL_L_X4Y151_SLICE_X4Y151_CO6;
  wire [0:0] CLBLL_L_X4Y151_SLICE_X4Y151_CQ;
  wire [0:0] CLBLL_L_X4Y151_SLICE_X4Y151_C_CY;
  wire [0:0] CLBLL_L_X4Y151_SLICE_X4Y151_C_XOR;
  wire [0:0] CLBLL_L_X4Y151_SLICE_X4Y151_D;
  wire [0:0] CLBLL_L_X4Y151_SLICE_X4Y151_D1;
  wire [0:0] CLBLL_L_X4Y151_SLICE_X4Y151_D2;
  wire [0:0] CLBLL_L_X4Y151_SLICE_X4Y151_D3;
  wire [0:0] CLBLL_L_X4Y151_SLICE_X4Y151_D4;
  wire [0:0] CLBLL_L_X4Y151_SLICE_X4Y151_D5;
  wire [0:0] CLBLL_L_X4Y151_SLICE_X4Y151_D6;
  wire [0:0] CLBLL_L_X4Y151_SLICE_X4Y151_DO5;
  wire [0:0] CLBLL_L_X4Y151_SLICE_X4Y151_DO6;
  wire [0:0] CLBLL_L_X4Y151_SLICE_X4Y151_DQ;
  wire [0:0] CLBLL_L_X4Y151_SLICE_X4Y151_D_CY;
  wire [0:0] CLBLL_L_X4Y151_SLICE_X4Y151_D_XOR;
  wire [0:0] CLBLL_L_X4Y151_SLICE_X5Y151_A;
  wire [0:0] CLBLL_L_X4Y151_SLICE_X5Y151_A1;
  wire [0:0] CLBLL_L_X4Y151_SLICE_X5Y151_A2;
  wire [0:0] CLBLL_L_X4Y151_SLICE_X5Y151_A3;
  wire [0:0] CLBLL_L_X4Y151_SLICE_X5Y151_A4;
  wire [0:0] CLBLL_L_X4Y151_SLICE_X5Y151_A5;
  wire [0:0] CLBLL_L_X4Y151_SLICE_X5Y151_A6;
  wire [0:0] CLBLL_L_X4Y151_SLICE_X5Y151_AO5;
  wire [0:0] CLBLL_L_X4Y151_SLICE_X5Y151_AO6;
  wire [0:0] CLBLL_L_X4Y151_SLICE_X5Y151_AQ;
  wire [0:0] CLBLL_L_X4Y151_SLICE_X5Y151_A_CY;
  wire [0:0] CLBLL_L_X4Y151_SLICE_X5Y151_A_XOR;
  wire [0:0] CLBLL_L_X4Y151_SLICE_X5Y151_B;
  wire [0:0] CLBLL_L_X4Y151_SLICE_X5Y151_B1;
  wire [0:0] CLBLL_L_X4Y151_SLICE_X5Y151_B2;
  wire [0:0] CLBLL_L_X4Y151_SLICE_X5Y151_B3;
  wire [0:0] CLBLL_L_X4Y151_SLICE_X5Y151_B4;
  wire [0:0] CLBLL_L_X4Y151_SLICE_X5Y151_B5;
  wire [0:0] CLBLL_L_X4Y151_SLICE_X5Y151_B5Q;
  wire [0:0] CLBLL_L_X4Y151_SLICE_X5Y151_B6;
  wire [0:0] CLBLL_L_X4Y151_SLICE_X5Y151_BMUX;
  wire [0:0] CLBLL_L_X4Y151_SLICE_X5Y151_BO5;
  wire [0:0] CLBLL_L_X4Y151_SLICE_X5Y151_BO6;
  wire [0:0] CLBLL_L_X4Y151_SLICE_X5Y151_BQ;
  wire [0:0] CLBLL_L_X4Y151_SLICE_X5Y151_B_CY;
  wire [0:0] CLBLL_L_X4Y151_SLICE_X5Y151_B_XOR;
  wire [0:0] CLBLL_L_X4Y151_SLICE_X5Y151_C;
  wire [0:0] CLBLL_L_X4Y151_SLICE_X5Y151_C1;
  wire [0:0] CLBLL_L_X4Y151_SLICE_X5Y151_C2;
  wire [0:0] CLBLL_L_X4Y151_SLICE_X5Y151_C3;
  wire [0:0] CLBLL_L_X4Y151_SLICE_X5Y151_C4;
  wire [0:0] CLBLL_L_X4Y151_SLICE_X5Y151_C5;
  wire [0:0] CLBLL_L_X4Y151_SLICE_X5Y151_C6;
  wire [0:0] CLBLL_L_X4Y151_SLICE_X5Y151_CLK;
  wire [0:0] CLBLL_L_X4Y151_SLICE_X5Y151_CO5;
  wire [0:0] CLBLL_L_X4Y151_SLICE_X5Y151_CO6;
  wire [0:0] CLBLL_L_X4Y151_SLICE_X5Y151_CQ;
  wire [0:0] CLBLL_L_X4Y151_SLICE_X5Y151_C_CY;
  wire [0:0] CLBLL_L_X4Y151_SLICE_X5Y151_C_XOR;
  wire [0:0] CLBLL_L_X4Y151_SLICE_X5Y151_D;
  wire [0:0] CLBLL_L_X4Y151_SLICE_X5Y151_D1;
  wire [0:0] CLBLL_L_X4Y151_SLICE_X5Y151_D2;
  wire [0:0] CLBLL_L_X4Y151_SLICE_X5Y151_D3;
  wire [0:0] CLBLL_L_X4Y151_SLICE_X5Y151_D4;
  wire [0:0] CLBLL_L_X4Y151_SLICE_X5Y151_D5;
  wire [0:0] CLBLL_L_X4Y151_SLICE_X5Y151_D5Q;
  wire [0:0] CLBLL_L_X4Y151_SLICE_X5Y151_D6;
  wire [0:0] CLBLL_L_X4Y151_SLICE_X5Y151_DMUX;
  wire [0:0] CLBLL_L_X4Y151_SLICE_X5Y151_DO5;
  wire [0:0] CLBLL_L_X4Y151_SLICE_X5Y151_DO6;
  wire [0:0] CLBLL_L_X4Y151_SLICE_X5Y151_DQ;
  wire [0:0] CLBLL_L_X4Y151_SLICE_X5Y151_D_CY;
  wire [0:0] CLBLL_L_X4Y151_SLICE_X5Y151_D_XOR;
  wire [0:0] CLBLL_L_X4Y152_SLICE_X4Y152_A;
  wire [0:0] CLBLL_L_X4Y152_SLICE_X4Y152_A1;
  wire [0:0] CLBLL_L_X4Y152_SLICE_X4Y152_A2;
  wire [0:0] CLBLL_L_X4Y152_SLICE_X4Y152_A3;
  wire [0:0] CLBLL_L_X4Y152_SLICE_X4Y152_A4;
  wire [0:0] CLBLL_L_X4Y152_SLICE_X4Y152_A5;
  wire [0:0] CLBLL_L_X4Y152_SLICE_X4Y152_A6;
  wire [0:0] CLBLL_L_X4Y152_SLICE_X4Y152_AO5;
  wire [0:0] CLBLL_L_X4Y152_SLICE_X4Y152_AO6;
  wire [0:0] CLBLL_L_X4Y152_SLICE_X4Y152_AQ;
  wire [0:0] CLBLL_L_X4Y152_SLICE_X4Y152_A_CY;
  wire [0:0] CLBLL_L_X4Y152_SLICE_X4Y152_A_XOR;
  wire [0:0] CLBLL_L_X4Y152_SLICE_X4Y152_B;
  wire [0:0] CLBLL_L_X4Y152_SLICE_X4Y152_B1;
  wire [0:0] CLBLL_L_X4Y152_SLICE_X4Y152_B2;
  wire [0:0] CLBLL_L_X4Y152_SLICE_X4Y152_B3;
  wire [0:0] CLBLL_L_X4Y152_SLICE_X4Y152_B4;
  wire [0:0] CLBLL_L_X4Y152_SLICE_X4Y152_B5;
  wire [0:0] CLBLL_L_X4Y152_SLICE_X4Y152_B5Q;
  wire [0:0] CLBLL_L_X4Y152_SLICE_X4Y152_B6;
  wire [0:0] CLBLL_L_X4Y152_SLICE_X4Y152_BMUX;
  wire [0:0] CLBLL_L_X4Y152_SLICE_X4Y152_BO5;
  wire [0:0] CLBLL_L_X4Y152_SLICE_X4Y152_BO6;
  wire [0:0] CLBLL_L_X4Y152_SLICE_X4Y152_BQ;
  wire [0:0] CLBLL_L_X4Y152_SLICE_X4Y152_B_CY;
  wire [0:0] CLBLL_L_X4Y152_SLICE_X4Y152_B_XOR;
  wire [0:0] CLBLL_L_X4Y152_SLICE_X4Y152_C;
  wire [0:0] CLBLL_L_X4Y152_SLICE_X4Y152_C1;
  wire [0:0] CLBLL_L_X4Y152_SLICE_X4Y152_C2;
  wire [0:0] CLBLL_L_X4Y152_SLICE_X4Y152_C3;
  wire [0:0] CLBLL_L_X4Y152_SLICE_X4Y152_C4;
  wire [0:0] CLBLL_L_X4Y152_SLICE_X4Y152_C5;
  wire [0:0] CLBLL_L_X4Y152_SLICE_X4Y152_C6;
  wire [0:0] CLBLL_L_X4Y152_SLICE_X4Y152_CLK;
  wire [0:0] CLBLL_L_X4Y152_SLICE_X4Y152_CO5;
  wire [0:0] CLBLL_L_X4Y152_SLICE_X4Y152_CO6;
  wire [0:0] CLBLL_L_X4Y152_SLICE_X4Y152_CQ;
  wire [0:0] CLBLL_L_X4Y152_SLICE_X4Y152_C_CY;
  wire [0:0] CLBLL_L_X4Y152_SLICE_X4Y152_C_XOR;
  wire [0:0] CLBLL_L_X4Y152_SLICE_X4Y152_D;
  wire [0:0] CLBLL_L_X4Y152_SLICE_X4Y152_D1;
  wire [0:0] CLBLL_L_X4Y152_SLICE_X4Y152_D2;
  wire [0:0] CLBLL_L_X4Y152_SLICE_X4Y152_D3;
  wire [0:0] CLBLL_L_X4Y152_SLICE_X4Y152_D4;
  wire [0:0] CLBLL_L_X4Y152_SLICE_X4Y152_D5;
  wire [0:0] CLBLL_L_X4Y152_SLICE_X4Y152_D6;
  wire [0:0] CLBLL_L_X4Y152_SLICE_X4Y152_DO5;
  wire [0:0] CLBLL_L_X4Y152_SLICE_X4Y152_DO6;
  wire [0:0] CLBLL_L_X4Y152_SLICE_X4Y152_DQ;
  wire [0:0] CLBLL_L_X4Y152_SLICE_X4Y152_D_CY;
  wire [0:0] CLBLL_L_X4Y152_SLICE_X4Y152_D_XOR;
  wire [0:0] CLBLL_L_X4Y152_SLICE_X5Y152_A;
  wire [0:0] CLBLL_L_X4Y152_SLICE_X5Y152_A1;
  wire [0:0] CLBLL_L_X4Y152_SLICE_X5Y152_A2;
  wire [0:0] CLBLL_L_X4Y152_SLICE_X5Y152_A3;
  wire [0:0] CLBLL_L_X4Y152_SLICE_X5Y152_A4;
  wire [0:0] CLBLL_L_X4Y152_SLICE_X5Y152_A5;
  wire [0:0] CLBLL_L_X4Y152_SLICE_X5Y152_A5Q;
  wire [0:0] CLBLL_L_X4Y152_SLICE_X5Y152_A6;
  wire [0:0] CLBLL_L_X4Y152_SLICE_X5Y152_AMUX;
  wire [0:0] CLBLL_L_X4Y152_SLICE_X5Y152_AO5;
  wire [0:0] CLBLL_L_X4Y152_SLICE_X5Y152_AO6;
  wire [0:0] CLBLL_L_X4Y152_SLICE_X5Y152_AQ;
  wire [0:0] CLBLL_L_X4Y152_SLICE_X5Y152_AX;
  wire [0:0] CLBLL_L_X4Y152_SLICE_X5Y152_A_CY;
  wire [0:0] CLBLL_L_X4Y152_SLICE_X5Y152_A_XOR;
  wire [0:0] CLBLL_L_X4Y152_SLICE_X5Y152_B;
  wire [0:0] CLBLL_L_X4Y152_SLICE_X5Y152_B1;
  wire [0:0] CLBLL_L_X4Y152_SLICE_X5Y152_B2;
  wire [0:0] CLBLL_L_X4Y152_SLICE_X5Y152_B3;
  wire [0:0] CLBLL_L_X4Y152_SLICE_X5Y152_B4;
  wire [0:0] CLBLL_L_X4Y152_SLICE_X5Y152_B5;
  wire [0:0] CLBLL_L_X4Y152_SLICE_X5Y152_B6;
  wire [0:0] CLBLL_L_X4Y152_SLICE_X5Y152_BO5;
  wire [0:0] CLBLL_L_X4Y152_SLICE_X5Y152_BO6;
  wire [0:0] CLBLL_L_X4Y152_SLICE_X5Y152_BQ;
  wire [0:0] CLBLL_L_X4Y152_SLICE_X5Y152_B_CY;
  wire [0:0] CLBLL_L_X4Y152_SLICE_X5Y152_B_XOR;
  wire [0:0] CLBLL_L_X4Y152_SLICE_X5Y152_C;
  wire [0:0] CLBLL_L_X4Y152_SLICE_X5Y152_C1;
  wire [0:0] CLBLL_L_X4Y152_SLICE_X5Y152_C2;
  wire [0:0] CLBLL_L_X4Y152_SLICE_X5Y152_C3;
  wire [0:0] CLBLL_L_X4Y152_SLICE_X5Y152_C4;
  wire [0:0] CLBLL_L_X4Y152_SLICE_X5Y152_C5;
  wire [0:0] CLBLL_L_X4Y152_SLICE_X5Y152_C6;
  wire [0:0] CLBLL_L_X4Y152_SLICE_X5Y152_CLK;
  wire [0:0] CLBLL_L_X4Y152_SLICE_X5Y152_CMUX;
  wire [0:0] CLBLL_L_X4Y152_SLICE_X5Y152_CO5;
  wire [0:0] CLBLL_L_X4Y152_SLICE_X5Y152_CO6;
  wire [0:0] CLBLL_L_X4Y152_SLICE_X5Y152_C_CY;
  wire [0:0] CLBLL_L_X4Y152_SLICE_X5Y152_C_XOR;
  wire [0:0] CLBLL_L_X4Y152_SLICE_X5Y152_D;
  wire [0:0] CLBLL_L_X4Y152_SLICE_X5Y152_D1;
  wire [0:0] CLBLL_L_X4Y152_SLICE_X5Y152_D2;
  wire [0:0] CLBLL_L_X4Y152_SLICE_X5Y152_D3;
  wire [0:0] CLBLL_L_X4Y152_SLICE_X5Y152_D4;
  wire [0:0] CLBLL_L_X4Y152_SLICE_X5Y152_D5;
  wire [0:0] CLBLL_L_X4Y152_SLICE_X5Y152_D6;
  wire [0:0] CLBLL_L_X4Y152_SLICE_X5Y152_DO5;
  wire [0:0] CLBLL_L_X4Y152_SLICE_X5Y152_DO6;
  wire [0:0] CLBLL_L_X4Y152_SLICE_X5Y152_D_CY;
  wire [0:0] CLBLL_L_X4Y152_SLICE_X5Y152_D_XOR;
  wire [0:0] CLBLL_L_X4Y153_SLICE_X4Y153_A;
  wire [0:0] CLBLL_L_X4Y153_SLICE_X4Y153_A1;
  wire [0:0] CLBLL_L_X4Y153_SLICE_X4Y153_A2;
  wire [0:0] CLBLL_L_X4Y153_SLICE_X4Y153_A3;
  wire [0:0] CLBLL_L_X4Y153_SLICE_X4Y153_A4;
  wire [0:0] CLBLL_L_X4Y153_SLICE_X4Y153_A5;
  wire [0:0] CLBLL_L_X4Y153_SLICE_X4Y153_A5Q;
  wire [0:0] CLBLL_L_X4Y153_SLICE_X4Y153_A6;
  wire [0:0] CLBLL_L_X4Y153_SLICE_X4Y153_AMUX;
  wire [0:0] CLBLL_L_X4Y153_SLICE_X4Y153_AO5;
  wire [0:0] CLBLL_L_X4Y153_SLICE_X4Y153_AO6;
  wire [0:0] CLBLL_L_X4Y153_SLICE_X4Y153_AQ;
  wire [0:0] CLBLL_L_X4Y153_SLICE_X4Y153_A_CY;
  wire [0:0] CLBLL_L_X4Y153_SLICE_X4Y153_A_XOR;
  wire [0:0] CLBLL_L_X4Y153_SLICE_X4Y153_B;
  wire [0:0] CLBLL_L_X4Y153_SLICE_X4Y153_B1;
  wire [0:0] CLBLL_L_X4Y153_SLICE_X4Y153_B2;
  wire [0:0] CLBLL_L_X4Y153_SLICE_X4Y153_B3;
  wire [0:0] CLBLL_L_X4Y153_SLICE_X4Y153_B4;
  wire [0:0] CLBLL_L_X4Y153_SLICE_X4Y153_B5;
  wire [0:0] CLBLL_L_X4Y153_SLICE_X4Y153_B5Q;
  wire [0:0] CLBLL_L_X4Y153_SLICE_X4Y153_B6;
  wire [0:0] CLBLL_L_X4Y153_SLICE_X4Y153_BMUX;
  wire [0:0] CLBLL_L_X4Y153_SLICE_X4Y153_BO5;
  wire [0:0] CLBLL_L_X4Y153_SLICE_X4Y153_BO6;
  wire [0:0] CLBLL_L_X4Y153_SLICE_X4Y153_BQ;
  wire [0:0] CLBLL_L_X4Y153_SLICE_X4Y153_B_CY;
  wire [0:0] CLBLL_L_X4Y153_SLICE_X4Y153_B_XOR;
  wire [0:0] CLBLL_L_X4Y153_SLICE_X4Y153_C;
  wire [0:0] CLBLL_L_X4Y153_SLICE_X4Y153_C1;
  wire [0:0] CLBLL_L_X4Y153_SLICE_X4Y153_C2;
  wire [0:0] CLBLL_L_X4Y153_SLICE_X4Y153_C3;
  wire [0:0] CLBLL_L_X4Y153_SLICE_X4Y153_C4;
  wire [0:0] CLBLL_L_X4Y153_SLICE_X4Y153_C5;
  wire [0:0] CLBLL_L_X4Y153_SLICE_X4Y153_C6;
  wire [0:0] CLBLL_L_X4Y153_SLICE_X4Y153_CLK;
  wire [0:0] CLBLL_L_X4Y153_SLICE_X4Y153_CMUX;
  wire [0:0] CLBLL_L_X4Y153_SLICE_X4Y153_CO5;
  wire [0:0] CLBLL_L_X4Y153_SLICE_X4Y153_CO6;
  wire [0:0] CLBLL_L_X4Y153_SLICE_X4Y153_C_CY;
  wire [0:0] CLBLL_L_X4Y153_SLICE_X4Y153_C_XOR;
  wire [0:0] CLBLL_L_X4Y153_SLICE_X4Y153_D;
  wire [0:0] CLBLL_L_X4Y153_SLICE_X4Y153_D1;
  wire [0:0] CLBLL_L_X4Y153_SLICE_X4Y153_D2;
  wire [0:0] CLBLL_L_X4Y153_SLICE_X4Y153_D3;
  wire [0:0] CLBLL_L_X4Y153_SLICE_X4Y153_D4;
  wire [0:0] CLBLL_L_X4Y153_SLICE_X4Y153_D5;
  wire [0:0] CLBLL_L_X4Y153_SLICE_X4Y153_D6;
  wire [0:0] CLBLL_L_X4Y153_SLICE_X4Y153_DMUX;
  wire [0:0] CLBLL_L_X4Y153_SLICE_X4Y153_DO5;
  wire [0:0] CLBLL_L_X4Y153_SLICE_X4Y153_DO6;
  wire [0:0] CLBLL_L_X4Y153_SLICE_X4Y153_D_CY;
  wire [0:0] CLBLL_L_X4Y153_SLICE_X4Y153_D_XOR;
  wire [0:0] CLBLL_L_X4Y153_SLICE_X5Y153_A;
  wire [0:0] CLBLL_L_X4Y153_SLICE_X5Y153_A1;
  wire [0:0] CLBLL_L_X4Y153_SLICE_X5Y153_A2;
  wire [0:0] CLBLL_L_X4Y153_SLICE_X5Y153_A3;
  wire [0:0] CLBLL_L_X4Y153_SLICE_X5Y153_A4;
  wire [0:0] CLBLL_L_X4Y153_SLICE_X5Y153_A5;
  wire [0:0] CLBLL_L_X4Y153_SLICE_X5Y153_A5Q;
  wire [0:0] CLBLL_L_X4Y153_SLICE_X5Y153_A6;
  wire [0:0] CLBLL_L_X4Y153_SLICE_X5Y153_AMUX;
  wire [0:0] CLBLL_L_X4Y153_SLICE_X5Y153_AO5;
  wire [0:0] CLBLL_L_X4Y153_SLICE_X5Y153_AO6;
  wire [0:0] CLBLL_L_X4Y153_SLICE_X5Y153_AQ;
  wire [0:0] CLBLL_L_X4Y153_SLICE_X5Y153_AX;
  wire [0:0] CLBLL_L_X4Y153_SLICE_X5Y153_A_CY;
  wire [0:0] CLBLL_L_X4Y153_SLICE_X5Y153_A_XOR;
  wire [0:0] CLBLL_L_X4Y153_SLICE_X5Y153_B;
  wire [0:0] CLBLL_L_X4Y153_SLICE_X5Y153_B1;
  wire [0:0] CLBLL_L_X4Y153_SLICE_X5Y153_B2;
  wire [0:0] CLBLL_L_X4Y153_SLICE_X5Y153_B3;
  wire [0:0] CLBLL_L_X4Y153_SLICE_X5Y153_B4;
  wire [0:0] CLBLL_L_X4Y153_SLICE_X5Y153_B5;
  wire [0:0] CLBLL_L_X4Y153_SLICE_X5Y153_B6;
  wire [0:0] CLBLL_L_X4Y153_SLICE_X5Y153_BMUX;
  wire [0:0] CLBLL_L_X4Y153_SLICE_X5Y153_BO5;
  wire [0:0] CLBLL_L_X4Y153_SLICE_X5Y153_BO6;
  wire [0:0] CLBLL_L_X4Y153_SLICE_X5Y153_B_CY;
  wire [0:0] CLBLL_L_X4Y153_SLICE_X5Y153_B_XOR;
  wire [0:0] CLBLL_L_X4Y153_SLICE_X5Y153_C;
  wire [0:0] CLBLL_L_X4Y153_SLICE_X5Y153_C1;
  wire [0:0] CLBLL_L_X4Y153_SLICE_X5Y153_C2;
  wire [0:0] CLBLL_L_X4Y153_SLICE_X5Y153_C3;
  wire [0:0] CLBLL_L_X4Y153_SLICE_X5Y153_C4;
  wire [0:0] CLBLL_L_X4Y153_SLICE_X5Y153_C5;
  wire [0:0] CLBLL_L_X4Y153_SLICE_X5Y153_C6;
  wire [0:0] CLBLL_L_X4Y153_SLICE_X5Y153_CLK;
  wire [0:0] CLBLL_L_X4Y153_SLICE_X5Y153_CO5;
  wire [0:0] CLBLL_L_X4Y153_SLICE_X5Y153_CO6;
  wire [0:0] CLBLL_L_X4Y153_SLICE_X5Y153_C_CY;
  wire [0:0] CLBLL_L_X4Y153_SLICE_X5Y153_C_XOR;
  wire [0:0] CLBLL_L_X4Y153_SLICE_X5Y153_D;
  wire [0:0] CLBLL_L_X4Y153_SLICE_X5Y153_D1;
  wire [0:0] CLBLL_L_X4Y153_SLICE_X5Y153_D2;
  wire [0:0] CLBLL_L_X4Y153_SLICE_X5Y153_D3;
  wire [0:0] CLBLL_L_X4Y153_SLICE_X5Y153_D4;
  wire [0:0] CLBLL_L_X4Y153_SLICE_X5Y153_D5;
  wire [0:0] CLBLL_L_X4Y153_SLICE_X5Y153_D6;
  wire [0:0] CLBLL_L_X4Y153_SLICE_X5Y153_DO5;
  wire [0:0] CLBLL_L_X4Y153_SLICE_X5Y153_DO6;
  wire [0:0] CLBLL_L_X4Y153_SLICE_X5Y153_D_CY;
  wire [0:0] CLBLL_L_X4Y153_SLICE_X5Y153_D_XOR;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X12Y142_A;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X12Y142_A1;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X12Y142_A2;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X12Y142_A3;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X12Y142_A4;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X12Y142_A5;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X12Y142_A6;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X12Y142_AO5;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X12Y142_AO6;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X12Y142_AQ;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X12Y142_A_CY;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X12Y142_A_XOR;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X12Y142_B;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X12Y142_B1;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X12Y142_B2;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X12Y142_B3;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X12Y142_B4;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X12Y142_B5;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X12Y142_B6;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X12Y142_BO5;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X12Y142_BO6;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X12Y142_B_CY;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X12Y142_B_XOR;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X12Y142_C;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X12Y142_C1;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X12Y142_C2;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X12Y142_C3;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X12Y142_C4;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X12Y142_C5;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X12Y142_C6;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X12Y142_CLK;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X12Y142_CO5;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X12Y142_CO6;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X12Y142_C_CY;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X12Y142_C_XOR;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X12Y142_D;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X12Y142_D1;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X12Y142_D2;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X12Y142_D3;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X12Y142_D4;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X12Y142_D5;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X12Y142_D6;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X12Y142_DO5;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X12Y142_DO6;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X12Y142_D_CY;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X12Y142_D_XOR;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X13Y142_A;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X13Y142_A1;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X13Y142_A2;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X13Y142_A3;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X13Y142_A4;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X13Y142_A5;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X13Y142_A6;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X13Y142_AO5;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X13Y142_AO6;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X13Y142_AQ;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X13Y142_A_CY;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X13Y142_A_XOR;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X13Y142_B;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X13Y142_B1;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X13Y142_B2;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X13Y142_B3;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X13Y142_B4;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X13Y142_B5;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X13Y142_B6;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X13Y142_BO5;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X13Y142_BO6;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X13Y142_B_CY;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X13Y142_B_XOR;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X13Y142_C;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X13Y142_C1;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X13Y142_C2;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X13Y142_C3;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X13Y142_C4;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X13Y142_C5;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X13Y142_C6;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X13Y142_CLK;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X13Y142_CO5;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X13Y142_CO6;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X13Y142_C_CY;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X13Y142_C_XOR;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X13Y142_D;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X13Y142_D1;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X13Y142_D2;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X13Y142_D3;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X13Y142_D4;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X13Y142_D5;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X13Y142_D6;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X13Y142_DO5;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X13Y142_DO6;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X13Y142_D_CY;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X13Y142_D_XOR;
  wire [0:0] CLBLM_L_X10Y143_SLICE_X12Y143_A;
  wire [0:0] CLBLM_L_X10Y143_SLICE_X12Y143_A1;
  wire [0:0] CLBLM_L_X10Y143_SLICE_X12Y143_A2;
  wire [0:0] CLBLM_L_X10Y143_SLICE_X12Y143_A3;
  wire [0:0] CLBLM_L_X10Y143_SLICE_X12Y143_A4;
  wire [0:0] CLBLM_L_X10Y143_SLICE_X12Y143_A5;
  wire [0:0] CLBLM_L_X10Y143_SLICE_X12Y143_A6;
  wire [0:0] CLBLM_L_X10Y143_SLICE_X12Y143_AO5;
  wire [0:0] CLBLM_L_X10Y143_SLICE_X12Y143_AO6;
  wire [0:0] CLBLM_L_X10Y143_SLICE_X12Y143_AQ;
  wire [0:0] CLBLM_L_X10Y143_SLICE_X12Y143_A_CY;
  wire [0:0] CLBLM_L_X10Y143_SLICE_X12Y143_A_XOR;
  wire [0:0] CLBLM_L_X10Y143_SLICE_X12Y143_B;
  wire [0:0] CLBLM_L_X10Y143_SLICE_X12Y143_B1;
  wire [0:0] CLBLM_L_X10Y143_SLICE_X12Y143_B2;
  wire [0:0] CLBLM_L_X10Y143_SLICE_X12Y143_B3;
  wire [0:0] CLBLM_L_X10Y143_SLICE_X12Y143_B4;
  wire [0:0] CLBLM_L_X10Y143_SLICE_X12Y143_B5;
  wire [0:0] CLBLM_L_X10Y143_SLICE_X12Y143_B6;
  wire [0:0] CLBLM_L_X10Y143_SLICE_X12Y143_BO5;
  wire [0:0] CLBLM_L_X10Y143_SLICE_X12Y143_BO6;
  wire [0:0] CLBLM_L_X10Y143_SLICE_X12Y143_BQ;
  wire [0:0] CLBLM_L_X10Y143_SLICE_X12Y143_B_CY;
  wire [0:0] CLBLM_L_X10Y143_SLICE_X12Y143_B_XOR;
  wire [0:0] CLBLM_L_X10Y143_SLICE_X12Y143_C;
  wire [0:0] CLBLM_L_X10Y143_SLICE_X12Y143_C1;
  wire [0:0] CLBLM_L_X10Y143_SLICE_X12Y143_C2;
  wire [0:0] CLBLM_L_X10Y143_SLICE_X12Y143_C3;
  wire [0:0] CLBLM_L_X10Y143_SLICE_X12Y143_C4;
  wire [0:0] CLBLM_L_X10Y143_SLICE_X12Y143_C5;
  wire [0:0] CLBLM_L_X10Y143_SLICE_X12Y143_C6;
  wire [0:0] CLBLM_L_X10Y143_SLICE_X12Y143_CLK;
  wire [0:0] CLBLM_L_X10Y143_SLICE_X12Y143_CMUX;
  wire [0:0] CLBLM_L_X10Y143_SLICE_X12Y143_CO5;
  wire [0:0] CLBLM_L_X10Y143_SLICE_X12Y143_CO6;
  wire [0:0] CLBLM_L_X10Y143_SLICE_X12Y143_C_CY;
  wire [0:0] CLBLM_L_X10Y143_SLICE_X12Y143_C_XOR;
  wire [0:0] CLBLM_L_X10Y143_SLICE_X12Y143_D;
  wire [0:0] CLBLM_L_X10Y143_SLICE_X12Y143_D1;
  wire [0:0] CLBLM_L_X10Y143_SLICE_X12Y143_D2;
  wire [0:0] CLBLM_L_X10Y143_SLICE_X12Y143_D3;
  wire [0:0] CLBLM_L_X10Y143_SLICE_X12Y143_D4;
  wire [0:0] CLBLM_L_X10Y143_SLICE_X12Y143_D5;
  wire [0:0] CLBLM_L_X10Y143_SLICE_X12Y143_D6;
  wire [0:0] CLBLM_L_X10Y143_SLICE_X12Y143_DO5;
  wire [0:0] CLBLM_L_X10Y143_SLICE_X12Y143_DO6;
  wire [0:0] CLBLM_L_X10Y143_SLICE_X12Y143_D_CY;
  wire [0:0] CLBLM_L_X10Y143_SLICE_X12Y143_D_XOR;
  wire [0:0] CLBLM_L_X10Y143_SLICE_X13Y143_A;
  wire [0:0] CLBLM_L_X10Y143_SLICE_X13Y143_A1;
  wire [0:0] CLBLM_L_X10Y143_SLICE_X13Y143_A2;
  wire [0:0] CLBLM_L_X10Y143_SLICE_X13Y143_A3;
  wire [0:0] CLBLM_L_X10Y143_SLICE_X13Y143_A4;
  wire [0:0] CLBLM_L_X10Y143_SLICE_X13Y143_A5;
  wire [0:0] CLBLM_L_X10Y143_SLICE_X13Y143_A6;
  wire [0:0] CLBLM_L_X10Y143_SLICE_X13Y143_AO5;
  wire [0:0] CLBLM_L_X10Y143_SLICE_X13Y143_AO6;
  wire [0:0] CLBLM_L_X10Y143_SLICE_X13Y143_AQ;
  wire [0:0] CLBLM_L_X10Y143_SLICE_X13Y143_A_CY;
  wire [0:0] CLBLM_L_X10Y143_SLICE_X13Y143_A_XOR;
  wire [0:0] CLBLM_L_X10Y143_SLICE_X13Y143_B;
  wire [0:0] CLBLM_L_X10Y143_SLICE_X13Y143_B1;
  wire [0:0] CLBLM_L_X10Y143_SLICE_X13Y143_B2;
  wire [0:0] CLBLM_L_X10Y143_SLICE_X13Y143_B3;
  wire [0:0] CLBLM_L_X10Y143_SLICE_X13Y143_B4;
  wire [0:0] CLBLM_L_X10Y143_SLICE_X13Y143_B5;
  wire [0:0] CLBLM_L_X10Y143_SLICE_X13Y143_B6;
  wire [0:0] CLBLM_L_X10Y143_SLICE_X13Y143_BO5;
  wire [0:0] CLBLM_L_X10Y143_SLICE_X13Y143_BO6;
  wire [0:0] CLBLM_L_X10Y143_SLICE_X13Y143_BQ;
  wire [0:0] CLBLM_L_X10Y143_SLICE_X13Y143_B_CY;
  wire [0:0] CLBLM_L_X10Y143_SLICE_X13Y143_B_XOR;
  wire [0:0] CLBLM_L_X10Y143_SLICE_X13Y143_C;
  wire [0:0] CLBLM_L_X10Y143_SLICE_X13Y143_C1;
  wire [0:0] CLBLM_L_X10Y143_SLICE_X13Y143_C2;
  wire [0:0] CLBLM_L_X10Y143_SLICE_X13Y143_C3;
  wire [0:0] CLBLM_L_X10Y143_SLICE_X13Y143_C4;
  wire [0:0] CLBLM_L_X10Y143_SLICE_X13Y143_C5;
  wire [0:0] CLBLM_L_X10Y143_SLICE_X13Y143_C5Q;
  wire [0:0] CLBLM_L_X10Y143_SLICE_X13Y143_C6;
  wire [0:0] CLBLM_L_X10Y143_SLICE_X13Y143_CLK;
  wire [0:0] CLBLM_L_X10Y143_SLICE_X13Y143_CMUX;
  wire [0:0] CLBLM_L_X10Y143_SLICE_X13Y143_CO5;
  wire [0:0] CLBLM_L_X10Y143_SLICE_X13Y143_CO6;
  wire [0:0] CLBLM_L_X10Y143_SLICE_X13Y143_CQ;
  wire [0:0] CLBLM_L_X10Y143_SLICE_X13Y143_C_CY;
  wire [0:0] CLBLM_L_X10Y143_SLICE_X13Y143_C_XOR;
  wire [0:0] CLBLM_L_X10Y143_SLICE_X13Y143_D;
  wire [0:0] CLBLM_L_X10Y143_SLICE_X13Y143_D1;
  wire [0:0] CLBLM_L_X10Y143_SLICE_X13Y143_D2;
  wire [0:0] CLBLM_L_X10Y143_SLICE_X13Y143_D3;
  wire [0:0] CLBLM_L_X10Y143_SLICE_X13Y143_D4;
  wire [0:0] CLBLM_L_X10Y143_SLICE_X13Y143_D5;
  wire [0:0] CLBLM_L_X10Y143_SLICE_X13Y143_D6;
  wire [0:0] CLBLM_L_X10Y143_SLICE_X13Y143_DMUX;
  wire [0:0] CLBLM_L_X10Y143_SLICE_X13Y143_DO5;
  wire [0:0] CLBLM_L_X10Y143_SLICE_X13Y143_DO6;
  wire [0:0] CLBLM_L_X10Y143_SLICE_X13Y143_D_CY;
  wire [0:0] CLBLM_L_X10Y143_SLICE_X13Y143_D_XOR;
  wire [0:0] CLBLM_L_X10Y144_SLICE_X12Y144_A;
  wire [0:0] CLBLM_L_X10Y144_SLICE_X12Y144_A1;
  wire [0:0] CLBLM_L_X10Y144_SLICE_X12Y144_A2;
  wire [0:0] CLBLM_L_X10Y144_SLICE_X12Y144_A3;
  wire [0:0] CLBLM_L_X10Y144_SLICE_X12Y144_A4;
  wire [0:0] CLBLM_L_X10Y144_SLICE_X12Y144_A5;
  wire [0:0] CLBLM_L_X10Y144_SLICE_X12Y144_A6;
  wire [0:0] CLBLM_L_X10Y144_SLICE_X12Y144_AMUX;
  wire [0:0] CLBLM_L_X10Y144_SLICE_X12Y144_AO5;
  wire [0:0] CLBLM_L_X10Y144_SLICE_X12Y144_AO6;
  wire [0:0] CLBLM_L_X10Y144_SLICE_X12Y144_AQ;
  wire [0:0] CLBLM_L_X10Y144_SLICE_X12Y144_AX;
  wire [0:0] CLBLM_L_X10Y144_SLICE_X12Y144_A_CY;
  wire [0:0] CLBLM_L_X10Y144_SLICE_X12Y144_A_XOR;
  wire [0:0] CLBLM_L_X10Y144_SLICE_X12Y144_B;
  wire [0:0] CLBLM_L_X10Y144_SLICE_X12Y144_B1;
  wire [0:0] CLBLM_L_X10Y144_SLICE_X12Y144_B2;
  wire [0:0] CLBLM_L_X10Y144_SLICE_X12Y144_B3;
  wire [0:0] CLBLM_L_X10Y144_SLICE_X12Y144_B4;
  wire [0:0] CLBLM_L_X10Y144_SLICE_X12Y144_B5;
  wire [0:0] CLBLM_L_X10Y144_SLICE_X12Y144_B6;
  wire [0:0] CLBLM_L_X10Y144_SLICE_X12Y144_BMUX;
  wire [0:0] CLBLM_L_X10Y144_SLICE_X12Y144_BO5;
  wire [0:0] CLBLM_L_X10Y144_SLICE_X12Y144_BO6;
  wire [0:0] CLBLM_L_X10Y144_SLICE_X12Y144_B_CY;
  wire [0:0] CLBLM_L_X10Y144_SLICE_X12Y144_B_XOR;
  wire [0:0] CLBLM_L_X10Y144_SLICE_X12Y144_C;
  wire [0:0] CLBLM_L_X10Y144_SLICE_X12Y144_C1;
  wire [0:0] CLBLM_L_X10Y144_SLICE_X12Y144_C2;
  wire [0:0] CLBLM_L_X10Y144_SLICE_X12Y144_C3;
  wire [0:0] CLBLM_L_X10Y144_SLICE_X12Y144_C4;
  wire [0:0] CLBLM_L_X10Y144_SLICE_X12Y144_C5;
  wire [0:0] CLBLM_L_X10Y144_SLICE_X12Y144_C6;
  wire [0:0] CLBLM_L_X10Y144_SLICE_X12Y144_CE;
  wire [0:0] CLBLM_L_X10Y144_SLICE_X12Y144_CLK;
  wire [0:0] CLBLM_L_X10Y144_SLICE_X12Y144_CO5;
  wire [0:0] CLBLM_L_X10Y144_SLICE_X12Y144_CO6;
  wire [0:0] CLBLM_L_X10Y144_SLICE_X12Y144_C_CY;
  wire [0:0] CLBLM_L_X10Y144_SLICE_X12Y144_C_XOR;
  wire [0:0] CLBLM_L_X10Y144_SLICE_X12Y144_D;
  wire [0:0] CLBLM_L_X10Y144_SLICE_X12Y144_D1;
  wire [0:0] CLBLM_L_X10Y144_SLICE_X12Y144_D2;
  wire [0:0] CLBLM_L_X10Y144_SLICE_X12Y144_D3;
  wire [0:0] CLBLM_L_X10Y144_SLICE_X12Y144_D4;
  wire [0:0] CLBLM_L_X10Y144_SLICE_X12Y144_D5;
  wire [0:0] CLBLM_L_X10Y144_SLICE_X12Y144_D6;
  wire [0:0] CLBLM_L_X10Y144_SLICE_X12Y144_DO5;
  wire [0:0] CLBLM_L_X10Y144_SLICE_X12Y144_DO6;
  wire [0:0] CLBLM_L_X10Y144_SLICE_X12Y144_D_CY;
  wire [0:0] CLBLM_L_X10Y144_SLICE_X12Y144_D_XOR;
  wire [0:0] CLBLM_L_X10Y144_SLICE_X13Y144_A;
  wire [0:0] CLBLM_L_X10Y144_SLICE_X13Y144_A1;
  wire [0:0] CLBLM_L_X10Y144_SLICE_X13Y144_A2;
  wire [0:0] CLBLM_L_X10Y144_SLICE_X13Y144_A3;
  wire [0:0] CLBLM_L_X10Y144_SLICE_X13Y144_A4;
  wire [0:0] CLBLM_L_X10Y144_SLICE_X13Y144_A5;
  wire [0:0] CLBLM_L_X10Y144_SLICE_X13Y144_A5Q;
  wire [0:0] CLBLM_L_X10Y144_SLICE_X13Y144_A6;
  wire [0:0] CLBLM_L_X10Y144_SLICE_X13Y144_AMUX;
  wire [0:0] CLBLM_L_X10Y144_SLICE_X13Y144_AO5;
  wire [0:0] CLBLM_L_X10Y144_SLICE_X13Y144_AO6;
  wire [0:0] CLBLM_L_X10Y144_SLICE_X13Y144_AQ;
  wire [0:0] CLBLM_L_X10Y144_SLICE_X13Y144_AX;
  wire [0:0] CLBLM_L_X10Y144_SLICE_X13Y144_A_CY;
  wire [0:0] CLBLM_L_X10Y144_SLICE_X13Y144_A_XOR;
  wire [0:0] CLBLM_L_X10Y144_SLICE_X13Y144_B;
  wire [0:0] CLBLM_L_X10Y144_SLICE_X13Y144_B1;
  wire [0:0] CLBLM_L_X10Y144_SLICE_X13Y144_B2;
  wire [0:0] CLBLM_L_X10Y144_SLICE_X13Y144_B3;
  wire [0:0] CLBLM_L_X10Y144_SLICE_X13Y144_B4;
  wire [0:0] CLBLM_L_X10Y144_SLICE_X13Y144_B5;
  wire [0:0] CLBLM_L_X10Y144_SLICE_X13Y144_B6;
  wire [0:0] CLBLM_L_X10Y144_SLICE_X13Y144_BO5;
  wire [0:0] CLBLM_L_X10Y144_SLICE_X13Y144_BO6;
  wire [0:0] CLBLM_L_X10Y144_SLICE_X13Y144_BQ;
  wire [0:0] CLBLM_L_X10Y144_SLICE_X13Y144_B_CY;
  wire [0:0] CLBLM_L_X10Y144_SLICE_X13Y144_B_XOR;
  wire [0:0] CLBLM_L_X10Y144_SLICE_X13Y144_C;
  wire [0:0] CLBLM_L_X10Y144_SLICE_X13Y144_C1;
  wire [0:0] CLBLM_L_X10Y144_SLICE_X13Y144_C2;
  wire [0:0] CLBLM_L_X10Y144_SLICE_X13Y144_C3;
  wire [0:0] CLBLM_L_X10Y144_SLICE_X13Y144_C4;
  wire [0:0] CLBLM_L_X10Y144_SLICE_X13Y144_C5;
  wire [0:0] CLBLM_L_X10Y144_SLICE_X13Y144_C5Q;
  wire [0:0] CLBLM_L_X10Y144_SLICE_X13Y144_C6;
  wire [0:0] CLBLM_L_X10Y144_SLICE_X13Y144_CLK;
  wire [0:0] CLBLM_L_X10Y144_SLICE_X13Y144_CMUX;
  wire [0:0] CLBLM_L_X10Y144_SLICE_X13Y144_CO5;
  wire [0:0] CLBLM_L_X10Y144_SLICE_X13Y144_CO6;
  wire [0:0] CLBLM_L_X10Y144_SLICE_X13Y144_CQ;
  wire [0:0] CLBLM_L_X10Y144_SLICE_X13Y144_C_CY;
  wire [0:0] CLBLM_L_X10Y144_SLICE_X13Y144_C_XOR;
  wire [0:0] CLBLM_L_X10Y144_SLICE_X13Y144_D;
  wire [0:0] CLBLM_L_X10Y144_SLICE_X13Y144_D1;
  wire [0:0] CLBLM_L_X10Y144_SLICE_X13Y144_D2;
  wire [0:0] CLBLM_L_X10Y144_SLICE_X13Y144_D3;
  wire [0:0] CLBLM_L_X10Y144_SLICE_X13Y144_D4;
  wire [0:0] CLBLM_L_X10Y144_SLICE_X13Y144_D5;
  wire [0:0] CLBLM_L_X10Y144_SLICE_X13Y144_D6;
  wire [0:0] CLBLM_L_X10Y144_SLICE_X13Y144_DO5;
  wire [0:0] CLBLM_L_X10Y144_SLICE_X13Y144_DO6;
  wire [0:0] CLBLM_L_X10Y144_SLICE_X13Y144_DQ;
  wire [0:0] CLBLM_L_X10Y144_SLICE_X13Y144_D_CY;
  wire [0:0] CLBLM_L_X10Y144_SLICE_X13Y144_D_XOR;
  wire [0:0] CLBLM_L_X10Y145_SLICE_X12Y145_A;
  wire [0:0] CLBLM_L_X10Y145_SLICE_X12Y145_A1;
  wire [0:0] CLBLM_L_X10Y145_SLICE_X12Y145_A2;
  wire [0:0] CLBLM_L_X10Y145_SLICE_X12Y145_A3;
  wire [0:0] CLBLM_L_X10Y145_SLICE_X12Y145_A4;
  wire [0:0] CLBLM_L_X10Y145_SLICE_X12Y145_A5;
  wire [0:0] CLBLM_L_X10Y145_SLICE_X12Y145_A5Q;
  wire [0:0] CLBLM_L_X10Y145_SLICE_X12Y145_A6;
  wire [0:0] CLBLM_L_X10Y145_SLICE_X12Y145_AMUX;
  wire [0:0] CLBLM_L_X10Y145_SLICE_X12Y145_AO5;
  wire [0:0] CLBLM_L_X10Y145_SLICE_X12Y145_AO6;
  wire [0:0] CLBLM_L_X10Y145_SLICE_X12Y145_AQ;
  wire [0:0] CLBLM_L_X10Y145_SLICE_X12Y145_A_CY;
  wire [0:0] CLBLM_L_X10Y145_SLICE_X12Y145_A_XOR;
  wire [0:0] CLBLM_L_X10Y145_SLICE_X12Y145_B;
  wire [0:0] CLBLM_L_X10Y145_SLICE_X12Y145_B1;
  wire [0:0] CLBLM_L_X10Y145_SLICE_X12Y145_B2;
  wire [0:0] CLBLM_L_X10Y145_SLICE_X12Y145_B3;
  wire [0:0] CLBLM_L_X10Y145_SLICE_X12Y145_B4;
  wire [0:0] CLBLM_L_X10Y145_SLICE_X12Y145_B5;
  wire [0:0] CLBLM_L_X10Y145_SLICE_X12Y145_B6;
  wire [0:0] CLBLM_L_X10Y145_SLICE_X12Y145_BO5;
  wire [0:0] CLBLM_L_X10Y145_SLICE_X12Y145_BO6;
  wire [0:0] CLBLM_L_X10Y145_SLICE_X12Y145_BQ;
  wire [0:0] CLBLM_L_X10Y145_SLICE_X12Y145_B_CY;
  wire [0:0] CLBLM_L_X10Y145_SLICE_X12Y145_B_XOR;
  wire [0:0] CLBLM_L_X10Y145_SLICE_X12Y145_C;
  wire [0:0] CLBLM_L_X10Y145_SLICE_X12Y145_C1;
  wire [0:0] CLBLM_L_X10Y145_SLICE_X12Y145_C2;
  wire [0:0] CLBLM_L_X10Y145_SLICE_X12Y145_C3;
  wire [0:0] CLBLM_L_X10Y145_SLICE_X12Y145_C4;
  wire [0:0] CLBLM_L_X10Y145_SLICE_X12Y145_C5;
  wire [0:0] CLBLM_L_X10Y145_SLICE_X12Y145_C6;
  wire [0:0] CLBLM_L_X10Y145_SLICE_X12Y145_CLK;
  wire [0:0] CLBLM_L_X10Y145_SLICE_X12Y145_CO5;
  wire [0:0] CLBLM_L_X10Y145_SLICE_X12Y145_CO6;
  wire [0:0] CLBLM_L_X10Y145_SLICE_X12Y145_C_CY;
  wire [0:0] CLBLM_L_X10Y145_SLICE_X12Y145_C_XOR;
  wire [0:0] CLBLM_L_X10Y145_SLICE_X12Y145_D;
  wire [0:0] CLBLM_L_X10Y145_SLICE_X12Y145_D1;
  wire [0:0] CLBLM_L_X10Y145_SLICE_X12Y145_D2;
  wire [0:0] CLBLM_L_X10Y145_SLICE_X12Y145_D3;
  wire [0:0] CLBLM_L_X10Y145_SLICE_X12Y145_D4;
  wire [0:0] CLBLM_L_X10Y145_SLICE_X12Y145_D5;
  wire [0:0] CLBLM_L_X10Y145_SLICE_X12Y145_D6;
  wire [0:0] CLBLM_L_X10Y145_SLICE_X12Y145_DO5;
  wire [0:0] CLBLM_L_X10Y145_SLICE_X12Y145_DO6;
  wire [0:0] CLBLM_L_X10Y145_SLICE_X12Y145_D_CY;
  wire [0:0] CLBLM_L_X10Y145_SLICE_X12Y145_D_XOR;
  wire [0:0] CLBLM_L_X10Y145_SLICE_X13Y145_A;
  wire [0:0] CLBLM_L_X10Y145_SLICE_X13Y145_A1;
  wire [0:0] CLBLM_L_X10Y145_SLICE_X13Y145_A2;
  wire [0:0] CLBLM_L_X10Y145_SLICE_X13Y145_A3;
  wire [0:0] CLBLM_L_X10Y145_SLICE_X13Y145_A4;
  wire [0:0] CLBLM_L_X10Y145_SLICE_X13Y145_A5;
  wire [0:0] CLBLM_L_X10Y145_SLICE_X13Y145_A6;
  wire [0:0] CLBLM_L_X10Y145_SLICE_X13Y145_AO5;
  wire [0:0] CLBLM_L_X10Y145_SLICE_X13Y145_AO6;
  wire [0:0] CLBLM_L_X10Y145_SLICE_X13Y145_AQ;
  wire [0:0] CLBLM_L_X10Y145_SLICE_X13Y145_A_CY;
  wire [0:0] CLBLM_L_X10Y145_SLICE_X13Y145_A_XOR;
  wire [0:0] CLBLM_L_X10Y145_SLICE_X13Y145_B;
  wire [0:0] CLBLM_L_X10Y145_SLICE_X13Y145_B1;
  wire [0:0] CLBLM_L_X10Y145_SLICE_X13Y145_B2;
  wire [0:0] CLBLM_L_X10Y145_SLICE_X13Y145_B3;
  wire [0:0] CLBLM_L_X10Y145_SLICE_X13Y145_B4;
  wire [0:0] CLBLM_L_X10Y145_SLICE_X13Y145_B5;
  wire [0:0] CLBLM_L_X10Y145_SLICE_X13Y145_B6;
  wire [0:0] CLBLM_L_X10Y145_SLICE_X13Y145_BO5;
  wire [0:0] CLBLM_L_X10Y145_SLICE_X13Y145_BO6;
  wire [0:0] CLBLM_L_X10Y145_SLICE_X13Y145_B_CY;
  wire [0:0] CLBLM_L_X10Y145_SLICE_X13Y145_B_XOR;
  wire [0:0] CLBLM_L_X10Y145_SLICE_X13Y145_C;
  wire [0:0] CLBLM_L_X10Y145_SLICE_X13Y145_C1;
  wire [0:0] CLBLM_L_X10Y145_SLICE_X13Y145_C2;
  wire [0:0] CLBLM_L_X10Y145_SLICE_X13Y145_C3;
  wire [0:0] CLBLM_L_X10Y145_SLICE_X13Y145_C4;
  wire [0:0] CLBLM_L_X10Y145_SLICE_X13Y145_C5;
  wire [0:0] CLBLM_L_X10Y145_SLICE_X13Y145_C6;
  wire [0:0] CLBLM_L_X10Y145_SLICE_X13Y145_CLK;
  wire [0:0] CLBLM_L_X10Y145_SLICE_X13Y145_CO5;
  wire [0:0] CLBLM_L_X10Y145_SLICE_X13Y145_CO6;
  wire [0:0] CLBLM_L_X10Y145_SLICE_X13Y145_C_CY;
  wire [0:0] CLBLM_L_X10Y145_SLICE_X13Y145_C_XOR;
  wire [0:0] CLBLM_L_X10Y145_SLICE_X13Y145_D;
  wire [0:0] CLBLM_L_X10Y145_SLICE_X13Y145_D1;
  wire [0:0] CLBLM_L_X10Y145_SLICE_X13Y145_D2;
  wire [0:0] CLBLM_L_X10Y145_SLICE_X13Y145_D3;
  wire [0:0] CLBLM_L_X10Y145_SLICE_X13Y145_D4;
  wire [0:0] CLBLM_L_X10Y145_SLICE_X13Y145_D5;
  wire [0:0] CLBLM_L_X10Y145_SLICE_X13Y145_D6;
  wire [0:0] CLBLM_L_X10Y145_SLICE_X13Y145_DO5;
  wire [0:0] CLBLM_L_X10Y145_SLICE_X13Y145_DO6;
  wire [0:0] CLBLM_L_X10Y145_SLICE_X13Y145_D_CY;
  wire [0:0] CLBLM_L_X10Y145_SLICE_X13Y145_D_XOR;
  wire [0:0] CLBLM_L_X10Y146_SLICE_X12Y146_A;
  wire [0:0] CLBLM_L_X10Y146_SLICE_X12Y146_A1;
  wire [0:0] CLBLM_L_X10Y146_SLICE_X12Y146_A2;
  wire [0:0] CLBLM_L_X10Y146_SLICE_X12Y146_A3;
  wire [0:0] CLBLM_L_X10Y146_SLICE_X12Y146_A4;
  wire [0:0] CLBLM_L_X10Y146_SLICE_X12Y146_A5;
  wire [0:0] CLBLM_L_X10Y146_SLICE_X12Y146_A6;
  wire [0:0] CLBLM_L_X10Y146_SLICE_X12Y146_AO5;
  wire [0:0] CLBLM_L_X10Y146_SLICE_X12Y146_AO6;
  wire [0:0] CLBLM_L_X10Y146_SLICE_X12Y146_AQ;
  wire [0:0] CLBLM_L_X10Y146_SLICE_X12Y146_A_CY;
  wire [0:0] CLBLM_L_X10Y146_SLICE_X12Y146_A_XOR;
  wire [0:0] CLBLM_L_X10Y146_SLICE_X12Y146_B;
  wire [0:0] CLBLM_L_X10Y146_SLICE_X12Y146_B1;
  wire [0:0] CLBLM_L_X10Y146_SLICE_X12Y146_B2;
  wire [0:0] CLBLM_L_X10Y146_SLICE_X12Y146_B3;
  wire [0:0] CLBLM_L_X10Y146_SLICE_X12Y146_B4;
  wire [0:0] CLBLM_L_X10Y146_SLICE_X12Y146_B5;
  wire [0:0] CLBLM_L_X10Y146_SLICE_X12Y146_B6;
  wire [0:0] CLBLM_L_X10Y146_SLICE_X12Y146_BO5;
  wire [0:0] CLBLM_L_X10Y146_SLICE_X12Y146_BO6;
  wire [0:0] CLBLM_L_X10Y146_SLICE_X12Y146_BQ;
  wire [0:0] CLBLM_L_X10Y146_SLICE_X12Y146_B_CY;
  wire [0:0] CLBLM_L_X10Y146_SLICE_X12Y146_B_XOR;
  wire [0:0] CLBLM_L_X10Y146_SLICE_X12Y146_C;
  wire [0:0] CLBLM_L_X10Y146_SLICE_X12Y146_C1;
  wire [0:0] CLBLM_L_X10Y146_SLICE_X12Y146_C2;
  wire [0:0] CLBLM_L_X10Y146_SLICE_X12Y146_C3;
  wire [0:0] CLBLM_L_X10Y146_SLICE_X12Y146_C4;
  wire [0:0] CLBLM_L_X10Y146_SLICE_X12Y146_C5;
  wire [0:0] CLBLM_L_X10Y146_SLICE_X12Y146_C6;
  wire [0:0] CLBLM_L_X10Y146_SLICE_X12Y146_CLK;
  wire [0:0] CLBLM_L_X10Y146_SLICE_X12Y146_CO5;
  wire [0:0] CLBLM_L_X10Y146_SLICE_X12Y146_CO6;
  wire [0:0] CLBLM_L_X10Y146_SLICE_X12Y146_CQ;
  wire [0:0] CLBLM_L_X10Y146_SLICE_X12Y146_C_CY;
  wire [0:0] CLBLM_L_X10Y146_SLICE_X12Y146_C_XOR;
  wire [0:0] CLBLM_L_X10Y146_SLICE_X12Y146_D;
  wire [0:0] CLBLM_L_X10Y146_SLICE_X12Y146_D1;
  wire [0:0] CLBLM_L_X10Y146_SLICE_X12Y146_D2;
  wire [0:0] CLBLM_L_X10Y146_SLICE_X12Y146_D3;
  wire [0:0] CLBLM_L_X10Y146_SLICE_X12Y146_D4;
  wire [0:0] CLBLM_L_X10Y146_SLICE_X12Y146_D5;
  wire [0:0] CLBLM_L_X10Y146_SLICE_X12Y146_D5Q;
  wire [0:0] CLBLM_L_X10Y146_SLICE_X12Y146_D6;
  wire [0:0] CLBLM_L_X10Y146_SLICE_X12Y146_DMUX;
  wire [0:0] CLBLM_L_X10Y146_SLICE_X12Y146_DO5;
  wire [0:0] CLBLM_L_X10Y146_SLICE_X12Y146_DO6;
  wire [0:0] CLBLM_L_X10Y146_SLICE_X12Y146_DQ;
  wire [0:0] CLBLM_L_X10Y146_SLICE_X12Y146_D_CY;
  wire [0:0] CLBLM_L_X10Y146_SLICE_X12Y146_D_XOR;
  wire [0:0] CLBLM_L_X10Y146_SLICE_X13Y146_A;
  wire [0:0] CLBLM_L_X10Y146_SLICE_X13Y146_A1;
  wire [0:0] CLBLM_L_X10Y146_SLICE_X13Y146_A2;
  wire [0:0] CLBLM_L_X10Y146_SLICE_X13Y146_A3;
  wire [0:0] CLBLM_L_X10Y146_SLICE_X13Y146_A4;
  wire [0:0] CLBLM_L_X10Y146_SLICE_X13Y146_A5;
  wire [0:0] CLBLM_L_X10Y146_SLICE_X13Y146_A6;
  wire [0:0] CLBLM_L_X10Y146_SLICE_X13Y146_AO5;
  wire [0:0] CLBLM_L_X10Y146_SLICE_X13Y146_AO6;
  wire [0:0] CLBLM_L_X10Y146_SLICE_X13Y146_AQ;
  wire [0:0] CLBLM_L_X10Y146_SLICE_X13Y146_A_CY;
  wire [0:0] CLBLM_L_X10Y146_SLICE_X13Y146_A_XOR;
  wire [0:0] CLBLM_L_X10Y146_SLICE_X13Y146_B;
  wire [0:0] CLBLM_L_X10Y146_SLICE_X13Y146_B1;
  wire [0:0] CLBLM_L_X10Y146_SLICE_X13Y146_B2;
  wire [0:0] CLBLM_L_X10Y146_SLICE_X13Y146_B3;
  wire [0:0] CLBLM_L_X10Y146_SLICE_X13Y146_B4;
  wire [0:0] CLBLM_L_X10Y146_SLICE_X13Y146_B5;
  wire [0:0] CLBLM_L_X10Y146_SLICE_X13Y146_B6;
  wire [0:0] CLBLM_L_X10Y146_SLICE_X13Y146_BO5;
  wire [0:0] CLBLM_L_X10Y146_SLICE_X13Y146_BO6;
  wire [0:0] CLBLM_L_X10Y146_SLICE_X13Y146_BQ;
  wire [0:0] CLBLM_L_X10Y146_SLICE_X13Y146_B_CY;
  wire [0:0] CLBLM_L_X10Y146_SLICE_X13Y146_B_XOR;
  wire [0:0] CLBLM_L_X10Y146_SLICE_X13Y146_C;
  wire [0:0] CLBLM_L_X10Y146_SLICE_X13Y146_C1;
  wire [0:0] CLBLM_L_X10Y146_SLICE_X13Y146_C2;
  wire [0:0] CLBLM_L_X10Y146_SLICE_X13Y146_C3;
  wire [0:0] CLBLM_L_X10Y146_SLICE_X13Y146_C4;
  wire [0:0] CLBLM_L_X10Y146_SLICE_X13Y146_C5;
  wire [0:0] CLBLM_L_X10Y146_SLICE_X13Y146_C6;
  wire [0:0] CLBLM_L_X10Y146_SLICE_X13Y146_CLK;
  wire [0:0] CLBLM_L_X10Y146_SLICE_X13Y146_CO5;
  wire [0:0] CLBLM_L_X10Y146_SLICE_X13Y146_CO6;
  wire [0:0] CLBLM_L_X10Y146_SLICE_X13Y146_CQ;
  wire [0:0] CLBLM_L_X10Y146_SLICE_X13Y146_C_CY;
  wire [0:0] CLBLM_L_X10Y146_SLICE_X13Y146_C_XOR;
  wire [0:0] CLBLM_L_X10Y146_SLICE_X13Y146_D;
  wire [0:0] CLBLM_L_X10Y146_SLICE_X13Y146_D1;
  wire [0:0] CLBLM_L_X10Y146_SLICE_X13Y146_D2;
  wire [0:0] CLBLM_L_X10Y146_SLICE_X13Y146_D3;
  wire [0:0] CLBLM_L_X10Y146_SLICE_X13Y146_D4;
  wire [0:0] CLBLM_L_X10Y146_SLICE_X13Y146_D5;
  wire [0:0] CLBLM_L_X10Y146_SLICE_X13Y146_D6;
  wire [0:0] CLBLM_L_X10Y146_SLICE_X13Y146_DMUX;
  wire [0:0] CLBLM_L_X10Y146_SLICE_X13Y146_DO5;
  wire [0:0] CLBLM_L_X10Y146_SLICE_X13Y146_DO6;
  wire [0:0] CLBLM_L_X10Y146_SLICE_X13Y146_D_CY;
  wire [0:0] CLBLM_L_X10Y146_SLICE_X13Y146_D_XOR;
  wire [0:0] CLBLM_L_X10Y147_SLICE_X12Y147_A;
  wire [0:0] CLBLM_L_X10Y147_SLICE_X12Y147_A1;
  wire [0:0] CLBLM_L_X10Y147_SLICE_X12Y147_A2;
  wire [0:0] CLBLM_L_X10Y147_SLICE_X12Y147_A3;
  wire [0:0] CLBLM_L_X10Y147_SLICE_X12Y147_A4;
  wire [0:0] CLBLM_L_X10Y147_SLICE_X12Y147_A5;
  wire [0:0] CLBLM_L_X10Y147_SLICE_X12Y147_A6;
  wire [0:0] CLBLM_L_X10Y147_SLICE_X12Y147_AMUX;
  wire [0:0] CLBLM_L_X10Y147_SLICE_X12Y147_AO5;
  wire [0:0] CLBLM_L_X10Y147_SLICE_X12Y147_AO6;
  wire [0:0] CLBLM_L_X10Y147_SLICE_X12Y147_AQ;
  wire [0:0] CLBLM_L_X10Y147_SLICE_X12Y147_AX;
  wire [0:0] CLBLM_L_X10Y147_SLICE_X12Y147_A_CY;
  wire [0:0] CLBLM_L_X10Y147_SLICE_X12Y147_A_XOR;
  wire [0:0] CLBLM_L_X10Y147_SLICE_X12Y147_B;
  wire [0:0] CLBLM_L_X10Y147_SLICE_X12Y147_B1;
  wire [0:0] CLBLM_L_X10Y147_SLICE_X12Y147_B2;
  wire [0:0] CLBLM_L_X10Y147_SLICE_X12Y147_B3;
  wire [0:0] CLBLM_L_X10Y147_SLICE_X12Y147_B4;
  wire [0:0] CLBLM_L_X10Y147_SLICE_X12Y147_B5;
  wire [0:0] CLBLM_L_X10Y147_SLICE_X12Y147_B6;
  wire [0:0] CLBLM_L_X10Y147_SLICE_X12Y147_BMUX;
  wire [0:0] CLBLM_L_X10Y147_SLICE_X12Y147_BO5;
  wire [0:0] CLBLM_L_X10Y147_SLICE_X12Y147_BO6;
  wire [0:0] CLBLM_L_X10Y147_SLICE_X12Y147_BQ;
  wire [0:0] CLBLM_L_X10Y147_SLICE_X12Y147_BX;
  wire [0:0] CLBLM_L_X10Y147_SLICE_X12Y147_B_CY;
  wire [0:0] CLBLM_L_X10Y147_SLICE_X12Y147_B_XOR;
  wire [0:0] CLBLM_L_X10Y147_SLICE_X12Y147_C;
  wire [0:0] CLBLM_L_X10Y147_SLICE_X12Y147_C1;
  wire [0:0] CLBLM_L_X10Y147_SLICE_X12Y147_C2;
  wire [0:0] CLBLM_L_X10Y147_SLICE_X12Y147_C3;
  wire [0:0] CLBLM_L_X10Y147_SLICE_X12Y147_C4;
  wire [0:0] CLBLM_L_X10Y147_SLICE_X12Y147_C5;
  wire [0:0] CLBLM_L_X10Y147_SLICE_X12Y147_C6;
  wire [0:0] CLBLM_L_X10Y147_SLICE_X12Y147_CE;
  wire [0:0] CLBLM_L_X10Y147_SLICE_X12Y147_CLK;
  wire [0:0] CLBLM_L_X10Y147_SLICE_X12Y147_CO5;
  wire [0:0] CLBLM_L_X10Y147_SLICE_X12Y147_CO6;
  wire [0:0] CLBLM_L_X10Y147_SLICE_X12Y147_CQ;
  wire [0:0] CLBLM_L_X10Y147_SLICE_X12Y147_CX;
  wire [0:0] CLBLM_L_X10Y147_SLICE_X12Y147_C_CY;
  wire [0:0] CLBLM_L_X10Y147_SLICE_X12Y147_C_XOR;
  wire [0:0] CLBLM_L_X10Y147_SLICE_X12Y147_D;
  wire [0:0] CLBLM_L_X10Y147_SLICE_X12Y147_D1;
  wire [0:0] CLBLM_L_X10Y147_SLICE_X12Y147_D2;
  wire [0:0] CLBLM_L_X10Y147_SLICE_X12Y147_D3;
  wire [0:0] CLBLM_L_X10Y147_SLICE_X12Y147_D4;
  wire [0:0] CLBLM_L_X10Y147_SLICE_X12Y147_D5;
  wire [0:0] CLBLM_L_X10Y147_SLICE_X12Y147_D6;
  wire [0:0] CLBLM_L_X10Y147_SLICE_X12Y147_DO5;
  wire [0:0] CLBLM_L_X10Y147_SLICE_X12Y147_DO6;
  wire [0:0] CLBLM_L_X10Y147_SLICE_X12Y147_D_CY;
  wire [0:0] CLBLM_L_X10Y147_SLICE_X12Y147_D_XOR;
  wire [0:0] CLBLM_L_X10Y147_SLICE_X13Y147_A;
  wire [0:0] CLBLM_L_X10Y147_SLICE_X13Y147_A1;
  wire [0:0] CLBLM_L_X10Y147_SLICE_X13Y147_A2;
  wire [0:0] CLBLM_L_X10Y147_SLICE_X13Y147_A3;
  wire [0:0] CLBLM_L_X10Y147_SLICE_X13Y147_A4;
  wire [0:0] CLBLM_L_X10Y147_SLICE_X13Y147_A5;
  wire [0:0] CLBLM_L_X10Y147_SLICE_X13Y147_A6;
  wire [0:0] CLBLM_L_X10Y147_SLICE_X13Y147_AO5;
  wire [0:0] CLBLM_L_X10Y147_SLICE_X13Y147_AO6;
  wire [0:0] CLBLM_L_X10Y147_SLICE_X13Y147_AQ;
  wire [0:0] CLBLM_L_X10Y147_SLICE_X13Y147_A_CY;
  wire [0:0] CLBLM_L_X10Y147_SLICE_X13Y147_A_XOR;
  wire [0:0] CLBLM_L_X10Y147_SLICE_X13Y147_B;
  wire [0:0] CLBLM_L_X10Y147_SLICE_X13Y147_B1;
  wire [0:0] CLBLM_L_X10Y147_SLICE_X13Y147_B2;
  wire [0:0] CLBLM_L_X10Y147_SLICE_X13Y147_B3;
  wire [0:0] CLBLM_L_X10Y147_SLICE_X13Y147_B4;
  wire [0:0] CLBLM_L_X10Y147_SLICE_X13Y147_B5;
  wire [0:0] CLBLM_L_X10Y147_SLICE_X13Y147_B6;
  wire [0:0] CLBLM_L_X10Y147_SLICE_X13Y147_BO5;
  wire [0:0] CLBLM_L_X10Y147_SLICE_X13Y147_BO6;
  wire [0:0] CLBLM_L_X10Y147_SLICE_X13Y147_B_CY;
  wire [0:0] CLBLM_L_X10Y147_SLICE_X13Y147_B_XOR;
  wire [0:0] CLBLM_L_X10Y147_SLICE_X13Y147_C;
  wire [0:0] CLBLM_L_X10Y147_SLICE_X13Y147_C1;
  wire [0:0] CLBLM_L_X10Y147_SLICE_X13Y147_C2;
  wire [0:0] CLBLM_L_X10Y147_SLICE_X13Y147_C3;
  wire [0:0] CLBLM_L_X10Y147_SLICE_X13Y147_C4;
  wire [0:0] CLBLM_L_X10Y147_SLICE_X13Y147_C5;
  wire [0:0] CLBLM_L_X10Y147_SLICE_X13Y147_C6;
  wire [0:0] CLBLM_L_X10Y147_SLICE_X13Y147_CLK;
  wire [0:0] CLBLM_L_X10Y147_SLICE_X13Y147_CO5;
  wire [0:0] CLBLM_L_X10Y147_SLICE_X13Y147_CO6;
  wire [0:0] CLBLM_L_X10Y147_SLICE_X13Y147_C_CY;
  wire [0:0] CLBLM_L_X10Y147_SLICE_X13Y147_C_XOR;
  wire [0:0] CLBLM_L_X10Y147_SLICE_X13Y147_D;
  wire [0:0] CLBLM_L_X10Y147_SLICE_X13Y147_D1;
  wire [0:0] CLBLM_L_X10Y147_SLICE_X13Y147_D2;
  wire [0:0] CLBLM_L_X10Y147_SLICE_X13Y147_D3;
  wire [0:0] CLBLM_L_X10Y147_SLICE_X13Y147_D4;
  wire [0:0] CLBLM_L_X10Y147_SLICE_X13Y147_D5;
  wire [0:0] CLBLM_L_X10Y147_SLICE_X13Y147_D6;
  wire [0:0] CLBLM_L_X10Y147_SLICE_X13Y147_DO5;
  wire [0:0] CLBLM_L_X10Y147_SLICE_X13Y147_DO6;
  wire [0:0] CLBLM_L_X10Y147_SLICE_X13Y147_D_CY;
  wire [0:0] CLBLM_L_X10Y147_SLICE_X13Y147_D_XOR;
  wire [0:0] CLBLM_L_X10Y148_SLICE_X12Y148_A;
  wire [0:0] CLBLM_L_X10Y148_SLICE_X12Y148_A1;
  wire [0:0] CLBLM_L_X10Y148_SLICE_X12Y148_A2;
  wire [0:0] CLBLM_L_X10Y148_SLICE_X12Y148_A3;
  wire [0:0] CLBLM_L_X10Y148_SLICE_X12Y148_A4;
  wire [0:0] CLBLM_L_X10Y148_SLICE_X12Y148_A5;
  wire [0:0] CLBLM_L_X10Y148_SLICE_X12Y148_A6;
  wire [0:0] CLBLM_L_X10Y148_SLICE_X12Y148_AMUX;
  wire [0:0] CLBLM_L_X10Y148_SLICE_X12Y148_AO5;
  wire [0:0] CLBLM_L_X10Y148_SLICE_X12Y148_AO6;
  wire [0:0] CLBLM_L_X10Y148_SLICE_X12Y148_AQ;
  wire [0:0] CLBLM_L_X10Y148_SLICE_X12Y148_AX;
  wire [0:0] CLBLM_L_X10Y148_SLICE_X12Y148_A_CY;
  wire [0:0] CLBLM_L_X10Y148_SLICE_X12Y148_A_XOR;
  wire [0:0] CLBLM_L_X10Y148_SLICE_X12Y148_B;
  wire [0:0] CLBLM_L_X10Y148_SLICE_X12Y148_B1;
  wire [0:0] CLBLM_L_X10Y148_SLICE_X12Y148_B2;
  wire [0:0] CLBLM_L_X10Y148_SLICE_X12Y148_B3;
  wire [0:0] CLBLM_L_X10Y148_SLICE_X12Y148_B4;
  wire [0:0] CLBLM_L_X10Y148_SLICE_X12Y148_B5;
  wire [0:0] CLBLM_L_X10Y148_SLICE_X12Y148_B6;
  wire [0:0] CLBLM_L_X10Y148_SLICE_X12Y148_BO5;
  wire [0:0] CLBLM_L_X10Y148_SLICE_X12Y148_BO6;
  wire [0:0] CLBLM_L_X10Y148_SLICE_X12Y148_B_CY;
  wire [0:0] CLBLM_L_X10Y148_SLICE_X12Y148_B_XOR;
  wire [0:0] CLBLM_L_X10Y148_SLICE_X12Y148_C;
  wire [0:0] CLBLM_L_X10Y148_SLICE_X12Y148_C1;
  wire [0:0] CLBLM_L_X10Y148_SLICE_X12Y148_C2;
  wire [0:0] CLBLM_L_X10Y148_SLICE_X12Y148_C3;
  wire [0:0] CLBLM_L_X10Y148_SLICE_X12Y148_C4;
  wire [0:0] CLBLM_L_X10Y148_SLICE_X12Y148_C5;
  wire [0:0] CLBLM_L_X10Y148_SLICE_X12Y148_C6;
  wire [0:0] CLBLM_L_X10Y148_SLICE_X12Y148_CLK;
  wire [0:0] CLBLM_L_X10Y148_SLICE_X12Y148_CO5;
  wire [0:0] CLBLM_L_X10Y148_SLICE_X12Y148_CO6;
  wire [0:0] CLBLM_L_X10Y148_SLICE_X12Y148_C_CY;
  wire [0:0] CLBLM_L_X10Y148_SLICE_X12Y148_C_XOR;
  wire [0:0] CLBLM_L_X10Y148_SLICE_X12Y148_D;
  wire [0:0] CLBLM_L_X10Y148_SLICE_X12Y148_D1;
  wire [0:0] CLBLM_L_X10Y148_SLICE_X12Y148_D2;
  wire [0:0] CLBLM_L_X10Y148_SLICE_X12Y148_D3;
  wire [0:0] CLBLM_L_X10Y148_SLICE_X12Y148_D4;
  wire [0:0] CLBLM_L_X10Y148_SLICE_X12Y148_D5;
  wire [0:0] CLBLM_L_X10Y148_SLICE_X12Y148_D6;
  wire [0:0] CLBLM_L_X10Y148_SLICE_X12Y148_DO5;
  wire [0:0] CLBLM_L_X10Y148_SLICE_X12Y148_DO6;
  wire [0:0] CLBLM_L_X10Y148_SLICE_X12Y148_D_CY;
  wire [0:0] CLBLM_L_X10Y148_SLICE_X12Y148_D_XOR;
  wire [0:0] CLBLM_L_X10Y148_SLICE_X13Y148_A;
  wire [0:0] CLBLM_L_X10Y148_SLICE_X13Y148_A1;
  wire [0:0] CLBLM_L_X10Y148_SLICE_X13Y148_A2;
  wire [0:0] CLBLM_L_X10Y148_SLICE_X13Y148_A3;
  wire [0:0] CLBLM_L_X10Y148_SLICE_X13Y148_A4;
  wire [0:0] CLBLM_L_X10Y148_SLICE_X13Y148_A5;
  wire [0:0] CLBLM_L_X10Y148_SLICE_X13Y148_A6;
  wire [0:0] CLBLM_L_X10Y148_SLICE_X13Y148_AO5;
  wire [0:0] CLBLM_L_X10Y148_SLICE_X13Y148_AO6;
  wire [0:0] CLBLM_L_X10Y148_SLICE_X13Y148_AQ;
  wire [0:0] CLBLM_L_X10Y148_SLICE_X13Y148_A_CY;
  wire [0:0] CLBLM_L_X10Y148_SLICE_X13Y148_A_XOR;
  wire [0:0] CLBLM_L_X10Y148_SLICE_X13Y148_B;
  wire [0:0] CLBLM_L_X10Y148_SLICE_X13Y148_B1;
  wire [0:0] CLBLM_L_X10Y148_SLICE_X13Y148_B2;
  wire [0:0] CLBLM_L_X10Y148_SLICE_X13Y148_B3;
  wire [0:0] CLBLM_L_X10Y148_SLICE_X13Y148_B4;
  wire [0:0] CLBLM_L_X10Y148_SLICE_X13Y148_B5;
  wire [0:0] CLBLM_L_X10Y148_SLICE_X13Y148_B6;
  wire [0:0] CLBLM_L_X10Y148_SLICE_X13Y148_BO5;
  wire [0:0] CLBLM_L_X10Y148_SLICE_X13Y148_BO6;
  wire [0:0] CLBLM_L_X10Y148_SLICE_X13Y148_BQ;
  wire [0:0] CLBLM_L_X10Y148_SLICE_X13Y148_B_CY;
  wire [0:0] CLBLM_L_X10Y148_SLICE_X13Y148_B_XOR;
  wire [0:0] CLBLM_L_X10Y148_SLICE_X13Y148_C;
  wire [0:0] CLBLM_L_X10Y148_SLICE_X13Y148_C1;
  wire [0:0] CLBLM_L_X10Y148_SLICE_X13Y148_C2;
  wire [0:0] CLBLM_L_X10Y148_SLICE_X13Y148_C3;
  wire [0:0] CLBLM_L_X10Y148_SLICE_X13Y148_C4;
  wire [0:0] CLBLM_L_X10Y148_SLICE_X13Y148_C5;
  wire [0:0] CLBLM_L_X10Y148_SLICE_X13Y148_C5Q;
  wire [0:0] CLBLM_L_X10Y148_SLICE_X13Y148_C6;
  wire [0:0] CLBLM_L_X10Y148_SLICE_X13Y148_CLK;
  wire [0:0] CLBLM_L_X10Y148_SLICE_X13Y148_CMUX;
  wire [0:0] CLBLM_L_X10Y148_SLICE_X13Y148_CO5;
  wire [0:0] CLBLM_L_X10Y148_SLICE_X13Y148_CO6;
  wire [0:0] CLBLM_L_X10Y148_SLICE_X13Y148_CQ;
  wire [0:0] CLBLM_L_X10Y148_SLICE_X13Y148_C_CY;
  wire [0:0] CLBLM_L_X10Y148_SLICE_X13Y148_C_XOR;
  wire [0:0] CLBLM_L_X10Y148_SLICE_X13Y148_D;
  wire [0:0] CLBLM_L_X10Y148_SLICE_X13Y148_D1;
  wire [0:0] CLBLM_L_X10Y148_SLICE_X13Y148_D2;
  wire [0:0] CLBLM_L_X10Y148_SLICE_X13Y148_D3;
  wire [0:0] CLBLM_L_X10Y148_SLICE_X13Y148_D4;
  wire [0:0] CLBLM_L_X10Y148_SLICE_X13Y148_D5;
  wire [0:0] CLBLM_L_X10Y148_SLICE_X13Y148_D6;
  wire [0:0] CLBLM_L_X10Y148_SLICE_X13Y148_DO5;
  wire [0:0] CLBLM_L_X10Y148_SLICE_X13Y148_DO6;
  wire [0:0] CLBLM_L_X10Y148_SLICE_X13Y148_D_CY;
  wire [0:0] CLBLM_L_X10Y148_SLICE_X13Y148_D_XOR;
  wire [0:0] CLBLM_L_X10Y149_SLICE_X12Y149_A;
  wire [0:0] CLBLM_L_X10Y149_SLICE_X12Y149_A1;
  wire [0:0] CLBLM_L_X10Y149_SLICE_X12Y149_A2;
  wire [0:0] CLBLM_L_X10Y149_SLICE_X12Y149_A3;
  wire [0:0] CLBLM_L_X10Y149_SLICE_X12Y149_A4;
  wire [0:0] CLBLM_L_X10Y149_SLICE_X12Y149_A5;
  wire [0:0] CLBLM_L_X10Y149_SLICE_X12Y149_A5Q;
  wire [0:0] CLBLM_L_X10Y149_SLICE_X12Y149_A6;
  wire [0:0] CLBLM_L_X10Y149_SLICE_X12Y149_AMUX;
  wire [0:0] CLBLM_L_X10Y149_SLICE_X12Y149_AO5;
  wire [0:0] CLBLM_L_X10Y149_SLICE_X12Y149_AO6;
  wire [0:0] CLBLM_L_X10Y149_SLICE_X12Y149_AQ;
  wire [0:0] CLBLM_L_X10Y149_SLICE_X12Y149_A_CY;
  wire [0:0] CLBLM_L_X10Y149_SLICE_X12Y149_A_XOR;
  wire [0:0] CLBLM_L_X10Y149_SLICE_X12Y149_B;
  wire [0:0] CLBLM_L_X10Y149_SLICE_X12Y149_B1;
  wire [0:0] CLBLM_L_X10Y149_SLICE_X12Y149_B2;
  wire [0:0] CLBLM_L_X10Y149_SLICE_X12Y149_B3;
  wire [0:0] CLBLM_L_X10Y149_SLICE_X12Y149_B4;
  wire [0:0] CLBLM_L_X10Y149_SLICE_X12Y149_B5;
  wire [0:0] CLBLM_L_X10Y149_SLICE_X12Y149_B6;
  wire [0:0] CLBLM_L_X10Y149_SLICE_X12Y149_BMUX;
  wire [0:0] CLBLM_L_X10Y149_SLICE_X12Y149_BO5;
  wire [0:0] CLBLM_L_X10Y149_SLICE_X12Y149_BO6;
  wire [0:0] CLBLM_L_X10Y149_SLICE_X12Y149_BQ;
  wire [0:0] CLBLM_L_X10Y149_SLICE_X12Y149_BX;
  wire [0:0] CLBLM_L_X10Y149_SLICE_X12Y149_B_CY;
  wire [0:0] CLBLM_L_X10Y149_SLICE_X12Y149_B_XOR;
  wire [0:0] CLBLM_L_X10Y149_SLICE_X12Y149_C;
  wire [0:0] CLBLM_L_X10Y149_SLICE_X12Y149_C1;
  wire [0:0] CLBLM_L_X10Y149_SLICE_X12Y149_C2;
  wire [0:0] CLBLM_L_X10Y149_SLICE_X12Y149_C3;
  wire [0:0] CLBLM_L_X10Y149_SLICE_X12Y149_C4;
  wire [0:0] CLBLM_L_X10Y149_SLICE_X12Y149_C5;
  wire [0:0] CLBLM_L_X10Y149_SLICE_X12Y149_C6;
  wire [0:0] CLBLM_L_X10Y149_SLICE_X12Y149_CLK;
  wire [0:0] CLBLM_L_X10Y149_SLICE_X12Y149_CMUX;
  wire [0:0] CLBLM_L_X10Y149_SLICE_X12Y149_CO5;
  wire [0:0] CLBLM_L_X10Y149_SLICE_X12Y149_CO6;
  wire [0:0] CLBLM_L_X10Y149_SLICE_X12Y149_C_CY;
  wire [0:0] CLBLM_L_X10Y149_SLICE_X12Y149_C_XOR;
  wire [0:0] CLBLM_L_X10Y149_SLICE_X12Y149_D;
  wire [0:0] CLBLM_L_X10Y149_SLICE_X12Y149_D1;
  wire [0:0] CLBLM_L_X10Y149_SLICE_X12Y149_D2;
  wire [0:0] CLBLM_L_X10Y149_SLICE_X12Y149_D3;
  wire [0:0] CLBLM_L_X10Y149_SLICE_X12Y149_D4;
  wire [0:0] CLBLM_L_X10Y149_SLICE_X12Y149_D5;
  wire [0:0] CLBLM_L_X10Y149_SLICE_X12Y149_D6;
  wire [0:0] CLBLM_L_X10Y149_SLICE_X12Y149_DO5;
  wire [0:0] CLBLM_L_X10Y149_SLICE_X12Y149_DO6;
  wire [0:0] CLBLM_L_X10Y149_SLICE_X12Y149_D_CY;
  wire [0:0] CLBLM_L_X10Y149_SLICE_X12Y149_D_XOR;
  wire [0:0] CLBLM_L_X10Y149_SLICE_X13Y149_A;
  wire [0:0] CLBLM_L_X10Y149_SLICE_X13Y149_A1;
  wire [0:0] CLBLM_L_X10Y149_SLICE_X13Y149_A2;
  wire [0:0] CLBLM_L_X10Y149_SLICE_X13Y149_A3;
  wire [0:0] CLBLM_L_X10Y149_SLICE_X13Y149_A4;
  wire [0:0] CLBLM_L_X10Y149_SLICE_X13Y149_A5;
  wire [0:0] CLBLM_L_X10Y149_SLICE_X13Y149_A6;
  wire [0:0] CLBLM_L_X10Y149_SLICE_X13Y149_AMUX;
  wire [0:0] CLBLM_L_X10Y149_SLICE_X13Y149_AO5;
  wire [0:0] CLBLM_L_X10Y149_SLICE_X13Y149_AO6;
  wire [0:0] CLBLM_L_X10Y149_SLICE_X13Y149_AQ;
  wire [0:0] CLBLM_L_X10Y149_SLICE_X13Y149_A_CY;
  wire [0:0] CLBLM_L_X10Y149_SLICE_X13Y149_A_XOR;
  wire [0:0] CLBLM_L_X10Y149_SLICE_X13Y149_B;
  wire [0:0] CLBLM_L_X10Y149_SLICE_X13Y149_B1;
  wire [0:0] CLBLM_L_X10Y149_SLICE_X13Y149_B2;
  wire [0:0] CLBLM_L_X10Y149_SLICE_X13Y149_B3;
  wire [0:0] CLBLM_L_X10Y149_SLICE_X13Y149_B4;
  wire [0:0] CLBLM_L_X10Y149_SLICE_X13Y149_B5;
  wire [0:0] CLBLM_L_X10Y149_SLICE_X13Y149_B6;
  wire [0:0] CLBLM_L_X10Y149_SLICE_X13Y149_BO5;
  wire [0:0] CLBLM_L_X10Y149_SLICE_X13Y149_BO6;
  wire [0:0] CLBLM_L_X10Y149_SLICE_X13Y149_B_CY;
  wire [0:0] CLBLM_L_X10Y149_SLICE_X13Y149_B_XOR;
  wire [0:0] CLBLM_L_X10Y149_SLICE_X13Y149_C;
  wire [0:0] CLBLM_L_X10Y149_SLICE_X13Y149_C1;
  wire [0:0] CLBLM_L_X10Y149_SLICE_X13Y149_C2;
  wire [0:0] CLBLM_L_X10Y149_SLICE_X13Y149_C3;
  wire [0:0] CLBLM_L_X10Y149_SLICE_X13Y149_C4;
  wire [0:0] CLBLM_L_X10Y149_SLICE_X13Y149_C5;
  wire [0:0] CLBLM_L_X10Y149_SLICE_X13Y149_C6;
  wire [0:0] CLBLM_L_X10Y149_SLICE_X13Y149_CLK;
  wire [0:0] CLBLM_L_X10Y149_SLICE_X13Y149_CO5;
  wire [0:0] CLBLM_L_X10Y149_SLICE_X13Y149_CO6;
  wire [0:0] CLBLM_L_X10Y149_SLICE_X13Y149_C_CY;
  wire [0:0] CLBLM_L_X10Y149_SLICE_X13Y149_C_XOR;
  wire [0:0] CLBLM_L_X10Y149_SLICE_X13Y149_D;
  wire [0:0] CLBLM_L_X10Y149_SLICE_X13Y149_D1;
  wire [0:0] CLBLM_L_X10Y149_SLICE_X13Y149_D2;
  wire [0:0] CLBLM_L_X10Y149_SLICE_X13Y149_D3;
  wire [0:0] CLBLM_L_X10Y149_SLICE_X13Y149_D4;
  wire [0:0] CLBLM_L_X10Y149_SLICE_X13Y149_D5;
  wire [0:0] CLBLM_L_X10Y149_SLICE_X13Y149_D6;
  wire [0:0] CLBLM_L_X10Y149_SLICE_X13Y149_DMUX;
  wire [0:0] CLBLM_L_X10Y149_SLICE_X13Y149_DO5;
  wire [0:0] CLBLM_L_X10Y149_SLICE_X13Y149_DO6;
  wire [0:0] CLBLM_L_X10Y149_SLICE_X13Y149_D_CY;
  wire [0:0] CLBLM_L_X10Y149_SLICE_X13Y149_D_XOR;
  wire [0:0] CLBLM_L_X10Y150_SLICE_X12Y150_A;
  wire [0:0] CLBLM_L_X10Y150_SLICE_X12Y150_A1;
  wire [0:0] CLBLM_L_X10Y150_SLICE_X12Y150_A2;
  wire [0:0] CLBLM_L_X10Y150_SLICE_X12Y150_A3;
  wire [0:0] CLBLM_L_X10Y150_SLICE_X12Y150_A4;
  wire [0:0] CLBLM_L_X10Y150_SLICE_X12Y150_A5;
  wire [0:0] CLBLM_L_X10Y150_SLICE_X12Y150_A6;
  wire [0:0] CLBLM_L_X10Y150_SLICE_X12Y150_AMUX;
  wire [0:0] CLBLM_L_X10Y150_SLICE_X12Y150_AO5;
  wire [0:0] CLBLM_L_X10Y150_SLICE_X12Y150_AO6;
  wire [0:0] CLBLM_L_X10Y150_SLICE_X12Y150_AQ;
  wire [0:0] CLBLM_L_X10Y150_SLICE_X12Y150_AX;
  wire [0:0] CLBLM_L_X10Y150_SLICE_X12Y150_A_CY;
  wire [0:0] CLBLM_L_X10Y150_SLICE_X12Y150_A_XOR;
  wire [0:0] CLBLM_L_X10Y150_SLICE_X12Y150_B;
  wire [0:0] CLBLM_L_X10Y150_SLICE_X12Y150_B1;
  wire [0:0] CLBLM_L_X10Y150_SLICE_X12Y150_B2;
  wire [0:0] CLBLM_L_X10Y150_SLICE_X12Y150_B3;
  wire [0:0] CLBLM_L_X10Y150_SLICE_X12Y150_B4;
  wire [0:0] CLBLM_L_X10Y150_SLICE_X12Y150_B5;
  wire [0:0] CLBLM_L_X10Y150_SLICE_X12Y150_B6;
  wire [0:0] CLBLM_L_X10Y150_SLICE_X12Y150_BMUX;
  wire [0:0] CLBLM_L_X10Y150_SLICE_X12Y150_BO5;
  wire [0:0] CLBLM_L_X10Y150_SLICE_X12Y150_BO6;
  wire [0:0] CLBLM_L_X10Y150_SLICE_X12Y150_B_CY;
  wire [0:0] CLBLM_L_X10Y150_SLICE_X12Y150_B_XOR;
  wire [0:0] CLBLM_L_X10Y150_SLICE_X12Y150_C;
  wire [0:0] CLBLM_L_X10Y150_SLICE_X12Y150_C1;
  wire [0:0] CLBLM_L_X10Y150_SLICE_X12Y150_C2;
  wire [0:0] CLBLM_L_X10Y150_SLICE_X12Y150_C3;
  wire [0:0] CLBLM_L_X10Y150_SLICE_X12Y150_C4;
  wire [0:0] CLBLM_L_X10Y150_SLICE_X12Y150_C5;
  wire [0:0] CLBLM_L_X10Y150_SLICE_X12Y150_C6;
  wire [0:0] CLBLM_L_X10Y150_SLICE_X12Y150_CE;
  wire [0:0] CLBLM_L_X10Y150_SLICE_X12Y150_CLK;
  wire [0:0] CLBLM_L_X10Y150_SLICE_X12Y150_CO5;
  wire [0:0] CLBLM_L_X10Y150_SLICE_X12Y150_CO6;
  wire [0:0] CLBLM_L_X10Y150_SLICE_X12Y150_C_CY;
  wire [0:0] CLBLM_L_X10Y150_SLICE_X12Y150_C_XOR;
  wire [0:0] CLBLM_L_X10Y150_SLICE_X12Y150_D;
  wire [0:0] CLBLM_L_X10Y150_SLICE_X12Y150_D1;
  wire [0:0] CLBLM_L_X10Y150_SLICE_X12Y150_D2;
  wire [0:0] CLBLM_L_X10Y150_SLICE_X12Y150_D3;
  wire [0:0] CLBLM_L_X10Y150_SLICE_X12Y150_D4;
  wire [0:0] CLBLM_L_X10Y150_SLICE_X12Y150_D5;
  wire [0:0] CLBLM_L_X10Y150_SLICE_X12Y150_D6;
  wire [0:0] CLBLM_L_X10Y150_SLICE_X12Y150_DO5;
  wire [0:0] CLBLM_L_X10Y150_SLICE_X12Y150_DO6;
  wire [0:0] CLBLM_L_X10Y150_SLICE_X12Y150_D_CY;
  wire [0:0] CLBLM_L_X10Y150_SLICE_X12Y150_D_XOR;
  wire [0:0] CLBLM_L_X10Y150_SLICE_X13Y150_A;
  wire [0:0] CLBLM_L_X10Y150_SLICE_X13Y150_A1;
  wire [0:0] CLBLM_L_X10Y150_SLICE_X13Y150_A2;
  wire [0:0] CLBLM_L_X10Y150_SLICE_X13Y150_A3;
  wire [0:0] CLBLM_L_X10Y150_SLICE_X13Y150_A4;
  wire [0:0] CLBLM_L_X10Y150_SLICE_X13Y150_A5;
  wire [0:0] CLBLM_L_X10Y150_SLICE_X13Y150_A6;
  wire [0:0] CLBLM_L_X10Y150_SLICE_X13Y150_AO5;
  wire [0:0] CLBLM_L_X10Y150_SLICE_X13Y150_AO6;
  wire [0:0] CLBLM_L_X10Y150_SLICE_X13Y150_AQ;
  wire [0:0] CLBLM_L_X10Y150_SLICE_X13Y150_A_CY;
  wire [0:0] CLBLM_L_X10Y150_SLICE_X13Y150_A_XOR;
  wire [0:0] CLBLM_L_X10Y150_SLICE_X13Y150_B;
  wire [0:0] CLBLM_L_X10Y150_SLICE_X13Y150_B1;
  wire [0:0] CLBLM_L_X10Y150_SLICE_X13Y150_B2;
  wire [0:0] CLBLM_L_X10Y150_SLICE_X13Y150_B3;
  wire [0:0] CLBLM_L_X10Y150_SLICE_X13Y150_B4;
  wire [0:0] CLBLM_L_X10Y150_SLICE_X13Y150_B5;
  wire [0:0] CLBLM_L_X10Y150_SLICE_X13Y150_B6;
  wire [0:0] CLBLM_L_X10Y150_SLICE_X13Y150_BMUX;
  wire [0:0] CLBLM_L_X10Y150_SLICE_X13Y150_BO5;
  wire [0:0] CLBLM_L_X10Y150_SLICE_X13Y150_BO6;
  wire [0:0] CLBLM_L_X10Y150_SLICE_X13Y150_B_CY;
  wire [0:0] CLBLM_L_X10Y150_SLICE_X13Y150_B_XOR;
  wire [0:0] CLBLM_L_X10Y150_SLICE_X13Y150_C;
  wire [0:0] CLBLM_L_X10Y150_SLICE_X13Y150_C1;
  wire [0:0] CLBLM_L_X10Y150_SLICE_X13Y150_C2;
  wire [0:0] CLBLM_L_X10Y150_SLICE_X13Y150_C3;
  wire [0:0] CLBLM_L_X10Y150_SLICE_X13Y150_C4;
  wire [0:0] CLBLM_L_X10Y150_SLICE_X13Y150_C5;
  wire [0:0] CLBLM_L_X10Y150_SLICE_X13Y150_C6;
  wire [0:0] CLBLM_L_X10Y150_SLICE_X13Y150_CLK;
  wire [0:0] CLBLM_L_X10Y150_SLICE_X13Y150_CO5;
  wire [0:0] CLBLM_L_X10Y150_SLICE_X13Y150_CO6;
  wire [0:0] CLBLM_L_X10Y150_SLICE_X13Y150_C_CY;
  wire [0:0] CLBLM_L_X10Y150_SLICE_X13Y150_C_XOR;
  wire [0:0] CLBLM_L_X10Y150_SLICE_X13Y150_D;
  wire [0:0] CLBLM_L_X10Y150_SLICE_X13Y150_D1;
  wire [0:0] CLBLM_L_X10Y150_SLICE_X13Y150_D2;
  wire [0:0] CLBLM_L_X10Y150_SLICE_X13Y150_D3;
  wire [0:0] CLBLM_L_X10Y150_SLICE_X13Y150_D4;
  wire [0:0] CLBLM_L_X10Y150_SLICE_X13Y150_D5;
  wire [0:0] CLBLM_L_X10Y150_SLICE_X13Y150_D6;
  wire [0:0] CLBLM_L_X10Y150_SLICE_X13Y150_DO5;
  wire [0:0] CLBLM_L_X10Y150_SLICE_X13Y150_DO6;
  wire [0:0] CLBLM_L_X10Y150_SLICE_X13Y150_D_CY;
  wire [0:0] CLBLM_L_X10Y150_SLICE_X13Y150_D_XOR;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X12Y151_A;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X12Y151_A1;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X12Y151_A2;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X12Y151_A3;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X12Y151_A4;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X12Y151_A5;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X12Y151_A6;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X12Y151_AO5;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X12Y151_AO6;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X12Y151_AQ;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X12Y151_A_CY;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X12Y151_A_XOR;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X12Y151_B;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X12Y151_B1;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X12Y151_B2;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X12Y151_B3;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X12Y151_B4;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X12Y151_B5;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X12Y151_B6;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X12Y151_BO5;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X12Y151_BO6;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X12Y151_BQ;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X12Y151_B_CY;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X12Y151_B_XOR;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X12Y151_C;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X12Y151_C1;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X12Y151_C2;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X12Y151_C3;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X12Y151_C4;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X12Y151_C5;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X12Y151_C6;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X12Y151_CLK;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X12Y151_CO5;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X12Y151_CO6;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X12Y151_CQ;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X12Y151_C_CY;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X12Y151_C_XOR;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X12Y151_D;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X12Y151_D1;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X12Y151_D2;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X12Y151_D3;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X12Y151_D4;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X12Y151_D5;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X12Y151_D6;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X12Y151_DO5;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X12Y151_DO6;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X12Y151_DQ;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X12Y151_D_CY;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X12Y151_D_XOR;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X13Y151_A;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X13Y151_A1;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X13Y151_A2;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X13Y151_A3;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X13Y151_A4;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X13Y151_A5;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X13Y151_A5Q;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X13Y151_A6;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X13Y151_AMUX;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X13Y151_AO5;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X13Y151_AO6;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X13Y151_AQ;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X13Y151_A_CY;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X13Y151_A_XOR;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X13Y151_B;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X13Y151_B1;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X13Y151_B2;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X13Y151_B3;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X13Y151_B4;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X13Y151_B5;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X13Y151_B6;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X13Y151_BMUX;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X13Y151_BO5;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X13Y151_BO6;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X13Y151_B_CY;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X13Y151_B_XOR;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X13Y151_C;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X13Y151_C1;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X13Y151_C2;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X13Y151_C3;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X13Y151_C4;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X13Y151_C5;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X13Y151_C6;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X13Y151_CLK;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X13Y151_CO5;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X13Y151_CO6;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X13Y151_C_CY;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X13Y151_C_XOR;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X13Y151_D;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X13Y151_D1;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X13Y151_D2;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X13Y151_D3;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X13Y151_D4;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X13Y151_D5;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X13Y151_D6;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X13Y151_DO5;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X13Y151_DO6;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X13Y151_D_CY;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X13Y151_D_XOR;
  wire [0:0] CLBLM_L_X10Y152_SLICE_X12Y152_A;
  wire [0:0] CLBLM_L_X10Y152_SLICE_X12Y152_A1;
  wire [0:0] CLBLM_L_X10Y152_SLICE_X12Y152_A2;
  wire [0:0] CLBLM_L_X10Y152_SLICE_X12Y152_A3;
  wire [0:0] CLBLM_L_X10Y152_SLICE_X12Y152_A4;
  wire [0:0] CLBLM_L_X10Y152_SLICE_X12Y152_A5;
  wire [0:0] CLBLM_L_X10Y152_SLICE_X12Y152_A6;
  wire [0:0] CLBLM_L_X10Y152_SLICE_X12Y152_AO5;
  wire [0:0] CLBLM_L_X10Y152_SLICE_X12Y152_AO6;
  wire [0:0] CLBLM_L_X10Y152_SLICE_X12Y152_AQ;
  wire [0:0] CLBLM_L_X10Y152_SLICE_X12Y152_A_CY;
  wire [0:0] CLBLM_L_X10Y152_SLICE_X12Y152_A_XOR;
  wire [0:0] CLBLM_L_X10Y152_SLICE_X12Y152_B;
  wire [0:0] CLBLM_L_X10Y152_SLICE_X12Y152_B1;
  wire [0:0] CLBLM_L_X10Y152_SLICE_X12Y152_B2;
  wire [0:0] CLBLM_L_X10Y152_SLICE_X12Y152_B3;
  wire [0:0] CLBLM_L_X10Y152_SLICE_X12Y152_B4;
  wire [0:0] CLBLM_L_X10Y152_SLICE_X12Y152_B5;
  wire [0:0] CLBLM_L_X10Y152_SLICE_X12Y152_B6;
  wire [0:0] CLBLM_L_X10Y152_SLICE_X12Y152_BO5;
  wire [0:0] CLBLM_L_X10Y152_SLICE_X12Y152_BO6;
  wire [0:0] CLBLM_L_X10Y152_SLICE_X12Y152_BQ;
  wire [0:0] CLBLM_L_X10Y152_SLICE_X12Y152_B_CY;
  wire [0:0] CLBLM_L_X10Y152_SLICE_X12Y152_B_XOR;
  wire [0:0] CLBLM_L_X10Y152_SLICE_X12Y152_C;
  wire [0:0] CLBLM_L_X10Y152_SLICE_X12Y152_C1;
  wire [0:0] CLBLM_L_X10Y152_SLICE_X12Y152_C2;
  wire [0:0] CLBLM_L_X10Y152_SLICE_X12Y152_C3;
  wire [0:0] CLBLM_L_X10Y152_SLICE_X12Y152_C4;
  wire [0:0] CLBLM_L_X10Y152_SLICE_X12Y152_C5;
  wire [0:0] CLBLM_L_X10Y152_SLICE_X12Y152_C6;
  wire [0:0] CLBLM_L_X10Y152_SLICE_X12Y152_CLK;
  wire [0:0] CLBLM_L_X10Y152_SLICE_X12Y152_CO5;
  wire [0:0] CLBLM_L_X10Y152_SLICE_X12Y152_CO6;
  wire [0:0] CLBLM_L_X10Y152_SLICE_X12Y152_CQ;
  wire [0:0] CLBLM_L_X10Y152_SLICE_X12Y152_C_CY;
  wire [0:0] CLBLM_L_X10Y152_SLICE_X12Y152_C_XOR;
  wire [0:0] CLBLM_L_X10Y152_SLICE_X12Y152_D;
  wire [0:0] CLBLM_L_X10Y152_SLICE_X12Y152_D1;
  wire [0:0] CLBLM_L_X10Y152_SLICE_X12Y152_D2;
  wire [0:0] CLBLM_L_X10Y152_SLICE_X12Y152_D3;
  wire [0:0] CLBLM_L_X10Y152_SLICE_X12Y152_D4;
  wire [0:0] CLBLM_L_X10Y152_SLICE_X12Y152_D5;
  wire [0:0] CLBLM_L_X10Y152_SLICE_X12Y152_D6;
  wire [0:0] CLBLM_L_X10Y152_SLICE_X12Y152_DO5;
  wire [0:0] CLBLM_L_X10Y152_SLICE_X12Y152_DO6;
  wire [0:0] CLBLM_L_X10Y152_SLICE_X12Y152_D_CY;
  wire [0:0] CLBLM_L_X10Y152_SLICE_X12Y152_D_XOR;
  wire [0:0] CLBLM_L_X10Y152_SLICE_X13Y152_A;
  wire [0:0] CLBLM_L_X10Y152_SLICE_X13Y152_A1;
  wire [0:0] CLBLM_L_X10Y152_SLICE_X13Y152_A2;
  wire [0:0] CLBLM_L_X10Y152_SLICE_X13Y152_A3;
  wire [0:0] CLBLM_L_X10Y152_SLICE_X13Y152_A4;
  wire [0:0] CLBLM_L_X10Y152_SLICE_X13Y152_A5;
  wire [0:0] CLBLM_L_X10Y152_SLICE_X13Y152_A6;
  wire [0:0] CLBLM_L_X10Y152_SLICE_X13Y152_AO5;
  wire [0:0] CLBLM_L_X10Y152_SLICE_X13Y152_AO6;
  wire [0:0] CLBLM_L_X10Y152_SLICE_X13Y152_AQ;
  wire [0:0] CLBLM_L_X10Y152_SLICE_X13Y152_A_CY;
  wire [0:0] CLBLM_L_X10Y152_SLICE_X13Y152_A_XOR;
  wire [0:0] CLBLM_L_X10Y152_SLICE_X13Y152_B;
  wire [0:0] CLBLM_L_X10Y152_SLICE_X13Y152_B1;
  wire [0:0] CLBLM_L_X10Y152_SLICE_X13Y152_B2;
  wire [0:0] CLBLM_L_X10Y152_SLICE_X13Y152_B3;
  wire [0:0] CLBLM_L_X10Y152_SLICE_X13Y152_B4;
  wire [0:0] CLBLM_L_X10Y152_SLICE_X13Y152_B5;
  wire [0:0] CLBLM_L_X10Y152_SLICE_X13Y152_B6;
  wire [0:0] CLBLM_L_X10Y152_SLICE_X13Y152_BO5;
  wire [0:0] CLBLM_L_X10Y152_SLICE_X13Y152_BO6;
  wire [0:0] CLBLM_L_X10Y152_SLICE_X13Y152_BQ;
  wire [0:0] CLBLM_L_X10Y152_SLICE_X13Y152_B_CY;
  wire [0:0] CLBLM_L_X10Y152_SLICE_X13Y152_B_XOR;
  wire [0:0] CLBLM_L_X10Y152_SLICE_X13Y152_C;
  wire [0:0] CLBLM_L_X10Y152_SLICE_X13Y152_C1;
  wire [0:0] CLBLM_L_X10Y152_SLICE_X13Y152_C2;
  wire [0:0] CLBLM_L_X10Y152_SLICE_X13Y152_C3;
  wire [0:0] CLBLM_L_X10Y152_SLICE_X13Y152_C4;
  wire [0:0] CLBLM_L_X10Y152_SLICE_X13Y152_C5;
  wire [0:0] CLBLM_L_X10Y152_SLICE_X13Y152_C6;
  wire [0:0] CLBLM_L_X10Y152_SLICE_X13Y152_CLK;
  wire [0:0] CLBLM_L_X10Y152_SLICE_X13Y152_CO5;
  wire [0:0] CLBLM_L_X10Y152_SLICE_X13Y152_CO6;
  wire [0:0] CLBLM_L_X10Y152_SLICE_X13Y152_CQ;
  wire [0:0] CLBLM_L_X10Y152_SLICE_X13Y152_C_CY;
  wire [0:0] CLBLM_L_X10Y152_SLICE_X13Y152_C_XOR;
  wire [0:0] CLBLM_L_X10Y152_SLICE_X13Y152_D;
  wire [0:0] CLBLM_L_X10Y152_SLICE_X13Y152_D1;
  wire [0:0] CLBLM_L_X10Y152_SLICE_X13Y152_D2;
  wire [0:0] CLBLM_L_X10Y152_SLICE_X13Y152_D3;
  wire [0:0] CLBLM_L_X10Y152_SLICE_X13Y152_D4;
  wire [0:0] CLBLM_L_X10Y152_SLICE_X13Y152_D5;
  wire [0:0] CLBLM_L_X10Y152_SLICE_X13Y152_D6;
  wire [0:0] CLBLM_L_X10Y152_SLICE_X13Y152_DMUX;
  wire [0:0] CLBLM_L_X10Y152_SLICE_X13Y152_DO5;
  wire [0:0] CLBLM_L_X10Y152_SLICE_X13Y152_DO6;
  wire [0:0] CLBLM_L_X10Y152_SLICE_X13Y152_D_CY;
  wire [0:0] CLBLM_L_X10Y152_SLICE_X13Y152_D_XOR;
  wire [0:0] CLBLM_L_X10Y153_SLICE_X12Y153_A;
  wire [0:0] CLBLM_L_X10Y153_SLICE_X12Y153_A1;
  wire [0:0] CLBLM_L_X10Y153_SLICE_X12Y153_A2;
  wire [0:0] CLBLM_L_X10Y153_SLICE_X12Y153_A3;
  wire [0:0] CLBLM_L_X10Y153_SLICE_X12Y153_A4;
  wire [0:0] CLBLM_L_X10Y153_SLICE_X12Y153_A5;
  wire [0:0] CLBLM_L_X10Y153_SLICE_X12Y153_A5Q;
  wire [0:0] CLBLM_L_X10Y153_SLICE_X12Y153_A6;
  wire [0:0] CLBLM_L_X10Y153_SLICE_X12Y153_AMUX;
  wire [0:0] CLBLM_L_X10Y153_SLICE_X12Y153_AO5;
  wire [0:0] CLBLM_L_X10Y153_SLICE_X12Y153_AO6;
  wire [0:0] CLBLM_L_X10Y153_SLICE_X12Y153_AQ;
  wire [0:0] CLBLM_L_X10Y153_SLICE_X12Y153_AX;
  wire [0:0] CLBLM_L_X10Y153_SLICE_X12Y153_A_CY;
  wire [0:0] CLBLM_L_X10Y153_SLICE_X12Y153_A_XOR;
  wire [0:0] CLBLM_L_X10Y153_SLICE_X12Y153_B;
  wire [0:0] CLBLM_L_X10Y153_SLICE_X12Y153_B1;
  wire [0:0] CLBLM_L_X10Y153_SLICE_X12Y153_B2;
  wire [0:0] CLBLM_L_X10Y153_SLICE_X12Y153_B3;
  wire [0:0] CLBLM_L_X10Y153_SLICE_X12Y153_B4;
  wire [0:0] CLBLM_L_X10Y153_SLICE_X12Y153_B5;
  wire [0:0] CLBLM_L_X10Y153_SLICE_X12Y153_B6;
  wire [0:0] CLBLM_L_X10Y153_SLICE_X12Y153_BO5;
  wire [0:0] CLBLM_L_X10Y153_SLICE_X12Y153_BO6;
  wire [0:0] CLBLM_L_X10Y153_SLICE_X12Y153_BQ;
  wire [0:0] CLBLM_L_X10Y153_SLICE_X12Y153_B_CY;
  wire [0:0] CLBLM_L_X10Y153_SLICE_X12Y153_B_XOR;
  wire [0:0] CLBLM_L_X10Y153_SLICE_X12Y153_C;
  wire [0:0] CLBLM_L_X10Y153_SLICE_X12Y153_C1;
  wire [0:0] CLBLM_L_X10Y153_SLICE_X12Y153_C2;
  wire [0:0] CLBLM_L_X10Y153_SLICE_X12Y153_C3;
  wire [0:0] CLBLM_L_X10Y153_SLICE_X12Y153_C4;
  wire [0:0] CLBLM_L_X10Y153_SLICE_X12Y153_C5;
  wire [0:0] CLBLM_L_X10Y153_SLICE_X12Y153_C6;
  wire [0:0] CLBLM_L_X10Y153_SLICE_X12Y153_CLK;
  wire [0:0] CLBLM_L_X10Y153_SLICE_X12Y153_CMUX;
  wire [0:0] CLBLM_L_X10Y153_SLICE_X12Y153_CO5;
  wire [0:0] CLBLM_L_X10Y153_SLICE_X12Y153_CO6;
  wire [0:0] CLBLM_L_X10Y153_SLICE_X12Y153_C_CY;
  wire [0:0] CLBLM_L_X10Y153_SLICE_X12Y153_C_XOR;
  wire [0:0] CLBLM_L_X10Y153_SLICE_X12Y153_D;
  wire [0:0] CLBLM_L_X10Y153_SLICE_X12Y153_D1;
  wire [0:0] CLBLM_L_X10Y153_SLICE_X12Y153_D2;
  wire [0:0] CLBLM_L_X10Y153_SLICE_X12Y153_D3;
  wire [0:0] CLBLM_L_X10Y153_SLICE_X12Y153_D4;
  wire [0:0] CLBLM_L_X10Y153_SLICE_X12Y153_D5;
  wire [0:0] CLBLM_L_X10Y153_SLICE_X12Y153_D6;
  wire [0:0] CLBLM_L_X10Y153_SLICE_X12Y153_DO5;
  wire [0:0] CLBLM_L_X10Y153_SLICE_X12Y153_DO6;
  wire [0:0] CLBLM_L_X10Y153_SLICE_X12Y153_D_CY;
  wire [0:0] CLBLM_L_X10Y153_SLICE_X12Y153_D_XOR;
  wire [0:0] CLBLM_L_X10Y153_SLICE_X13Y153_A;
  wire [0:0] CLBLM_L_X10Y153_SLICE_X13Y153_A1;
  wire [0:0] CLBLM_L_X10Y153_SLICE_X13Y153_A2;
  wire [0:0] CLBLM_L_X10Y153_SLICE_X13Y153_A3;
  wire [0:0] CLBLM_L_X10Y153_SLICE_X13Y153_A4;
  wire [0:0] CLBLM_L_X10Y153_SLICE_X13Y153_A5;
  wire [0:0] CLBLM_L_X10Y153_SLICE_X13Y153_A5Q;
  wire [0:0] CLBLM_L_X10Y153_SLICE_X13Y153_A6;
  wire [0:0] CLBLM_L_X10Y153_SLICE_X13Y153_AMUX;
  wire [0:0] CLBLM_L_X10Y153_SLICE_X13Y153_AO5;
  wire [0:0] CLBLM_L_X10Y153_SLICE_X13Y153_AO6;
  wire [0:0] CLBLM_L_X10Y153_SLICE_X13Y153_AQ;
  wire [0:0] CLBLM_L_X10Y153_SLICE_X13Y153_AX;
  wire [0:0] CLBLM_L_X10Y153_SLICE_X13Y153_A_CY;
  wire [0:0] CLBLM_L_X10Y153_SLICE_X13Y153_A_XOR;
  wire [0:0] CLBLM_L_X10Y153_SLICE_X13Y153_B;
  wire [0:0] CLBLM_L_X10Y153_SLICE_X13Y153_B1;
  wire [0:0] CLBLM_L_X10Y153_SLICE_X13Y153_B2;
  wire [0:0] CLBLM_L_X10Y153_SLICE_X13Y153_B3;
  wire [0:0] CLBLM_L_X10Y153_SLICE_X13Y153_B4;
  wire [0:0] CLBLM_L_X10Y153_SLICE_X13Y153_B5;
  wire [0:0] CLBLM_L_X10Y153_SLICE_X13Y153_B6;
  wire [0:0] CLBLM_L_X10Y153_SLICE_X13Y153_BO5;
  wire [0:0] CLBLM_L_X10Y153_SLICE_X13Y153_BO6;
  wire [0:0] CLBLM_L_X10Y153_SLICE_X13Y153_BQ;
  wire [0:0] CLBLM_L_X10Y153_SLICE_X13Y153_B_CY;
  wire [0:0] CLBLM_L_X10Y153_SLICE_X13Y153_B_XOR;
  wire [0:0] CLBLM_L_X10Y153_SLICE_X13Y153_C;
  wire [0:0] CLBLM_L_X10Y153_SLICE_X13Y153_C1;
  wire [0:0] CLBLM_L_X10Y153_SLICE_X13Y153_C2;
  wire [0:0] CLBLM_L_X10Y153_SLICE_X13Y153_C3;
  wire [0:0] CLBLM_L_X10Y153_SLICE_X13Y153_C4;
  wire [0:0] CLBLM_L_X10Y153_SLICE_X13Y153_C5;
  wire [0:0] CLBLM_L_X10Y153_SLICE_X13Y153_C6;
  wire [0:0] CLBLM_L_X10Y153_SLICE_X13Y153_CLK;
  wire [0:0] CLBLM_L_X10Y153_SLICE_X13Y153_CO5;
  wire [0:0] CLBLM_L_X10Y153_SLICE_X13Y153_CO6;
  wire [0:0] CLBLM_L_X10Y153_SLICE_X13Y153_CQ;
  wire [0:0] CLBLM_L_X10Y153_SLICE_X13Y153_C_CY;
  wire [0:0] CLBLM_L_X10Y153_SLICE_X13Y153_C_XOR;
  wire [0:0] CLBLM_L_X10Y153_SLICE_X13Y153_D;
  wire [0:0] CLBLM_L_X10Y153_SLICE_X13Y153_D1;
  wire [0:0] CLBLM_L_X10Y153_SLICE_X13Y153_D2;
  wire [0:0] CLBLM_L_X10Y153_SLICE_X13Y153_D3;
  wire [0:0] CLBLM_L_X10Y153_SLICE_X13Y153_D4;
  wire [0:0] CLBLM_L_X10Y153_SLICE_X13Y153_D5;
  wire [0:0] CLBLM_L_X10Y153_SLICE_X13Y153_D6;
  wire [0:0] CLBLM_L_X10Y153_SLICE_X13Y153_DMUX;
  wire [0:0] CLBLM_L_X10Y153_SLICE_X13Y153_DO5;
  wire [0:0] CLBLM_L_X10Y153_SLICE_X13Y153_DO6;
  wire [0:0] CLBLM_L_X10Y153_SLICE_X13Y153_D_CY;
  wire [0:0] CLBLM_L_X10Y153_SLICE_X13Y153_D_XOR;
  wire [0:0] CLBLM_L_X10Y154_SLICE_X12Y154_A;
  wire [0:0] CLBLM_L_X10Y154_SLICE_X12Y154_A1;
  wire [0:0] CLBLM_L_X10Y154_SLICE_X12Y154_A2;
  wire [0:0] CLBLM_L_X10Y154_SLICE_X12Y154_A3;
  wire [0:0] CLBLM_L_X10Y154_SLICE_X12Y154_A4;
  wire [0:0] CLBLM_L_X10Y154_SLICE_X12Y154_A5;
  wire [0:0] CLBLM_L_X10Y154_SLICE_X12Y154_A5Q;
  wire [0:0] CLBLM_L_X10Y154_SLICE_X12Y154_A6;
  wire [0:0] CLBLM_L_X10Y154_SLICE_X12Y154_AMUX;
  wire [0:0] CLBLM_L_X10Y154_SLICE_X12Y154_AO5;
  wire [0:0] CLBLM_L_X10Y154_SLICE_X12Y154_AO6;
  wire [0:0] CLBLM_L_X10Y154_SLICE_X12Y154_AQ;
  wire [0:0] CLBLM_L_X10Y154_SLICE_X12Y154_AX;
  wire [0:0] CLBLM_L_X10Y154_SLICE_X12Y154_A_CY;
  wire [0:0] CLBLM_L_X10Y154_SLICE_X12Y154_A_XOR;
  wire [0:0] CLBLM_L_X10Y154_SLICE_X12Y154_B;
  wire [0:0] CLBLM_L_X10Y154_SLICE_X12Y154_B1;
  wire [0:0] CLBLM_L_X10Y154_SLICE_X12Y154_B2;
  wire [0:0] CLBLM_L_X10Y154_SLICE_X12Y154_B3;
  wire [0:0] CLBLM_L_X10Y154_SLICE_X12Y154_B4;
  wire [0:0] CLBLM_L_X10Y154_SLICE_X12Y154_B5;
  wire [0:0] CLBLM_L_X10Y154_SLICE_X12Y154_B5Q;
  wire [0:0] CLBLM_L_X10Y154_SLICE_X12Y154_B6;
  wire [0:0] CLBLM_L_X10Y154_SLICE_X12Y154_BMUX;
  wire [0:0] CLBLM_L_X10Y154_SLICE_X12Y154_BO5;
  wire [0:0] CLBLM_L_X10Y154_SLICE_X12Y154_BO6;
  wire [0:0] CLBLM_L_X10Y154_SLICE_X12Y154_BQ;
  wire [0:0] CLBLM_L_X10Y154_SLICE_X12Y154_BX;
  wire [0:0] CLBLM_L_X10Y154_SLICE_X12Y154_B_CY;
  wire [0:0] CLBLM_L_X10Y154_SLICE_X12Y154_B_XOR;
  wire [0:0] CLBLM_L_X10Y154_SLICE_X12Y154_C;
  wire [0:0] CLBLM_L_X10Y154_SLICE_X12Y154_C1;
  wire [0:0] CLBLM_L_X10Y154_SLICE_X12Y154_C2;
  wire [0:0] CLBLM_L_X10Y154_SLICE_X12Y154_C3;
  wire [0:0] CLBLM_L_X10Y154_SLICE_X12Y154_C4;
  wire [0:0] CLBLM_L_X10Y154_SLICE_X12Y154_C5;
  wire [0:0] CLBLM_L_X10Y154_SLICE_X12Y154_C6;
  wire [0:0] CLBLM_L_X10Y154_SLICE_X12Y154_CLK;
  wire [0:0] CLBLM_L_X10Y154_SLICE_X12Y154_CMUX;
  wire [0:0] CLBLM_L_X10Y154_SLICE_X12Y154_CO5;
  wire [0:0] CLBLM_L_X10Y154_SLICE_X12Y154_CO6;
  wire [0:0] CLBLM_L_X10Y154_SLICE_X12Y154_C_CY;
  wire [0:0] CLBLM_L_X10Y154_SLICE_X12Y154_C_XOR;
  wire [0:0] CLBLM_L_X10Y154_SLICE_X12Y154_D;
  wire [0:0] CLBLM_L_X10Y154_SLICE_X12Y154_D1;
  wire [0:0] CLBLM_L_X10Y154_SLICE_X12Y154_D2;
  wire [0:0] CLBLM_L_X10Y154_SLICE_X12Y154_D3;
  wire [0:0] CLBLM_L_X10Y154_SLICE_X12Y154_D4;
  wire [0:0] CLBLM_L_X10Y154_SLICE_X12Y154_D5;
  wire [0:0] CLBLM_L_X10Y154_SLICE_X12Y154_D6;
  wire [0:0] CLBLM_L_X10Y154_SLICE_X12Y154_DMUX;
  wire [0:0] CLBLM_L_X10Y154_SLICE_X12Y154_DO5;
  wire [0:0] CLBLM_L_X10Y154_SLICE_X12Y154_DO6;
  wire [0:0] CLBLM_L_X10Y154_SLICE_X12Y154_D_CY;
  wire [0:0] CLBLM_L_X10Y154_SLICE_X12Y154_D_XOR;
  wire [0:0] CLBLM_L_X10Y154_SLICE_X13Y154_A;
  wire [0:0] CLBLM_L_X10Y154_SLICE_X13Y154_A1;
  wire [0:0] CLBLM_L_X10Y154_SLICE_X13Y154_A2;
  wire [0:0] CLBLM_L_X10Y154_SLICE_X13Y154_A3;
  wire [0:0] CLBLM_L_X10Y154_SLICE_X13Y154_A4;
  wire [0:0] CLBLM_L_X10Y154_SLICE_X13Y154_A5;
  wire [0:0] CLBLM_L_X10Y154_SLICE_X13Y154_A6;
  wire [0:0] CLBLM_L_X10Y154_SLICE_X13Y154_AO5;
  wire [0:0] CLBLM_L_X10Y154_SLICE_X13Y154_AO6;
  wire [0:0] CLBLM_L_X10Y154_SLICE_X13Y154_AQ;
  wire [0:0] CLBLM_L_X10Y154_SLICE_X13Y154_A_CY;
  wire [0:0] CLBLM_L_X10Y154_SLICE_X13Y154_A_XOR;
  wire [0:0] CLBLM_L_X10Y154_SLICE_X13Y154_B;
  wire [0:0] CLBLM_L_X10Y154_SLICE_X13Y154_B1;
  wire [0:0] CLBLM_L_X10Y154_SLICE_X13Y154_B2;
  wire [0:0] CLBLM_L_X10Y154_SLICE_X13Y154_B3;
  wire [0:0] CLBLM_L_X10Y154_SLICE_X13Y154_B4;
  wire [0:0] CLBLM_L_X10Y154_SLICE_X13Y154_B5;
  wire [0:0] CLBLM_L_X10Y154_SLICE_X13Y154_B6;
  wire [0:0] CLBLM_L_X10Y154_SLICE_X13Y154_BMUX;
  wire [0:0] CLBLM_L_X10Y154_SLICE_X13Y154_BO5;
  wire [0:0] CLBLM_L_X10Y154_SLICE_X13Y154_BO6;
  wire [0:0] CLBLM_L_X10Y154_SLICE_X13Y154_B_CY;
  wire [0:0] CLBLM_L_X10Y154_SLICE_X13Y154_B_XOR;
  wire [0:0] CLBLM_L_X10Y154_SLICE_X13Y154_C;
  wire [0:0] CLBLM_L_X10Y154_SLICE_X13Y154_C1;
  wire [0:0] CLBLM_L_X10Y154_SLICE_X13Y154_C2;
  wire [0:0] CLBLM_L_X10Y154_SLICE_X13Y154_C3;
  wire [0:0] CLBLM_L_X10Y154_SLICE_X13Y154_C4;
  wire [0:0] CLBLM_L_X10Y154_SLICE_X13Y154_C5;
  wire [0:0] CLBLM_L_X10Y154_SLICE_X13Y154_C6;
  wire [0:0] CLBLM_L_X10Y154_SLICE_X13Y154_CLK;
  wire [0:0] CLBLM_L_X10Y154_SLICE_X13Y154_CMUX;
  wire [0:0] CLBLM_L_X10Y154_SLICE_X13Y154_CO5;
  wire [0:0] CLBLM_L_X10Y154_SLICE_X13Y154_CO6;
  wire [0:0] CLBLM_L_X10Y154_SLICE_X13Y154_C_CY;
  wire [0:0] CLBLM_L_X10Y154_SLICE_X13Y154_C_XOR;
  wire [0:0] CLBLM_L_X10Y154_SLICE_X13Y154_D;
  wire [0:0] CLBLM_L_X10Y154_SLICE_X13Y154_D1;
  wire [0:0] CLBLM_L_X10Y154_SLICE_X13Y154_D2;
  wire [0:0] CLBLM_L_X10Y154_SLICE_X13Y154_D3;
  wire [0:0] CLBLM_L_X10Y154_SLICE_X13Y154_D4;
  wire [0:0] CLBLM_L_X10Y154_SLICE_X13Y154_D5;
  wire [0:0] CLBLM_L_X10Y154_SLICE_X13Y154_D6;
  wire [0:0] CLBLM_L_X10Y154_SLICE_X13Y154_DO5;
  wire [0:0] CLBLM_L_X10Y154_SLICE_X13Y154_DO6;
  wire [0:0] CLBLM_L_X10Y154_SLICE_X13Y154_D_CY;
  wire [0:0] CLBLM_L_X10Y154_SLICE_X13Y154_D_XOR;
  wire [0:0] CLBLM_L_X10Y155_SLICE_X12Y155_A;
  wire [0:0] CLBLM_L_X10Y155_SLICE_X12Y155_A1;
  wire [0:0] CLBLM_L_X10Y155_SLICE_X12Y155_A2;
  wire [0:0] CLBLM_L_X10Y155_SLICE_X12Y155_A3;
  wire [0:0] CLBLM_L_X10Y155_SLICE_X12Y155_A4;
  wire [0:0] CLBLM_L_X10Y155_SLICE_X12Y155_A5;
  wire [0:0] CLBLM_L_X10Y155_SLICE_X12Y155_A6;
  wire [0:0] CLBLM_L_X10Y155_SLICE_X12Y155_AO5;
  wire [0:0] CLBLM_L_X10Y155_SLICE_X12Y155_AO6;
  wire [0:0] CLBLM_L_X10Y155_SLICE_X12Y155_AQ;
  wire [0:0] CLBLM_L_X10Y155_SLICE_X12Y155_A_CY;
  wire [0:0] CLBLM_L_X10Y155_SLICE_X12Y155_A_XOR;
  wire [0:0] CLBLM_L_X10Y155_SLICE_X12Y155_B;
  wire [0:0] CLBLM_L_X10Y155_SLICE_X12Y155_B1;
  wire [0:0] CLBLM_L_X10Y155_SLICE_X12Y155_B2;
  wire [0:0] CLBLM_L_X10Y155_SLICE_X12Y155_B3;
  wire [0:0] CLBLM_L_X10Y155_SLICE_X12Y155_B4;
  wire [0:0] CLBLM_L_X10Y155_SLICE_X12Y155_B5;
  wire [0:0] CLBLM_L_X10Y155_SLICE_X12Y155_B6;
  wire [0:0] CLBLM_L_X10Y155_SLICE_X12Y155_BMUX;
  wire [0:0] CLBLM_L_X10Y155_SLICE_X12Y155_BO5;
  wire [0:0] CLBLM_L_X10Y155_SLICE_X12Y155_BO6;
  wire [0:0] CLBLM_L_X10Y155_SLICE_X12Y155_B_CY;
  wire [0:0] CLBLM_L_X10Y155_SLICE_X12Y155_B_XOR;
  wire [0:0] CLBLM_L_X10Y155_SLICE_X12Y155_C;
  wire [0:0] CLBLM_L_X10Y155_SLICE_X12Y155_C1;
  wire [0:0] CLBLM_L_X10Y155_SLICE_X12Y155_C2;
  wire [0:0] CLBLM_L_X10Y155_SLICE_X12Y155_C3;
  wire [0:0] CLBLM_L_X10Y155_SLICE_X12Y155_C4;
  wire [0:0] CLBLM_L_X10Y155_SLICE_X12Y155_C5;
  wire [0:0] CLBLM_L_X10Y155_SLICE_X12Y155_C6;
  wire [0:0] CLBLM_L_X10Y155_SLICE_X12Y155_CLK;
  wire [0:0] CLBLM_L_X10Y155_SLICE_X12Y155_CO5;
  wire [0:0] CLBLM_L_X10Y155_SLICE_X12Y155_CO6;
  wire [0:0] CLBLM_L_X10Y155_SLICE_X12Y155_C_CY;
  wire [0:0] CLBLM_L_X10Y155_SLICE_X12Y155_C_XOR;
  wire [0:0] CLBLM_L_X10Y155_SLICE_X12Y155_D;
  wire [0:0] CLBLM_L_X10Y155_SLICE_X12Y155_D1;
  wire [0:0] CLBLM_L_X10Y155_SLICE_X12Y155_D2;
  wire [0:0] CLBLM_L_X10Y155_SLICE_X12Y155_D3;
  wire [0:0] CLBLM_L_X10Y155_SLICE_X12Y155_D4;
  wire [0:0] CLBLM_L_X10Y155_SLICE_X12Y155_D5;
  wire [0:0] CLBLM_L_X10Y155_SLICE_X12Y155_D6;
  wire [0:0] CLBLM_L_X10Y155_SLICE_X12Y155_DO5;
  wire [0:0] CLBLM_L_X10Y155_SLICE_X12Y155_DO6;
  wire [0:0] CLBLM_L_X10Y155_SLICE_X12Y155_D_CY;
  wire [0:0] CLBLM_L_X10Y155_SLICE_X12Y155_D_XOR;
  wire [0:0] CLBLM_L_X10Y155_SLICE_X13Y155_A;
  wire [0:0] CLBLM_L_X10Y155_SLICE_X13Y155_A1;
  wire [0:0] CLBLM_L_X10Y155_SLICE_X13Y155_A2;
  wire [0:0] CLBLM_L_X10Y155_SLICE_X13Y155_A3;
  wire [0:0] CLBLM_L_X10Y155_SLICE_X13Y155_A4;
  wire [0:0] CLBLM_L_X10Y155_SLICE_X13Y155_A5;
  wire [0:0] CLBLM_L_X10Y155_SLICE_X13Y155_A6;
  wire [0:0] CLBLM_L_X10Y155_SLICE_X13Y155_AMUX;
  wire [0:0] CLBLM_L_X10Y155_SLICE_X13Y155_AO5;
  wire [0:0] CLBLM_L_X10Y155_SLICE_X13Y155_AO6;
  wire [0:0] CLBLM_L_X10Y155_SLICE_X13Y155_A_CY;
  wire [0:0] CLBLM_L_X10Y155_SLICE_X13Y155_A_XOR;
  wire [0:0] CLBLM_L_X10Y155_SLICE_X13Y155_B;
  wire [0:0] CLBLM_L_X10Y155_SLICE_X13Y155_B1;
  wire [0:0] CLBLM_L_X10Y155_SLICE_X13Y155_B2;
  wire [0:0] CLBLM_L_X10Y155_SLICE_X13Y155_B3;
  wire [0:0] CLBLM_L_X10Y155_SLICE_X13Y155_B4;
  wire [0:0] CLBLM_L_X10Y155_SLICE_X13Y155_B5;
  wire [0:0] CLBLM_L_X10Y155_SLICE_X13Y155_B6;
  wire [0:0] CLBLM_L_X10Y155_SLICE_X13Y155_BO5;
  wire [0:0] CLBLM_L_X10Y155_SLICE_X13Y155_BO6;
  wire [0:0] CLBLM_L_X10Y155_SLICE_X13Y155_B_CY;
  wire [0:0] CLBLM_L_X10Y155_SLICE_X13Y155_B_XOR;
  wire [0:0] CLBLM_L_X10Y155_SLICE_X13Y155_C;
  wire [0:0] CLBLM_L_X10Y155_SLICE_X13Y155_C1;
  wire [0:0] CLBLM_L_X10Y155_SLICE_X13Y155_C2;
  wire [0:0] CLBLM_L_X10Y155_SLICE_X13Y155_C3;
  wire [0:0] CLBLM_L_X10Y155_SLICE_X13Y155_C4;
  wire [0:0] CLBLM_L_X10Y155_SLICE_X13Y155_C5;
  wire [0:0] CLBLM_L_X10Y155_SLICE_X13Y155_C6;
  wire [0:0] CLBLM_L_X10Y155_SLICE_X13Y155_CO5;
  wire [0:0] CLBLM_L_X10Y155_SLICE_X13Y155_CO6;
  wire [0:0] CLBLM_L_X10Y155_SLICE_X13Y155_C_CY;
  wire [0:0] CLBLM_L_X10Y155_SLICE_X13Y155_C_XOR;
  wire [0:0] CLBLM_L_X10Y155_SLICE_X13Y155_D;
  wire [0:0] CLBLM_L_X10Y155_SLICE_X13Y155_D1;
  wire [0:0] CLBLM_L_X10Y155_SLICE_X13Y155_D2;
  wire [0:0] CLBLM_L_X10Y155_SLICE_X13Y155_D3;
  wire [0:0] CLBLM_L_X10Y155_SLICE_X13Y155_D4;
  wire [0:0] CLBLM_L_X10Y155_SLICE_X13Y155_D5;
  wire [0:0] CLBLM_L_X10Y155_SLICE_X13Y155_D6;
  wire [0:0] CLBLM_L_X10Y155_SLICE_X13Y155_DO5;
  wire [0:0] CLBLM_L_X10Y155_SLICE_X13Y155_DO6;
  wire [0:0] CLBLM_L_X10Y155_SLICE_X13Y155_D_CY;
  wire [0:0] CLBLM_L_X10Y155_SLICE_X13Y155_D_XOR;
  wire [0:0] CLBLM_L_X12Y145_SLICE_X16Y145_A;
  wire [0:0] CLBLM_L_X12Y145_SLICE_X16Y145_A1;
  wire [0:0] CLBLM_L_X12Y145_SLICE_X16Y145_A2;
  wire [0:0] CLBLM_L_X12Y145_SLICE_X16Y145_A3;
  wire [0:0] CLBLM_L_X12Y145_SLICE_X16Y145_A4;
  wire [0:0] CLBLM_L_X12Y145_SLICE_X16Y145_A5;
  wire [0:0] CLBLM_L_X12Y145_SLICE_X16Y145_A6;
  wire [0:0] CLBLM_L_X12Y145_SLICE_X16Y145_AMUX;
  wire [0:0] CLBLM_L_X12Y145_SLICE_X16Y145_AO5;
  wire [0:0] CLBLM_L_X12Y145_SLICE_X16Y145_AO6;
  wire [0:0] CLBLM_L_X12Y145_SLICE_X16Y145_AQ;
  wire [0:0] CLBLM_L_X12Y145_SLICE_X16Y145_AX;
  wire [0:0] CLBLM_L_X12Y145_SLICE_X16Y145_A_CY;
  wire [0:0] CLBLM_L_X12Y145_SLICE_X16Y145_A_XOR;
  wire [0:0] CLBLM_L_X12Y145_SLICE_X16Y145_B;
  wire [0:0] CLBLM_L_X12Y145_SLICE_X16Y145_B1;
  wire [0:0] CLBLM_L_X12Y145_SLICE_X16Y145_B2;
  wire [0:0] CLBLM_L_X12Y145_SLICE_X16Y145_B3;
  wire [0:0] CLBLM_L_X12Y145_SLICE_X16Y145_B4;
  wire [0:0] CLBLM_L_X12Y145_SLICE_X16Y145_B5;
  wire [0:0] CLBLM_L_X12Y145_SLICE_X16Y145_B6;
  wire [0:0] CLBLM_L_X12Y145_SLICE_X16Y145_BO5;
  wire [0:0] CLBLM_L_X12Y145_SLICE_X16Y145_BO6;
  wire [0:0] CLBLM_L_X12Y145_SLICE_X16Y145_B_CY;
  wire [0:0] CLBLM_L_X12Y145_SLICE_X16Y145_B_XOR;
  wire [0:0] CLBLM_L_X12Y145_SLICE_X16Y145_C;
  wire [0:0] CLBLM_L_X12Y145_SLICE_X16Y145_C1;
  wire [0:0] CLBLM_L_X12Y145_SLICE_X16Y145_C2;
  wire [0:0] CLBLM_L_X12Y145_SLICE_X16Y145_C3;
  wire [0:0] CLBLM_L_X12Y145_SLICE_X16Y145_C4;
  wire [0:0] CLBLM_L_X12Y145_SLICE_X16Y145_C5;
  wire [0:0] CLBLM_L_X12Y145_SLICE_X16Y145_C6;
  wire [0:0] CLBLM_L_X12Y145_SLICE_X16Y145_CE;
  wire [0:0] CLBLM_L_X12Y145_SLICE_X16Y145_CLK;
  wire [0:0] CLBLM_L_X12Y145_SLICE_X16Y145_CO5;
  wire [0:0] CLBLM_L_X12Y145_SLICE_X16Y145_CO6;
  wire [0:0] CLBLM_L_X12Y145_SLICE_X16Y145_C_CY;
  wire [0:0] CLBLM_L_X12Y145_SLICE_X16Y145_C_XOR;
  wire [0:0] CLBLM_L_X12Y145_SLICE_X16Y145_D;
  wire [0:0] CLBLM_L_X12Y145_SLICE_X16Y145_D1;
  wire [0:0] CLBLM_L_X12Y145_SLICE_X16Y145_D2;
  wire [0:0] CLBLM_L_X12Y145_SLICE_X16Y145_D3;
  wire [0:0] CLBLM_L_X12Y145_SLICE_X16Y145_D4;
  wire [0:0] CLBLM_L_X12Y145_SLICE_X16Y145_D5;
  wire [0:0] CLBLM_L_X12Y145_SLICE_X16Y145_D6;
  wire [0:0] CLBLM_L_X12Y145_SLICE_X16Y145_DO5;
  wire [0:0] CLBLM_L_X12Y145_SLICE_X16Y145_DO6;
  wire [0:0] CLBLM_L_X12Y145_SLICE_X16Y145_D_CY;
  wire [0:0] CLBLM_L_X12Y145_SLICE_X16Y145_D_XOR;
  wire [0:0] CLBLM_L_X12Y145_SLICE_X17Y145_A;
  wire [0:0] CLBLM_L_X12Y145_SLICE_X17Y145_A1;
  wire [0:0] CLBLM_L_X12Y145_SLICE_X17Y145_A2;
  wire [0:0] CLBLM_L_X12Y145_SLICE_X17Y145_A3;
  wire [0:0] CLBLM_L_X12Y145_SLICE_X17Y145_A4;
  wire [0:0] CLBLM_L_X12Y145_SLICE_X17Y145_A5;
  wire [0:0] CLBLM_L_X12Y145_SLICE_X17Y145_A6;
  wire [0:0] CLBLM_L_X12Y145_SLICE_X17Y145_AMUX;
  wire [0:0] CLBLM_L_X12Y145_SLICE_X17Y145_AO5;
  wire [0:0] CLBLM_L_X12Y145_SLICE_X17Y145_AO6;
  wire [0:0] CLBLM_L_X12Y145_SLICE_X17Y145_A_CY;
  wire [0:0] CLBLM_L_X12Y145_SLICE_X17Y145_A_XOR;
  wire [0:0] CLBLM_L_X12Y145_SLICE_X17Y145_B;
  wire [0:0] CLBLM_L_X12Y145_SLICE_X17Y145_B1;
  wire [0:0] CLBLM_L_X12Y145_SLICE_X17Y145_B2;
  wire [0:0] CLBLM_L_X12Y145_SLICE_X17Y145_B3;
  wire [0:0] CLBLM_L_X12Y145_SLICE_X17Y145_B4;
  wire [0:0] CLBLM_L_X12Y145_SLICE_X17Y145_B5;
  wire [0:0] CLBLM_L_X12Y145_SLICE_X17Y145_B6;
  wire [0:0] CLBLM_L_X12Y145_SLICE_X17Y145_BO5;
  wire [0:0] CLBLM_L_X12Y145_SLICE_X17Y145_BO6;
  wire [0:0] CLBLM_L_X12Y145_SLICE_X17Y145_B_CY;
  wire [0:0] CLBLM_L_X12Y145_SLICE_X17Y145_B_XOR;
  wire [0:0] CLBLM_L_X12Y145_SLICE_X17Y145_C;
  wire [0:0] CLBLM_L_X12Y145_SLICE_X17Y145_C1;
  wire [0:0] CLBLM_L_X12Y145_SLICE_X17Y145_C2;
  wire [0:0] CLBLM_L_X12Y145_SLICE_X17Y145_C3;
  wire [0:0] CLBLM_L_X12Y145_SLICE_X17Y145_C4;
  wire [0:0] CLBLM_L_X12Y145_SLICE_X17Y145_C5;
  wire [0:0] CLBLM_L_X12Y145_SLICE_X17Y145_C6;
  wire [0:0] CLBLM_L_X12Y145_SLICE_X17Y145_CMUX;
  wire [0:0] CLBLM_L_X12Y145_SLICE_X17Y145_CO5;
  wire [0:0] CLBLM_L_X12Y145_SLICE_X17Y145_CO6;
  wire [0:0] CLBLM_L_X12Y145_SLICE_X17Y145_C_CY;
  wire [0:0] CLBLM_L_X12Y145_SLICE_X17Y145_C_XOR;
  wire [0:0] CLBLM_L_X12Y145_SLICE_X17Y145_D;
  wire [0:0] CLBLM_L_X12Y145_SLICE_X17Y145_D1;
  wire [0:0] CLBLM_L_X12Y145_SLICE_X17Y145_D2;
  wire [0:0] CLBLM_L_X12Y145_SLICE_X17Y145_D3;
  wire [0:0] CLBLM_L_X12Y145_SLICE_X17Y145_D4;
  wire [0:0] CLBLM_L_X12Y145_SLICE_X17Y145_D5;
  wire [0:0] CLBLM_L_X12Y145_SLICE_X17Y145_D6;
  wire [0:0] CLBLM_L_X12Y145_SLICE_X17Y145_DO5;
  wire [0:0] CLBLM_L_X12Y145_SLICE_X17Y145_DO6;
  wire [0:0] CLBLM_L_X12Y145_SLICE_X17Y145_D_CY;
  wire [0:0] CLBLM_L_X12Y145_SLICE_X17Y145_D_XOR;
  wire [0:0] CLBLM_L_X12Y146_SLICE_X16Y146_A;
  wire [0:0] CLBLM_L_X12Y146_SLICE_X16Y146_A1;
  wire [0:0] CLBLM_L_X12Y146_SLICE_X16Y146_A2;
  wire [0:0] CLBLM_L_X12Y146_SLICE_X16Y146_A3;
  wire [0:0] CLBLM_L_X12Y146_SLICE_X16Y146_A4;
  wire [0:0] CLBLM_L_X12Y146_SLICE_X16Y146_A5;
  wire [0:0] CLBLM_L_X12Y146_SLICE_X16Y146_A6;
  wire [0:0] CLBLM_L_X12Y146_SLICE_X16Y146_AMUX;
  wire [0:0] CLBLM_L_X12Y146_SLICE_X16Y146_AO5;
  wire [0:0] CLBLM_L_X12Y146_SLICE_X16Y146_AO6;
  wire [0:0] CLBLM_L_X12Y146_SLICE_X16Y146_AQ;
  wire [0:0] CLBLM_L_X12Y146_SLICE_X16Y146_AX;
  wire [0:0] CLBLM_L_X12Y146_SLICE_X16Y146_A_CY;
  wire [0:0] CLBLM_L_X12Y146_SLICE_X16Y146_A_XOR;
  wire [0:0] CLBLM_L_X12Y146_SLICE_X16Y146_B;
  wire [0:0] CLBLM_L_X12Y146_SLICE_X16Y146_B1;
  wire [0:0] CLBLM_L_X12Y146_SLICE_X16Y146_B2;
  wire [0:0] CLBLM_L_X12Y146_SLICE_X16Y146_B3;
  wire [0:0] CLBLM_L_X12Y146_SLICE_X16Y146_B4;
  wire [0:0] CLBLM_L_X12Y146_SLICE_X16Y146_B5;
  wire [0:0] CLBLM_L_X12Y146_SLICE_X16Y146_B6;
  wire [0:0] CLBLM_L_X12Y146_SLICE_X16Y146_BO5;
  wire [0:0] CLBLM_L_X12Y146_SLICE_X16Y146_BO6;
  wire [0:0] CLBLM_L_X12Y146_SLICE_X16Y146_BQ;
  wire [0:0] CLBLM_L_X12Y146_SLICE_X16Y146_BX;
  wire [0:0] CLBLM_L_X12Y146_SLICE_X16Y146_B_CY;
  wire [0:0] CLBLM_L_X12Y146_SLICE_X16Y146_B_XOR;
  wire [0:0] CLBLM_L_X12Y146_SLICE_X16Y146_C;
  wire [0:0] CLBLM_L_X12Y146_SLICE_X16Y146_C1;
  wire [0:0] CLBLM_L_X12Y146_SLICE_X16Y146_C2;
  wire [0:0] CLBLM_L_X12Y146_SLICE_X16Y146_C3;
  wire [0:0] CLBLM_L_X12Y146_SLICE_X16Y146_C4;
  wire [0:0] CLBLM_L_X12Y146_SLICE_X16Y146_C5;
  wire [0:0] CLBLM_L_X12Y146_SLICE_X16Y146_C6;
  wire [0:0] CLBLM_L_X12Y146_SLICE_X16Y146_CE;
  wire [0:0] CLBLM_L_X12Y146_SLICE_X16Y146_CLK;
  wire [0:0] CLBLM_L_X12Y146_SLICE_X16Y146_CO5;
  wire [0:0] CLBLM_L_X12Y146_SLICE_X16Y146_CO6;
  wire [0:0] CLBLM_L_X12Y146_SLICE_X16Y146_CQ;
  wire [0:0] CLBLM_L_X12Y146_SLICE_X16Y146_CX;
  wire [0:0] CLBLM_L_X12Y146_SLICE_X16Y146_C_CY;
  wire [0:0] CLBLM_L_X12Y146_SLICE_X16Y146_C_XOR;
  wire [0:0] CLBLM_L_X12Y146_SLICE_X16Y146_D;
  wire [0:0] CLBLM_L_X12Y146_SLICE_X16Y146_D1;
  wire [0:0] CLBLM_L_X12Y146_SLICE_X16Y146_D2;
  wire [0:0] CLBLM_L_X12Y146_SLICE_X16Y146_D3;
  wire [0:0] CLBLM_L_X12Y146_SLICE_X16Y146_D4;
  wire [0:0] CLBLM_L_X12Y146_SLICE_X16Y146_D5;
  wire [0:0] CLBLM_L_X12Y146_SLICE_X16Y146_D6;
  wire [0:0] CLBLM_L_X12Y146_SLICE_X16Y146_DO5;
  wire [0:0] CLBLM_L_X12Y146_SLICE_X16Y146_DO6;
  wire [0:0] CLBLM_L_X12Y146_SLICE_X16Y146_DQ;
  wire [0:0] CLBLM_L_X12Y146_SLICE_X16Y146_DX;
  wire [0:0] CLBLM_L_X12Y146_SLICE_X16Y146_D_CY;
  wire [0:0] CLBLM_L_X12Y146_SLICE_X16Y146_D_XOR;
  wire [0:0] CLBLM_L_X12Y146_SLICE_X17Y146_A;
  wire [0:0] CLBLM_L_X12Y146_SLICE_X17Y146_A1;
  wire [0:0] CLBLM_L_X12Y146_SLICE_X17Y146_A2;
  wire [0:0] CLBLM_L_X12Y146_SLICE_X17Y146_A3;
  wire [0:0] CLBLM_L_X12Y146_SLICE_X17Y146_A4;
  wire [0:0] CLBLM_L_X12Y146_SLICE_X17Y146_A5;
  wire [0:0] CLBLM_L_X12Y146_SLICE_X17Y146_A6;
  wire [0:0] CLBLM_L_X12Y146_SLICE_X17Y146_AO5;
  wire [0:0] CLBLM_L_X12Y146_SLICE_X17Y146_AO6;
  wire [0:0] CLBLM_L_X12Y146_SLICE_X17Y146_AQ;
  wire [0:0] CLBLM_L_X12Y146_SLICE_X17Y146_A_CY;
  wire [0:0] CLBLM_L_X12Y146_SLICE_X17Y146_A_XOR;
  wire [0:0] CLBLM_L_X12Y146_SLICE_X17Y146_B;
  wire [0:0] CLBLM_L_X12Y146_SLICE_X17Y146_B1;
  wire [0:0] CLBLM_L_X12Y146_SLICE_X17Y146_B2;
  wire [0:0] CLBLM_L_X12Y146_SLICE_X17Y146_B3;
  wire [0:0] CLBLM_L_X12Y146_SLICE_X17Y146_B4;
  wire [0:0] CLBLM_L_X12Y146_SLICE_X17Y146_B5;
  wire [0:0] CLBLM_L_X12Y146_SLICE_X17Y146_B6;
  wire [0:0] CLBLM_L_X12Y146_SLICE_X17Y146_BO5;
  wire [0:0] CLBLM_L_X12Y146_SLICE_X17Y146_BO6;
  wire [0:0] CLBLM_L_X12Y146_SLICE_X17Y146_B_CY;
  wire [0:0] CLBLM_L_X12Y146_SLICE_X17Y146_B_XOR;
  wire [0:0] CLBLM_L_X12Y146_SLICE_X17Y146_C;
  wire [0:0] CLBLM_L_X12Y146_SLICE_X17Y146_C1;
  wire [0:0] CLBLM_L_X12Y146_SLICE_X17Y146_C2;
  wire [0:0] CLBLM_L_X12Y146_SLICE_X17Y146_C3;
  wire [0:0] CLBLM_L_X12Y146_SLICE_X17Y146_C4;
  wire [0:0] CLBLM_L_X12Y146_SLICE_X17Y146_C5;
  wire [0:0] CLBLM_L_X12Y146_SLICE_X17Y146_C6;
  wire [0:0] CLBLM_L_X12Y146_SLICE_X17Y146_CLK;
  wire [0:0] CLBLM_L_X12Y146_SLICE_X17Y146_CMUX;
  wire [0:0] CLBLM_L_X12Y146_SLICE_X17Y146_CO5;
  wire [0:0] CLBLM_L_X12Y146_SLICE_X17Y146_CO6;
  wire [0:0] CLBLM_L_X12Y146_SLICE_X17Y146_C_CY;
  wire [0:0] CLBLM_L_X12Y146_SLICE_X17Y146_C_XOR;
  wire [0:0] CLBLM_L_X12Y146_SLICE_X17Y146_D;
  wire [0:0] CLBLM_L_X12Y146_SLICE_X17Y146_D1;
  wire [0:0] CLBLM_L_X12Y146_SLICE_X17Y146_D2;
  wire [0:0] CLBLM_L_X12Y146_SLICE_X17Y146_D3;
  wire [0:0] CLBLM_L_X12Y146_SLICE_X17Y146_D4;
  wire [0:0] CLBLM_L_X12Y146_SLICE_X17Y146_D5;
  wire [0:0] CLBLM_L_X12Y146_SLICE_X17Y146_D6;
  wire [0:0] CLBLM_L_X12Y146_SLICE_X17Y146_DO5;
  wire [0:0] CLBLM_L_X12Y146_SLICE_X17Y146_DO6;
  wire [0:0] CLBLM_L_X12Y146_SLICE_X17Y146_D_CY;
  wire [0:0] CLBLM_L_X12Y146_SLICE_X17Y146_D_XOR;
  wire [0:0] CLBLM_L_X12Y147_SLICE_X16Y147_A;
  wire [0:0] CLBLM_L_X12Y147_SLICE_X16Y147_A1;
  wire [0:0] CLBLM_L_X12Y147_SLICE_X16Y147_A2;
  wire [0:0] CLBLM_L_X12Y147_SLICE_X16Y147_A3;
  wire [0:0] CLBLM_L_X12Y147_SLICE_X16Y147_A4;
  wire [0:0] CLBLM_L_X12Y147_SLICE_X16Y147_A5;
  wire [0:0] CLBLM_L_X12Y147_SLICE_X16Y147_A6;
  wire [0:0] CLBLM_L_X12Y147_SLICE_X16Y147_AMUX;
  wire [0:0] CLBLM_L_X12Y147_SLICE_X16Y147_AO5;
  wire [0:0] CLBLM_L_X12Y147_SLICE_X16Y147_AO6;
  wire [0:0] CLBLM_L_X12Y147_SLICE_X16Y147_A_CY;
  wire [0:0] CLBLM_L_X12Y147_SLICE_X16Y147_A_XOR;
  wire [0:0] CLBLM_L_X12Y147_SLICE_X16Y147_B;
  wire [0:0] CLBLM_L_X12Y147_SLICE_X16Y147_B1;
  wire [0:0] CLBLM_L_X12Y147_SLICE_X16Y147_B2;
  wire [0:0] CLBLM_L_X12Y147_SLICE_X16Y147_B3;
  wire [0:0] CLBLM_L_X12Y147_SLICE_X16Y147_B4;
  wire [0:0] CLBLM_L_X12Y147_SLICE_X16Y147_B5;
  wire [0:0] CLBLM_L_X12Y147_SLICE_X16Y147_B6;
  wire [0:0] CLBLM_L_X12Y147_SLICE_X16Y147_BO5;
  wire [0:0] CLBLM_L_X12Y147_SLICE_X16Y147_BO6;
  wire [0:0] CLBLM_L_X12Y147_SLICE_X16Y147_B_CY;
  wire [0:0] CLBLM_L_X12Y147_SLICE_X16Y147_B_XOR;
  wire [0:0] CLBLM_L_X12Y147_SLICE_X16Y147_C;
  wire [0:0] CLBLM_L_X12Y147_SLICE_X16Y147_C1;
  wire [0:0] CLBLM_L_X12Y147_SLICE_X16Y147_C2;
  wire [0:0] CLBLM_L_X12Y147_SLICE_X16Y147_C3;
  wire [0:0] CLBLM_L_X12Y147_SLICE_X16Y147_C4;
  wire [0:0] CLBLM_L_X12Y147_SLICE_X16Y147_C5;
  wire [0:0] CLBLM_L_X12Y147_SLICE_X16Y147_C6;
  wire [0:0] CLBLM_L_X12Y147_SLICE_X16Y147_CMUX;
  wire [0:0] CLBLM_L_X12Y147_SLICE_X16Y147_CO5;
  wire [0:0] CLBLM_L_X12Y147_SLICE_X16Y147_CO6;
  wire [0:0] CLBLM_L_X12Y147_SLICE_X16Y147_C_CY;
  wire [0:0] CLBLM_L_X12Y147_SLICE_X16Y147_C_XOR;
  wire [0:0] CLBLM_L_X12Y147_SLICE_X16Y147_D;
  wire [0:0] CLBLM_L_X12Y147_SLICE_X16Y147_D1;
  wire [0:0] CLBLM_L_X12Y147_SLICE_X16Y147_D2;
  wire [0:0] CLBLM_L_X12Y147_SLICE_X16Y147_D3;
  wire [0:0] CLBLM_L_X12Y147_SLICE_X16Y147_D4;
  wire [0:0] CLBLM_L_X12Y147_SLICE_X16Y147_D5;
  wire [0:0] CLBLM_L_X12Y147_SLICE_X16Y147_D6;
  wire [0:0] CLBLM_L_X12Y147_SLICE_X16Y147_DMUX;
  wire [0:0] CLBLM_L_X12Y147_SLICE_X16Y147_DO5;
  wire [0:0] CLBLM_L_X12Y147_SLICE_X16Y147_DO6;
  wire [0:0] CLBLM_L_X12Y147_SLICE_X16Y147_D_CY;
  wire [0:0] CLBLM_L_X12Y147_SLICE_X16Y147_D_XOR;
  wire [0:0] CLBLM_L_X12Y147_SLICE_X17Y147_A;
  wire [0:0] CLBLM_L_X12Y147_SLICE_X17Y147_A1;
  wire [0:0] CLBLM_L_X12Y147_SLICE_X17Y147_A2;
  wire [0:0] CLBLM_L_X12Y147_SLICE_X17Y147_A3;
  wire [0:0] CLBLM_L_X12Y147_SLICE_X17Y147_A4;
  wire [0:0] CLBLM_L_X12Y147_SLICE_X17Y147_A5;
  wire [0:0] CLBLM_L_X12Y147_SLICE_X17Y147_A6;
  wire [0:0] CLBLM_L_X12Y147_SLICE_X17Y147_AMUX;
  wire [0:0] CLBLM_L_X12Y147_SLICE_X17Y147_AO5;
  wire [0:0] CLBLM_L_X12Y147_SLICE_X17Y147_AO6;
  wire [0:0] CLBLM_L_X12Y147_SLICE_X17Y147_A_CY;
  wire [0:0] CLBLM_L_X12Y147_SLICE_X17Y147_A_XOR;
  wire [0:0] CLBLM_L_X12Y147_SLICE_X17Y147_B;
  wire [0:0] CLBLM_L_X12Y147_SLICE_X17Y147_B1;
  wire [0:0] CLBLM_L_X12Y147_SLICE_X17Y147_B2;
  wire [0:0] CLBLM_L_X12Y147_SLICE_X17Y147_B3;
  wire [0:0] CLBLM_L_X12Y147_SLICE_X17Y147_B4;
  wire [0:0] CLBLM_L_X12Y147_SLICE_X17Y147_B5;
  wire [0:0] CLBLM_L_X12Y147_SLICE_X17Y147_B6;
  wire [0:0] CLBLM_L_X12Y147_SLICE_X17Y147_BO5;
  wire [0:0] CLBLM_L_X12Y147_SLICE_X17Y147_BO6;
  wire [0:0] CLBLM_L_X12Y147_SLICE_X17Y147_B_CY;
  wire [0:0] CLBLM_L_X12Y147_SLICE_X17Y147_B_XOR;
  wire [0:0] CLBLM_L_X12Y147_SLICE_X17Y147_C;
  wire [0:0] CLBLM_L_X12Y147_SLICE_X17Y147_C1;
  wire [0:0] CLBLM_L_X12Y147_SLICE_X17Y147_C2;
  wire [0:0] CLBLM_L_X12Y147_SLICE_X17Y147_C3;
  wire [0:0] CLBLM_L_X12Y147_SLICE_X17Y147_C4;
  wire [0:0] CLBLM_L_X12Y147_SLICE_X17Y147_C5;
  wire [0:0] CLBLM_L_X12Y147_SLICE_X17Y147_C6;
  wire [0:0] CLBLM_L_X12Y147_SLICE_X17Y147_CO5;
  wire [0:0] CLBLM_L_X12Y147_SLICE_X17Y147_CO6;
  wire [0:0] CLBLM_L_X12Y147_SLICE_X17Y147_C_CY;
  wire [0:0] CLBLM_L_X12Y147_SLICE_X17Y147_C_XOR;
  wire [0:0] CLBLM_L_X12Y147_SLICE_X17Y147_D;
  wire [0:0] CLBLM_L_X12Y147_SLICE_X17Y147_D1;
  wire [0:0] CLBLM_L_X12Y147_SLICE_X17Y147_D2;
  wire [0:0] CLBLM_L_X12Y147_SLICE_X17Y147_D3;
  wire [0:0] CLBLM_L_X12Y147_SLICE_X17Y147_D4;
  wire [0:0] CLBLM_L_X12Y147_SLICE_X17Y147_D5;
  wire [0:0] CLBLM_L_X12Y147_SLICE_X17Y147_D6;
  wire [0:0] CLBLM_L_X12Y147_SLICE_X17Y147_DO5;
  wire [0:0] CLBLM_L_X12Y147_SLICE_X17Y147_DO6;
  wire [0:0] CLBLM_L_X12Y147_SLICE_X17Y147_D_CY;
  wire [0:0] CLBLM_L_X12Y147_SLICE_X17Y147_D_XOR;
  wire [0:0] CLBLM_L_X12Y148_SLICE_X16Y148_A;
  wire [0:0] CLBLM_L_X12Y148_SLICE_X16Y148_A1;
  wire [0:0] CLBLM_L_X12Y148_SLICE_X16Y148_A2;
  wire [0:0] CLBLM_L_X12Y148_SLICE_X16Y148_A3;
  wire [0:0] CLBLM_L_X12Y148_SLICE_X16Y148_A4;
  wire [0:0] CLBLM_L_X12Y148_SLICE_X16Y148_A5;
  wire [0:0] CLBLM_L_X12Y148_SLICE_X16Y148_A6;
  wire [0:0] CLBLM_L_X12Y148_SLICE_X16Y148_AMUX;
  wire [0:0] CLBLM_L_X12Y148_SLICE_X16Y148_AO5;
  wire [0:0] CLBLM_L_X12Y148_SLICE_X16Y148_AO6;
  wire [0:0] CLBLM_L_X12Y148_SLICE_X16Y148_A_CY;
  wire [0:0] CLBLM_L_X12Y148_SLICE_X16Y148_A_XOR;
  wire [0:0] CLBLM_L_X12Y148_SLICE_X16Y148_B;
  wire [0:0] CLBLM_L_X12Y148_SLICE_X16Y148_B1;
  wire [0:0] CLBLM_L_X12Y148_SLICE_X16Y148_B2;
  wire [0:0] CLBLM_L_X12Y148_SLICE_X16Y148_B3;
  wire [0:0] CLBLM_L_X12Y148_SLICE_X16Y148_B4;
  wire [0:0] CLBLM_L_X12Y148_SLICE_X16Y148_B5;
  wire [0:0] CLBLM_L_X12Y148_SLICE_X16Y148_B6;
  wire [0:0] CLBLM_L_X12Y148_SLICE_X16Y148_BO5;
  wire [0:0] CLBLM_L_X12Y148_SLICE_X16Y148_BO6;
  wire [0:0] CLBLM_L_X12Y148_SLICE_X16Y148_B_CY;
  wire [0:0] CLBLM_L_X12Y148_SLICE_X16Y148_B_XOR;
  wire [0:0] CLBLM_L_X12Y148_SLICE_X16Y148_C;
  wire [0:0] CLBLM_L_X12Y148_SLICE_X16Y148_C1;
  wire [0:0] CLBLM_L_X12Y148_SLICE_X16Y148_C2;
  wire [0:0] CLBLM_L_X12Y148_SLICE_X16Y148_C3;
  wire [0:0] CLBLM_L_X12Y148_SLICE_X16Y148_C4;
  wire [0:0] CLBLM_L_X12Y148_SLICE_X16Y148_C5;
  wire [0:0] CLBLM_L_X12Y148_SLICE_X16Y148_C6;
  wire [0:0] CLBLM_L_X12Y148_SLICE_X16Y148_CO5;
  wire [0:0] CLBLM_L_X12Y148_SLICE_X16Y148_CO6;
  wire [0:0] CLBLM_L_X12Y148_SLICE_X16Y148_C_CY;
  wire [0:0] CLBLM_L_X12Y148_SLICE_X16Y148_C_XOR;
  wire [0:0] CLBLM_L_X12Y148_SLICE_X16Y148_D;
  wire [0:0] CLBLM_L_X12Y148_SLICE_X16Y148_D1;
  wire [0:0] CLBLM_L_X12Y148_SLICE_X16Y148_D2;
  wire [0:0] CLBLM_L_X12Y148_SLICE_X16Y148_D3;
  wire [0:0] CLBLM_L_X12Y148_SLICE_X16Y148_D4;
  wire [0:0] CLBLM_L_X12Y148_SLICE_X16Y148_D5;
  wire [0:0] CLBLM_L_X12Y148_SLICE_X16Y148_D6;
  wire [0:0] CLBLM_L_X12Y148_SLICE_X16Y148_DO5;
  wire [0:0] CLBLM_L_X12Y148_SLICE_X16Y148_DO6;
  wire [0:0] CLBLM_L_X12Y148_SLICE_X16Y148_D_CY;
  wire [0:0] CLBLM_L_X12Y148_SLICE_X16Y148_D_XOR;
  wire [0:0] CLBLM_L_X12Y148_SLICE_X17Y148_A;
  wire [0:0] CLBLM_L_X12Y148_SLICE_X17Y148_A1;
  wire [0:0] CLBLM_L_X12Y148_SLICE_X17Y148_A2;
  wire [0:0] CLBLM_L_X12Y148_SLICE_X17Y148_A3;
  wire [0:0] CLBLM_L_X12Y148_SLICE_X17Y148_A4;
  wire [0:0] CLBLM_L_X12Y148_SLICE_X17Y148_A5;
  wire [0:0] CLBLM_L_X12Y148_SLICE_X17Y148_A6;
  wire [0:0] CLBLM_L_X12Y148_SLICE_X17Y148_AO5;
  wire [0:0] CLBLM_L_X12Y148_SLICE_X17Y148_AO6;
  wire [0:0] CLBLM_L_X12Y148_SLICE_X17Y148_A_CY;
  wire [0:0] CLBLM_L_X12Y148_SLICE_X17Y148_A_XOR;
  wire [0:0] CLBLM_L_X12Y148_SLICE_X17Y148_B;
  wire [0:0] CLBLM_L_X12Y148_SLICE_X17Y148_B1;
  wire [0:0] CLBLM_L_X12Y148_SLICE_X17Y148_B2;
  wire [0:0] CLBLM_L_X12Y148_SLICE_X17Y148_B3;
  wire [0:0] CLBLM_L_X12Y148_SLICE_X17Y148_B4;
  wire [0:0] CLBLM_L_X12Y148_SLICE_X17Y148_B5;
  wire [0:0] CLBLM_L_X12Y148_SLICE_X17Y148_B6;
  wire [0:0] CLBLM_L_X12Y148_SLICE_X17Y148_BO5;
  wire [0:0] CLBLM_L_X12Y148_SLICE_X17Y148_BO6;
  wire [0:0] CLBLM_L_X12Y148_SLICE_X17Y148_B_CY;
  wire [0:0] CLBLM_L_X12Y148_SLICE_X17Y148_B_XOR;
  wire [0:0] CLBLM_L_X12Y148_SLICE_X17Y148_C;
  wire [0:0] CLBLM_L_X12Y148_SLICE_X17Y148_C1;
  wire [0:0] CLBLM_L_X12Y148_SLICE_X17Y148_C2;
  wire [0:0] CLBLM_L_X12Y148_SLICE_X17Y148_C3;
  wire [0:0] CLBLM_L_X12Y148_SLICE_X17Y148_C4;
  wire [0:0] CLBLM_L_X12Y148_SLICE_X17Y148_C5;
  wire [0:0] CLBLM_L_X12Y148_SLICE_X17Y148_C6;
  wire [0:0] CLBLM_L_X12Y148_SLICE_X17Y148_CO5;
  wire [0:0] CLBLM_L_X12Y148_SLICE_X17Y148_CO6;
  wire [0:0] CLBLM_L_X12Y148_SLICE_X17Y148_C_CY;
  wire [0:0] CLBLM_L_X12Y148_SLICE_X17Y148_C_XOR;
  wire [0:0] CLBLM_L_X12Y148_SLICE_X17Y148_D;
  wire [0:0] CLBLM_L_X12Y148_SLICE_X17Y148_D1;
  wire [0:0] CLBLM_L_X12Y148_SLICE_X17Y148_D2;
  wire [0:0] CLBLM_L_X12Y148_SLICE_X17Y148_D3;
  wire [0:0] CLBLM_L_X12Y148_SLICE_X17Y148_D4;
  wire [0:0] CLBLM_L_X12Y148_SLICE_X17Y148_D5;
  wire [0:0] CLBLM_L_X12Y148_SLICE_X17Y148_D6;
  wire [0:0] CLBLM_L_X12Y148_SLICE_X17Y148_DO5;
  wire [0:0] CLBLM_L_X12Y148_SLICE_X17Y148_DO6;
  wire [0:0] CLBLM_L_X12Y148_SLICE_X17Y148_D_CY;
  wire [0:0] CLBLM_L_X12Y148_SLICE_X17Y148_D_XOR;
  wire [0:0] CLBLM_L_X12Y149_SLICE_X16Y149_A;
  wire [0:0] CLBLM_L_X12Y149_SLICE_X16Y149_A1;
  wire [0:0] CLBLM_L_X12Y149_SLICE_X16Y149_A2;
  wire [0:0] CLBLM_L_X12Y149_SLICE_X16Y149_A3;
  wire [0:0] CLBLM_L_X12Y149_SLICE_X16Y149_A4;
  wire [0:0] CLBLM_L_X12Y149_SLICE_X16Y149_A5;
  wire [0:0] CLBLM_L_X12Y149_SLICE_X16Y149_A6;
  wire [0:0] CLBLM_L_X12Y149_SLICE_X16Y149_AO5;
  wire [0:0] CLBLM_L_X12Y149_SLICE_X16Y149_AO6;
  wire [0:0] CLBLM_L_X12Y149_SLICE_X16Y149_A_CY;
  wire [0:0] CLBLM_L_X12Y149_SLICE_X16Y149_A_XOR;
  wire [0:0] CLBLM_L_X12Y149_SLICE_X16Y149_B;
  wire [0:0] CLBLM_L_X12Y149_SLICE_X16Y149_B1;
  wire [0:0] CLBLM_L_X12Y149_SLICE_X16Y149_B2;
  wire [0:0] CLBLM_L_X12Y149_SLICE_X16Y149_B3;
  wire [0:0] CLBLM_L_X12Y149_SLICE_X16Y149_B4;
  wire [0:0] CLBLM_L_X12Y149_SLICE_X16Y149_B5;
  wire [0:0] CLBLM_L_X12Y149_SLICE_X16Y149_B6;
  wire [0:0] CLBLM_L_X12Y149_SLICE_X16Y149_BO5;
  wire [0:0] CLBLM_L_X12Y149_SLICE_X16Y149_BO6;
  wire [0:0] CLBLM_L_X12Y149_SLICE_X16Y149_B_CY;
  wire [0:0] CLBLM_L_X12Y149_SLICE_X16Y149_B_XOR;
  wire [0:0] CLBLM_L_X12Y149_SLICE_X16Y149_C;
  wire [0:0] CLBLM_L_X12Y149_SLICE_X16Y149_C1;
  wire [0:0] CLBLM_L_X12Y149_SLICE_X16Y149_C2;
  wire [0:0] CLBLM_L_X12Y149_SLICE_X16Y149_C3;
  wire [0:0] CLBLM_L_X12Y149_SLICE_X16Y149_C4;
  wire [0:0] CLBLM_L_X12Y149_SLICE_X16Y149_C5;
  wire [0:0] CLBLM_L_X12Y149_SLICE_X16Y149_C6;
  wire [0:0] CLBLM_L_X12Y149_SLICE_X16Y149_CO5;
  wire [0:0] CLBLM_L_X12Y149_SLICE_X16Y149_CO6;
  wire [0:0] CLBLM_L_X12Y149_SLICE_X16Y149_C_CY;
  wire [0:0] CLBLM_L_X12Y149_SLICE_X16Y149_C_XOR;
  wire [0:0] CLBLM_L_X12Y149_SLICE_X16Y149_D;
  wire [0:0] CLBLM_L_X12Y149_SLICE_X16Y149_D1;
  wire [0:0] CLBLM_L_X12Y149_SLICE_X16Y149_D2;
  wire [0:0] CLBLM_L_X12Y149_SLICE_X16Y149_D3;
  wire [0:0] CLBLM_L_X12Y149_SLICE_X16Y149_D4;
  wire [0:0] CLBLM_L_X12Y149_SLICE_X16Y149_D5;
  wire [0:0] CLBLM_L_X12Y149_SLICE_X16Y149_D6;
  wire [0:0] CLBLM_L_X12Y149_SLICE_X16Y149_DO5;
  wire [0:0] CLBLM_L_X12Y149_SLICE_X16Y149_DO6;
  wire [0:0] CLBLM_L_X12Y149_SLICE_X16Y149_D_CY;
  wire [0:0] CLBLM_L_X12Y149_SLICE_X16Y149_D_XOR;
  wire [0:0] CLBLM_L_X12Y149_SLICE_X17Y149_A;
  wire [0:0] CLBLM_L_X12Y149_SLICE_X17Y149_A1;
  wire [0:0] CLBLM_L_X12Y149_SLICE_X17Y149_A2;
  wire [0:0] CLBLM_L_X12Y149_SLICE_X17Y149_A3;
  wire [0:0] CLBLM_L_X12Y149_SLICE_X17Y149_A4;
  wire [0:0] CLBLM_L_X12Y149_SLICE_X17Y149_A5;
  wire [0:0] CLBLM_L_X12Y149_SLICE_X17Y149_A6;
  wire [0:0] CLBLM_L_X12Y149_SLICE_X17Y149_AMUX;
  wire [0:0] CLBLM_L_X12Y149_SLICE_X17Y149_AO5;
  wire [0:0] CLBLM_L_X12Y149_SLICE_X17Y149_AO6;
  wire [0:0] CLBLM_L_X12Y149_SLICE_X17Y149_A_CY;
  wire [0:0] CLBLM_L_X12Y149_SLICE_X17Y149_A_XOR;
  wire [0:0] CLBLM_L_X12Y149_SLICE_X17Y149_B;
  wire [0:0] CLBLM_L_X12Y149_SLICE_X17Y149_B1;
  wire [0:0] CLBLM_L_X12Y149_SLICE_X17Y149_B2;
  wire [0:0] CLBLM_L_X12Y149_SLICE_X17Y149_B3;
  wire [0:0] CLBLM_L_X12Y149_SLICE_X17Y149_B4;
  wire [0:0] CLBLM_L_X12Y149_SLICE_X17Y149_B5;
  wire [0:0] CLBLM_L_X12Y149_SLICE_X17Y149_B6;
  wire [0:0] CLBLM_L_X12Y149_SLICE_X17Y149_BMUX;
  wire [0:0] CLBLM_L_X12Y149_SLICE_X17Y149_BO5;
  wire [0:0] CLBLM_L_X12Y149_SLICE_X17Y149_BO6;
  wire [0:0] CLBLM_L_X12Y149_SLICE_X17Y149_B_CY;
  wire [0:0] CLBLM_L_X12Y149_SLICE_X17Y149_B_XOR;
  wire [0:0] CLBLM_L_X12Y149_SLICE_X17Y149_C;
  wire [0:0] CLBLM_L_X12Y149_SLICE_X17Y149_C1;
  wire [0:0] CLBLM_L_X12Y149_SLICE_X17Y149_C2;
  wire [0:0] CLBLM_L_X12Y149_SLICE_X17Y149_C3;
  wire [0:0] CLBLM_L_X12Y149_SLICE_X17Y149_C4;
  wire [0:0] CLBLM_L_X12Y149_SLICE_X17Y149_C5;
  wire [0:0] CLBLM_L_X12Y149_SLICE_X17Y149_C6;
  wire [0:0] CLBLM_L_X12Y149_SLICE_X17Y149_CO5;
  wire [0:0] CLBLM_L_X12Y149_SLICE_X17Y149_CO6;
  wire [0:0] CLBLM_L_X12Y149_SLICE_X17Y149_C_CY;
  wire [0:0] CLBLM_L_X12Y149_SLICE_X17Y149_C_XOR;
  wire [0:0] CLBLM_L_X12Y149_SLICE_X17Y149_D;
  wire [0:0] CLBLM_L_X12Y149_SLICE_X17Y149_D1;
  wire [0:0] CLBLM_L_X12Y149_SLICE_X17Y149_D2;
  wire [0:0] CLBLM_L_X12Y149_SLICE_X17Y149_D3;
  wire [0:0] CLBLM_L_X12Y149_SLICE_X17Y149_D4;
  wire [0:0] CLBLM_L_X12Y149_SLICE_X17Y149_D5;
  wire [0:0] CLBLM_L_X12Y149_SLICE_X17Y149_D6;
  wire [0:0] CLBLM_L_X12Y149_SLICE_X17Y149_DMUX;
  wire [0:0] CLBLM_L_X12Y149_SLICE_X17Y149_DO5;
  wire [0:0] CLBLM_L_X12Y149_SLICE_X17Y149_DO6;
  wire [0:0] CLBLM_L_X12Y149_SLICE_X17Y149_D_CY;
  wire [0:0] CLBLM_L_X12Y149_SLICE_X17Y149_D_XOR;
  wire [0:0] CLBLM_L_X12Y150_SLICE_X16Y150_A;
  wire [0:0] CLBLM_L_X12Y150_SLICE_X16Y150_A1;
  wire [0:0] CLBLM_L_X12Y150_SLICE_X16Y150_A2;
  wire [0:0] CLBLM_L_X12Y150_SLICE_X16Y150_A3;
  wire [0:0] CLBLM_L_X12Y150_SLICE_X16Y150_A4;
  wire [0:0] CLBLM_L_X12Y150_SLICE_X16Y150_A5;
  wire [0:0] CLBLM_L_X12Y150_SLICE_X16Y150_A6;
  wire [0:0] CLBLM_L_X12Y150_SLICE_X16Y150_AMUX;
  wire [0:0] CLBLM_L_X12Y150_SLICE_X16Y150_AO5;
  wire [0:0] CLBLM_L_X12Y150_SLICE_X16Y150_AO6;
  wire [0:0] CLBLM_L_X12Y150_SLICE_X16Y150_A_CY;
  wire [0:0] CLBLM_L_X12Y150_SLICE_X16Y150_A_XOR;
  wire [0:0] CLBLM_L_X12Y150_SLICE_X16Y150_B;
  wire [0:0] CLBLM_L_X12Y150_SLICE_X16Y150_B1;
  wire [0:0] CLBLM_L_X12Y150_SLICE_X16Y150_B2;
  wire [0:0] CLBLM_L_X12Y150_SLICE_X16Y150_B3;
  wire [0:0] CLBLM_L_X12Y150_SLICE_X16Y150_B4;
  wire [0:0] CLBLM_L_X12Y150_SLICE_X16Y150_B5;
  wire [0:0] CLBLM_L_X12Y150_SLICE_X16Y150_B6;
  wire [0:0] CLBLM_L_X12Y150_SLICE_X16Y150_BO5;
  wire [0:0] CLBLM_L_X12Y150_SLICE_X16Y150_BO6;
  wire [0:0] CLBLM_L_X12Y150_SLICE_X16Y150_B_CY;
  wire [0:0] CLBLM_L_X12Y150_SLICE_X16Y150_B_XOR;
  wire [0:0] CLBLM_L_X12Y150_SLICE_X16Y150_C;
  wire [0:0] CLBLM_L_X12Y150_SLICE_X16Y150_C1;
  wire [0:0] CLBLM_L_X12Y150_SLICE_X16Y150_C2;
  wire [0:0] CLBLM_L_X12Y150_SLICE_X16Y150_C3;
  wire [0:0] CLBLM_L_X12Y150_SLICE_X16Y150_C4;
  wire [0:0] CLBLM_L_X12Y150_SLICE_X16Y150_C5;
  wire [0:0] CLBLM_L_X12Y150_SLICE_X16Y150_C6;
  wire [0:0] CLBLM_L_X12Y150_SLICE_X16Y150_CO5;
  wire [0:0] CLBLM_L_X12Y150_SLICE_X16Y150_CO6;
  wire [0:0] CLBLM_L_X12Y150_SLICE_X16Y150_C_CY;
  wire [0:0] CLBLM_L_X12Y150_SLICE_X16Y150_C_XOR;
  wire [0:0] CLBLM_L_X12Y150_SLICE_X16Y150_D;
  wire [0:0] CLBLM_L_X12Y150_SLICE_X16Y150_D1;
  wire [0:0] CLBLM_L_X12Y150_SLICE_X16Y150_D2;
  wire [0:0] CLBLM_L_X12Y150_SLICE_X16Y150_D3;
  wire [0:0] CLBLM_L_X12Y150_SLICE_X16Y150_D4;
  wire [0:0] CLBLM_L_X12Y150_SLICE_X16Y150_D5;
  wire [0:0] CLBLM_L_X12Y150_SLICE_X16Y150_D6;
  wire [0:0] CLBLM_L_X12Y150_SLICE_X16Y150_DO5;
  wire [0:0] CLBLM_L_X12Y150_SLICE_X16Y150_DO6;
  wire [0:0] CLBLM_L_X12Y150_SLICE_X16Y150_D_CY;
  wire [0:0] CLBLM_L_X12Y150_SLICE_X16Y150_D_XOR;
  wire [0:0] CLBLM_L_X12Y150_SLICE_X17Y150_A;
  wire [0:0] CLBLM_L_X12Y150_SLICE_X17Y150_A1;
  wire [0:0] CLBLM_L_X12Y150_SLICE_X17Y150_A2;
  wire [0:0] CLBLM_L_X12Y150_SLICE_X17Y150_A3;
  wire [0:0] CLBLM_L_X12Y150_SLICE_X17Y150_A4;
  wire [0:0] CLBLM_L_X12Y150_SLICE_X17Y150_A5;
  wire [0:0] CLBLM_L_X12Y150_SLICE_X17Y150_A6;
  wire [0:0] CLBLM_L_X12Y150_SLICE_X17Y150_AO5;
  wire [0:0] CLBLM_L_X12Y150_SLICE_X17Y150_AO6;
  wire [0:0] CLBLM_L_X12Y150_SLICE_X17Y150_A_CY;
  wire [0:0] CLBLM_L_X12Y150_SLICE_X17Y150_A_XOR;
  wire [0:0] CLBLM_L_X12Y150_SLICE_X17Y150_B;
  wire [0:0] CLBLM_L_X12Y150_SLICE_X17Y150_B1;
  wire [0:0] CLBLM_L_X12Y150_SLICE_X17Y150_B2;
  wire [0:0] CLBLM_L_X12Y150_SLICE_X17Y150_B3;
  wire [0:0] CLBLM_L_X12Y150_SLICE_X17Y150_B4;
  wire [0:0] CLBLM_L_X12Y150_SLICE_X17Y150_B5;
  wire [0:0] CLBLM_L_X12Y150_SLICE_X17Y150_B6;
  wire [0:0] CLBLM_L_X12Y150_SLICE_X17Y150_BO5;
  wire [0:0] CLBLM_L_X12Y150_SLICE_X17Y150_BO6;
  wire [0:0] CLBLM_L_X12Y150_SLICE_X17Y150_B_CY;
  wire [0:0] CLBLM_L_X12Y150_SLICE_X17Y150_B_XOR;
  wire [0:0] CLBLM_L_X12Y150_SLICE_X17Y150_C;
  wire [0:0] CLBLM_L_X12Y150_SLICE_X17Y150_C1;
  wire [0:0] CLBLM_L_X12Y150_SLICE_X17Y150_C2;
  wire [0:0] CLBLM_L_X12Y150_SLICE_X17Y150_C3;
  wire [0:0] CLBLM_L_X12Y150_SLICE_X17Y150_C4;
  wire [0:0] CLBLM_L_X12Y150_SLICE_X17Y150_C5;
  wire [0:0] CLBLM_L_X12Y150_SLICE_X17Y150_C6;
  wire [0:0] CLBLM_L_X12Y150_SLICE_X17Y150_CO5;
  wire [0:0] CLBLM_L_X12Y150_SLICE_X17Y150_CO6;
  wire [0:0] CLBLM_L_X12Y150_SLICE_X17Y150_C_CY;
  wire [0:0] CLBLM_L_X12Y150_SLICE_X17Y150_C_XOR;
  wire [0:0] CLBLM_L_X12Y150_SLICE_X17Y150_D;
  wire [0:0] CLBLM_L_X12Y150_SLICE_X17Y150_D1;
  wire [0:0] CLBLM_L_X12Y150_SLICE_X17Y150_D2;
  wire [0:0] CLBLM_L_X12Y150_SLICE_X17Y150_D3;
  wire [0:0] CLBLM_L_X12Y150_SLICE_X17Y150_D4;
  wire [0:0] CLBLM_L_X12Y150_SLICE_X17Y150_D5;
  wire [0:0] CLBLM_L_X12Y150_SLICE_X17Y150_D6;
  wire [0:0] CLBLM_L_X12Y150_SLICE_X17Y150_DO5;
  wire [0:0] CLBLM_L_X12Y150_SLICE_X17Y150_DO6;
  wire [0:0] CLBLM_L_X12Y150_SLICE_X17Y150_D_CY;
  wire [0:0] CLBLM_L_X12Y150_SLICE_X17Y150_D_XOR;
  wire [0:0] CLBLM_L_X12Y151_SLICE_X16Y151_A;
  wire [0:0] CLBLM_L_X12Y151_SLICE_X16Y151_A1;
  wire [0:0] CLBLM_L_X12Y151_SLICE_X16Y151_A2;
  wire [0:0] CLBLM_L_X12Y151_SLICE_X16Y151_A3;
  wire [0:0] CLBLM_L_X12Y151_SLICE_X16Y151_A4;
  wire [0:0] CLBLM_L_X12Y151_SLICE_X16Y151_A5;
  wire [0:0] CLBLM_L_X12Y151_SLICE_X16Y151_A6;
  wire [0:0] CLBLM_L_X12Y151_SLICE_X16Y151_AMUX;
  wire [0:0] CLBLM_L_X12Y151_SLICE_X16Y151_AO5;
  wire [0:0] CLBLM_L_X12Y151_SLICE_X16Y151_AO6;
  wire [0:0] CLBLM_L_X12Y151_SLICE_X16Y151_AQ;
  wire [0:0] CLBLM_L_X12Y151_SLICE_X16Y151_A_CY;
  wire [0:0] CLBLM_L_X12Y151_SLICE_X16Y151_A_XOR;
  wire [0:0] CLBLM_L_X12Y151_SLICE_X16Y151_B;
  wire [0:0] CLBLM_L_X12Y151_SLICE_X16Y151_B1;
  wire [0:0] CLBLM_L_X12Y151_SLICE_X16Y151_B2;
  wire [0:0] CLBLM_L_X12Y151_SLICE_X16Y151_B3;
  wire [0:0] CLBLM_L_X12Y151_SLICE_X16Y151_B4;
  wire [0:0] CLBLM_L_X12Y151_SLICE_X16Y151_B5;
  wire [0:0] CLBLM_L_X12Y151_SLICE_X16Y151_B6;
  wire [0:0] CLBLM_L_X12Y151_SLICE_X16Y151_BMUX;
  wire [0:0] CLBLM_L_X12Y151_SLICE_X16Y151_BO5;
  wire [0:0] CLBLM_L_X12Y151_SLICE_X16Y151_BO6;
  wire [0:0] CLBLM_L_X12Y151_SLICE_X16Y151_B_CY;
  wire [0:0] CLBLM_L_X12Y151_SLICE_X16Y151_B_XOR;
  wire [0:0] CLBLM_L_X12Y151_SLICE_X16Y151_C;
  wire [0:0] CLBLM_L_X12Y151_SLICE_X16Y151_C1;
  wire [0:0] CLBLM_L_X12Y151_SLICE_X16Y151_C2;
  wire [0:0] CLBLM_L_X12Y151_SLICE_X16Y151_C3;
  wire [0:0] CLBLM_L_X12Y151_SLICE_X16Y151_C4;
  wire [0:0] CLBLM_L_X12Y151_SLICE_X16Y151_C5;
  wire [0:0] CLBLM_L_X12Y151_SLICE_X16Y151_C6;
  wire [0:0] CLBLM_L_X12Y151_SLICE_X16Y151_CLK;
  wire [0:0] CLBLM_L_X12Y151_SLICE_X16Y151_CO5;
  wire [0:0] CLBLM_L_X12Y151_SLICE_X16Y151_CO6;
  wire [0:0] CLBLM_L_X12Y151_SLICE_X16Y151_C_CY;
  wire [0:0] CLBLM_L_X12Y151_SLICE_X16Y151_C_XOR;
  wire [0:0] CLBLM_L_X12Y151_SLICE_X16Y151_D;
  wire [0:0] CLBLM_L_X12Y151_SLICE_X16Y151_D1;
  wire [0:0] CLBLM_L_X12Y151_SLICE_X16Y151_D2;
  wire [0:0] CLBLM_L_X12Y151_SLICE_X16Y151_D3;
  wire [0:0] CLBLM_L_X12Y151_SLICE_X16Y151_D4;
  wire [0:0] CLBLM_L_X12Y151_SLICE_X16Y151_D5;
  wire [0:0] CLBLM_L_X12Y151_SLICE_X16Y151_D6;
  wire [0:0] CLBLM_L_X12Y151_SLICE_X16Y151_DO5;
  wire [0:0] CLBLM_L_X12Y151_SLICE_X16Y151_DO6;
  wire [0:0] CLBLM_L_X12Y151_SLICE_X16Y151_D_CY;
  wire [0:0] CLBLM_L_X12Y151_SLICE_X16Y151_D_XOR;
  wire [0:0] CLBLM_L_X12Y151_SLICE_X17Y151_A;
  wire [0:0] CLBLM_L_X12Y151_SLICE_X17Y151_A1;
  wire [0:0] CLBLM_L_X12Y151_SLICE_X17Y151_A2;
  wire [0:0] CLBLM_L_X12Y151_SLICE_X17Y151_A3;
  wire [0:0] CLBLM_L_X12Y151_SLICE_X17Y151_A4;
  wire [0:0] CLBLM_L_X12Y151_SLICE_X17Y151_A5;
  wire [0:0] CLBLM_L_X12Y151_SLICE_X17Y151_A6;
  wire [0:0] CLBLM_L_X12Y151_SLICE_X17Y151_AO5;
  wire [0:0] CLBLM_L_X12Y151_SLICE_X17Y151_AO6;
  wire [0:0] CLBLM_L_X12Y151_SLICE_X17Y151_A_CY;
  wire [0:0] CLBLM_L_X12Y151_SLICE_X17Y151_A_XOR;
  wire [0:0] CLBLM_L_X12Y151_SLICE_X17Y151_B;
  wire [0:0] CLBLM_L_X12Y151_SLICE_X17Y151_B1;
  wire [0:0] CLBLM_L_X12Y151_SLICE_X17Y151_B2;
  wire [0:0] CLBLM_L_X12Y151_SLICE_X17Y151_B3;
  wire [0:0] CLBLM_L_X12Y151_SLICE_X17Y151_B4;
  wire [0:0] CLBLM_L_X12Y151_SLICE_X17Y151_B5;
  wire [0:0] CLBLM_L_X12Y151_SLICE_X17Y151_B6;
  wire [0:0] CLBLM_L_X12Y151_SLICE_X17Y151_BO5;
  wire [0:0] CLBLM_L_X12Y151_SLICE_X17Y151_BO6;
  wire [0:0] CLBLM_L_X12Y151_SLICE_X17Y151_B_CY;
  wire [0:0] CLBLM_L_X12Y151_SLICE_X17Y151_B_XOR;
  wire [0:0] CLBLM_L_X12Y151_SLICE_X17Y151_C;
  wire [0:0] CLBLM_L_X12Y151_SLICE_X17Y151_C1;
  wire [0:0] CLBLM_L_X12Y151_SLICE_X17Y151_C2;
  wire [0:0] CLBLM_L_X12Y151_SLICE_X17Y151_C3;
  wire [0:0] CLBLM_L_X12Y151_SLICE_X17Y151_C4;
  wire [0:0] CLBLM_L_X12Y151_SLICE_X17Y151_C5;
  wire [0:0] CLBLM_L_X12Y151_SLICE_X17Y151_C6;
  wire [0:0] CLBLM_L_X12Y151_SLICE_X17Y151_CO5;
  wire [0:0] CLBLM_L_X12Y151_SLICE_X17Y151_CO6;
  wire [0:0] CLBLM_L_X12Y151_SLICE_X17Y151_C_CY;
  wire [0:0] CLBLM_L_X12Y151_SLICE_X17Y151_C_XOR;
  wire [0:0] CLBLM_L_X12Y151_SLICE_X17Y151_D;
  wire [0:0] CLBLM_L_X12Y151_SLICE_X17Y151_D1;
  wire [0:0] CLBLM_L_X12Y151_SLICE_X17Y151_D2;
  wire [0:0] CLBLM_L_X12Y151_SLICE_X17Y151_D3;
  wire [0:0] CLBLM_L_X12Y151_SLICE_X17Y151_D4;
  wire [0:0] CLBLM_L_X12Y151_SLICE_X17Y151_D5;
  wire [0:0] CLBLM_L_X12Y151_SLICE_X17Y151_D6;
  wire [0:0] CLBLM_L_X12Y151_SLICE_X17Y151_DO5;
  wire [0:0] CLBLM_L_X12Y151_SLICE_X17Y151_DO6;
  wire [0:0] CLBLM_L_X12Y151_SLICE_X17Y151_D_CY;
  wire [0:0] CLBLM_L_X12Y151_SLICE_X17Y151_D_XOR;
  wire [0:0] CLBLM_L_X12Y152_SLICE_X16Y152_A;
  wire [0:0] CLBLM_L_X12Y152_SLICE_X16Y152_A1;
  wire [0:0] CLBLM_L_X12Y152_SLICE_X16Y152_A2;
  wire [0:0] CLBLM_L_X12Y152_SLICE_X16Y152_A3;
  wire [0:0] CLBLM_L_X12Y152_SLICE_X16Y152_A4;
  wire [0:0] CLBLM_L_X12Y152_SLICE_X16Y152_A5;
  wire [0:0] CLBLM_L_X12Y152_SLICE_X16Y152_A6;
  wire [0:0] CLBLM_L_X12Y152_SLICE_X16Y152_AMUX;
  wire [0:0] CLBLM_L_X12Y152_SLICE_X16Y152_AO5;
  wire [0:0] CLBLM_L_X12Y152_SLICE_X16Y152_AO6;
  wire [0:0] CLBLM_L_X12Y152_SLICE_X16Y152_A_CY;
  wire [0:0] CLBLM_L_X12Y152_SLICE_X16Y152_A_XOR;
  wire [0:0] CLBLM_L_X12Y152_SLICE_X16Y152_B;
  wire [0:0] CLBLM_L_X12Y152_SLICE_X16Y152_B1;
  wire [0:0] CLBLM_L_X12Y152_SLICE_X16Y152_B2;
  wire [0:0] CLBLM_L_X12Y152_SLICE_X16Y152_B3;
  wire [0:0] CLBLM_L_X12Y152_SLICE_X16Y152_B4;
  wire [0:0] CLBLM_L_X12Y152_SLICE_X16Y152_B5;
  wire [0:0] CLBLM_L_X12Y152_SLICE_X16Y152_B6;
  wire [0:0] CLBLM_L_X12Y152_SLICE_X16Y152_BO5;
  wire [0:0] CLBLM_L_X12Y152_SLICE_X16Y152_BO6;
  wire [0:0] CLBLM_L_X12Y152_SLICE_X16Y152_B_CY;
  wire [0:0] CLBLM_L_X12Y152_SLICE_X16Y152_B_XOR;
  wire [0:0] CLBLM_L_X12Y152_SLICE_X16Y152_C;
  wire [0:0] CLBLM_L_X12Y152_SLICE_X16Y152_C1;
  wire [0:0] CLBLM_L_X12Y152_SLICE_X16Y152_C2;
  wire [0:0] CLBLM_L_X12Y152_SLICE_X16Y152_C3;
  wire [0:0] CLBLM_L_X12Y152_SLICE_X16Y152_C4;
  wire [0:0] CLBLM_L_X12Y152_SLICE_X16Y152_C5;
  wire [0:0] CLBLM_L_X12Y152_SLICE_X16Y152_C6;
  wire [0:0] CLBLM_L_X12Y152_SLICE_X16Y152_CO5;
  wire [0:0] CLBLM_L_X12Y152_SLICE_X16Y152_CO6;
  wire [0:0] CLBLM_L_X12Y152_SLICE_X16Y152_C_CY;
  wire [0:0] CLBLM_L_X12Y152_SLICE_X16Y152_C_XOR;
  wire [0:0] CLBLM_L_X12Y152_SLICE_X16Y152_D;
  wire [0:0] CLBLM_L_X12Y152_SLICE_X16Y152_D1;
  wire [0:0] CLBLM_L_X12Y152_SLICE_X16Y152_D2;
  wire [0:0] CLBLM_L_X12Y152_SLICE_X16Y152_D3;
  wire [0:0] CLBLM_L_X12Y152_SLICE_X16Y152_D4;
  wire [0:0] CLBLM_L_X12Y152_SLICE_X16Y152_D5;
  wire [0:0] CLBLM_L_X12Y152_SLICE_X16Y152_D6;
  wire [0:0] CLBLM_L_X12Y152_SLICE_X16Y152_DO5;
  wire [0:0] CLBLM_L_X12Y152_SLICE_X16Y152_DO6;
  wire [0:0] CLBLM_L_X12Y152_SLICE_X16Y152_D_CY;
  wire [0:0] CLBLM_L_X12Y152_SLICE_X16Y152_D_XOR;
  wire [0:0] CLBLM_L_X12Y152_SLICE_X17Y152_A;
  wire [0:0] CLBLM_L_X12Y152_SLICE_X17Y152_A1;
  wire [0:0] CLBLM_L_X12Y152_SLICE_X17Y152_A2;
  wire [0:0] CLBLM_L_X12Y152_SLICE_X17Y152_A3;
  wire [0:0] CLBLM_L_X12Y152_SLICE_X17Y152_A4;
  wire [0:0] CLBLM_L_X12Y152_SLICE_X17Y152_A5;
  wire [0:0] CLBLM_L_X12Y152_SLICE_X17Y152_A6;
  wire [0:0] CLBLM_L_X12Y152_SLICE_X17Y152_AO5;
  wire [0:0] CLBLM_L_X12Y152_SLICE_X17Y152_AO6;
  wire [0:0] CLBLM_L_X12Y152_SLICE_X17Y152_A_CY;
  wire [0:0] CLBLM_L_X12Y152_SLICE_X17Y152_A_XOR;
  wire [0:0] CLBLM_L_X12Y152_SLICE_X17Y152_B;
  wire [0:0] CLBLM_L_X12Y152_SLICE_X17Y152_B1;
  wire [0:0] CLBLM_L_X12Y152_SLICE_X17Y152_B2;
  wire [0:0] CLBLM_L_X12Y152_SLICE_X17Y152_B3;
  wire [0:0] CLBLM_L_X12Y152_SLICE_X17Y152_B4;
  wire [0:0] CLBLM_L_X12Y152_SLICE_X17Y152_B5;
  wire [0:0] CLBLM_L_X12Y152_SLICE_X17Y152_B6;
  wire [0:0] CLBLM_L_X12Y152_SLICE_X17Y152_BO5;
  wire [0:0] CLBLM_L_X12Y152_SLICE_X17Y152_BO6;
  wire [0:0] CLBLM_L_X12Y152_SLICE_X17Y152_B_CY;
  wire [0:0] CLBLM_L_X12Y152_SLICE_X17Y152_B_XOR;
  wire [0:0] CLBLM_L_X12Y152_SLICE_X17Y152_C;
  wire [0:0] CLBLM_L_X12Y152_SLICE_X17Y152_C1;
  wire [0:0] CLBLM_L_X12Y152_SLICE_X17Y152_C2;
  wire [0:0] CLBLM_L_X12Y152_SLICE_X17Y152_C3;
  wire [0:0] CLBLM_L_X12Y152_SLICE_X17Y152_C4;
  wire [0:0] CLBLM_L_X12Y152_SLICE_X17Y152_C5;
  wire [0:0] CLBLM_L_X12Y152_SLICE_X17Y152_C6;
  wire [0:0] CLBLM_L_X12Y152_SLICE_X17Y152_CO5;
  wire [0:0] CLBLM_L_X12Y152_SLICE_X17Y152_CO6;
  wire [0:0] CLBLM_L_X12Y152_SLICE_X17Y152_C_CY;
  wire [0:0] CLBLM_L_X12Y152_SLICE_X17Y152_C_XOR;
  wire [0:0] CLBLM_L_X12Y152_SLICE_X17Y152_D;
  wire [0:0] CLBLM_L_X12Y152_SLICE_X17Y152_D1;
  wire [0:0] CLBLM_L_X12Y152_SLICE_X17Y152_D2;
  wire [0:0] CLBLM_L_X12Y152_SLICE_X17Y152_D3;
  wire [0:0] CLBLM_L_X12Y152_SLICE_X17Y152_D4;
  wire [0:0] CLBLM_L_X12Y152_SLICE_X17Y152_D5;
  wire [0:0] CLBLM_L_X12Y152_SLICE_X17Y152_D6;
  wire [0:0] CLBLM_L_X12Y152_SLICE_X17Y152_DO5;
  wire [0:0] CLBLM_L_X12Y152_SLICE_X17Y152_DO6;
  wire [0:0] CLBLM_L_X12Y152_SLICE_X17Y152_D_CY;
  wire [0:0] CLBLM_L_X12Y152_SLICE_X17Y152_D_XOR;
  wire [0:0] CLBLM_L_X12Y153_SLICE_X16Y153_A;
  wire [0:0] CLBLM_L_X12Y153_SLICE_X16Y153_A1;
  wire [0:0] CLBLM_L_X12Y153_SLICE_X16Y153_A2;
  wire [0:0] CLBLM_L_X12Y153_SLICE_X16Y153_A3;
  wire [0:0] CLBLM_L_X12Y153_SLICE_X16Y153_A4;
  wire [0:0] CLBLM_L_X12Y153_SLICE_X16Y153_A5;
  wire [0:0] CLBLM_L_X12Y153_SLICE_X16Y153_A6;
  wire [0:0] CLBLM_L_X12Y153_SLICE_X16Y153_AMUX;
  wire [0:0] CLBLM_L_X12Y153_SLICE_X16Y153_AO5;
  wire [0:0] CLBLM_L_X12Y153_SLICE_X16Y153_AO6;
  wire [0:0] CLBLM_L_X12Y153_SLICE_X16Y153_A_CY;
  wire [0:0] CLBLM_L_X12Y153_SLICE_X16Y153_A_XOR;
  wire [0:0] CLBLM_L_X12Y153_SLICE_X16Y153_B;
  wire [0:0] CLBLM_L_X12Y153_SLICE_X16Y153_B1;
  wire [0:0] CLBLM_L_X12Y153_SLICE_X16Y153_B2;
  wire [0:0] CLBLM_L_X12Y153_SLICE_X16Y153_B3;
  wire [0:0] CLBLM_L_X12Y153_SLICE_X16Y153_B4;
  wire [0:0] CLBLM_L_X12Y153_SLICE_X16Y153_B5;
  wire [0:0] CLBLM_L_X12Y153_SLICE_X16Y153_B6;
  wire [0:0] CLBLM_L_X12Y153_SLICE_X16Y153_BO5;
  wire [0:0] CLBLM_L_X12Y153_SLICE_X16Y153_BO6;
  wire [0:0] CLBLM_L_X12Y153_SLICE_X16Y153_B_CY;
  wire [0:0] CLBLM_L_X12Y153_SLICE_X16Y153_B_XOR;
  wire [0:0] CLBLM_L_X12Y153_SLICE_X16Y153_C;
  wire [0:0] CLBLM_L_X12Y153_SLICE_X16Y153_C1;
  wire [0:0] CLBLM_L_X12Y153_SLICE_X16Y153_C2;
  wire [0:0] CLBLM_L_X12Y153_SLICE_X16Y153_C3;
  wire [0:0] CLBLM_L_X12Y153_SLICE_X16Y153_C4;
  wire [0:0] CLBLM_L_X12Y153_SLICE_X16Y153_C5;
  wire [0:0] CLBLM_L_X12Y153_SLICE_X16Y153_C6;
  wire [0:0] CLBLM_L_X12Y153_SLICE_X16Y153_CO5;
  wire [0:0] CLBLM_L_X12Y153_SLICE_X16Y153_CO6;
  wire [0:0] CLBLM_L_X12Y153_SLICE_X16Y153_C_CY;
  wire [0:0] CLBLM_L_X12Y153_SLICE_X16Y153_C_XOR;
  wire [0:0] CLBLM_L_X12Y153_SLICE_X16Y153_D;
  wire [0:0] CLBLM_L_X12Y153_SLICE_X16Y153_D1;
  wire [0:0] CLBLM_L_X12Y153_SLICE_X16Y153_D2;
  wire [0:0] CLBLM_L_X12Y153_SLICE_X16Y153_D3;
  wire [0:0] CLBLM_L_X12Y153_SLICE_X16Y153_D4;
  wire [0:0] CLBLM_L_X12Y153_SLICE_X16Y153_D5;
  wire [0:0] CLBLM_L_X12Y153_SLICE_X16Y153_D6;
  wire [0:0] CLBLM_L_X12Y153_SLICE_X16Y153_DO5;
  wire [0:0] CLBLM_L_X12Y153_SLICE_X16Y153_DO6;
  wire [0:0] CLBLM_L_X12Y153_SLICE_X16Y153_D_CY;
  wire [0:0] CLBLM_L_X12Y153_SLICE_X16Y153_D_XOR;
  wire [0:0] CLBLM_L_X12Y153_SLICE_X17Y153_A;
  wire [0:0] CLBLM_L_X12Y153_SLICE_X17Y153_A1;
  wire [0:0] CLBLM_L_X12Y153_SLICE_X17Y153_A2;
  wire [0:0] CLBLM_L_X12Y153_SLICE_X17Y153_A3;
  wire [0:0] CLBLM_L_X12Y153_SLICE_X17Y153_A4;
  wire [0:0] CLBLM_L_X12Y153_SLICE_X17Y153_A5;
  wire [0:0] CLBLM_L_X12Y153_SLICE_X17Y153_A6;
  wire [0:0] CLBLM_L_X12Y153_SLICE_X17Y153_AO5;
  wire [0:0] CLBLM_L_X12Y153_SLICE_X17Y153_AO6;
  wire [0:0] CLBLM_L_X12Y153_SLICE_X17Y153_A_CY;
  wire [0:0] CLBLM_L_X12Y153_SLICE_X17Y153_A_XOR;
  wire [0:0] CLBLM_L_X12Y153_SLICE_X17Y153_B;
  wire [0:0] CLBLM_L_X12Y153_SLICE_X17Y153_B1;
  wire [0:0] CLBLM_L_X12Y153_SLICE_X17Y153_B2;
  wire [0:0] CLBLM_L_X12Y153_SLICE_X17Y153_B3;
  wire [0:0] CLBLM_L_X12Y153_SLICE_X17Y153_B4;
  wire [0:0] CLBLM_L_X12Y153_SLICE_X17Y153_B5;
  wire [0:0] CLBLM_L_X12Y153_SLICE_X17Y153_B6;
  wire [0:0] CLBLM_L_X12Y153_SLICE_X17Y153_BO5;
  wire [0:0] CLBLM_L_X12Y153_SLICE_X17Y153_BO6;
  wire [0:0] CLBLM_L_X12Y153_SLICE_X17Y153_B_CY;
  wire [0:0] CLBLM_L_X12Y153_SLICE_X17Y153_B_XOR;
  wire [0:0] CLBLM_L_X12Y153_SLICE_X17Y153_C;
  wire [0:0] CLBLM_L_X12Y153_SLICE_X17Y153_C1;
  wire [0:0] CLBLM_L_X12Y153_SLICE_X17Y153_C2;
  wire [0:0] CLBLM_L_X12Y153_SLICE_X17Y153_C3;
  wire [0:0] CLBLM_L_X12Y153_SLICE_X17Y153_C4;
  wire [0:0] CLBLM_L_X12Y153_SLICE_X17Y153_C5;
  wire [0:0] CLBLM_L_X12Y153_SLICE_X17Y153_C6;
  wire [0:0] CLBLM_L_X12Y153_SLICE_X17Y153_CO5;
  wire [0:0] CLBLM_L_X12Y153_SLICE_X17Y153_CO6;
  wire [0:0] CLBLM_L_X12Y153_SLICE_X17Y153_C_CY;
  wire [0:0] CLBLM_L_X12Y153_SLICE_X17Y153_C_XOR;
  wire [0:0] CLBLM_L_X12Y153_SLICE_X17Y153_D;
  wire [0:0] CLBLM_L_X12Y153_SLICE_X17Y153_D1;
  wire [0:0] CLBLM_L_X12Y153_SLICE_X17Y153_D2;
  wire [0:0] CLBLM_L_X12Y153_SLICE_X17Y153_D3;
  wire [0:0] CLBLM_L_X12Y153_SLICE_X17Y153_D4;
  wire [0:0] CLBLM_L_X12Y153_SLICE_X17Y153_D5;
  wire [0:0] CLBLM_L_X12Y153_SLICE_X17Y153_D6;
  wire [0:0] CLBLM_L_X12Y153_SLICE_X17Y153_DO5;
  wire [0:0] CLBLM_L_X12Y153_SLICE_X17Y153_DO6;
  wire [0:0] CLBLM_L_X12Y153_SLICE_X17Y153_D_CY;
  wire [0:0] CLBLM_L_X12Y153_SLICE_X17Y153_D_XOR;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X10Y142_A;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X10Y142_A1;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X10Y142_A2;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X10Y142_A3;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X10Y142_A4;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X10Y142_A5;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X10Y142_A5Q;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X10Y142_A6;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X10Y142_AMUX;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X10Y142_AO5;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X10Y142_AO6;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X10Y142_AQ;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X10Y142_AX;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X10Y142_A_CY;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X10Y142_A_XOR;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X10Y142_B;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X10Y142_B1;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X10Y142_B2;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X10Y142_B3;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X10Y142_B4;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X10Y142_B5;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X10Y142_B6;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X10Y142_BO5;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X10Y142_BO6;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X10Y142_BQ;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X10Y142_B_CY;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X10Y142_B_XOR;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X10Y142_C;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X10Y142_C1;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X10Y142_C2;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X10Y142_C3;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X10Y142_C4;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X10Y142_C5;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X10Y142_C6;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X10Y142_CLK;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X10Y142_CO5;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X10Y142_CO6;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X10Y142_CQ;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X10Y142_C_CY;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X10Y142_C_XOR;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X10Y142_D;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X10Y142_D1;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X10Y142_D2;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X10Y142_D3;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X10Y142_D4;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X10Y142_D5;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X10Y142_D6;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X10Y142_DO5;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X10Y142_DO6;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X10Y142_D_CY;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X10Y142_D_XOR;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X11Y142_A;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X11Y142_A1;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X11Y142_A2;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X11Y142_A3;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X11Y142_A4;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X11Y142_A5;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X11Y142_A6;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X11Y142_AO5;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X11Y142_AO6;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X11Y142_AQ;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X11Y142_A_CY;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X11Y142_A_XOR;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X11Y142_B;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X11Y142_B1;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X11Y142_B2;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X11Y142_B3;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X11Y142_B4;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X11Y142_B5;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X11Y142_B6;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X11Y142_BO5;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X11Y142_BO6;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X11Y142_BQ;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X11Y142_B_CY;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X11Y142_B_XOR;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X11Y142_C;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X11Y142_C1;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X11Y142_C2;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X11Y142_C3;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X11Y142_C4;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X11Y142_C5;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X11Y142_C6;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X11Y142_CLK;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X11Y142_CMUX;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X11Y142_CO5;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X11Y142_CO6;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X11Y142_C_CY;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X11Y142_C_XOR;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X11Y142_D;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X11Y142_D1;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X11Y142_D2;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X11Y142_D3;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X11Y142_D4;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X11Y142_D5;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X11Y142_D6;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X11Y142_DMUX;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X11Y142_DO5;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X11Y142_DO6;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X11Y142_D_CY;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X11Y142_D_XOR;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X10Y143_A;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X10Y143_A1;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X10Y143_A2;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X10Y143_A3;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X10Y143_A4;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X10Y143_A5;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X10Y143_A6;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X10Y143_AO5;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X10Y143_AO6;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X10Y143_AQ;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X10Y143_A_CY;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X10Y143_A_XOR;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X10Y143_B;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X10Y143_B1;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X10Y143_B2;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X10Y143_B3;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X10Y143_B4;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X10Y143_B5;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X10Y143_B6;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X10Y143_BO5;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X10Y143_BO6;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X10Y143_BQ;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X10Y143_B_CY;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X10Y143_B_XOR;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X10Y143_C;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X10Y143_C1;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X10Y143_C2;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X10Y143_C3;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X10Y143_C4;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X10Y143_C5;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X10Y143_C6;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X10Y143_CLK;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X10Y143_CO5;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X10Y143_CO6;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X10Y143_CQ;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X10Y143_C_CY;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X10Y143_C_XOR;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X10Y143_D;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X10Y143_D1;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X10Y143_D2;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X10Y143_D3;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X10Y143_D4;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X10Y143_D5;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X10Y143_D6;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X10Y143_DO5;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X10Y143_DO6;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X10Y143_DQ;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X10Y143_D_CY;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X10Y143_D_XOR;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X11Y143_A;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X11Y143_A1;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X11Y143_A2;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X11Y143_A3;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X11Y143_A4;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X11Y143_A5;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X11Y143_A6;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X11Y143_AO5;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X11Y143_AO6;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X11Y143_AQ;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X11Y143_A_CY;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X11Y143_A_XOR;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X11Y143_B;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X11Y143_B1;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X11Y143_B2;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X11Y143_B3;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X11Y143_B4;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X11Y143_B5;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X11Y143_B6;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X11Y143_BO5;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X11Y143_BO6;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X11Y143_BQ;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X11Y143_B_CY;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X11Y143_B_XOR;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X11Y143_C;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X11Y143_C1;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X11Y143_C2;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X11Y143_C3;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X11Y143_C4;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X11Y143_C5;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X11Y143_C6;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X11Y143_CLK;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X11Y143_CO5;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X11Y143_CO6;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X11Y143_CQ;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X11Y143_C_CY;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X11Y143_C_XOR;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X11Y143_D;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X11Y143_D1;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X11Y143_D2;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X11Y143_D3;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X11Y143_D4;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X11Y143_D5;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X11Y143_D5Q;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X11Y143_D6;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X11Y143_DMUX;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X11Y143_DO5;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X11Y143_DO6;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X11Y143_DQ;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X11Y143_D_CY;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X11Y143_D_XOR;
  wire [0:0] CLBLM_L_X8Y144_SLICE_X10Y144_A;
  wire [0:0] CLBLM_L_X8Y144_SLICE_X10Y144_A1;
  wire [0:0] CLBLM_L_X8Y144_SLICE_X10Y144_A2;
  wire [0:0] CLBLM_L_X8Y144_SLICE_X10Y144_A3;
  wire [0:0] CLBLM_L_X8Y144_SLICE_X10Y144_A4;
  wire [0:0] CLBLM_L_X8Y144_SLICE_X10Y144_A5;
  wire [0:0] CLBLM_L_X8Y144_SLICE_X10Y144_A6;
  wire [0:0] CLBLM_L_X8Y144_SLICE_X10Y144_AMUX;
  wire [0:0] CLBLM_L_X8Y144_SLICE_X10Y144_AO5;
  wire [0:0] CLBLM_L_X8Y144_SLICE_X10Y144_AO6;
  wire [0:0] CLBLM_L_X8Y144_SLICE_X10Y144_AQ;
  wire [0:0] CLBLM_L_X8Y144_SLICE_X10Y144_AX;
  wire [0:0] CLBLM_L_X8Y144_SLICE_X10Y144_A_CY;
  wire [0:0] CLBLM_L_X8Y144_SLICE_X10Y144_A_XOR;
  wire [0:0] CLBLM_L_X8Y144_SLICE_X10Y144_B;
  wire [0:0] CLBLM_L_X8Y144_SLICE_X10Y144_B1;
  wire [0:0] CLBLM_L_X8Y144_SLICE_X10Y144_B2;
  wire [0:0] CLBLM_L_X8Y144_SLICE_X10Y144_B3;
  wire [0:0] CLBLM_L_X8Y144_SLICE_X10Y144_B4;
  wire [0:0] CLBLM_L_X8Y144_SLICE_X10Y144_B5;
  wire [0:0] CLBLM_L_X8Y144_SLICE_X10Y144_B6;
  wire [0:0] CLBLM_L_X8Y144_SLICE_X10Y144_BMUX;
  wire [0:0] CLBLM_L_X8Y144_SLICE_X10Y144_BO5;
  wire [0:0] CLBLM_L_X8Y144_SLICE_X10Y144_BO6;
  wire [0:0] CLBLM_L_X8Y144_SLICE_X10Y144_BQ;
  wire [0:0] CLBLM_L_X8Y144_SLICE_X10Y144_BX;
  wire [0:0] CLBLM_L_X8Y144_SLICE_X10Y144_B_CY;
  wire [0:0] CLBLM_L_X8Y144_SLICE_X10Y144_B_XOR;
  wire [0:0] CLBLM_L_X8Y144_SLICE_X10Y144_C;
  wire [0:0] CLBLM_L_X8Y144_SLICE_X10Y144_C1;
  wire [0:0] CLBLM_L_X8Y144_SLICE_X10Y144_C2;
  wire [0:0] CLBLM_L_X8Y144_SLICE_X10Y144_C3;
  wire [0:0] CLBLM_L_X8Y144_SLICE_X10Y144_C4;
  wire [0:0] CLBLM_L_X8Y144_SLICE_X10Y144_C5;
  wire [0:0] CLBLM_L_X8Y144_SLICE_X10Y144_C6;
  wire [0:0] CLBLM_L_X8Y144_SLICE_X10Y144_CE;
  wire [0:0] CLBLM_L_X8Y144_SLICE_X10Y144_CLK;
  wire [0:0] CLBLM_L_X8Y144_SLICE_X10Y144_CO5;
  wire [0:0] CLBLM_L_X8Y144_SLICE_X10Y144_CO6;
  wire [0:0] CLBLM_L_X8Y144_SLICE_X10Y144_C_CY;
  wire [0:0] CLBLM_L_X8Y144_SLICE_X10Y144_C_XOR;
  wire [0:0] CLBLM_L_X8Y144_SLICE_X10Y144_D;
  wire [0:0] CLBLM_L_X8Y144_SLICE_X10Y144_D1;
  wire [0:0] CLBLM_L_X8Y144_SLICE_X10Y144_D2;
  wire [0:0] CLBLM_L_X8Y144_SLICE_X10Y144_D3;
  wire [0:0] CLBLM_L_X8Y144_SLICE_X10Y144_D4;
  wire [0:0] CLBLM_L_X8Y144_SLICE_X10Y144_D5;
  wire [0:0] CLBLM_L_X8Y144_SLICE_X10Y144_D6;
  wire [0:0] CLBLM_L_X8Y144_SLICE_X10Y144_DO5;
  wire [0:0] CLBLM_L_X8Y144_SLICE_X10Y144_DO6;
  wire [0:0] CLBLM_L_X8Y144_SLICE_X10Y144_D_CY;
  wire [0:0] CLBLM_L_X8Y144_SLICE_X10Y144_D_XOR;
  wire [0:0] CLBLM_L_X8Y144_SLICE_X11Y144_A;
  wire [0:0] CLBLM_L_X8Y144_SLICE_X11Y144_A1;
  wire [0:0] CLBLM_L_X8Y144_SLICE_X11Y144_A2;
  wire [0:0] CLBLM_L_X8Y144_SLICE_X11Y144_A3;
  wire [0:0] CLBLM_L_X8Y144_SLICE_X11Y144_A4;
  wire [0:0] CLBLM_L_X8Y144_SLICE_X11Y144_A5;
  wire [0:0] CLBLM_L_X8Y144_SLICE_X11Y144_A6;
  wire [0:0] CLBLM_L_X8Y144_SLICE_X11Y144_AO5;
  wire [0:0] CLBLM_L_X8Y144_SLICE_X11Y144_AO6;
  wire [0:0] CLBLM_L_X8Y144_SLICE_X11Y144_AQ;
  wire [0:0] CLBLM_L_X8Y144_SLICE_X11Y144_A_CY;
  wire [0:0] CLBLM_L_X8Y144_SLICE_X11Y144_A_XOR;
  wire [0:0] CLBLM_L_X8Y144_SLICE_X11Y144_B;
  wire [0:0] CLBLM_L_X8Y144_SLICE_X11Y144_B1;
  wire [0:0] CLBLM_L_X8Y144_SLICE_X11Y144_B2;
  wire [0:0] CLBLM_L_X8Y144_SLICE_X11Y144_B3;
  wire [0:0] CLBLM_L_X8Y144_SLICE_X11Y144_B4;
  wire [0:0] CLBLM_L_X8Y144_SLICE_X11Y144_B5;
  wire [0:0] CLBLM_L_X8Y144_SLICE_X11Y144_B5Q;
  wire [0:0] CLBLM_L_X8Y144_SLICE_X11Y144_B6;
  wire [0:0] CLBLM_L_X8Y144_SLICE_X11Y144_BMUX;
  wire [0:0] CLBLM_L_X8Y144_SLICE_X11Y144_BO5;
  wire [0:0] CLBLM_L_X8Y144_SLICE_X11Y144_BO6;
  wire [0:0] CLBLM_L_X8Y144_SLICE_X11Y144_BQ;
  wire [0:0] CLBLM_L_X8Y144_SLICE_X11Y144_B_CY;
  wire [0:0] CLBLM_L_X8Y144_SLICE_X11Y144_B_XOR;
  wire [0:0] CLBLM_L_X8Y144_SLICE_X11Y144_C;
  wire [0:0] CLBLM_L_X8Y144_SLICE_X11Y144_C1;
  wire [0:0] CLBLM_L_X8Y144_SLICE_X11Y144_C2;
  wire [0:0] CLBLM_L_X8Y144_SLICE_X11Y144_C3;
  wire [0:0] CLBLM_L_X8Y144_SLICE_X11Y144_C4;
  wire [0:0] CLBLM_L_X8Y144_SLICE_X11Y144_C5;
  wire [0:0] CLBLM_L_X8Y144_SLICE_X11Y144_C6;
  wire [0:0] CLBLM_L_X8Y144_SLICE_X11Y144_CLK;
  wire [0:0] CLBLM_L_X8Y144_SLICE_X11Y144_CO5;
  wire [0:0] CLBLM_L_X8Y144_SLICE_X11Y144_CO6;
  wire [0:0] CLBLM_L_X8Y144_SLICE_X11Y144_CQ;
  wire [0:0] CLBLM_L_X8Y144_SLICE_X11Y144_C_CY;
  wire [0:0] CLBLM_L_X8Y144_SLICE_X11Y144_C_XOR;
  wire [0:0] CLBLM_L_X8Y144_SLICE_X11Y144_D;
  wire [0:0] CLBLM_L_X8Y144_SLICE_X11Y144_D1;
  wire [0:0] CLBLM_L_X8Y144_SLICE_X11Y144_D2;
  wire [0:0] CLBLM_L_X8Y144_SLICE_X11Y144_D3;
  wire [0:0] CLBLM_L_X8Y144_SLICE_X11Y144_D4;
  wire [0:0] CLBLM_L_X8Y144_SLICE_X11Y144_D5;
  wire [0:0] CLBLM_L_X8Y144_SLICE_X11Y144_D6;
  wire [0:0] CLBLM_L_X8Y144_SLICE_X11Y144_DO5;
  wire [0:0] CLBLM_L_X8Y144_SLICE_X11Y144_DO6;
  wire [0:0] CLBLM_L_X8Y144_SLICE_X11Y144_DQ;
  wire [0:0] CLBLM_L_X8Y144_SLICE_X11Y144_D_CY;
  wire [0:0] CLBLM_L_X8Y144_SLICE_X11Y144_D_XOR;
  wire [0:0] CLBLM_L_X8Y145_SLICE_X10Y145_A;
  wire [0:0] CLBLM_L_X8Y145_SLICE_X10Y145_A1;
  wire [0:0] CLBLM_L_X8Y145_SLICE_X10Y145_A2;
  wire [0:0] CLBLM_L_X8Y145_SLICE_X10Y145_A3;
  wire [0:0] CLBLM_L_X8Y145_SLICE_X10Y145_A4;
  wire [0:0] CLBLM_L_X8Y145_SLICE_X10Y145_A5;
  wire [0:0] CLBLM_L_X8Y145_SLICE_X10Y145_A5Q;
  wire [0:0] CLBLM_L_X8Y145_SLICE_X10Y145_A6;
  wire [0:0] CLBLM_L_X8Y145_SLICE_X10Y145_AMUX;
  wire [0:0] CLBLM_L_X8Y145_SLICE_X10Y145_AO5;
  wire [0:0] CLBLM_L_X8Y145_SLICE_X10Y145_AO6;
  wire [0:0] CLBLM_L_X8Y145_SLICE_X10Y145_AQ;
  wire [0:0] CLBLM_L_X8Y145_SLICE_X10Y145_A_CY;
  wire [0:0] CLBLM_L_X8Y145_SLICE_X10Y145_A_XOR;
  wire [0:0] CLBLM_L_X8Y145_SLICE_X10Y145_B;
  wire [0:0] CLBLM_L_X8Y145_SLICE_X10Y145_B1;
  wire [0:0] CLBLM_L_X8Y145_SLICE_X10Y145_B2;
  wire [0:0] CLBLM_L_X8Y145_SLICE_X10Y145_B3;
  wire [0:0] CLBLM_L_X8Y145_SLICE_X10Y145_B4;
  wire [0:0] CLBLM_L_X8Y145_SLICE_X10Y145_B5;
  wire [0:0] CLBLM_L_X8Y145_SLICE_X10Y145_B6;
  wire [0:0] CLBLM_L_X8Y145_SLICE_X10Y145_BO5;
  wire [0:0] CLBLM_L_X8Y145_SLICE_X10Y145_BO6;
  wire [0:0] CLBLM_L_X8Y145_SLICE_X10Y145_B_CY;
  wire [0:0] CLBLM_L_X8Y145_SLICE_X10Y145_B_XOR;
  wire [0:0] CLBLM_L_X8Y145_SLICE_X10Y145_C;
  wire [0:0] CLBLM_L_X8Y145_SLICE_X10Y145_C1;
  wire [0:0] CLBLM_L_X8Y145_SLICE_X10Y145_C2;
  wire [0:0] CLBLM_L_X8Y145_SLICE_X10Y145_C3;
  wire [0:0] CLBLM_L_X8Y145_SLICE_X10Y145_C4;
  wire [0:0] CLBLM_L_X8Y145_SLICE_X10Y145_C5;
  wire [0:0] CLBLM_L_X8Y145_SLICE_X10Y145_C6;
  wire [0:0] CLBLM_L_X8Y145_SLICE_X10Y145_CLK;
  wire [0:0] CLBLM_L_X8Y145_SLICE_X10Y145_CO5;
  wire [0:0] CLBLM_L_X8Y145_SLICE_X10Y145_CO6;
  wire [0:0] CLBLM_L_X8Y145_SLICE_X10Y145_C_CY;
  wire [0:0] CLBLM_L_X8Y145_SLICE_X10Y145_C_XOR;
  wire [0:0] CLBLM_L_X8Y145_SLICE_X10Y145_D;
  wire [0:0] CLBLM_L_X8Y145_SLICE_X10Y145_D1;
  wire [0:0] CLBLM_L_X8Y145_SLICE_X10Y145_D2;
  wire [0:0] CLBLM_L_X8Y145_SLICE_X10Y145_D3;
  wire [0:0] CLBLM_L_X8Y145_SLICE_X10Y145_D4;
  wire [0:0] CLBLM_L_X8Y145_SLICE_X10Y145_D5;
  wire [0:0] CLBLM_L_X8Y145_SLICE_X10Y145_D6;
  wire [0:0] CLBLM_L_X8Y145_SLICE_X10Y145_DO5;
  wire [0:0] CLBLM_L_X8Y145_SLICE_X10Y145_DO6;
  wire [0:0] CLBLM_L_X8Y145_SLICE_X10Y145_D_CY;
  wire [0:0] CLBLM_L_X8Y145_SLICE_X10Y145_D_XOR;
  wire [0:0] CLBLM_L_X8Y145_SLICE_X11Y145_A;
  wire [0:0] CLBLM_L_X8Y145_SLICE_X11Y145_A1;
  wire [0:0] CLBLM_L_X8Y145_SLICE_X11Y145_A2;
  wire [0:0] CLBLM_L_X8Y145_SLICE_X11Y145_A3;
  wire [0:0] CLBLM_L_X8Y145_SLICE_X11Y145_A4;
  wire [0:0] CLBLM_L_X8Y145_SLICE_X11Y145_A5;
  wire [0:0] CLBLM_L_X8Y145_SLICE_X11Y145_A6;
  wire [0:0] CLBLM_L_X8Y145_SLICE_X11Y145_AO5;
  wire [0:0] CLBLM_L_X8Y145_SLICE_X11Y145_AO6;
  wire [0:0] CLBLM_L_X8Y145_SLICE_X11Y145_AQ;
  wire [0:0] CLBLM_L_X8Y145_SLICE_X11Y145_A_CY;
  wire [0:0] CLBLM_L_X8Y145_SLICE_X11Y145_A_XOR;
  wire [0:0] CLBLM_L_X8Y145_SLICE_X11Y145_B;
  wire [0:0] CLBLM_L_X8Y145_SLICE_X11Y145_B1;
  wire [0:0] CLBLM_L_X8Y145_SLICE_X11Y145_B2;
  wire [0:0] CLBLM_L_X8Y145_SLICE_X11Y145_B3;
  wire [0:0] CLBLM_L_X8Y145_SLICE_X11Y145_B4;
  wire [0:0] CLBLM_L_X8Y145_SLICE_X11Y145_B5;
  wire [0:0] CLBLM_L_X8Y145_SLICE_X11Y145_B6;
  wire [0:0] CLBLM_L_X8Y145_SLICE_X11Y145_BO5;
  wire [0:0] CLBLM_L_X8Y145_SLICE_X11Y145_BO6;
  wire [0:0] CLBLM_L_X8Y145_SLICE_X11Y145_BQ;
  wire [0:0] CLBLM_L_X8Y145_SLICE_X11Y145_B_CY;
  wire [0:0] CLBLM_L_X8Y145_SLICE_X11Y145_B_XOR;
  wire [0:0] CLBLM_L_X8Y145_SLICE_X11Y145_C;
  wire [0:0] CLBLM_L_X8Y145_SLICE_X11Y145_C1;
  wire [0:0] CLBLM_L_X8Y145_SLICE_X11Y145_C2;
  wire [0:0] CLBLM_L_X8Y145_SLICE_X11Y145_C3;
  wire [0:0] CLBLM_L_X8Y145_SLICE_X11Y145_C4;
  wire [0:0] CLBLM_L_X8Y145_SLICE_X11Y145_C5;
  wire [0:0] CLBLM_L_X8Y145_SLICE_X11Y145_C5Q;
  wire [0:0] CLBLM_L_X8Y145_SLICE_X11Y145_C6;
  wire [0:0] CLBLM_L_X8Y145_SLICE_X11Y145_CLK;
  wire [0:0] CLBLM_L_X8Y145_SLICE_X11Y145_CMUX;
  wire [0:0] CLBLM_L_X8Y145_SLICE_X11Y145_CO5;
  wire [0:0] CLBLM_L_X8Y145_SLICE_X11Y145_CO6;
  wire [0:0] CLBLM_L_X8Y145_SLICE_X11Y145_CQ;
  wire [0:0] CLBLM_L_X8Y145_SLICE_X11Y145_C_CY;
  wire [0:0] CLBLM_L_X8Y145_SLICE_X11Y145_C_XOR;
  wire [0:0] CLBLM_L_X8Y145_SLICE_X11Y145_D;
  wire [0:0] CLBLM_L_X8Y145_SLICE_X11Y145_D1;
  wire [0:0] CLBLM_L_X8Y145_SLICE_X11Y145_D2;
  wire [0:0] CLBLM_L_X8Y145_SLICE_X11Y145_D3;
  wire [0:0] CLBLM_L_X8Y145_SLICE_X11Y145_D4;
  wire [0:0] CLBLM_L_X8Y145_SLICE_X11Y145_D5;
  wire [0:0] CLBLM_L_X8Y145_SLICE_X11Y145_D6;
  wire [0:0] CLBLM_L_X8Y145_SLICE_X11Y145_DO5;
  wire [0:0] CLBLM_L_X8Y145_SLICE_X11Y145_DO6;
  wire [0:0] CLBLM_L_X8Y145_SLICE_X11Y145_DQ;
  wire [0:0] CLBLM_L_X8Y145_SLICE_X11Y145_D_CY;
  wire [0:0] CLBLM_L_X8Y145_SLICE_X11Y145_D_XOR;
  wire [0:0] CLBLM_L_X8Y146_SLICE_X10Y146_A;
  wire [0:0] CLBLM_L_X8Y146_SLICE_X10Y146_A1;
  wire [0:0] CLBLM_L_X8Y146_SLICE_X10Y146_A2;
  wire [0:0] CLBLM_L_X8Y146_SLICE_X10Y146_A3;
  wire [0:0] CLBLM_L_X8Y146_SLICE_X10Y146_A4;
  wire [0:0] CLBLM_L_X8Y146_SLICE_X10Y146_A5;
  wire [0:0] CLBLM_L_X8Y146_SLICE_X10Y146_A6;
  wire [0:0] CLBLM_L_X8Y146_SLICE_X10Y146_AMUX;
  wire [0:0] CLBLM_L_X8Y146_SLICE_X10Y146_AO5;
  wire [0:0] CLBLM_L_X8Y146_SLICE_X10Y146_AO6;
  wire [0:0] CLBLM_L_X8Y146_SLICE_X10Y146_AQ;
  wire [0:0] CLBLM_L_X8Y146_SLICE_X10Y146_AX;
  wire [0:0] CLBLM_L_X8Y146_SLICE_X10Y146_A_CY;
  wire [0:0] CLBLM_L_X8Y146_SLICE_X10Y146_A_XOR;
  wire [0:0] CLBLM_L_X8Y146_SLICE_X10Y146_B;
  wire [0:0] CLBLM_L_X8Y146_SLICE_X10Y146_B1;
  wire [0:0] CLBLM_L_X8Y146_SLICE_X10Y146_B2;
  wire [0:0] CLBLM_L_X8Y146_SLICE_X10Y146_B3;
  wire [0:0] CLBLM_L_X8Y146_SLICE_X10Y146_B4;
  wire [0:0] CLBLM_L_X8Y146_SLICE_X10Y146_B5;
  wire [0:0] CLBLM_L_X8Y146_SLICE_X10Y146_B6;
  wire [0:0] CLBLM_L_X8Y146_SLICE_X10Y146_BMUX;
  wire [0:0] CLBLM_L_X8Y146_SLICE_X10Y146_BO5;
  wire [0:0] CLBLM_L_X8Y146_SLICE_X10Y146_BO6;
  wire [0:0] CLBLM_L_X8Y146_SLICE_X10Y146_BQ;
  wire [0:0] CLBLM_L_X8Y146_SLICE_X10Y146_BX;
  wire [0:0] CLBLM_L_X8Y146_SLICE_X10Y146_B_CY;
  wire [0:0] CLBLM_L_X8Y146_SLICE_X10Y146_B_XOR;
  wire [0:0] CLBLM_L_X8Y146_SLICE_X10Y146_C;
  wire [0:0] CLBLM_L_X8Y146_SLICE_X10Y146_C1;
  wire [0:0] CLBLM_L_X8Y146_SLICE_X10Y146_C2;
  wire [0:0] CLBLM_L_X8Y146_SLICE_X10Y146_C3;
  wire [0:0] CLBLM_L_X8Y146_SLICE_X10Y146_C4;
  wire [0:0] CLBLM_L_X8Y146_SLICE_X10Y146_C5;
  wire [0:0] CLBLM_L_X8Y146_SLICE_X10Y146_C6;
  wire [0:0] CLBLM_L_X8Y146_SLICE_X10Y146_CE;
  wire [0:0] CLBLM_L_X8Y146_SLICE_X10Y146_CLK;
  wire [0:0] CLBLM_L_X8Y146_SLICE_X10Y146_CMUX;
  wire [0:0] CLBLM_L_X8Y146_SLICE_X10Y146_CO5;
  wire [0:0] CLBLM_L_X8Y146_SLICE_X10Y146_CO6;
  wire [0:0] CLBLM_L_X8Y146_SLICE_X10Y146_C_CY;
  wire [0:0] CLBLM_L_X8Y146_SLICE_X10Y146_C_XOR;
  wire [0:0] CLBLM_L_X8Y146_SLICE_X10Y146_D;
  wire [0:0] CLBLM_L_X8Y146_SLICE_X10Y146_D1;
  wire [0:0] CLBLM_L_X8Y146_SLICE_X10Y146_D2;
  wire [0:0] CLBLM_L_X8Y146_SLICE_X10Y146_D3;
  wire [0:0] CLBLM_L_X8Y146_SLICE_X10Y146_D4;
  wire [0:0] CLBLM_L_X8Y146_SLICE_X10Y146_D5;
  wire [0:0] CLBLM_L_X8Y146_SLICE_X10Y146_D6;
  wire [0:0] CLBLM_L_X8Y146_SLICE_X10Y146_DO5;
  wire [0:0] CLBLM_L_X8Y146_SLICE_X10Y146_DO6;
  wire [0:0] CLBLM_L_X8Y146_SLICE_X10Y146_D_CY;
  wire [0:0] CLBLM_L_X8Y146_SLICE_X10Y146_D_XOR;
  wire [0:0] CLBLM_L_X8Y146_SLICE_X11Y146_A;
  wire [0:0] CLBLM_L_X8Y146_SLICE_X11Y146_A1;
  wire [0:0] CLBLM_L_X8Y146_SLICE_X11Y146_A2;
  wire [0:0] CLBLM_L_X8Y146_SLICE_X11Y146_A3;
  wire [0:0] CLBLM_L_X8Y146_SLICE_X11Y146_A4;
  wire [0:0] CLBLM_L_X8Y146_SLICE_X11Y146_A5;
  wire [0:0] CLBLM_L_X8Y146_SLICE_X11Y146_A6;
  wire [0:0] CLBLM_L_X8Y146_SLICE_X11Y146_AO5;
  wire [0:0] CLBLM_L_X8Y146_SLICE_X11Y146_AO6;
  wire [0:0] CLBLM_L_X8Y146_SLICE_X11Y146_AQ;
  wire [0:0] CLBLM_L_X8Y146_SLICE_X11Y146_A_CY;
  wire [0:0] CLBLM_L_X8Y146_SLICE_X11Y146_A_XOR;
  wire [0:0] CLBLM_L_X8Y146_SLICE_X11Y146_B;
  wire [0:0] CLBLM_L_X8Y146_SLICE_X11Y146_B1;
  wire [0:0] CLBLM_L_X8Y146_SLICE_X11Y146_B2;
  wire [0:0] CLBLM_L_X8Y146_SLICE_X11Y146_B3;
  wire [0:0] CLBLM_L_X8Y146_SLICE_X11Y146_B4;
  wire [0:0] CLBLM_L_X8Y146_SLICE_X11Y146_B5;
  wire [0:0] CLBLM_L_X8Y146_SLICE_X11Y146_B5Q;
  wire [0:0] CLBLM_L_X8Y146_SLICE_X11Y146_B6;
  wire [0:0] CLBLM_L_X8Y146_SLICE_X11Y146_BMUX;
  wire [0:0] CLBLM_L_X8Y146_SLICE_X11Y146_BO5;
  wire [0:0] CLBLM_L_X8Y146_SLICE_X11Y146_BO6;
  wire [0:0] CLBLM_L_X8Y146_SLICE_X11Y146_BQ;
  wire [0:0] CLBLM_L_X8Y146_SLICE_X11Y146_B_CY;
  wire [0:0] CLBLM_L_X8Y146_SLICE_X11Y146_B_XOR;
  wire [0:0] CLBLM_L_X8Y146_SLICE_X11Y146_C;
  wire [0:0] CLBLM_L_X8Y146_SLICE_X11Y146_C1;
  wire [0:0] CLBLM_L_X8Y146_SLICE_X11Y146_C2;
  wire [0:0] CLBLM_L_X8Y146_SLICE_X11Y146_C3;
  wire [0:0] CLBLM_L_X8Y146_SLICE_X11Y146_C4;
  wire [0:0] CLBLM_L_X8Y146_SLICE_X11Y146_C5;
  wire [0:0] CLBLM_L_X8Y146_SLICE_X11Y146_C5Q;
  wire [0:0] CLBLM_L_X8Y146_SLICE_X11Y146_C6;
  wire [0:0] CLBLM_L_X8Y146_SLICE_X11Y146_CLK;
  wire [0:0] CLBLM_L_X8Y146_SLICE_X11Y146_CMUX;
  wire [0:0] CLBLM_L_X8Y146_SLICE_X11Y146_CO5;
  wire [0:0] CLBLM_L_X8Y146_SLICE_X11Y146_CO6;
  wire [0:0] CLBLM_L_X8Y146_SLICE_X11Y146_CQ;
  wire [0:0] CLBLM_L_X8Y146_SLICE_X11Y146_C_CY;
  wire [0:0] CLBLM_L_X8Y146_SLICE_X11Y146_C_XOR;
  wire [0:0] CLBLM_L_X8Y146_SLICE_X11Y146_D;
  wire [0:0] CLBLM_L_X8Y146_SLICE_X11Y146_D1;
  wire [0:0] CLBLM_L_X8Y146_SLICE_X11Y146_D2;
  wire [0:0] CLBLM_L_X8Y146_SLICE_X11Y146_D3;
  wire [0:0] CLBLM_L_X8Y146_SLICE_X11Y146_D4;
  wire [0:0] CLBLM_L_X8Y146_SLICE_X11Y146_D5;
  wire [0:0] CLBLM_L_X8Y146_SLICE_X11Y146_D5Q;
  wire [0:0] CLBLM_L_X8Y146_SLICE_X11Y146_D6;
  wire [0:0] CLBLM_L_X8Y146_SLICE_X11Y146_DMUX;
  wire [0:0] CLBLM_L_X8Y146_SLICE_X11Y146_DO5;
  wire [0:0] CLBLM_L_X8Y146_SLICE_X11Y146_DO6;
  wire [0:0] CLBLM_L_X8Y146_SLICE_X11Y146_DQ;
  wire [0:0] CLBLM_L_X8Y146_SLICE_X11Y146_D_CY;
  wire [0:0] CLBLM_L_X8Y146_SLICE_X11Y146_D_XOR;
  wire [0:0] CLBLM_L_X8Y147_SLICE_X10Y147_A;
  wire [0:0] CLBLM_L_X8Y147_SLICE_X10Y147_A1;
  wire [0:0] CLBLM_L_X8Y147_SLICE_X10Y147_A2;
  wire [0:0] CLBLM_L_X8Y147_SLICE_X10Y147_A3;
  wire [0:0] CLBLM_L_X8Y147_SLICE_X10Y147_A4;
  wire [0:0] CLBLM_L_X8Y147_SLICE_X10Y147_A5;
  wire [0:0] CLBLM_L_X8Y147_SLICE_X10Y147_A6;
  wire [0:0] CLBLM_L_X8Y147_SLICE_X10Y147_AO5;
  wire [0:0] CLBLM_L_X8Y147_SLICE_X10Y147_AO6;
  wire [0:0] CLBLM_L_X8Y147_SLICE_X10Y147_AQ;
  wire [0:0] CLBLM_L_X8Y147_SLICE_X10Y147_A_CY;
  wire [0:0] CLBLM_L_X8Y147_SLICE_X10Y147_A_XOR;
  wire [0:0] CLBLM_L_X8Y147_SLICE_X10Y147_B;
  wire [0:0] CLBLM_L_X8Y147_SLICE_X10Y147_B1;
  wire [0:0] CLBLM_L_X8Y147_SLICE_X10Y147_B2;
  wire [0:0] CLBLM_L_X8Y147_SLICE_X10Y147_B3;
  wire [0:0] CLBLM_L_X8Y147_SLICE_X10Y147_B4;
  wire [0:0] CLBLM_L_X8Y147_SLICE_X10Y147_B5;
  wire [0:0] CLBLM_L_X8Y147_SLICE_X10Y147_B6;
  wire [0:0] CLBLM_L_X8Y147_SLICE_X10Y147_BO5;
  wire [0:0] CLBLM_L_X8Y147_SLICE_X10Y147_BO6;
  wire [0:0] CLBLM_L_X8Y147_SLICE_X10Y147_BQ;
  wire [0:0] CLBLM_L_X8Y147_SLICE_X10Y147_B_CY;
  wire [0:0] CLBLM_L_X8Y147_SLICE_X10Y147_B_XOR;
  wire [0:0] CLBLM_L_X8Y147_SLICE_X10Y147_C;
  wire [0:0] CLBLM_L_X8Y147_SLICE_X10Y147_C1;
  wire [0:0] CLBLM_L_X8Y147_SLICE_X10Y147_C2;
  wire [0:0] CLBLM_L_X8Y147_SLICE_X10Y147_C3;
  wire [0:0] CLBLM_L_X8Y147_SLICE_X10Y147_C4;
  wire [0:0] CLBLM_L_X8Y147_SLICE_X10Y147_C5;
  wire [0:0] CLBLM_L_X8Y147_SLICE_X10Y147_C5Q;
  wire [0:0] CLBLM_L_X8Y147_SLICE_X10Y147_C6;
  wire [0:0] CLBLM_L_X8Y147_SLICE_X10Y147_CLK;
  wire [0:0] CLBLM_L_X8Y147_SLICE_X10Y147_CMUX;
  wire [0:0] CLBLM_L_X8Y147_SLICE_X10Y147_CO5;
  wire [0:0] CLBLM_L_X8Y147_SLICE_X10Y147_CO6;
  wire [0:0] CLBLM_L_X8Y147_SLICE_X10Y147_CQ;
  wire [0:0] CLBLM_L_X8Y147_SLICE_X10Y147_C_CY;
  wire [0:0] CLBLM_L_X8Y147_SLICE_X10Y147_C_XOR;
  wire [0:0] CLBLM_L_X8Y147_SLICE_X10Y147_D;
  wire [0:0] CLBLM_L_X8Y147_SLICE_X10Y147_D1;
  wire [0:0] CLBLM_L_X8Y147_SLICE_X10Y147_D2;
  wire [0:0] CLBLM_L_X8Y147_SLICE_X10Y147_D3;
  wire [0:0] CLBLM_L_X8Y147_SLICE_X10Y147_D4;
  wire [0:0] CLBLM_L_X8Y147_SLICE_X10Y147_D5;
  wire [0:0] CLBLM_L_X8Y147_SLICE_X10Y147_D6;
  wire [0:0] CLBLM_L_X8Y147_SLICE_X10Y147_DO5;
  wire [0:0] CLBLM_L_X8Y147_SLICE_X10Y147_DO6;
  wire [0:0] CLBLM_L_X8Y147_SLICE_X10Y147_D_CY;
  wire [0:0] CLBLM_L_X8Y147_SLICE_X10Y147_D_XOR;
  wire [0:0] CLBLM_L_X8Y147_SLICE_X11Y147_A;
  wire [0:0] CLBLM_L_X8Y147_SLICE_X11Y147_A1;
  wire [0:0] CLBLM_L_X8Y147_SLICE_X11Y147_A2;
  wire [0:0] CLBLM_L_X8Y147_SLICE_X11Y147_A3;
  wire [0:0] CLBLM_L_X8Y147_SLICE_X11Y147_A4;
  wire [0:0] CLBLM_L_X8Y147_SLICE_X11Y147_A5;
  wire [0:0] CLBLM_L_X8Y147_SLICE_X11Y147_A6;
  wire [0:0] CLBLM_L_X8Y147_SLICE_X11Y147_AO5;
  wire [0:0] CLBLM_L_X8Y147_SLICE_X11Y147_AO6;
  wire [0:0] CLBLM_L_X8Y147_SLICE_X11Y147_AQ;
  wire [0:0] CLBLM_L_X8Y147_SLICE_X11Y147_A_CY;
  wire [0:0] CLBLM_L_X8Y147_SLICE_X11Y147_A_XOR;
  wire [0:0] CLBLM_L_X8Y147_SLICE_X11Y147_B;
  wire [0:0] CLBLM_L_X8Y147_SLICE_X11Y147_B1;
  wire [0:0] CLBLM_L_X8Y147_SLICE_X11Y147_B2;
  wire [0:0] CLBLM_L_X8Y147_SLICE_X11Y147_B3;
  wire [0:0] CLBLM_L_X8Y147_SLICE_X11Y147_B4;
  wire [0:0] CLBLM_L_X8Y147_SLICE_X11Y147_B5;
  wire [0:0] CLBLM_L_X8Y147_SLICE_X11Y147_B6;
  wire [0:0] CLBLM_L_X8Y147_SLICE_X11Y147_BO5;
  wire [0:0] CLBLM_L_X8Y147_SLICE_X11Y147_BO6;
  wire [0:0] CLBLM_L_X8Y147_SLICE_X11Y147_BQ;
  wire [0:0] CLBLM_L_X8Y147_SLICE_X11Y147_B_CY;
  wire [0:0] CLBLM_L_X8Y147_SLICE_X11Y147_B_XOR;
  wire [0:0] CLBLM_L_X8Y147_SLICE_X11Y147_C;
  wire [0:0] CLBLM_L_X8Y147_SLICE_X11Y147_C1;
  wire [0:0] CLBLM_L_X8Y147_SLICE_X11Y147_C2;
  wire [0:0] CLBLM_L_X8Y147_SLICE_X11Y147_C3;
  wire [0:0] CLBLM_L_X8Y147_SLICE_X11Y147_C4;
  wire [0:0] CLBLM_L_X8Y147_SLICE_X11Y147_C5;
  wire [0:0] CLBLM_L_X8Y147_SLICE_X11Y147_C5Q;
  wire [0:0] CLBLM_L_X8Y147_SLICE_X11Y147_C6;
  wire [0:0] CLBLM_L_X8Y147_SLICE_X11Y147_CLK;
  wire [0:0] CLBLM_L_X8Y147_SLICE_X11Y147_CMUX;
  wire [0:0] CLBLM_L_X8Y147_SLICE_X11Y147_CO5;
  wire [0:0] CLBLM_L_X8Y147_SLICE_X11Y147_CO6;
  wire [0:0] CLBLM_L_X8Y147_SLICE_X11Y147_CQ;
  wire [0:0] CLBLM_L_X8Y147_SLICE_X11Y147_C_CY;
  wire [0:0] CLBLM_L_X8Y147_SLICE_X11Y147_C_XOR;
  wire [0:0] CLBLM_L_X8Y147_SLICE_X11Y147_D;
  wire [0:0] CLBLM_L_X8Y147_SLICE_X11Y147_D1;
  wire [0:0] CLBLM_L_X8Y147_SLICE_X11Y147_D2;
  wire [0:0] CLBLM_L_X8Y147_SLICE_X11Y147_D3;
  wire [0:0] CLBLM_L_X8Y147_SLICE_X11Y147_D4;
  wire [0:0] CLBLM_L_X8Y147_SLICE_X11Y147_D5;
  wire [0:0] CLBLM_L_X8Y147_SLICE_X11Y147_D6;
  wire [0:0] CLBLM_L_X8Y147_SLICE_X11Y147_DO5;
  wire [0:0] CLBLM_L_X8Y147_SLICE_X11Y147_DO6;
  wire [0:0] CLBLM_L_X8Y147_SLICE_X11Y147_DQ;
  wire [0:0] CLBLM_L_X8Y147_SLICE_X11Y147_D_CY;
  wire [0:0] CLBLM_L_X8Y147_SLICE_X11Y147_D_XOR;
  wire [0:0] CLBLM_L_X8Y148_SLICE_X10Y148_A;
  wire [0:0] CLBLM_L_X8Y148_SLICE_X10Y148_A1;
  wire [0:0] CLBLM_L_X8Y148_SLICE_X10Y148_A2;
  wire [0:0] CLBLM_L_X8Y148_SLICE_X10Y148_A3;
  wire [0:0] CLBLM_L_X8Y148_SLICE_X10Y148_A4;
  wire [0:0] CLBLM_L_X8Y148_SLICE_X10Y148_A5;
  wire [0:0] CLBLM_L_X8Y148_SLICE_X10Y148_A6;
  wire [0:0] CLBLM_L_X8Y148_SLICE_X10Y148_AO5;
  wire [0:0] CLBLM_L_X8Y148_SLICE_X10Y148_AO6;
  wire [0:0] CLBLM_L_X8Y148_SLICE_X10Y148_AQ;
  wire [0:0] CLBLM_L_X8Y148_SLICE_X10Y148_A_CY;
  wire [0:0] CLBLM_L_X8Y148_SLICE_X10Y148_A_XOR;
  wire [0:0] CLBLM_L_X8Y148_SLICE_X10Y148_B;
  wire [0:0] CLBLM_L_X8Y148_SLICE_X10Y148_B1;
  wire [0:0] CLBLM_L_X8Y148_SLICE_X10Y148_B2;
  wire [0:0] CLBLM_L_X8Y148_SLICE_X10Y148_B3;
  wire [0:0] CLBLM_L_X8Y148_SLICE_X10Y148_B4;
  wire [0:0] CLBLM_L_X8Y148_SLICE_X10Y148_B5;
  wire [0:0] CLBLM_L_X8Y148_SLICE_X10Y148_B5Q;
  wire [0:0] CLBLM_L_X8Y148_SLICE_X10Y148_B6;
  wire [0:0] CLBLM_L_X8Y148_SLICE_X10Y148_BMUX;
  wire [0:0] CLBLM_L_X8Y148_SLICE_X10Y148_BO5;
  wire [0:0] CLBLM_L_X8Y148_SLICE_X10Y148_BO6;
  wire [0:0] CLBLM_L_X8Y148_SLICE_X10Y148_BQ;
  wire [0:0] CLBLM_L_X8Y148_SLICE_X10Y148_B_CY;
  wire [0:0] CLBLM_L_X8Y148_SLICE_X10Y148_B_XOR;
  wire [0:0] CLBLM_L_X8Y148_SLICE_X10Y148_C;
  wire [0:0] CLBLM_L_X8Y148_SLICE_X10Y148_C1;
  wire [0:0] CLBLM_L_X8Y148_SLICE_X10Y148_C2;
  wire [0:0] CLBLM_L_X8Y148_SLICE_X10Y148_C3;
  wire [0:0] CLBLM_L_X8Y148_SLICE_X10Y148_C4;
  wire [0:0] CLBLM_L_X8Y148_SLICE_X10Y148_C5;
  wire [0:0] CLBLM_L_X8Y148_SLICE_X10Y148_C6;
  wire [0:0] CLBLM_L_X8Y148_SLICE_X10Y148_CLK;
  wire [0:0] CLBLM_L_X8Y148_SLICE_X10Y148_CO5;
  wire [0:0] CLBLM_L_X8Y148_SLICE_X10Y148_CO6;
  wire [0:0] CLBLM_L_X8Y148_SLICE_X10Y148_C_CY;
  wire [0:0] CLBLM_L_X8Y148_SLICE_X10Y148_C_XOR;
  wire [0:0] CLBLM_L_X8Y148_SLICE_X10Y148_D;
  wire [0:0] CLBLM_L_X8Y148_SLICE_X10Y148_D1;
  wire [0:0] CLBLM_L_X8Y148_SLICE_X10Y148_D2;
  wire [0:0] CLBLM_L_X8Y148_SLICE_X10Y148_D3;
  wire [0:0] CLBLM_L_X8Y148_SLICE_X10Y148_D4;
  wire [0:0] CLBLM_L_X8Y148_SLICE_X10Y148_D5;
  wire [0:0] CLBLM_L_X8Y148_SLICE_X10Y148_D6;
  wire [0:0] CLBLM_L_X8Y148_SLICE_X10Y148_DO5;
  wire [0:0] CLBLM_L_X8Y148_SLICE_X10Y148_DO6;
  wire [0:0] CLBLM_L_X8Y148_SLICE_X10Y148_D_CY;
  wire [0:0] CLBLM_L_X8Y148_SLICE_X10Y148_D_XOR;
  wire [0:0] CLBLM_L_X8Y148_SLICE_X11Y148_A;
  wire [0:0] CLBLM_L_X8Y148_SLICE_X11Y148_A1;
  wire [0:0] CLBLM_L_X8Y148_SLICE_X11Y148_A2;
  wire [0:0] CLBLM_L_X8Y148_SLICE_X11Y148_A3;
  wire [0:0] CLBLM_L_X8Y148_SLICE_X11Y148_A4;
  wire [0:0] CLBLM_L_X8Y148_SLICE_X11Y148_A5;
  wire [0:0] CLBLM_L_X8Y148_SLICE_X11Y148_A6;
  wire [0:0] CLBLM_L_X8Y148_SLICE_X11Y148_AO5;
  wire [0:0] CLBLM_L_X8Y148_SLICE_X11Y148_AO6;
  wire [0:0] CLBLM_L_X8Y148_SLICE_X11Y148_AQ;
  wire [0:0] CLBLM_L_X8Y148_SLICE_X11Y148_A_CY;
  wire [0:0] CLBLM_L_X8Y148_SLICE_X11Y148_A_XOR;
  wire [0:0] CLBLM_L_X8Y148_SLICE_X11Y148_B;
  wire [0:0] CLBLM_L_X8Y148_SLICE_X11Y148_B1;
  wire [0:0] CLBLM_L_X8Y148_SLICE_X11Y148_B2;
  wire [0:0] CLBLM_L_X8Y148_SLICE_X11Y148_B3;
  wire [0:0] CLBLM_L_X8Y148_SLICE_X11Y148_B4;
  wire [0:0] CLBLM_L_X8Y148_SLICE_X11Y148_B5;
  wire [0:0] CLBLM_L_X8Y148_SLICE_X11Y148_B5Q;
  wire [0:0] CLBLM_L_X8Y148_SLICE_X11Y148_B6;
  wire [0:0] CLBLM_L_X8Y148_SLICE_X11Y148_BMUX;
  wire [0:0] CLBLM_L_X8Y148_SLICE_X11Y148_BO5;
  wire [0:0] CLBLM_L_X8Y148_SLICE_X11Y148_BO6;
  wire [0:0] CLBLM_L_X8Y148_SLICE_X11Y148_BQ;
  wire [0:0] CLBLM_L_X8Y148_SLICE_X11Y148_B_CY;
  wire [0:0] CLBLM_L_X8Y148_SLICE_X11Y148_B_XOR;
  wire [0:0] CLBLM_L_X8Y148_SLICE_X11Y148_C;
  wire [0:0] CLBLM_L_X8Y148_SLICE_X11Y148_C1;
  wire [0:0] CLBLM_L_X8Y148_SLICE_X11Y148_C2;
  wire [0:0] CLBLM_L_X8Y148_SLICE_X11Y148_C3;
  wire [0:0] CLBLM_L_X8Y148_SLICE_X11Y148_C4;
  wire [0:0] CLBLM_L_X8Y148_SLICE_X11Y148_C5;
  wire [0:0] CLBLM_L_X8Y148_SLICE_X11Y148_C6;
  wire [0:0] CLBLM_L_X8Y148_SLICE_X11Y148_CLK;
  wire [0:0] CLBLM_L_X8Y148_SLICE_X11Y148_CO5;
  wire [0:0] CLBLM_L_X8Y148_SLICE_X11Y148_CO6;
  wire [0:0] CLBLM_L_X8Y148_SLICE_X11Y148_C_CY;
  wire [0:0] CLBLM_L_X8Y148_SLICE_X11Y148_C_XOR;
  wire [0:0] CLBLM_L_X8Y148_SLICE_X11Y148_D;
  wire [0:0] CLBLM_L_X8Y148_SLICE_X11Y148_D1;
  wire [0:0] CLBLM_L_X8Y148_SLICE_X11Y148_D2;
  wire [0:0] CLBLM_L_X8Y148_SLICE_X11Y148_D3;
  wire [0:0] CLBLM_L_X8Y148_SLICE_X11Y148_D4;
  wire [0:0] CLBLM_L_X8Y148_SLICE_X11Y148_D5;
  wire [0:0] CLBLM_L_X8Y148_SLICE_X11Y148_D6;
  wire [0:0] CLBLM_L_X8Y148_SLICE_X11Y148_DO5;
  wire [0:0] CLBLM_L_X8Y148_SLICE_X11Y148_DO6;
  wire [0:0] CLBLM_L_X8Y148_SLICE_X11Y148_D_CY;
  wire [0:0] CLBLM_L_X8Y148_SLICE_X11Y148_D_XOR;
  wire [0:0] CLBLM_L_X8Y149_SLICE_X10Y149_A;
  wire [0:0] CLBLM_L_X8Y149_SLICE_X10Y149_A1;
  wire [0:0] CLBLM_L_X8Y149_SLICE_X10Y149_A2;
  wire [0:0] CLBLM_L_X8Y149_SLICE_X10Y149_A3;
  wire [0:0] CLBLM_L_X8Y149_SLICE_X10Y149_A4;
  wire [0:0] CLBLM_L_X8Y149_SLICE_X10Y149_A5;
  wire [0:0] CLBLM_L_X8Y149_SLICE_X10Y149_A6;
  wire [0:0] CLBLM_L_X8Y149_SLICE_X10Y149_AO5;
  wire [0:0] CLBLM_L_X8Y149_SLICE_X10Y149_AO6;
  wire [0:0] CLBLM_L_X8Y149_SLICE_X10Y149_AQ;
  wire [0:0] CLBLM_L_X8Y149_SLICE_X10Y149_AX;
  wire [0:0] CLBLM_L_X8Y149_SLICE_X10Y149_A_CY;
  wire [0:0] CLBLM_L_X8Y149_SLICE_X10Y149_A_XOR;
  wire [0:0] CLBLM_L_X8Y149_SLICE_X10Y149_B;
  wire [0:0] CLBLM_L_X8Y149_SLICE_X10Y149_B1;
  wire [0:0] CLBLM_L_X8Y149_SLICE_X10Y149_B2;
  wire [0:0] CLBLM_L_X8Y149_SLICE_X10Y149_B3;
  wire [0:0] CLBLM_L_X8Y149_SLICE_X10Y149_B4;
  wire [0:0] CLBLM_L_X8Y149_SLICE_X10Y149_B5;
  wire [0:0] CLBLM_L_X8Y149_SLICE_X10Y149_B6;
  wire [0:0] CLBLM_L_X8Y149_SLICE_X10Y149_BO5;
  wire [0:0] CLBLM_L_X8Y149_SLICE_X10Y149_BO6;
  wire [0:0] CLBLM_L_X8Y149_SLICE_X10Y149_B_CY;
  wire [0:0] CLBLM_L_X8Y149_SLICE_X10Y149_B_XOR;
  wire [0:0] CLBLM_L_X8Y149_SLICE_X10Y149_C;
  wire [0:0] CLBLM_L_X8Y149_SLICE_X10Y149_C1;
  wire [0:0] CLBLM_L_X8Y149_SLICE_X10Y149_C2;
  wire [0:0] CLBLM_L_X8Y149_SLICE_X10Y149_C3;
  wire [0:0] CLBLM_L_X8Y149_SLICE_X10Y149_C4;
  wire [0:0] CLBLM_L_X8Y149_SLICE_X10Y149_C5;
  wire [0:0] CLBLM_L_X8Y149_SLICE_X10Y149_C6;
  wire [0:0] CLBLM_L_X8Y149_SLICE_X10Y149_CE;
  wire [0:0] CLBLM_L_X8Y149_SLICE_X10Y149_CLK;
  wire [0:0] CLBLM_L_X8Y149_SLICE_X10Y149_CO5;
  wire [0:0] CLBLM_L_X8Y149_SLICE_X10Y149_CO6;
  wire [0:0] CLBLM_L_X8Y149_SLICE_X10Y149_C_CY;
  wire [0:0] CLBLM_L_X8Y149_SLICE_X10Y149_C_XOR;
  wire [0:0] CLBLM_L_X8Y149_SLICE_X10Y149_D;
  wire [0:0] CLBLM_L_X8Y149_SLICE_X10Y149_D1;
  wire [0:0] CLBLM_L_X8Y149_SLICE_X10Y149_D2;
  wire [0:0] CLBLM_L_X8Y149_SLICE_X10Y149_D3;
  wire [0:0] CLBLM_L_X8Y149_SLICE_X10Y149_D4;
  wire [0:0] CLBLM_L_X8Y149_SLICE_X10Y149_D5;
  wire [0:0] CLBLM_L_X8Y149_SLICE_X10Y149_D6;
  wire [0:0] CLBLM_L_X8Y149_SLICE_X10Y149_DO5;
  wire [0:0] CLBLM_L_X8Y149_SLICE_X10Y149_DO6;
  wire [0:0] CLBLM_L_X8Y149_SLICE_X10Y149_D_CY;
  wire [0:0] CLBLM_L_X8Y149_SLICE_X10Y149_D_XOR;
  wire [0:0] CLBLM_L_X8Y149_SLICE_X11Y149_A;
  wire [0:0] CLBLM_L_X8Y149_SLICE_X11Y149_A1;
  wire [0:0] CLBLM_L_X8Y149_SLICE_X11Y149_A2;
  wire [0:0] CLBLM_L_X8Y149_SLICE_X11Y149_A3;
  wire [0:0] CLBLM_L_X8Y149_SLICE_X11Y149_A4;
  wire [0:0] CLBLM_L_X8Y149_SLICE_X11Y149_A5;
  wire [0:0] CLBLM_L_X8Y149_SLICE_X11Y149_A5Q;
  wire [0:0] CLBLM_L_X8Y149_SLICE_X11Y149_A6;
  wire [0:0] CLBLM_L_X8Y149_SLICE_X11Y149_AMUX;
  wire [0:0] CLBLM_L_X8Y149_SLICE_X11Y149_AO5;
  wire [0:0] CLBLM_L_X8Y149_SLICE_X11Y149_AO6;
  wire [0:0] CLBLM_L_X8Y149_SLICE_X11Y149_AQ;
  wire [0:0] CLBLM_L_X8Y149_SLICE_X11Y149_A_CY;
  wire [0:0] CLBLM_L_X8Y149_SLICE_X11Y149_A_XOR;
  wire [0:0] CLBLM_L_X8Y149_SLICE_X11Y149_B;
  wire [0:0] CLBLM_L_X8Y149_SLICE_X11Y149_B1;
  wire [0:0] CLBLM_L_X8Y149_SLICE_X11Y149_B2;
  wire [0:0] CLBLM_L_X8Y149_SLICE_X11Y149_B3;
  wire [0:0] CLBLM_L_X8Y149_SLICE_X11Y149_B4;
  wire [0:0] CLBLM_L_X8Y149_SLICE_X11Y149_B5;
  wire [0:0] CLBLM_L_X8Y149_SLICE_X11Y149_B6;
  wire [0:0] CLBLM_L_X8Y149_SLICE_X11Y149_BO5;
  wire [0:0] CLBLM_L_X8Y149_SLICE_X11Y149_BO6;
  wire [0:0] CLBLM_L_X8Y149_SLICE_X11Y149_B_CY;
  wire [0:0] CLBLM_L_X8Y149_SLICE_X11Y149_B_XOR;
  wire [0:0] CLBLM_L_X8Y149_SLICE_X11Y149_C;
  wire [0:0] CLBLM_L_X8Y149_SLICE_X11Y149_C1;
  wire [0:0] CLBLM_L_X8Y149_SLICE_X11Y149_C2;
  wire [0:0] CLBLM_L_X8Y149_SLICE_X11Y149_C3;
  wire [0:0] CLBLM_L_X8Y149_SLICE_X11Y149_C4;
  wire [0:0] CLBLM_L_X8Y149_SLICE_X11Y149_C5;
  wire [0:0] CLBLM_L_X8Y149_SLICE_X11Y149_C6;
  wire [0:0] CLBLM_L_X8Y149_SLICE_X11Y149_CLK;
  wire [0:0] CLBLM_L_X8Y149_SLICE_X11Y149_CO5;
  wire [0:0] CLBLM_L_X8Y149_SLICE_X11Y149_CO6;
  wire [0:0] CLBLM_L_X8Y149_SLICE_X11Y149_C_CY;
  wire [0:0] CLBLM_L_X8Y149_SLICE_X11Y149_C_XOR;
  wire [0:0] CLBLM_L_X8Y149_SLICE_X11Y149_D;
  wire [0:0] CLBLM_L_X8Y149_SLICE_X11Y149_D1;
  wire [0:0] CLBLM_L_X8Y149_SLICE_X11Y149_D2;
  wire [0:0] CLBLM_L_X8Y149_SLICE_X11Y149_D3;
  wire [0:0] CLBLM_L_X8Y149_SLICE_X11Y149_D4;
  wire [0:0] CLBLM_L_X8Y149_SLICE_X11Y149_D5;
  wire [0:0] CLBLM_L_X8Y149_SLICE_X11Y149_D6;
  wire [0:0] CLBLM_L_X8Y149_SLICE_X11Y149_DO5;
  wire [0:0] CLBLM_L_X8Y149_SLICE_X11Y149_DO6;
  wire [0:0] CLBLM_L_X8Y149_SLICE_X11Y149_D_CY;
  wire [0:0] CLBLM_L_X8Y149_SLICE_X11Y149_D_XOR;
  wire [0:0] CLBLM_L_X8Y150_SLICE_X10Y150_A;
  wire [0:0] CLBLM_L_X8Y150_SLICE_X10Y150_A1;
  wire [0:0] CLBLM_L_X8Y150_SLICE_X10Y150_A2;
  wire [0:0] CLBLM_L_X8Y150_SLICE_X10Y150_A3;
  wire [0:0] CLBLM_L_X8Y150_SLICE_X10Y150_A4;
  wire [0:0] CLBLM_L_X8Y150_SLICE_X10Y150_A5;
  wire [0:0] CLBLM_L_X8Y150_SLICE_X10Y150_A6;
  wire [0:0] CLBLM_L_X8Y150_SLICE_X10Y150_AO5;
  wire [0:0] CLBLM_L_X8Y150_SLICE_X10Y150_AO6;
  wire [0:0] CLBLM_L_X8Y150_SLICE_X10Y150_AQ;
  wire [0:0] CLBLM_L_X8Y150_SLICE_X10Y150_A_CY;
  wire [0:0] CLBLM_L_X8Y150_SLICE_X10Y150_A_XOR;
  wire [0:0] CLBLM_L_X8Y150_SLICE_X10Y150_B;
  wire [0:0] CLBLM_L_X8Y150_SLICE_X10Y150_B1;
  wire [0:0] CLBLM_L_X8Y150_SLICE_X10Y150_B2;
  wire [0:0] CLBLM_L_X8Y150_SLICE_X10Y150_B3;
  wire [0:0] CLBLM_L_X8Y150_SLICE_X10Y150_B4;
  wire [0:0] CLBLM_L_X8Y150_SLICE_X10Y150_B5;
  wire [0:0] CLBLM_L_X8Y150_SLICE_X10Y150_B6;
  wire [0:0] CLBLM_L_X8Y150_SLICE_X10Y150_BMUX;
  wire [0:0] CLBLM_L_X8Y150_SLICE_X10Y150_BO5;
  wire [0:0] CLBLM_L_X8Y150_SLICE_X10Y150_BO6;
  wire [0:0] CLBLM_L_X8Y150_SLICE_X10Y150_B_CY;
  wire [0:0] CLBLM_L_X8Y150_SLICE_X10Y150_B_XOR;
  wire [0:0] CLBLM_L_X8Y150_SLICE_X10Y150_C;
  wire [0:0] CLBLM_L_X8Y150_SLICE_X10Y150_C1;
  wire [0:0] CLBLM_L_X8Y150_SLICE_X10Y150_C2;
  wire [0:0] CLBLM_L_X8Y150_SLICE_X10Y150_C3;
  wire [0:0] CLBLM_L_X8Y150_SLICE_X10Y150_C4;
  wire [0:0] CLBLM_L_X8Y150_SLICE_X10Y150_C5;
  wire [0:0] CLBLM_L_X8Y150_SLICE_X10Y150_C6;
  wire [0:0] CLBLM_L_X8Y150_SLICE_X10Y150_CLK;
  wire [0:0] CLBLM_L_X8Y150_SLICE_X10Y150_CMUX;
  wire [0:0] CLBLM_L_X8Y150_SLICE_X10Y150_CO5;
  wire [0:0] CLBLM_L_X8Y150_SLICE_X10Y150_CO6;
  wire [0:0] CLBLM_L_X8Y150_SLICE_X10Y150_C_CY;
  wire [0:0] CLBLM_L_X8Y150_SLICE_X10Y150_C_XOR;
  wire [0:0] CLBLM_L_X8Y150_SLICE_X10Y150_D;
  wire [0:0] CLBLM_L_X8Y150_SLICE_X10Y150_D1;
  wire [0:0] CLBLM_L_X8Y150_SLICE_X10Y150_D2;
  wire [0:0] CLBLM_L_X8Y150_SLICE_X10Y150_D3;
  wire [0:0] CLBLM_L_X8Y150_SLICE_X10Y150_D4;
  wire [0:0] CLBLM_L_X8Y150_SLICE_X10Y150_D5;
  wire [0:0] CLBLM_L_X8Y150_SLICE_X10Y150_D6;
  wire [0:0] CLBLM_L_X8Y150_SLICE_X10Y150_DO5;
  wire [0:0] CLBLM_L_X8Y150_SLICE_X10Y150_DO6;
  wire [0:0] CLBLM_L_X8Y150_SLICE_X10Y150_D_CY;
  wire [0:0] CLBLM_L_X8Y150_SLICE_X10Y150_D_XOR;
  wire [0:0] CLBLM_L_X8Y150_SLICE_X11Y150_A;
  wire [0:0] CLBLM_L_X8Y150_SLICE_X11Y150_A1;
  wire [0:0] CLBLM_L_X8Y150_SLICE_X11Y150_A2;
  wire [0:0] CLBLM_L_X8Y150_SLICE_X11Y150_A3;
  wire [0:0] CLBLM_L_X8Y150_SLICE_X11Y150_A4;
  wire [0:0] CLBLM_L_X8Y150_SLICE_X11Y150_A5;
  wire [0:0] CLBLM_L_X8Y150_SLICE_X11Y150_A6;
  wire [0:0] CLBLM_L_X8Y150_SLICE_X11Y150_AO5;
  wire [0:0] CLBLM_L_X8Y150_SLICE_X11Y150_AO6;
  wire [0:0] CLBLM_L_X8Y150_SLICE_X11Y150_AQ;
  wire [0:0] CLBLM_L_X8Y150_SLICE_X11Y150_A_CY;
  wire [0:0] CLBLM_L_X8Y150_SLICE_X11Y150_A_XOR;
  wire [0:0] CLBLM_L_X8Y150_SLICE_X11Y150_B;
  wire [0:0] CLBLM_L_X8Y150_SLICE_X11Y150_B1;
  wire [0:0] CLBLM_L_X8Y150_SLICE_X11Y150_B2;
  wire [0:0] CLBLM_L_X8Y150_SLICE_X11Y150_B3;
  wire [0:0] CLBLM_L_X8Y150_SLICE_X11Y150_B4;
  wire [0:0] CLBLM_L_X8Y150_SLICE_X11Y150_B5;
  wire [0:0] CLBLM_L_X8Y150_SLICE_X11Y150_B6;
  wire [0:0] CLBLM_L_X8Y150_SLICE_X11Y150_BMUX;
  wire [0:0] CLBLM_L_X8Y150_SLICE_X11Y150_BO5;
  wire [0:0] CLBLM_L_X8Y150_SLICE_X11Y150_BO6;
  wire [0:0] CLBLM_L_X8Y150_SLICE_X11Y150_B_CY;
  wire [0:0] CLBLM_L_X8Y150_SLICE_X11Y150_B_XOR;
  wire [0:0] CLBLM_L_X8Y150_SLICE_X11Y150_C;
  wire [0:0] CLBLM_L_X8Y150_SLICE_X11Y150_C1;
  wire [0:0] CLBLM_L_X8Y150_SLICE_X11Y150_C2;
  wire [0:0] CLBLM_L_X8Y150_SLICE_X11Y150_C3;
  wire [0:0] CLBLM_L_X8Y150_SLICE_X11Y150_C4;
  wire [0:0] CLBLM_L_X8Y150_SLICE_X11Y150_C5;
  wire [0:0] CLBLM_L_X8Y150_SLICE_X11Y150_C6;
  wire [0:0] CLBLM_L_X8Y150_SLICE_X11Y150_CLK;
  wire [0:0] CLBLM_L_X8Y150_SLICE_X11Y150_CO5;
  wire [0:0] CLBLM_L_X8Y150_SLICE_X11Y150_CO6;
  wire [0:0] CLBLM_L_X8Y150_SLICE_X11Y150_C_CY;
  wire [0:0] CLBLM_L_X8Y150_SLICE_X11Y150_C_XOR;
  wire [0:0] CLBLM_L_X8Y150_SLICE_X11Y150_D;
  wire [0:0] CLBLM_L_X8Y150_SLICE_X11Y150_D1;
  wire [0:0] CLBLM_L_X8Y150_SLICE_X11Y150_D2;
  wire [0:0] CLBLM_L_X8Y150_SLICE_X11Y150_D3;
  wire [0:0] CLBLM_L_X8Y150_SLICE_X11Y150_D4;
  wire [0:0] CLBLM_L_X8Y150_SLICE_X11Y150_D5;
  wire [0:0] CLBLM_L_X8Y150_SLICE_X11Y150_D6;
  wire [0:0] CLBLM_L_X8Y150_SLICE_X11Y150_DO5;
  wire [0:0] CLBLM_L_X8Y150_SLICE_X11Y150_DO6;
  wire [0:0] CLBLM_L_X8Y150_SLICE_X11Y150_D_CY;
  wire [0:0] CLBLM_L_X8Y150_SLICE_X11Y150_D_XOR;
  wire [0:0] CLBLM_L_X8Y151_SLICE_X10Y151_A;
  wire [0:0] CLBLM_L_X8Y151_SLICE_X10Y151_A1;
  wire [0:0] CLBLM_L_X8Y151_SLICE_X10Y151_A2;
  wire [0:0] CLBLM_L_X8Y151_SLICE_X10Y151_A3;
  wire [0:0] CLBLM_L_X8Y151_SLICE_X10Y151_A4;
  wire [0:0] CLBLM_L_X8Y151_SLICE_X10Y151_A5;
  wire [0:0] CLBLM_L_X8Y151_SLICE_X10Y151_A5Q;
  wire [0:0] CLBLM_L_X8Y151_SLICE_X10Y151_A6;
  wire [0:0] CLBLM_L_X8Y151_SLICE_X10Y151_AMUX;
  wire [0:0] CLBLM_L_X8Y151_SLICE_X10Y151_AO5;
  wire [0:0] CLBLM_L_X8Y151_SLICE_X10Y151_AO6;
  wire [0:0] CLBLM_L_X8Y151_SLICE_X10Y151_AQ;
  wire [0:0] CLBLM_L_X8Y151_SLICE_X10Y151_A_CY;
  wire [0:0] CLBLM_L_X8Y151_SLICE_X10Y151_A_XOR;
  wire [0:0] CLBLM_L_X8Y151_SLICE_X10Y151_B;
  wire [0:0] CLBLM_L_X8Y151_SLICE_X10Y151_B1;
  wire [0:0] CLBLM_L_X8Y151_SLICE_X10Y151_B2;
  wire [0:0] CLBLM_L_X8Y151_SLICE_X10Y151_B3;
  wire [0:0] CLBLM_L_X8Y151_SLICE_X10Y151_B4;
  wire [0:0] CLBLM_L_X8Y151_SLICE_X10Y151_B5;
  wire [0:0] CLBLM_L_X8Y151_SLICE_X10Y151_B5Q;
  wire [0:0] CLBLM_L_X8Y151_SLICE_X10Y151_B6;
  wire [0:0] CLBLM_L_X8Y151_SLICE_X10Y151_BMUX;
  wire [0:0] CLBLM_L_X8Y151_SLICE_X10Y151_BO5;
  wire [0:0] CLBLM_L_X8Y151_SLICE_X10Y151_BO6;
  wire [0:0] CLBLM_L_X8Y151_SLICE_X10Y151_BQ;
  wire [0:0] CLBLM_L_X8Y151_SLICE_X10Y151_B_CY;
  wire [0:0] CLBLM_L_X8Y151_SLICE_X10Y151_B_XOR;
  wire [0:0] CLBLM_L_X8Y151_SLICE_X10Y151_C;
  wire [0:0] CLBLM_L_X8Y151_SLICE_X10Y151_C1;
  wire [0:0] CLBLM_L_X8Y151_SLICE_X10Y151_C2;
  wire [0:0] CLBLM_L_X8Y151_SLICE_X10Y151_C3;
  wire [0:0] CLBLM_L_X8Y151_SLICE_X10Y151_C4;
  wire [0:0] CLBLM_L_X8Y151_SLICE_X10Y151_C5;
  wire [0:0] CLBLM_L_X8Y151_SLICE_X10Y151_C5Q;
  wire [0:0] CLBLM_L_X8Y151_SLICE_X10Y151_C6;
  wire [0:0] CLBLM_L_X8Y151_SLICE_X10Y151_CLK;
  wire [0:0] CLBLM_L_X8Y151_SLICE_X10Y151_CMUX;
  wire [0:0] CLBLM_L_X8Y151_SLICE_X10Y151_CO5;
  wire [0:0] CLBLM_L_X8Y151_SLICE_X10Y151_CO6;
  wire [0:0] CLBLM_L_X8Y151_SLICE_X10Y151_CQ;
  wire [0:0] CLBLM_L_X8Y151_SLICE_X10Y151_C_CY;
  wire [0:0] CLBLM_L_X8Y151_SLICE_X10Y151_C_XOR;
  wire [0:0] CLBLM_L_X8Y151_SLICE_X10Y151_D;
  wire [0:0] CLBLM_L_X8Y151_SLICE_X10Y151_D1;
  wire [0:0] CLBLM_L_X8Y151_SLICE_X10Y151_D2;
  wire [0:0] CLBLM_L_X8Y151_SLICE_X10Y151_D3;
  wire [0:0] CLBLM_L_X8Y151_SLICE_X10Y151_D4;
  wire [0:0] CLBLM_L_X8Y151_SLICE_X10Y151_D5;
  wire [0:0] CLBLM_L_X8Y151_SLICE_X10Y151_D6;
  wire [0:0] CLBLM_L_X8Y151_SLICE_X10Y151_DO5;
  wire [0:0] CLBLM_L_X8Y151_SLICE_X10Y151_DO6;
  wire [0:0] CLBLM_L_X8Y151_SLICE_X10Y151_D_CY;
  wire [0:0] CLBLM_L_X8Y151_SLICE_X10Y151_D_XOR;
  wire [0:0] CLBLM_L_X8Y151_SLICE_X11Y151_A;
  wire [0:0] CLBLM_L_X8Y151_SLICE_X11Y151_A1;
  wire [0:0] CLBLM_L_X8Y151_SLICE_X11Y151_A2;
  wire [0:0] CLBLM_L_X8Y151_SLICE_X11Y151_A3;
  wire [0:0] CLBLM_L_X8Y151_SLICE_X11Y151_A4;
  wire [0:0] CLBLM_L_X8Y151_SLICE_X11Y151_A5;
  wire [0:0] CLBLM_L_X8Y151_SLICE_X11Y151_A6;
  wire [0:0] CLBLM_L_X8Y151_SLICE_X11Y151_AO5;
  wire [0:0] CLBLM_L_X8Y151_SLICE_X11Y151_AO6;
  wire [0:0] CLBLM_L_X8Y151_SLICE_X11Y151_AQ;
  wire [0:0] CLBLM_L_X8Y151_SLICE_X11Y151_A_CY;
  wire [0:0] CLBLM_L_X8Y151_SLICE_X11Y151_A_XOR;
  wire [0:0] CLBLM_L_X8Y151_SLICE_X11Y151_B;
  wire [0:0] CLBLM_L_X8Y151_SLICE_X11Y151_B1;
  wire [0:0] CLBLM_L_X8Y151_SLICE_X11Y151_B2;
  wire [0:0] CLBLM_L_X8Y151_SLICE_X11Y151_B3;
  wire [0:0] CLBLM_L_X8Y151_SLICE_X11Y151_B4;
  wire [0:0] CLBLM_L_X8Y151_SLICE_X11Y151_B5;
  wire [0:0] CLBLM_L_X8Y151_SLICE_X11Y151_B6;
  wire [0:0] CLBLM_L_X8Y151_SLICE_X11Y151_BO5;
  wire [0:0] CLBLM_L_X8Y151_SLICE_X11Y151_BO6;
  wire [0:0] CLBLM_L_X8Y151_SLICE_X11Y151_B_CY;
  wire [0:0] CLBLM_L_X8Y151_SLICE_X11Y151_B_XOR;
  wire [0:0] CLBLM_L_X8Y151_SLICE_X11Y151_C;
  wire [0:0] CLBLM_L_X8Y151_SLICE_X11Y151_C1;
  wire [0:0] CLBLM_L_X8Y151_SLICE_X11Y151_C2;
  wire [0:0] CLBLM_L_X8Y151_SLICE_X11Y151_C3;
  wire [0:0] CLBLM_L_X8Y151_SLICE_X11Y151_C4;
  wire [0:0] CLBLM_L_X8Y151_SLICE_X11Y151_C5;
  wire [0:0] CLBLM_L_X8Y151_SLICE_X11Y151_C6;
  wire [0:0] CLBLM_L_X8Y151_SLICE_X11Y151_CLK;
  wire [0:0] CLBLM_L_X8Y151_SLICE_X11Y151_CO5;
  wire [0:0] CLBLM_L_X8Y151_SLICE_X11Y151_CO6;
  wire [0:0] CLBLM_L_X8Y151_SLICE_X11Y151_C_CY;
  wire [0:0] CLBLM_L_X8Y151_SLICE_X11Y151_C_XOR;
  wire [0:0] CLBLM_L_X8Y151_SLICE_X11Y151_D;
  wire [0:0] CLBLM_L_X8Y151_SLICE_X11Y151_D1;
  wire [0:0] CLBLM_L_X8Y151_SLICE_X11Y151_D2;
  wire [0:0] CLBLM_L_X8Y151_SLICE_X11Y151_D3;
  wire [0:0] CLBLM_L_X8Y151_SLICE_X11Y151_D4;
  wire [0:0] CLBLM_L_X8Y151_SLICE_X11Y151_D5;
  wire [0:0] CLBLM_L_X8Y151_SLICE_X11Y151_D6;
  wire [0:0] CLBLM_L_X8Y151_SLICE_X11Y151_DO5;
  wire [0:0] CLBLM_L_X8Y151_SLICE_X11Y151_DO6;
  wire [0:0] CLBLM_L_X8Y151_SLICE_X11Y151_D_CY;
  wire [0:0] CLBLM_L_X8Y151_SLICE_X11Y151_D_XOR;
  wire [0:0] CLBLM_L_X8Y152_SLICE_X10Y152_A;
  wire [0:0] CLBLM_L_X8Y152_SLICE_X10Y152_A1;
  wire [0:0] CLBLM_L_X8Y152_SLICE_X10Y152_A2;
  wire [0:0] CLBLM_L_X8Y152_SLICE_X10Y152_A3;
  wire [0:0] CLBLM_L_X8Y152_SLICE_X10Y152_A4;
  wire [0:0] CLBLM_L_X8Y152_SLICE_X10Y152_A5;
  wire [0:0] CLBLM_L_X8Y152_SLICE_X10Y152_A5Q;
  wire [0:0] CLBLM_L_X8Y152_SLICE_X10Y152_A6;
  wire [0:0] CLBLM_L_X8Y152_SLICE_X10Y152_AMUX;
  wire [0:0] CLBLM_L_X8Y152_SLICE_X10Y152_AO5;
  wire [0:0] CLBLM_L_X8Y152_SLICE_X10Y152_AO6;
  wire [0:0] CLBLM_L_X8Y152_SLICE_X10Y152_AQ;
  wire [0:0] CLBLM_L_X8Y152_SLICE_X10Y152_AX;
  wire [0:0] CLBLM_L_X8Y152_SLICE_X10Y152_A_CY;
  wire [0:0] CLBLM_L_X8Y152_SLICE_X10Y152_A_XOR;
  wire [0:0] CLBLM_L_X8Y152_SLICE_X10Y152_B;
  wire [0:0] CLBLM_L_X8Y152_SLICE_X10Y152_B1;
  wire [0:0] CLBLM_L_X8Y152_SLICE_X10Y152_B2;
  wire [0:0] CLBLM_L_X8Y152_SLICE_X10Y152_B3;
  wire [0:0] CLBLM_L_X8Y152_SLICE_X10Y152_B4;
  wire [0:0] CLBLM_L_X8Y152_SLICE_X10Y152_B5;
  wire [0:0] CLBLM_L_X8Y152_SLICE_X10Y152_B6;
  wire [0:0] CLBLM_L_X8Y152_SLICE_X10Y152_BO5;
  wire [0:0] CLBLM_L_X8Y152_SLICE_X10Y152_BO6;
  wire [0:0] CLBLM_L_X8Y152_SLICE_X10Y152_BQ;
  wire [0:0] CLBLM_L_X8Y152_SLICE_X10Y152_B_CY;
  wire [0:0] CLBLM_L_X8Y152_SLICE_X10Y152_B_XOR;
  wire [0:0] CLBLM_L_X8Y152_SLICE_X10Y152_C;
  wire [0:0] CLBLM_L_X8Y152_SLICE_X10Y152_C1;
  wire [0:0] CLBLM_L_X8Y152_SLICE_X10Y152_C2;
  wire [0:0] CLBLM_L_X8Y152_SLICE_X10Y152_C3;
  wire [0:0] CLBLM_L_X8Y152_SLICE_X10Y152_C4;
  wire [0:0] CLBLM_L_X8Y152_SLICE_X10Y152_C5;
  wire [0:0] CLBLM_L_X8Y152_SLICE_X10Y152_C5Q;
  wire [0:0] CLBLM_L_X8Y152_SLICE_X10Y152_C6;
  wire [0:0] CLBLM_L_X8Y152_SLICE_X10Y152_CLK;
  wire [0:0] CLBLM_L_X8Y152_SLICE_X10Y152_CMUX;
  wire [0:0] CLBLM_L_X8Y152_SLICE_X10Y152_CO5;
  wire [0:0] CLBLM_L_X8Y152_SLICE_X10Y152_CO6;
  wire [0:0] CLBLM_L_X8Y152_SLICE_X10Y152_CQ;
  wire [0:0] CLBLM_L_X8Y152_SLICE_X10Y152_C_CY;
  wire [0:0] CLBLM_L_X8Y152_SLICE_X10Y152_C_XOR;
  wire [0:0] CLBLM_L_X8Y152_SLICE_X10Y152_D;
  wire [0:0] CLBLM_L_X8Y152_SLICE_X10Y152_D1;
  wire [0:0] CLBLM_L_X8Y152_SLICE_X10Y152_D2;
  wire [0:0] CLBLM_L_X8Y152_SLICE_X10Y152_D3;
  wire [0:0] CLBLM_L_X8Y152_SLICE_X10Y152_D4;
  wire [0:0] CLBLM_L_X8Y152_SLICE_X10Y152_D5;
  wire [0:0] CLBLM_L_X8Y152_SLICE_X10Y152_D6;
  wire [0:0] CLBLM_L_X8Y152_SLICE_X10Y152_DO5;
  wire [0:0] CLBLM_L_X8Y152_SLICE_X10Y152_DO6;
  wire [0:0] CLBLM_L_X8Y152_SLICE_X10Y152_DQ;
  wire [0:0] CLBLM_L_X8Y152_SLICE_X10Y152_D_CY;
  wire [0:0] CLBLM_L_X8Y152_SLICE_X10Y152_D_XOR;
  wire [0:0] CLBLM_L_X8Y152_SLICE_X11Y152_A;
  wire [0:0] CLBLM_L_X8Y152_SLICE_X11Y152_A1;
  wire [0:0] CLBLM_L_X8Y152_SLICE_X11Y152_A2;
  wire [0:0] CLBLM_L_X8Y152_SLICE_X11Y152_A3;
  wire [0:0] CLBLM_L_X8Y152_SLICE_X11Y152_A4;
  wire [0:0] CLBLM_L_X8Y152_SLICE_X11Y152_A5;
  wire [0:0] CLBLM_L_X8Y152_SLICE_X11Y152_A6;
  wire [0:0] CLBLM_L_X8Y152_SLICE_X11Y152_AO5;
  wire [0:0] CLBLM_L_X8Y152_SLICE_X11Y152_AO6;
  wire [0:0] CLBLM_L_X8Y152_SLICE_X11Y152_AQ;
  wire [0:0] CLBLM_L_X8Y152_SLICE_X11Y152_A_CY;
  wire [0:0] CLBLM_L_X8Y152_SLICE_X11Y152_A_XOR;
  wire [0:0] CLBLM_L_X8Y152_SLICE_X11Y152_B;
  wire [0:0] CLBLM_L_X8Y152_SLICE_X11Y152_B1;
  wire [0:0] CLBLM_L_X8Y152_SLICE_X11Y152_B2;
  wire [0:0] CLBLM_L_X8Y152_SLICE_X11Y152_B3;
  wire [0:0] CLBLM_L_X8Y152_SLICE_X11Y152_B4;
  wire [0:0] CLBLM_L_X8Y152_SLICE_X11Y152_B5;
  wire [0:0] CLBLM_L_X8Y152_SLICE_X11Y152_B6;
  wire [0:0] CLBLM_L_X8Y152_SLICE_X11Y152_BO5;
  wire [0:0] CLBLM_L_X8Y152_SLICE_X11Y152_BO6;
  wire [0:0] CLBLM_L_X8Y152_SLICE_X11Y152_BQ;
  wire [0:0] CLBLM_L_X8Y152_SLICE_X11Y152_B_CY;
  wire [0:0] CLBLM_L_X8Y152_SLICE_X11Y152_B_XOR;
  wire [0:0] CLBLM_L_X8Y152_SLICE_X11Y152_C;
  wire [0:0] CLBLM_L_X8Y152_SLICE_X11Y152_C1;
  wire [0:0] CLBLM_L_X8Y152_SLICE_X11Y152_C2;
  wire [0:0] CLBLM_L_X8Y152_SLICE_X11Y152_C3;
  wire [0:0] CLBLM_L_X8Y152_SLICE_X11Y152_C4;
  wire [0:0] CLBLM_L_X8Y152_SLICE_X11Y152_C5;
  wire [0:0] CLBLM_L_X8Y152_SLICE_X11Y152_C6;
  wire [0:0] CLBLM_L_X8Y152_SLICE_X11Y152_CLK;
  wire [0:0] CLBLM_L_X8Y152_SLICE_X11Y152_CO5;
  wire [0:0] CLBLM_L_X8Y152_SLICE_X11Y152_CO6;
  wire [0:0] CLBLM_L_X8Y152_SLICE_X11Y152_CQ;
  wire [0:0] CLBLM_L_X8Y152_SLICE_X11Y152_C_CY;
  wire [0:0] CLBLM_L_X8Y152_SLICE_X11Y152_C_XOR;
  wire [0:0] CLBLM_L_X8Y152_SLICE_X11Y152_D;
  wire [0:0] CLBLM_L_X8Y152_SLICE_X11Y152_D1;
  wire [0:0] CLBLM_L_X8Y152_SLICE_X11Y152_D2;
  wire [0:0] CLBLM_L_X8Y152_SLICE_X11Y152_D3;
  wire [0:0] CLBLM_L_X8Y152_SLICE_X11Y152_D4;
  wire [0:0] CLBLM_L_X8Y152_SLICE_X11Y152_D5;
  wire [0:0] CLBLM_L_X8Y152_SLICE_X11Y152_D5Q;
  wire [0:0] CLBLM_L_X8Y152_SLICE_X11Y152_D6;
  wire [0:0] CLBLM_L_X8Y152_SLICE_X11Y152_DMUX;
  wire [0:0] CLBLM_L_X8Y152_SLICE_X11Y152_DO5;
  wire [0:0] CLBLM_L_X8Y152_SLICE_X11Y152_DO6;
  wire [0:0] CLBLM_L_X8Y152_SLICE_X11Y152_DQ;
  wire [0:0] CLBLM_L_X8Y152_SLICE_X11Y152_D_CY;
  wire [0:0] CLBLM_L_X8Y152_SLICE_X11Y152_D_XOR;
  wire [0:0] CLBLM_L_X8Y153_SLICE_X10Y153_A;
  wire [0:0] CLBLM_L_X8Y153_SLICE_X10Y153_A1;
  wire [0:0] CLBLM_L_X8Y153_SLICE_X10Y153_A2;
  wire [0:0] CLBLM_L_X8Y153_SLICE_X10Y153_A3;
  wire [0:0] CLBLM_L_X8Y153_SLICE_X10Y153_A4;
  wire [0:0] CLBLM_L_X8Y153_SLICE_X10Y153_A5;
  wire [0:0] CLBLM_L_X8Y153_SLICE_X10Y153_A5Q;
  wire [0:0] CLBLM_L_X8Y153_SLICE_X10Y153_A6;
  wire [0:0] CLBLM_L_X8Y153_SLICE_X10Y153_AMUX;
  wire [0:0] CLBLM_L_X8Y153_SLICE_X10Y153_AO5;
  wire [0:0] CLBLM_L_X8Y153_SLICE_X10Y153_AO6;
  wire [0:0] CLBLM_L_X8Y153_SLICE_X10Y153_AQ;
  wire [0:0] CLBLM_L_X8Y153_SLICE_X10Y153_A_CY;
  wire [0:0] CLBLM_L_X8Y153_SLICE_X10Y153_A_XOR;
  wire [0:0] CLBLM_L_X8Y153_SLICE_X10Y153_B;
  wire [0:0] CLBLM_L_X8Y153_SLICE_X10Y153_B1;
  wire [0:0] CLBLM_L_X8Y153_SLICE_X10Y153_B2;
  wire [0:0] CLBLM_L_X8Y153_SLICE_X10Y153_B3;
  wire [0:0] CLBLM_L_X8Y153_SLICE_X10Y153_B4;
  wire [0:0] CLBLM_L_X8Y153_SLICE_X10Y153_B5;
  wire [0:0] CLBLM_L_X8Y153_SLICE_X10Y153_B5Q;
  wire [0:0] CLBLM_L_X8Y153_SLICE_X10Y153_B6;
  wire [0:0] CLBLM_L_X8Y153_SLICE_X10Y153_BMUX;
  wire [0:0] CLBLM_L_X8Y153_SLICE_X10Y153_BO5;
  wire [0:0] CLBLM_L_X8Y153_SLICE_X10Y153_BO6;
  wire [0:0] CLBLM_L_X8Y153_SLICE_X10Y153_BQ;
  wire [0:0] CLBLM_L_X8Y153_SLICE_X10Y153_B_CY;
  wire [0:0] CLBLM_L_X8Y153_SLICE_X10Y153_B_XOR;
  wire [0:0] CLBLM_L_X8Y153_SLICE_X10Y153_C;
  wire [0:0] CLBLM_L_X8Y153_SLICE_X10Y153_C1;
  wire [0:0] CLBLM_L_X8Y153_SLICE_X10Y153_C2;
  wire [0:0] CLBLM_L_X8Y153_SLICE_X10Y153_C3;
  wire [0:0] CLBLM_L_X8Y153_SLICE_X10Y153_C4;
  wire [0:0] CLBLM_L_X8Y153_SLICE_X10Y153_C5;
  wire [0:0] CLBLM_L_X8Y153_SLICE_X10Y153_C5Q;
  wire [0:0] CLBLM_L_X8Y153_SLICE_X10Y153_C6;
  wire [0:0] CLBLM_L_X8Y153_SLICE_X10Y153_CLK;
  wire [0:0] CLBLM_L_X8Y153_SLICE_X10Y153_CMUX;
  wire [0:0] CLBLM_L_X8Y153_SLICE_X10Y153_CO5;
  wire [0:0] CLBLM_L_X8Y153_SLICE_X10Y153_CO6;
  wire [0:0] CLBLM_L_X8Y153_SLICE_X10Y153_CQ;
  wire [0:0] CLBLM_L_X8Y153_SLICE_X10Y153_C_CY;
  wire [0:0] CLBLM_L_X8Y153_SLICE_X10Y153_C_XOR;
  wire [0:0] CLBLM_L_X8Y153_SLICE_X10Y153_D;
  wire [0:0] CLBLM_L_X8Y153_SLICE_X10Y153_D1;
  wire [0:0] CLBLM_L_X8Y153_SLICE_X10Y153_D2;
  wire [0:0] CLBLM_L_X8Y153_SLICE_X10Y153_D3;
  wire [0:0] CLBLM_L_X8Y153_SLICE_X10Y153_D4;
  wire [0:0] CLBLM_L_X8Y153_SLICE_X10Y153_D5;
  wire [0:0] CLBLM_L_X8Y153_SLICE_X10Y153_D5Q;
  wire [0:0] CLBLM_L_X8Y153_SLICE_X10Y153_D6;
  wire [0:0] CLBLM_L_X8Y153_SLICE_X10Y153_DMUX;
  wire [0:0] CLBLM_L_X8Y153_SLICE_X10Y153_DO5;
  wire [0:0] CLBLM_L_X8Y153_SLICE_X10Y153_DO6;
  wire [0:0] CLBLM_L_X8Y153_SLICE_X10Y153_DQ;
  wire [0:0] CLBLM_L_X8Y153_SLICE_X10Y153_D_CY;
  wire [0:0] CLBLM_L_X8Y153_SLICE_X10Y153_D_XOR;
  wire [0:0] CLBLM_L_X8Y153_SLICE_X11Y153_A;
  wire [0:0] CLBLM_L_X8Y153_SLICE_X11Y153_A1;
  wire [0:0] CLBLM_L_X8Y153_SLICE_X11Y153_A2;
  wire [0:0] CLBLM_L_X8Y153_SLICE_X11Y153_A3;
  wire [0:0] CLBLM_L_X8Y153_SLICE_X11Y153_A4;
  wire [0:0] CLBLM_L_X8Y153_SLICE_X11Y153_A5;
  wire [0:0] CLBLM_L_X8Y153_SLICE_X11Y153_A6;
  wire [0:0] CLBLM_L_X8Y153_SLICE_X11Y153_AO5;
  wire [0:0] CLBLM_L_X8Y153_SLICE_X11Y153_AO6;
  wire [0:0] CLBLM_L_X8Y153_SLICE_X11Y153_AQ;
  wire [0:0] CLBLM_L_X8Y153_SLICE_X11Y153_A_CY;
  wire [0:0] CLBLM_L_X8Y153_SLICE_X11Y153_A_XOR;
  wire [0:0] CLBLM_L_X8Y153_SLICE_X11Y153_B;
  wire [0:0] CLBLM_L_X8Y153_SLICE_X11Y153_B1;
  wire [0:0] CLBLM_L_X8Y153_SLICE_X11Y153_B2;
  wire [0:0] CLBLM_L_X8Y153_SLICE_X11Y153_B3;
  wire [0:0] CLBLM_L_X8Y153_SLICE_X11Y153_B4;
  wire [0:0] CLBLM_L_X8Y153_SLICE_X11Y153_B5;
  wire [0:0] CLBLM_L_X8Y153_SLICE_X11Y153_B6;
  wire [0:0] CLBLM_L_X8Y153_SLICE_X11Y153_BO5;
  wire [0:0] CLBLM_L_X8Y153_SLICE_X11Y153_BO6;
  wire [0:0] CLBLM_L_X8Y153_SLICE_X11Y153_BQ;
  wire [0:0] CLBLM_L_X8Y153_SLICE_X11Y153_B_CY;
  wire [0:0] CLBLM_L_X8Y153_SLICE_X11Y153_B_XOR;
  wire [0:0] CLBLM_L_X8Y153_SLICE_X11Y153_C;
  wire [0:0] CLBLM_L_X8Y153_SLICE_X11Y153_C1;
  wire [0:0] CLBLM_L_X8Y153_SLICE_X11Y153_C2;
  wire [0:0] CLBLM_L_X8Y153_SLICE_X11Y153_C3;
  wire [0:0] CLBLM_L_X8Y153_SLICE_X11Y153_C4;
  wire [0:0] CLBLM_L_X8Y153_SLICE_X11Y153_C5;
  wire [0:0] CLBLM_L_X8Y153_SLICE_X11Y153_C6;
  wire [0:0] CLBLM_L_X8Y153_SLICE_X11Y153_CLK;
  wire [0:0] CLBLM_L_X8Y153_SLICE_X11Y153_CO5;
  wire [0:0] CLBLM_L_X8Y153_SLICE_X11Y153_CO6;
  wire [0:0] CLBLM_L_X8Y153_SLICE_X11Y153_C_CY;
  wire [0:0] CLBLM_L_X8Y153_SLICE_X11Y153_C_XOR;
  wire [0:0] CLBLM_L_X8Y153_SLICE_X11Y153_D;
  wire [0:0] CLBLM_L_X8Y153_SLICE_X11Y153_D1;
  wire [0:0] CLBLM_L_X8Y153_SLICE_X11Y153_D2;
  wire [0:0] CLBLM_L_X8Y153_SLICE_X11Y153_D3;
  wire [0:0] CLBLM_L_X8Y153_SLICE_X11Y153_D4;
  wire [0:0] CLBLM_L_X8Y153_SLICE_X11Y153_D5;
  wire [0:0] CLBLM_L_X8Y153_SLICE_X11Y153_D6;
  wire [0:0] CLBLM_L_X8Y153_SLICE_X11Y153_DO5;
  wire [0:0] CLBLM_L_X8Y153_SLICE_X11Y153_DO6;
  wire [0:0] CLBLM_L_X8Y153_SLICE_X11Y153_D_CY;
  wire [0:0] CLBLM_L_X8Y153_SLICE_X11Y153_D_XOR;
  wire [0:0] CLBLM_L_X8Y154_SLICE_X10Y154_A;
  wire [0:0] CLBLM_L_X8Y154_SLICE_X10Y154_A1;
  wire [0:0] CLBLM_L_X8Y154_SLICE_X10Y154_A2;
  wire [0:0] CLBLM_L_X8Y154_SLICE_X10Y154_A3;
  wire [0:0] CLBLM_L_X8Y154_SLICE_X10Y154_A4;
  wire [0:0] CLBLM_L_X8Y154_SLICE_X10Y154_A5;
  wire [0:0] CLBLM_L_X8Y154_SLICE_X10Y154_A6;
  wire [0:0] CLBLM_L_X8Y154_SLICE_X10Y154_AO5;
  wire [0:0] CLBLM_L_X8Y154_SLICE_X10Y154_AO6;
  wire [0:0] CLBLM_L_X8Y154_SLICE_X10Y154_AQ;
  wire [0:0] CLBLM_L_X8Y154_SLICE_X10Y154_A_CY;
  wire [0:0] CLBLM_L_X8Y154_SLICE_X10Y154_A_XOR;
  wire [0:0] CLBLM_L_X8Y154_SLICE_X10Y154_B;
  wire [0:0] CLBLM_L_X8Y154_SLICE_X10Y154_B1;
  wire [0:0] CLBLM_L_X8Y154_SLICE_X10Y154_B2;
  wire [0:0] CLBLM_L_X8Y154_SLICE_X10Y154_B3;
  wire [0:0] CLBLM_L_X8Y154_SLICE_X10Y154_B4;
  wire [0:0] CLBLM_L_X8Y154_SLICE_X10Y154_B5;
  wire [0:0] CLBLM_L_X8Y154_SLICE_X10Y154_B6;
  wire [0:0] CLBLM_L_X8Y154_SLICE_X10Y154_BMUX;
  wire [0:0] CLBLM_L_X8Y154_SLICE_X10Y154_BO5;
  wire [0:0] CLBLM_L_X8Y154_SLICE_X10Y154_BO6;
  wire [0:0] CLBLM_L_X8Y154_SLICE_X10Y154_B_CY;
  wire [0:0] CLBLM_L_X8Y154_SLICE_X10Y154_B_XOR;
  wire [0:0] CLBLM_L_X8Y154_SLICE_X10Y154_C;
  wire [0:0] CLBLM_L_X8Y154_SLICE_X10Y154_C1;
  wire [0:0] CLBLM_L_X8Y154_SLICE_X10Y154_C2;
  wire [0:0] CLBLM_L_X8Y154_SLICE_X10Y154_C3;
  wire [0:0] CLBLM_L_X8Y154_SLICE_X10Y154_C4;
  wire [0:0] CLBLM_L_X8Y154_SLICE_X10Y154_C5;
  wire [0:0] CLBLM_L_X8Y154_SLICE_X10Y154_C6;
  wire [0:0] CLBLM_L_X8Y154_SLICE_X10Y154_CLK;
  wire [0:0] CLBLM_L_X8Y154_SLICE_X10Y154_CO5;
  wire [0:0] CLBLM_L_X8Y154_SLICE_X10Y154_CO6;
  wire [0:0] CLBLM_L_X8Y154_SLICE_X10Y154_C_CY;
  wire [0:0] CLBLM_L_X8Y154_SLICE_X10Y154_C_XOR;
  wire [0:0] CLBLM_L_X8Y154_SLICE_X10Y154_D;
  wire [0:0] CLBLM_L_X8Y154_SLICE_X10Y154_D1;
  wire [0:0] CLBLM_L_X8Y154_SLICE_X10Y154_D2;
  wire [0:0] CLBLM_L_X8Y154_SLICE_X10Y154_D3;
  wire [0:0] CLBLM_L_X8Y154_SLICE_X10Y154_D4;
  wire [0:0] CLBLM_L_X8Y154_SLICE_X10Y154_D5;
  wire [0:0] CLBLM_L_X8Y154_SLICE_X10Y154_D6;
  wire [0:0] CLBLM_L_X8Y154_SLICE_X10Y154_DO5;
  wire [0:0] CLBLM_L_X8Y154_SLICE_X10Y154_DO6;
  wire [0:0] CLBLM_L_X8Y154_SLICE_X10Y154_D_CY;
  wire [0:0] CLBLM_L_X8Y154_SLICE_X10Y154_D_XOR;
  wire [0:0] CLBLM_L_X8Y154_SLICE_X11Y154_A;
  wire [0:0] CLBLM_L_X8Y154_SLICE_X11Y154_A1;
  wire [0:0] CLBLM_L_X8Y154_SLICE_X11Y154_A2;
  wire [0:0] CLBLM_L_X8Y154_SLICE_X11Y154_A3;
  wire [0:0] CLBLM_L_X8Y154_SLICE_X11Y154_A4;
  wire [0:0] CLBLM_L_X8Y154_SLICE_X11Y154_A5;
  wire [0:0] CLBLM_L_X8Y154_SLICE_X11Y154_A6;
  wire [0:0] CLBLM_L_X8Y154_SLICE_X11Y154_AO5;
  wire [0:0] CLBLM_L_X8Y154_SLICE_X11Y154_AO6;
  wire [0:0] CLBLM_L_X8Y154_SLICE_X11Y154_AQ;
  wire [0:0] CLBLM_L_X8Y154_SLICE_X11Y154_A_CY;
  wire [0:0] CLBLM_L_X8Y154_SLICE_X11Y154_A_XOR;
  wire [0:0] CLBLM_L_X8Y154_SLICE_X11Y154_B;
  wire [0:0] CLBLM_L_X8Y154_SLICE_X11Y154_B1;
  wire [0:0] CLBLM_L_X8Y154_SLICE_X11Y154_B2;
  wire [0:0] CLBLM_L_X8Y154_SLICE_X11Y154_B3;
  wire [0:0] CLBLM_L_X8Y154_SLICE_X11Y154_B4;
  wire [0:0] CLBLM_L_X8Y154_SLICE_X11Y154_B5;
  wire [0:0] CLBLM_L_X8Y154_SLICE_X11Y154_B6;
  wire [0:0] CLBLM_L_X8Y154_SLICE_X11Y154_BO5;
  wire [0:0] CLBLM_L_X8Y154_SLICE_X11Y154_BO6;
  wire [0:0] CLBLM_L_X8Y154_SLICE_X11Y154_B_CY;
  wire [0:0] CLBLM_L_X8Y154_SLICE_X11Y154_B_XOR;
  wire [0:0] CLBLM_L_X8Y154_SLICE_X11Y154_C;
  wire [0:0] CLBLM_L_X8Y154_SLICE_X11Y154_C1;
  wire [0:0] CLBLM_L_X8Y154_SLICE_X11Y154_C2;
  wire [0:0] CLBLM_L_X8Y154_SLICE_X11Y154_C3;
  wire [0:0] CLBLM_L_X8Y154_SLICE_X11Y154_C4;
  wire [0:0] CLBLM_L_X8Y154_SLICE_X11Y154_C5;
  wire [0:0] CLBLM_L_X8Y154_SLICE_X11Y154_C6;
  wire [0:0] CLBLM_L_X8Y154_SLICE_X11Y154_CLK;
  wire [0:0] CLBLM_L_X8Y154_SLICE_X11Y154_CO5;
  wire [0:0] CLBLM_L_X8Y154_SLICE_X11Y154_CO6;
  wire [0:0] CLBLM_L_X8Y154_SLICE_X11Y154_C_CY;
  wire [0:0] CLBLM_L_X8Y154_SLICE_X11Y154_C_XOR;
  wire [0:0] CLBLM_L_X8Y154_SLICE_X11Y154_D;
  wire [0:0] CLBLM_L_X8Y154_SLICE_X11Y154_D1;
  wire [0:0] CLBLM_L_X8Y154_SLICE_X11Y154_D2;
  wire [0:0] CLBLM_L_X8Y154_SLICE_X11Y154_D3;
  wire [0:0] CLBLM_L_X8Y154_SLICE_X11Y154_D4;
  wire [0:0] CLBLM_L_X8Y154_SLICE_X11Y154_D5;
  wire [0:0] CLBLM_L_X8Y154_SLICE_X11Y154_D6;
  wire [0:0] CLBLM_L_X8Y154_SLICE_X11Y154_DO5;
  wire [0:0] CLBLM_L_X8Y154_SLICE_X11Y154_DO6;
  wire [0:0] CLBLM_L_X8Y154_SLICE_X11Y154_D_CY;
  wire [0:0] CLBLM_L_X8Y154_SLICE_X11Y154_D_XOR;
  wire [0:0] CLBLM_R_X103Y178_SLICE_X162Y178_A;
  wire [0:0] CLBLM_R_X103Y178_SLICE_X162Y178_A1;
  wire [0:0] CLBLM_R_X103Y178_SLICE_X162Y178_A2;
  wire [0:0] CLBLM_R_X103Y178_SLICE_X162Y178_A3;
  wire [0:0] CLBLM_R_X103Y178_SLICE_X162Y178_A4;
  wire [0:0] CLBLM_R_X103Y178_SLICE_X162Y178_A5;
  wire [0:0] CLBLM_R_X103Y178_SLICE_X162Y178_A6;
  wire [0:0] CLBLM_R_X103Y178_SLICE_X162Y178_AO5;
  wire [0:0] CLBLM_R_X103Y178_SLICE_X162Y178_AO6;
  wire [0:0] CLBLM_R_X103Y178_SLICE_X162Y178_A_CY;
  wire [0:0] CLBLM_R_X103Y178_SLICE_X162Y178_A_XOR;
  wire [0:0] CLBLM_R_X103Y178_SLICE_X162Y178_B;
  wire [0:0] CLBLM_R_X103Y178_SLICE_X162Y178_B1;
  wire [0:0] CLBLM_R_X103Y178_SLICE_X162Y178_B2;
  wire [0:0] CLBLM_R_X103Y178_SLICE_X162Y178_B3;
  wire [0:0] CLBLM_R_X103Y178_SLICE_X162Y178_B4;
  wire [0:0] CLBLM_R_X103Y178_SLICE_X162Y178_B5;
  wire [0:0] CLBLM_R_X103Y178_SLICE_X162Y178_B6;
  wire [0:0] CLBLM_R_X103Y178_SLICE_X162Y178_BO5;
  wire [0:0] CLBLM_R_X103Y178_SLICE_X162Y178_BO6;
  wire [0:0] CLBLM_R_X103Y178_SLICE_X162Y178_B_CY;
  wire [0:0] CLBLM_R_X103Y178_SLICE_X162Y178_B_XOR;
  wire [0:0] CLBLM_R_X103Y178_SLICE_X162Y178_C;
  wire [0:0] CLBLM_R_X103Y178_SLICE_X162Y178_C1;
  wire [0:0] CLBLM_R_X103Y178_SLICE_X162Y178_C2;
  wire [0:0] CLBLM_R_X103Y178_SLICE_X162Y178_C3;
  wire [0:0] CLBLM_R_X103Y178_SLICE_X162Y178_C4;
  wire [0:0] CLBLM_R_X103Y178_SLICE_X162Y178_C5;
  wire [0:0] CLBLM_R_X103Y178_SLICE_X162Y178_C6;
  wire [0:0] CLBLM_R_X103Y178_SLICE_X162Y178_CO5;
  wire [0:0] CLBLM_R_X103Y178_SLICE_X162Y178_CO6;
  wire [0:0] CLBLM_R_X103Y178_SLICE_X162Y178_C_CY;
  wire [0:0] CLBLM_R_X103Y178_SLICE_X162Y178_C_XOR;
  wire [0:0] CLBLM_R_X103Y178_SLICE_X162Y178_D;
  wire [0:0] CLBLM_R_X103Y178_SLICE_X162Y178_D1;
  wire [0:0] CLBLM_R_X103Y178_SLICE_X162Y178_D2;
  wire [0:0] CLBLM_R_X103Y178_SLICE_X162Y178_D3;
  wire [0:0] CLBLM_R_X103Y178_SLICE_X162Y178_D4;
  wire [0:0] CLBLM_R_X103Y178_SLICE_X162Y178_D5;
  wire [0:0] CLBLM_R_X103Y178_SLICE_X162Y178_D6;
  wire [0:0] CLBLM_R_X103Y178_SLICE_X162Y178_DO5;
  wire [0:0] CLBLM_R_X103Y178_SLICE_X162Y178_DO6;
  wire [0:0] CLBLM_R_X103Y178_SLICE_X162Y178_D_CY;
  wire [0:0] CLBLM_R_X103Y178_SLICE_X162Y178_D_XOR;
  wire [0:0] CLBLM_R_X103Y178_SLICE_X163Y178_A;
  wire [0:0] CLBLM_R_X103Y178_SLICE_X163Y178_A1;
  wire [0:0] CLBLM_R_X103Y178_SLICE_X163Y178_A2;
  wire [0:0] CLBLM_R_X103Y178_SLICE_X163Y178_A3;
  wire [0:0] CLBLM_R_X103Y178_SLICE_X163Y178_A4;
  wire [0:0] CLBLM_R_X103Y178_SLICE_X163Y178_A5;
  wire [0:0] CLBLM_R_X103Y178_SLICE_X163Y178_A6;
  wire [0:0] CLBLM_R_X103Y178_SLICE_X163Y178_AO5;
  wire [0:0] CLBLM_R_X103Y178_SLICE_X163Y178_AO6;
  wire [0:0] CLBLM_R_X103Y178_SLICE_X163Y178_A_CY;
  wire [0:0] CLBLM_R_X103Y178_SLICE_X163Y178_A_XOR;
  wire [0:0] CLBLM_R_X103Y178_SLICE_X163Y178_B;
  wire [0:0] CLBLM_R_X103Y178_SLICE_X163Y178_B1;
  wire [0:0] CLBLM_R_X103Y178_SLICE_X163Y178_B2;
  wire [0:0] CLBLM_R_X103Y178_SLICE_X163Y178_B3;
  wire [0:0] CLBLM_R_X103Y178_SLICE_X163Y178_B4;
  wire [0:0] CLBLM_R_X103Y178_SLICE_X163Y178_B5;
  wire [0:0] CLBLM_R_X103Y178_SLICE_X163Y178_B6;
  wire [0:0] CLBLM_R_X103Y178_SLICE_X163Y178_BO5;
  wire [0:0] CLBLM_R_X103Y178_SLICE_X163Y178_BO6;
  wire [0:0] CLBLM_R_X103Y178_SLICE_X163Y178_B_CY;
  wire [0:0] CLBLM_R_X103Y178_SLICE_X163Y178_B_XOR;
  wire [0:0] CLBLM_R_X103Y178_SLICE_X163Y178_C;
  wire [0:0] CLBLM_R_X103Y178_SLICE_X163Y178_C1;
  wire [0:0] CLBLM_R_X103Y178_SLICE_X163Y178_C2;
  wire [0:0] CLBLM_R_X103Y178_SLICE_X163Y178_C3;
  wire [0:0] CLBLM_R_X103Y178_SLICE_X163Y178_C4;
  wire [0:0] CLBLM_R_X103Y178_SLICE_X163Y178_C5;
  wire [0:0] CLBLM_R_X103Y178_SLICE_X163Y178_C6;
  wire [0:0] CLBLM_R_X103Y178_SLICE_X163Y178_CO5;
  wire [0:0] CLBLM_R_X103Y178_SLICE_X163Y178_CO6;
  wire [0:0] CLBLM_R_X103Y178_SLICE_X163Y178_C_CY;
  wire [0:0] CLBLM_R_X103Y178_SLICE_X163Y178_C_XOR;
  wire [0:0] CLBLM_R_X103Y178_SLICE_X163Y178_D;
  wire [0:0] CLBLM_R_X103Y178_SLICE_X163Y178_D1;
  wire [0:0] CLBLM_R_X103Y178_SLICE_X163Y178_D2;
  wire [0:0] CLBLM_R_X103Y178_SLICE_X163Y178_D3;
  wire [0:0] CLBLM_R_X103Y178_SLICE_X163Y178_D4;
  wire [0:0] CLBLM_R_X103Y178_SLICE_X163Y178_D5;
  wire [0:0] CLBLM_R_X103Y178_SLICE_X163Y178_D6;
  wire [0:0] CLBLM_R_X103Y178_SLICE_X163Y178_DO5;
  wire [0:0] CLBLM_R_X103Y178_SLICE_X163Y178_DO6;
  wire [0:0] CLBLM_R_X103Y178_SLICE_X163Y178_D_CY;
  wire [0:0] CLBLM_R_X103Y178_SLICE_X163Y178_D_XOR;
  wire [0:0] CLBLM_R_X11Y144_SLICE_X14Y144_A;
  wire [0:0] CLBLM_R_X11Y144_SLICE_X14Y144_A1;
  wire [0:0] CLBLM_R_X11Y144_SLICE_X14Y144_A2;
  wire [0:0] CLBLM_R_X11Y144_SLICE_X14Y144_A3;
  wire [0:0] CLBLM_R_X11Y144_SLICE_X14Y144_A4;
  wire [0:0] CLBLM_R_X11Y144_SLICE_X14Y144_A5;
  wire [0:0] CLBLM_R_X11Y144_SLICE_X14Y144_A6;
  wire [0:0] CLBLM_R_X11Y144_SLICE_X14Y144_AO5;
  wire [0:0] CLBLM_R_X11Y144_SLICE_X14Y144_AO6;
  wire [0:0] CLBLM_R_X11Y144_SLICE_X14Y144_A_CY;
  wire [0:0] CLBLM_R_X11Y144_SLICE_X14Y144_A_XOR;
  wire [0:0] CLBLM_R_X11Y144_SLICE_X14Y144_B;
  wire [0:0] CLBLM_R_X11Y144_SLICE_X14Y144_B1;
  wire [0:0] CLBLM_R_X11Y144_SLICE_X14Y144_B2;
  wire [0:0] CLBLM_R_X11Y144_SLICE_X14Y144_B3;
  wire [0:0] CLBLM_R_X11Y144_SLICE_X14Y144_B4;
  wire [0:0] CLBLM_R_X11Y144_SLICE_X14Y144_B5;
  wire [0:0] CLBLM_R_X11Y144_SLICE_X14Y144_B6;
  wire [0:0] CLBLM_R_X11Y144_SLICE_X14Y144_BO5;
  wire [0:0] CLBLM_R_X11Y144_SLICE_X14Y144_BO6;
  wire [0:0] CLBLM_R_X11Y144_SLICE_X14Y144_B_CY;
  wire [0:0] CLBLM_R_X11Y144_SLICE_X14Y144_B_XOR;
  wire [0:0] CLBLM_R_X11Y144_SLICE_X14Y144_C;
  wire [0:0] CLBLM_R_X11Y144_SLICE_X14Y144_C1;
  wire [0:0] CLBLM_R_X11Y144_SLICE_X14Y144_C2;
  wire [0:0] CLBLM_R_X11Y144_SLICE_X14Y144_C3;
  wire [0:0] CLBLM_R_X11Y144_SLICE_X14Y144_C4;
  wire [0:0] CLBLM_R_X11Y144_SLICE_X14Y144_C5;
  wire [0:0] CLBLM_R_X11Y144_SLICE_X14Y144_C6;
  wire [0:0] CLBLM_R_X11Y144_SLICE_X14Y144_CO5;
  wire [0:0] CLBLM_R_X11Y144_SLICE_X14Y144_CO6;
  wire [0:0] CLBLM_R_X11Y144_SLICE_X14Y144_C_CY;
  wire [0:0] CLBLM_R_X11Y144_SLICE_X14Y144_C_XOR;
  wire [0:0] CLBLM_R_X11Y144_SLICE_X14Y144_D;
  wire [0:0] CLBLM_R_X11Y144_SLICE_X14Y144_D1;
  wire [0:0] CLBLM_R_X11Y144_SLICE_X14Y144_D2;
  wire [0:0] CLBLM_R_X11Y144_SLICE_X14Y144_D3;
  wire [0:0] CLBLM_R_X11Y144_SLICE_X14Y144_D4;
  wire [0:0] CLBLM_R_X11Y144_SLICE_X14Y144_D5;
  wire [0:0] CLBLM_R_X11Y144_SLICE_X14Y144_D6;
  wire [0:0] CLBLM_R_X11Y144_SLICE_X14Y144_DO5;
  wire [0:0] CLBLM_R_X11Y144_SLICE_X14Y144_DO6;
  wire [0:0] CLBLM_R_X11Y144_SLICE_X14Y144_D_CY;
  wire [0:0] CLBLM_R_X11Y144_SLICE_X14Y144_D_XOR;
  wire [0:0] CLBLM_R_X11Y144_SLICE_X15Y144_A;
  wire [0:0] CLBLM_R_X11Y144_SLICE_X15Y144_A1;
  wire [0:0] CLBLM_R_X11Y144_SLICE_X15Y144_A2;
  wire [0:0] CLBLM_R_X11Y144_SLICE_X15Y144_A3;
  wire [0:0] CLBLM_R_X11Y144_SLICE_X15Y144_A4;
  wire [0:0] CLBLM_R_X11Y144_SLICE_X15Y144_A5;
  wire [0:0] CLBLM_R_X11Y144_SLICE_X15Y144_A6;
  wire [0:0] CLBLM_R_X11Y144_SLICE_X15Y144_AO5;
  wire [0:0] CLBLM_R_X11Y144_SLICE_X15Y144_AO6;
  wire [0:0] CLBLM_R_X11Y144_SLICE_X15Y144_A_CY;
  wire [0:0] CLBLM_R_X11Y144_SLICE_X15Y144_A_XOR;
  wire [0:0] CLBLM_R_X11Y144_SLICE_X15Y144_B;
  wire [0:0] CLBLM_R_X11Y144_SLICE_X15Y144_B1;
  wire [0:0] CLBLM_R_X11Y144_SLICE_X15Y144_B2;
  wire [0:0] CLBLM_R_X11Y144_SLICE_X15Y144_B3;
  wire [0:0] CLBLM_R_X11Y144_SLICE_X15Y144_B4;
  wire [0:0] CLBLM_R_X11Y144_SLICE_X15Y144_B5;
  wire [0:0] CLBLM_R_X11Y144_SLICE_X15Y144_B6;
  wire [0:0] CLBLM_R_X11Y144_SLICE_X15Y144_BO5;
  wire [0:0] CLBLM_R_X11Y144_SLICE_X15Y144_BO6;
  wire [0:0] CLBLM_R_X11Y144_SLICE_X15Y144_B_CY;
  wire [0:0] CLBLM_R_X11Y144_SLICE_X15Y144_B_XOR;
  wire [0:0] CLBLM_R_X11Y144_SLICE_X15Y144_C;
  wire [0:0] CLBLM_R_X11Y144_SLICE_X15Y144_C1;
  wire [0:0] CLBLM_R_X11Y144_SLICE_X15Y144_C2;
  wire [0:0] CLBLM_R_X11Y144_SLICE_X15Y144_C3;
  wire [0:0] CLBLM_R_X11Y144_SLICE_X15Y144_C4;
  wire [0:0] CLBLM_R_X11Y144_SLICE_X15Y144_C5;
  wire [0:0] CLBLM_R_X11Y144_SLICE_X15Y144_C6;
  wire [0:0] CLBLM_R_X11Y144_SLICE_X15Y144_CO5;
  wire [0:0] CLBLM_R_X11Y144_SLICE_X15Y144_CO6;
  wire [0:0] CLBLM_R_X11Y144_SLICE_X15Y144_C_CY;
  wire [0:0] CLBLM_R_X11Y144_SLICE_X15Y144_C_XOR;
  wire [0:0] CLBLM_R_X11Y144_SLICE_X15Y144_D;
  wire [0:0] CLBLM_R_X11Y144_SLICE_X15Y144_D1;
  wire [0:0] CLBLM_R_X11Y144_SLICE_X15Y144_D2;
  wire [0:0] CLBLM_R_X11Y144_SLICE_X15Y144_D3;
  wire [0:0] CLBLM_R_X11Y144_SLICE_X15Y144_D4;
  wire [0:0] CLBLM_R_X11Y144_SLICE_X15Y144_D5;
  wire [0:0] CLBLM_R_X11Y144_SLICE_X15Y144_D6;
  wire [0:0] CLBLM_R_X11Y144_SLICE_X15Y144_DO5;
  wire [0:0] CLBLM_R_X11Y144_SLICE_X15Y144_DO6;
  wire [0:0] CLBLM_R_X11Y144_SLICE_X15Y144_D_CY;
  wire [0:0] CLBLM_R_X11Y144_SLICE_X15Y144_D_XOR;
  wire [0:0] CLBLM_R_X11Y145_SLICE_X14Y145_A;
  wire [0:0] CLBLM_R_X11Y145_SLICE_X14Y145_A1;
  wire [0:0] CLBLM_R_X11Y145_SLICE_X14Y145_A2;
  wire [0:0] CLBLM_R_X11Y145_SLICE_X14Y145_A3;
  wire [0:0] CLBLM_R_X11Y145_SLICE_X14Y145_A4;
  wire [0:0] CLBLM_R_X11Y145_SLICE_X14Y145_A5;
  wire [0:0] CLBLM_R_X11Y145_SLICE_X14Y145_A6;
  wire [0:0] CLBLM_R_X11Y145_SLICE_X14Y145_AO5;
  wire [0:0] CLBLM_R_X11Y145_SLICE_X14Y145_AO6;
  wire [0:0] CLBLM_R_X11Y145_SLICE_X14Y145_A_CY;
  wire [0:0] CLBLM_R_X11Y145_SLICE_X14Y145_A_XOR;
  wire [0:0] CLBLM_R_X11Y145_SLICE_X14Y145_B;
  wire [0:0] CLBLM_R_X11Y145_SLICE_X14Y145_B1;
  wire [0:0] CLBLM_R_X11Y145_SLICE_X14Y145_B2;
  wire [0:0] CLBLM_R_X11Y145_SLICE_X14Y145_B3;
  wire [0:0] CLBLM_R_X11Y145_SLICE_X14Y145_B4;
  wire [0:0] CLBLM_R_X11Y145_SLICE_X14Y145_B5;
  wire [0:0] CLBLM_R_X11Y145_SLICE_X14Y145_B6;
  wire [0:0] CLBLM_R_X11Y145_SLICE_X14Y145_BO5;
  wire [0:0] CLBLM_R_X11Y145_SLICE_X14Y145_BO6;
  wire [0:0] CLBLM_R_X11Y145_SLICE_X14Y145_B_CY;
  wire [0:0] CLBLM_R_X11Y145_SLICE_X14Y145_B_XOR;
  wire [0:0] CLBLM_R_X11Y145_SLICE_X14Y145_C;
  wire [0:0] CLBLM_R_X11Y145_SLICE_X14Y145_C1;
  wire [0:0] CLBLM_R_X11Y145_SLICE_X14Y145_C2;
  wire [0:0] CLBLM_R_X11Y145_SLICE_X14Y145_C3;
  wire [0:0] CLBLM_R_X11Y145_SLICE_X14Y145_C4;
  wire [0:0] CLBLM_R_X11Y145_SLICE_X14Y145_C5;
  wire [0:0] CLBLM_R_X11Y145_SLICE_X14Y145_C6;
  wire [0:0] CLBLM_R_X11Y145_SLICE_X14Y145_CO5;
  wire [0:0] CLBLM_R_X11Y145_SLICE_X14Y145_CO6;
  wire [0:0] CLBLM_R_X11Y145_SLICE_X14Y145_C_CY;
  wire [0:0] CLBLM_R_X11Y145_SLICE_X14Y145_C_XOR;
  wire [0:0] CLBLM_R_X11Y145_SLICE_X14Y145_D;
  wire [0:0] CLBLM_R_X11Y145_SLICE_X14Y145_D1;
  wire [0:0] CLBLM_R_X11Y145_SLICE_X14Y145_D2;
  wire [0:0] CLBLM_R_X11Y145_SLICE_X14Y145_D3;
  wire [0:0] CLBLM_R_X11Y145_SLICE_X14Y145_D4;
  wire [0:0] CLBLM_R_X11Y145_SLICE_X14Y145_D5;
  wire [0:0] CLBLM_R_X11Y145_SLICE_X14Y145_D6;
  wire [0:0] CLBLM_R_X11Y145_SLICE_X14Y145_DO5;
  wire [0:0] CLBLM_R_X11Y145_SLICE_X14Y145_DO6;
  wire [0:0] CLBLM_R_X11Y145_SLICE_X14Y145_D_CY;
  wire [0:0] CLBLM_R_X11Y145_SLICE_X14Y145_D_XOR;
  wire [0:0] CLBLM_R_X11Y145_SLICE_X15Y145_A;
  wire [0:0] CLBLM_R_X11Y145_SLICE_X15Y145_A1;
  wire [0:0] CLBLM_R_X11Y145_SLICE_X15Y145_A2;
  wire [0:0] CLBLM_R_X11Y145_SLICE_X15Y145_A3;
  wire [0:0] CLBLM_R_X11Y145_SLICE_X15Y145_A4;
  wire [0:0] CLBLM_R_X11Y145_SLICE_X15Y145_A5;
  wire [0:0] CLBLM_R_X11Y145_SLICE_X15Y145_A6;
  wire [0:0] CLBLM_R_X11Y145_SLICE_X15Y145_AO5;
  wire [0:0] CLBLM_R_X11Y145_SLICE_X15Y145_AO6;
  wire [0:0] CLBLM_R_X11Y145_SLICE_X15Y145_AQ;
  wire [0:0] CLBLM_R_X11Y145_SLICE_X15Y145_A_CY;
  wire [0:0] CLBLM_R_X11Y145_SLICE_X15Y145_A_XOR;
  wire [0:0] CLBLM_R_X11Y145_SLICE_X15Y145_B;
  wire [0:0] CLBLM_R_X11Y145_SLICE_X15Y145_B1;
  wire [0:0] CLBLM_R_X11Y145_SLICE_X15Y145_B2;
  wire [0:0] CLBLM_R_X11Y145_SLICE_X15Y145_B3;
  wire [0:0] CLBLM_R_X11Y145_SLICE_X15Y145_B4;
  wire [0:0] CLBLM_R_X11Y145_SLICE_X15Y145_B5;
  wire [0:0] CLBLM_R_X11Y145_SLICE_X15Y145_B6;
  wire [0:0] CLBLM_R_X11Y145_SLICE_X15Y145_BMUX;
  wire [0:0] CLBLM_R_X11Y145_SLICE_X15Y145_BO5;
  wire [0:0] CLBLM_R_X11Y145_SLICE_X15Y145_BO6;
  wire [0:0] CLBLM_R_X11Y145_SLICE_X15Y145_B_CY;
  wire [0:0] CLBLM_R_X11Y145_SLICE_X15Y145_B_XOR;
  wire [0:0] CLBLM_R_X11Y145_SLICE_X15Y145_C;
  wire [0:0] CLBLM_R_X11Y145_SLICE_X15Y145_C1;
  wire [0:0] CLBLM_R_X11Y145_SLICE_X15Y145_C2;
  wire [0:0] CLBLM_R_X11Y145_SLICE_X15Y145_C3;
  wire [0:0] CLBLM_R_X11Y145_SLICE_X15Y145_C4;
  wire [0:0] CLBLM_R_X11Y145_SLICE_X15Y145_C5;
  wire [0:0] CLBLM_R_X11Y145_SLICE_X15Y145_C6;
  wire [0:0] CLBLM_R_X11Y145_SLICE_X15Y145_CLK;
  wire [0:0] CLBLM_R_X11Y145_SLICE_X15Y145_CO5;
  wire [0:0] CLBLM_R_X11Y145_SLICE_X15Y145_CO6;
  wire [0:0] CLBLM_R_X11Y145_SLICE_X15Y145_C_CY;
  wire [0:0] CLBLM_R_X11Y145_SLICE_X15Y145_C_XOR;
  wire [0:0] CLBLM_R_X11Y145_SLICE_X15Y145_D;
  wire [0:0] CLBLM_R_X11Y145_SLICE_X15Y145_D1;
  wire [0:0] CLBLM_R_X11Y145_SLICE_X15Y145_D2;
  wire [0:0] CLBLM_R_X11Y145_SLICE_X15Y145_D3;
  wire [0:0] CLBLM_R_X11Y145_SLICE_X15Y145_D4;
  wire [0:0] CLBLM_R_X11Y145_SLICE_X15Y145_D5;
  wire [0:0] CLBLM_R_X11Y145_SLICE_X15Y145_D6;
  wire [0:0] CLBLM_R_X11Y145_SLICE_X15Y145_DO5;
  wire [0:0] CLBLM_R_X11Y145_SLICE_X15Y145_DO6;
  wire [0:0] CLBLM_R_X11Y145_SLICE_X15Y145_D_CY;
  wire [0:0] CLBLM_R_X11Y145_SLICE_X15Y145_D_XOR;
  wire [0:0] CLBLM_R_X11Y146_SLICE_X14Y146_A;
  wire [0:0] CLBLM_R_X11Y146_SLICE_X14Y146_A1;
  wire [0:0] CLBLM_R_X11Y146_SLICE_X14Y146_A2;
  wire [0:0] CLBLM_R_X11Y146_SLICE_X14Y146_A3;
  wire [0:0] CLBLM_R_X11Y146_SLICE_X14Y146_A4;
  wire [0:0] CLBLM_R_X11Y146_SLICE_X14Y146_A5;
  wire [0:0] CLBLM_R_X11Y146_SLICE_X14Y146_A6;
  wire [0:0] CLBLM_R_X11Y146_SLICE_X14Y146_AO5;
  wire [0:0] CLBLM_R_X11Y146_SLICE_X14Y146_AO6;
  wire [0:0] CLBLM_R_X11Y146_SLICE_X14Y146_AQ;
  wire [0:0] CLBLM_R_X11Y146_SLICE_X14Y146_A_CY;
  wire [0:0] CLBLM_R_X11Y146_SLICE_X14Y146_A_XOR;
  wire [0:0] CLBLM_R_X11Y146_SLICE_X14Y146_B;
  wire [0:0] CLBLM_R_X11Y146_SLICE_X14Y146_B1;
  wire [0:0] CLBLM_R_X11Y146_SLICE_X14Y146_B2;
  wire [0:0] CLBLM_R_X11Y146_SLICE_X14Y146_B3;
  wire [0:0] CLBLM_R_X11Y146_SLICE_X14Y146_B4;
  wire [0:0] CLBLM_R_X11Y146_SLICE_X14Y146_B5;
  wire [0:0] CLBLM_R_X11Y146_SLICE_X14Y146_B6;
  wire [0:0] CLBLM_R_X11Y146_SLICE_X14Y146_BMUX;
  wire [0:0] CLBLM_R_X11Y146_SLICE_X14Y146_BO5;
  wire [0:0] CLBLM_R_X11Y146_SLICE_X14Y146_BO6;
  wire [0:0] CLBLM_R_X11Y146_SLICE_X14Y146_B_CY;
  wire [0:0] CLBLM_R_X11Y146_SLICE_X14Y146_B_XOR;
  wire [0:0] CLBLM_R_X11Y146_SLICE_X14Y146_C;
  wire [0:0] CLBLM_R_X11Y146_SLICE_X14Y146_C1;
  wire [0:0] CLBLM_R_X11Y146_SLICE_X14Y146_C2;
  wire [0:0] CLBLM_R_X11Y146_SLICE_X14Y146_C3;
  wire [0:0] CLBLM_R_X11Y146_SLICE_X14Y146_C4;
  wire [0:0] CLBLM_R_X11Y146_SLICE_X14Y146_C5;
  wire [0:0] CLBLM_R_X11Y146_SLICE_X14Y146_C6;
  wire [0:0] CLBLM_R_X11Y146_SLICE_X14Y146_CLK;
  wire [0:0] CLBLM_R_X11Y146_SLICE_X14Y146_CMUX;
  wire [0:0] CLBLM_R_X11Y146_SLICE_X14Y146_CO5;
  wire [0:0] CLBLM_R_X11Y146_SLICE_X14Y146_CO6;
  wire [0:0] CLBLM_R_X11Y146_SLICE_X14Y146_C_CY;
  wire [0:0] CLBLM_R_X11Y146_SLICE_X14Y146_C_XOR;
  wire [0:0] CLBLM_R_X11Y146_SLICE_X14Y146_D;
  wire [0:0] CLBLM_R_X11Y146_SLICE_X14Y146_D1;
  wire [0:0] CLBLM_R_X11Y146_SLICE_X14Y146_D2;
  wire [0:0] CLBLM_R_X11Y146_SLICE_X14Y146_D3;
  wire [0:0] CLBLM_R_X11Y146_SLICE_X14Y146_D4;
  wire [0:0] CLBLM_R_X11Y146_SLICE_X14Y146_D5;
  wire [0:0] CLBLM_R_X11Y146_SLICE_X14Y146_D6;
  wire [0:0] CLBLM_R_X11Y146_SLICE_X14Y146_DO5;
  wire [0:0] CLBLM_R_X11Y146_SLICE_X14Y146_DO6;
  wire [0:0] CLBLM_R_X11Y146_SLICE_X14Y146_D_CY;
  wire [0:0] CLBLM_R_X11Y146_SLICE_X14Y146_D_XOR;
  wire [0:0] CLBLM_R_X11Y146_SLICE_X15Y146_A;
  wire [0:0] CLBLM_R_X11Y146_SLICE_X15Y146_A1;
  wire [0:0] CLBLM_R_X11Y146_SLICE_X15Y146_A2;
  wire [0:0] CLBLM_R_X11Y146_SLICE_X15Y146_A3;
  wire [0:0] CLBLM_R_X11Y146_SLICE_X15Y146_A4;
  wire [0:0] CLBLM_R_X11Y146_SLICE_X15Y146_A5;
  wire [0:0] CLBLM_R_X11Y146_SLICE_X15Y146_A6;
  wire [0:0] CLBLM_R_X11Y146_SLICE_X15Y146_AMUX;
  wire [0:0] CLBLM_R_X11Y146_SLICE_X15Y146_AO5;
  wire [0:0] CLBLM_R_X11Y146_SLICE_X15Y146_AO6;
  wire [0:0] CLBLM_R_X11Y146_SLICE_X15Y146_A_CY;
  wire [0:0] CLBLM_R_X11Y146_SLICE_X15Y146_A_XOR;
  wire [0:0] CLBLM_R_X11Y146_SLICE_X15Y146_B;
  wire [0:0] CLBLM_R_X11Y146_SLICE_X15Y146_B1;
  wire [0:0] CLBLM_R_X11Y146_SLICE_X15Y146_B2;
  wire [0:0] CLBLM_R_X11Y146_SLICE_X15Y146_B3;
  wire [0:0] CLBLM_R_X11Y146_SLICE_X15Y146_B4;
  wire [0:0] CLBLM_R_X11Y146_SLICE_X15Y146_B5;
  wire [0:0] CLBLM_R_X11Y146_SLICE_X15Y146_B6;
  wire [0:0] CLBLM_R_X11Y146_SLICE_X15Y146_BMUX;
  wire [0:0] CLBLM_R_X11Y146_SLICE_X15Y146_BO5;
  wire [0:0] CLBLM_R_X11Y146_SLICE_X15Y146_BO6;
  wire [0:0] CLBLM_R_X11Y146_SLICE_X15Y146_B_CY;
  wire [0:0] CLBLM_R_X11Y146_SLICE_X15Y146_B_XOR;
  wire [0:0] CLBLM_R_X11Y146_SLICE_X15Y146_C;
  wire [0:0] CLBLM_R_X11Y146_SLICE_X15Y146_C1;
  wire [0:0] CLBLM_R_X11Y146_SLICE_X15Y146_C2;
  wire [0:0] CLBLM_R_X11Y146_SLICE_X15Y146_C3;
  wire [0:0] CLBLM_R_X11Y146_SLICE_X15Y146_C4;
  wire [0:0] CLBLM_R_X11Y146_SLICE_X15Y146_C5;
  wire [0:0] CLBLM_R_X11Y146_SLICE_X15Y146_C6;
  wire [0:0] CLBLM_R_X11Y146_SLICE_X15Y146_CO5;
  wire [0:0] CLBLM_R_X11Y146_SLICE_X15Y146_CO6;
  wire [0:0] CLBLM_R_X11Y146_SLICE_X15Y146_C_CY;
  wire [0:0] CLBLM_R_X11Y146_SLICE_X15Y146_C_XOR;
  wire [0:0] CLBLM_R_X11Y146_SLICE_X15Y146_D;
  wire [0:0] CLBLM_R_X11Y146_SLICE_X15Y146_D1;
  wire [0:0] CLBLM_R_X11Y146_SLICE_X15Y146_D2;
  wire [0:0] CLBLM_R_X11Y146_SLICE_X15Y146_D3;
  wire [0:0] CLBLM_R_X11Y146_SLICE_X15Y146_D4;
  wire [0:0] CLBLM_R_X11Y146_SLICE_X15Y146_D5;
  wire [0:0] CLBLM_R_X11Y146_SLICE_X15Y146_D6;
  wire [0:0] CLBLM_R_X11Y146_SLICE_X15Y146_DO5;
  wire [0:0] CLBLM_R_X11Y146_SLICE_X15Y146_DO6;
  wire [0:0] CLBLM_R_X11Y146_SLICE_X15Y146_D_CY;
  wire [0:0] CLBLM_R_X11Y146_SLICE_X15Y146_D_XOR;
  wire [0:0] CLBLM_R_X11Y147_SLICE_X14Y147_A;
  wire [0:0] CLBLM_R_X11Y147_SLICE_X14Y147_A1;
  wire [0:0] CLBLM_R_X11Y147_SLICE_X14Y147_A2;
  wire [0:0] CLBLM_R_X11Y147_SLICE_X14Y147_A3;
  wire [0:0] CLBLM_R_X11Y147_SLICE_X14Y147_A4;
  wire [0:0] CLBLM_R_X11Y147_SLICE_X14Y147_A5;
  wire [0:0] CLBLM_R_X11Y147_SLICE_X14Y147_A6;
  wire [0:0] CLBLM_R_X11Y147_SLICE_X14Y147_AMUX;
  wire [0:0] CLBLM_R_X11Y147_SLICE_X14Y147_AO5;
  wire [0:0] CLBLM_R_X11Y147_SLICE_X14Y147_AO6;
  wire [0:0] CLBLM_R_X11Y147_SLICE_X14Y147_A_CY;
  wire [0:0] CLBLM_R_X11Y147_SLICE_X14Y147_A_XOR;
  wire [0:0] CLBLM_R_X11Y147_SLICE_X14Y147_B;
  wire [0:0] CLBLM_R_X11Y147_SLICE_X14Y147_B1;
  wire [0:0] CLBLM_R_X11Y147_SLICE_X14Y147_B2;
  wire [0:0] CLBLM_R_X11Y147_SLICE_X14Y147_B3;
  wire [0:0] CLBLM_R_X11Y147_SLICE_X14Y147_B4;
  wire [0:0] CLBLM_R_X11Y147_SLICE_X14Y147_B5;
  wire [0:0] CLBLM_R_X11Y147_SLICE_X14Y147_B6;
  wire [0:0] CLBLM_R_X11Y147_SLICE_X14Y147_BMUX;
  wire [0:0] CLBLM_R_X11Y147_SLICE_X14Y147_BO5;
  wire [0:0] CLBLM_R_X11Y147_SLICE_X14Y147_BO6;
  wire [0:0] CLBLM_R_X11Y147_SLICE_X14Y147_B_CY;
  wire [0:0] CLBLM_R_X11Y147_SLICE_X14Y147_B_XOR;
  wire [0:0] CLBLM_R_X11Y147_SLICE_X14Y147_C;
  wire [0:0] CLBLM_R_X11Y147_SLICE_X14Y147_C1;
  wire [0:0] CLBLM_R_X11Y147_SLICE_X14Y147_C2;
  wire [0:0] CLBLM_R_X11Y147_SLICE_X14Y147_C3;
  wire [0:0] CLBLM_R_X11Y147_SLICE_X14Y147_C4;
  wire [0:0] CLBLM_R_X11Y147_SLICE_X14Y147_C5;
  wire [0:0] CLBLM_R_X11Y147_SLICE_X14Y147_C6;
  wire [0:0] CLBLM_R_X11Y147_SLICE_X14Y147_CO5;
  wire [0:0] CLBLM_R_X11Y147_SLICE_X14Y147_CO6;
  wire [0:0] CLBLM_R_X11Y147_SLICE_X14Y147_C_CY;
  wire [0:0] CLBLM_R_X11Y147_SLICE_X14Y147_C_XOR;
  wire [0:0] CLBLM_R_X11Y147_SLICE_X14Y147_D;
  wire [0:0] CLBLM_R_X11Y147_SLICE_X14Y147_D1;
  wire [0:0] CLBLM_R_X11Y147_SLICE_X14Y147_D2;
  wire [0:0] CLBLM_R_X11Y147_SLICE_X14Y147_D3;
  wire [0:0] CLBLM_R_X11Y147_SLICE_X14Y147_D4;
  wire [0:0] CLBLM_R_X11Y147_SLICE_X14Y147_D5;
  wire [0:0] CLBLM_R_X11Y147_SLICE_X14Y147_D6;
  wire [0:0] CLBLM_R_X11Y147_SLICE_X14Y147_DO5;
  wire [0:0] CLBLM_R_X11Y147_SLICE_X14Y147_DO6;
  wire [0:0] CLBLM_R_X11Y147_SLICE_X14Y147_D_CY;
  wire [0:0] CLBLM_R_X11Y147_SLICE_X14Y147_D_XOR;
  wire [0:0] CLBLM_R_X11Y147_SLICE_X15Y147_A;
  wire [0:0] CLBLM_R_X11Y147_SLICE_X15Y147_A1;
  wire [0:0] CLBLM_R_X11Y147_SLICE_X15Y147_A2;
  wire [0:0] CLBLM_R_X11Y147_SLICE_X15Y147_A3;
  wire [0:0] CLBLM_R_X11Y147_SLICE_X15Y147_A4;
  wire [0:0] CLBLM_R_X11Y147_SLICE_X15Y147_A5;
  wire [0:0] CLBLM_R_X11Y147_SLICE_X15Y147_A6;
  wire [0:0] CLBLM_R_X11Y147_SLICE_X15Y147_AO5;
  wire [0:0] CLBLM_R_X11Y147_SLICE_X15Y147_AO6;
  wire [0:0] CLBLM_R_X11Y147_SLICE_X15Y147_A_CY;
  wire [0:0] CLBLM_R_X11Y147_SLICE_X15Y147_A_XOR;
  wire [0:0] CLBLM_R_X11Y147_SLICE_X15Y147_B;
  wire [0:0] CLBLM_R_X11Y147_SLICE_X15Y147_B1;
  wire [0:0] CLBLM_R_X11Y147_SLICE_X15Y147_B2;
  wire [0:0] CLBLM_R_X11Y147_SLICE_X15Y147_B3;
  wire [0:0] CLBLM_R_X11Y147_SLICE_X15Y147_B4;
  wire [0:0] CLBLM_R_X11Y147_SLICE_X15Y147_B5;
  wire [0:0] CLBLM_R_X11Y147_SLICE_X15Y147_B6;
  wire [0:0] CLBLM_R_X11Y147_SLICE_X15Y147_BO5;
  wire [0:0] CLBLM_R_X11Y147_SLICE_X15Y147_BO6;
  wire [0:0] CLBLM_R_X11Y147_SLICE_X15Y147_B_CY;
  wire [0:0] CLBLM_R_X11Y147_SLICE_X15Y147_B_XOR;
  wire [0:0] CLBLM_R_X11Y147_SLICE_X15Y147_C;
  wire [0:0] CLBLM_R_X11Y147_SLICE_X15Y147_C1;
  wire [0:0] CLBLM_R_X11Y147_SLICE_X15Y147_C2;
  wire [0:0] CLBLM_R_X11Y147_SLICE_X15Y147_C3;
  wire [0:0] CLBLM_R_X11Y147_SLICE_X15Y147_C4;
  wire [0:0] CLBLM_R_X11Y147_SLICE_X15Y147_C5;
  wire [0:0] CLBLM_R_X11Y147_SLICE_X15Y147_C6;
  wire [0:0] CLBLM_R_X11Y147_SLICE_X15Y147_CO5;
  wire [0:0] CLBLM_R_X11Y147_SLICE_X15Y147_CO6;
  wire [0:0] CLBLM_R_X11Y147_SLICE_X15Y147_C_CY;
  wire [0:0] CLBLM_R_X11Y147_SLICE_X15Y147_C_XOR;
  wire [0:0] CLBLM_R_X11Y147_SLICE_X15Y147_D;
  wire [0:0] CLBLM_R_X11Y147_SLICE_X15Y147_D1;
  wire [0:0] CLBLM_R_X11Y147_SLICE_X15Y147_D2;
  wire [0:0] CLBLM_R_X11Y147_SLICE_X15Y147_D3;
  wire [0:0] CLBLM_R_X11Y147_SLICE_X15Y147_D4;
  wire [0:0] CLBLM_R_X11Y147_SLICE_X15Y147_D5;
  wire [0:0] CLBLM_R_X11Y147_SLICE_X15Y147_D6;
  wire [0:0] CLBLM_R_X11Y147_SLICE_X15Y147_DO5;
  wire [0:0] CLBLM_R_X11Y147_SLICE_X15Y147_DO6;
  wire [0:0] CLBLM_R_X11Y147_SLICE_X15Y147_D_CY;
  wire [0:0] CLBLM_R_X11Y147_SLICE_X15Y147_D_XOR;
  wire [0:0] CLBLM_R_X11Y148_SLICE_X14Y148_A;
  wire [0:0] CLBLM_R_X11Y148_SLICE_X14Y148_A1;
  wire [0:0] CLBLM_R_X11Y148_SLICE_X14Y148_A2;
  wire [0:0] CLBLM_R_X11Y148_SLICE_X14Y148_A3;
  wire [0:0] CLBLM_R_X11Y148_SLICE_X14Y148_A4;
  wire [0:0] CLBLM_R_X11Y148_SLICE_X14Y148_A5;
  wire [0:0] CLBLM_R_X11Y148_SLICE_X14Y148_A6;
  wire [0:0] CLBLM_R_X11Y148_SLICE_X14Y148_AO5;
  wire [0:0] CLBLM_R_X11Y148_SLICE_X14Y148_AO6;
  wire [0:0] CLBLM_R_X11Y148_SLICE_X14Y148_A_CY;
  wire [0:0] CLBLM_R_X11Y148_SLICE_X14Y148_A_XOR;
  wire [0:0] CLBLM_R_X11Y148_SLICE_X14Y148_B;
  wire [0:0] CLBLM_R_X11Y148_SLICE_X14Y148_B1;
  wire [0:0] CLBLM_R_X11Y148_SLICE_X14Y148_B2;
  wire [0:0] CLBLM_R_X11Y148_SLICE_X14Y148_B3;
  wire [0:0] CLBLM_R_X11Y148_SLICE_X14Y148_B4;
  wire [0:0] CLBLM_R_X11Y148_SLICE_X14Y148_B5;
  wire [0:0] CLBLM_R_X11Y148_SLICE_X14Y148_B6;
  wire [0:0] CLBLM_R_X11Y148_SLICE_X14Y148_BO5;
  wire [0:0] CLBLM_R_X11Y148_SLICE_X14Y148_BO6;
  wire [0:0] CLBLM_R_X11Y148_SLICE_X14Y148_B_CY;
  wire [0:0] CLBLM_R_X11Y148_SLICE_X14Y148_B_XOR;
  wire [0:0] CLBLM_R_X11Y148_SLICE_X14Y148_C;
  wire [0:0] CLBLM_R_X11Y148_SLICE_X14Y148_C1;
  wire [0:0] CLBLM_R_X11Y148_SLICE_X14Y148_C2;
  wire [0:0] CLBLM_R_X11Y148_SLICE_X14Y148_C3;
  wire [0:0] CLBLM_R_X11Y148_SLICE_X14Y148_C4;
  wire [0:0] CLBLM_R_X11Y148_SLICE_X14Y148_C5;
  wire [0:0] CLBLM_R_X11Y148_SLICE_X14Y148_C6;
  wire [0:0] CLBLM_R_X11Y148_SLICE_X14Y148_CO5;
  wire [0:0] CLBLM_R_X11Y148_SLICE_X14Y148_CO6;
  wire [0:0] CLBLM_R_X11Y148_SLICE_X14Y148_C_CY;
  wire [0:0] CLBLM_R_X11Y148_SLICE_X14Y148_C_XOR;
  wire [0:0] CLBLM_R_X11Y148_SLICE_X14Y148_D;
  wire [0:0] CLBLM_R_X11Y148_SLICE_X14Y148_D1;
  wire [0:0] CLBLM_R_X11Y148_SLICE_X14Y148_D2;
  wire [0:0] CLBLM_R_X11Y148_SLICE_X14Y148_D3;
  wire [0:0] CLBLM_R_X11Y148_SLICE_X14Y148_D4;
  wire [0:0] CLBLM_R_X11Y148_SLICE_X14Y148_D5;
  wire [0:0] CLBLM_R_X11Y148_SLICE_X14Y148_D6;
  wire [0:0] CLBLM_R_X11Y148_SLICE_X14Y148_DO5;
  wire [0:0] CLBLM_R_X11Y148_SLICE_X14Y148_DO6;
  wire [0:0] CLBLM_R_X11Y148_SLICE_X14Y148_D_CY;
  wire [0:0] CLBLM_R_X11Y148_SLICE_X14Y148_D_XOR;
  wire [0:0] CLBLM_R_X11Y148_SLICE_X15Y148_A;
  wire [0:0] CLBLM_R_X11Y148_SLICE_X15Y148_A1;
  wire [0:0] CLBLM_R_X11Y148_SLICE_X15Y148_A2;
  wire [0:0] CLBLM_R_X11Y148_SLICE_X15Y148_A3;
  wire [0:0] CLBLM_R_X11Y148_SLICE_X15Y148_A4;
  wire [0:0] CLBLM_R_X11Y148_SLICE_X15Y148_A5;
  wire [0:0] CLBLM_R_X11Y148_SLICE_X15Y148_A6;
  wire [0:0] CLBLM_R_X11Y148_SLICE_X15Y148_AO5;
  wire [0:0] CLBLM_R_X11Y148_SLICE_X15Y148_AO6;
  wire [0:0] CLBLM_R_X11Y148_SLICE_X15Y148_A_CY;
  wire [0:0] CLBLM_R_X11Y148_SLICE_X15Y148_A_XOR;
  wire [0:0] CLBLM_R_X11Y148_SLICE_X15Y148_B;
  wire [0:0] CLBLM_R_X11Y148_SLICE_X15Y148_B1;
  wire [0:0] CLBLM_R_X11Y148_SLICE_X15Y148_B2;
  wire [0:0] CLBLM_R_X11Y148_SLICE_X15Y148_B3;
  wire [0:0] CLBLM_R_X11Y148_SLICE_X15Y148_B4;
  wire [0:0] CLBLM_R_X11Y148_SLICE_X15Y148_B5;
  wire [0:0] CLBLM_R_X11Y148_SLICE_X15Y148_B6;
  wire [0:0] CLBLM_R_X11Y148_SLICE_X15Y148_BMUX;
  wire [0:0] CLBLM_R_X11Y148_SLICE_X15Y148_BO5;
  wire [0:0] CLBLM_R_X11Y148_SLICE_X15Y148_BO6;
  wire [0:0] CLBLM_R_X11Y148_SLICE_X15Y148_B_CY;
  wire [0:0] CLBLM_R_X11Y148_SLICE_X15Y148_B_XOR;
  wire [0:0] CLBLM_R_X11Y148_SLICE_X15Y148_C;
  wire [0:0] CLBLM_R_X11Y148_SLICE_X15Y148_C1;
  wire [0:0] CLBLM_R_X11Y148_SLICE_X15Y148_C2;
  wire [0:0] CLBLM_R_X11Y148_SLICE_X15Y148_C3;
  wire [0:0] CLBLM_R_X11Y148_SLICE_X15Y148_C4;
  wire [0:0] CLBLM_R_X11Y148_SLICE_X15Y148_C5;
  wire [0:0] CLBLM_R_X11Y148_SLICE_X15Y148_C6;
  wire [0:0] CLBLM_R_X11Y148_SLICE_X15Y148_CMUX;
  wire [0:0] CLBLM_R_X11Y148_SLICE_X15Y148_CO5;
  wire [0:0] CLBLM_R_X11Y148_SLICE_X15Y148_CO6;
  wire [0:0] CLBLM_R_X11Y148_SLICE_X15Y148_C_CY;
  wire [0:0] CLBLM_R_X11Y148_SLICE_X15Y148_C_XOR;
  wire [0:0] CLBLM_R_X11Y148_SLICE_X15Y148_D;
  wire [0:0] CLBLM_R_X11Y148_SLICE_X15Y148_D1;
  wire [0:0] CLBLM_R_X11Y148_SLICE_X15Y148_D2;
  wire [0:0] CLBLM_R_X11Y148_SLICE_X15Y148_D3;
  wire [0:0] CLBLM_R_X11Y148_SLICE_X15Y148_D4;
  wire [0:0] CLBLM_R_X11Y148_SLICE_X15Y148_D5;
  wire [0:0] CLBLM_R_X11Y148_SLICE_X15Y148_D6;
  wire [0:0] CLBLM_R_X11Y148_SLICE_X15Y148_DO5;
  wire [0:0] CLBLM_R_X11Y148_SLICE_X15Y148_DO6;
  wire [0:0] CLBLM_R_X11Y148_SLICE_X15Y148_D_CY;
  wire [0:0] CLBLM_R_X11Y148_SLICE_X15Y148_D_XOR;
  wire [0:0] CLBLM_R_X11Y149_SLICE_X14Y149_A;
  wire [0:0] CLBLM_R_X11Y149_SLICE_X14Y149_A1;
  wire [0:0] CLBLM_R_X11Y149_SLICE_X14Y149_A2;
  wire [0:0] CLBLM_R_X11Y149_SLICE_X14Y149_A3;
  wire [0:0] CLBLM_R_X11Y149_SLICE_X14Y149_A4;
  wire [0:0] CLBLM_R_X11Y149_SLICE_X14Y149_A5;
  wire [0:0] CLBLM_R_X11Y149_SLICE_X14Y149_A6;
  wire [0:0] CLBLM_R_X11Y149_SLICE_X14Y149_AO5;
  wire [0:0] CLBLM_R_X11Y149_SLICE_X14Y149_AO6;
  wire [0:0] CLBLM_R_X11Y149_SLICE_X14Y149_A_CY;
  wire [0:0] CLBLM_R_X11Y149_SLICE_X14Y149_A_XOR;
  wire [0:0] CLBLM_R_X11Y149_SLICE_X14Y149_B;
  wire [0:0] CLBLM_R_X11Y149_SLICE_X14Y149_B1;
  wire [0:0] CLBLM_R_X11Y149_SLICE_X14Y149_B2;
  wire [0:0] CLBLM_R_X11Y149_SLICE_X14Y149_B3;
  wire [0:0] CLBLM_R_X11Y149_SLICE_X14Y149_B4;
  wire [0:0] CLBLM_R_X11Y149_SLICE_X14Y149_B5;
  wire [0:0] CLBLM_R_X11Y149_SLICE_X14Y149_B6;
  wire [0:0] CLBLM_R_X11Y149_SLICE_X14Y149_BO5;
  wire [0:0] CLBLM_R_X11Y149_SLICE_X14Y149_BO6;
  wire [0:0] CLBLM_R_X11Y149_SLICE_X14Y149_B_CY;
  wire [0:0] CLBLM_R_X11Y149_SLICE_X14Y149_B_XOR;
  wire [0:0] CLBLM_R_X11Y149_SLICE_X14Y149_C;
  wire [0:0] CLBLM_R_X11Y149_SLICE_X14Y149_C1;
  wire [0:0] CLBLM_R_X11Y149_SLICE_X14Y149_C2;
  wire [0:0] CLBLM_R_X11Y149_SLICE_X14Y149_C3;
  wire [0:0] CLBLM_R_X11Y149_SLICE_X14Y149_C4;
  wire [0:0] CLBLM_R_X11Y149_SLICE_X14Y149_C5;
  wire [0:0] CLBLM_R_X11Y149_SLICE_X14Y149_C6;
  wire [0:0] CLBLM_R_X11Y149_SLICE_X14Y149_CO5;
  wire [0:0] CLBLM_R_X11Y149_SLICE_X14Y149_CO6;
  wire [0:0] CLBLM_R_X11Y149_SLICE_X14Y149_C_CY;
  wire [0:0] CLBLM_R_X11Y149_SLICE_X14Y149_C_XOR;
  wire [0:0] CLBLM_R_X11Y149_SLICE_X14Y149_D;
  wire [0:0] CLBLM_R_X11Y149_SLICE_X14Y149_D1;
  wire [0:0] CLBLM_R_X11Y149_SLICE_X14Y149_D2;
  wire [0:0] CLBLM_R_X11Y149_SLICE_X14Y149_D3;
  wire [0:0] CLBLM_R_X11Y149_SLICE_X14Y149_D4;
  wire [0:0] CLBLM_R_X11Y149_SLICE_X14Y149_D5;
  wire [0:0] CLBLM_R_X11Y149_SLICE_X14Y149_D6;
  wire [0:0] CLBLM_R_X11Y149_SLICE_X14Y149_DMUX;
  wire [0:0] CLBLM_R_X11Y149_SLICE_X14Y149_DO5;
  wire [0:0] CLBLM_R_X11Y149_SLICE_X14Y149_DO6;
  wire [0:0] CLBLM_R_X11Y149_SLICE_X14Y149_D_CY;
  wire [0:0] CLBLM_R_X11Y149_SLICE_X14Y149_D_XOR;
  wire [0:0] CLBLM_R_X11Y149_SLICE_X15Y149_A;
  wire [0:0] CLBLM_R_X11Y149_SLICE_X15Y149_A1;
  wire [0:0] CLBLM_R_X11Y149_SLICE_X15Y149_A2;
  wire [0:0] CLBLM_R_X11Y149_SLICE_X15Y149_A3;
  wire [0:0] CLBLM_R_X11Y149_SLICE_X15Y149_A4;
  wire [0:0] CLBLM_R_X11Y149_SLICE_X15Y149_A5;
  wire [0:0] CLBLM_R_X11Y149_SLICE_X15Y149_A6;
  wire [0:0] CLBLM_R_X11Y149_SLICE_X15Y149_AO5;
  wire [0:0] CLBLM_R_X11Y149_SLICE_X15Y149_AO6;
  wire [0:0] CLBLM_R_X11Y149_SLICE_X15Y149_A_CY;
  wire [0:0] CLBLM_R_X11Y149_SLICE_X15Y149_A_XOR;
  wire [0:0] CLBLM_R_X11Y149_SLICE_X15Y149_B;
  wire [0:0] CLBLM_R_X11Y149_SLICE_X15Y149_B1;
  wire [0:0] CLBLM_R_X11Y149_SLICE_X15Y149_B2;
  wire [0:0] CLBLM_R_X11Y149_SLICE_X15Y149_B3;
  wire [0:0] CLBLM_R_X11Y149_SLICE_X15Y149_B4;
  wire [0:0] CLBLM_R_X11Y149_SLICE_X15Y149_B5;
  wire [0:0] CLBLM_R_X11Y149_SLICE_X15Y149_B6;
  wire [0:0] CLBLM_R_X11Y149_SLICE_X15Y149_BO5;
  wire [0:0] CLBLM_R_X11Y149_SLICE_X15Y149_BO6;
  wire [0:0] CLBLM_R_X11Y149_SLICE_X15Y149_B_CY;
  wire [0:0] CLBLM_R_X11Y149_SLICE_X15Y149_B_XOR;
  wire [0:0] CLBLM_R_X11Y149_SLICE_X15Y149_C;
  wire [0:0] CLBLM_R_X11Y149_SLICE_X15Y149_C1;
  wire [0:0] CLBLM_R_X11Y149_SLICE_X15Y149_C2;
  wire [0:0] CLBLM_R_X11Y149_SLICE_X15Y149_C3;
  wire [0:0] CLBLM_R_X11Y149_SLICE_X15Y149_C4;
  wire [0:0] CLBLM_R_X11Y149_SLICE_X15Y149_C5;
  wire [0:0] CLBLM_R_X11Y149_SLICE_X15Y149_C6;
  wire [0:0] CLBLM_R_X11Y149_SLICE_X15Y149_CO5;
  wire [0:0] CLBLM_R_X11Y149_SLICE_X15Y149_CO6;
  wire [0:0] CLBLM_R_X11Y149_SLICE_X15Y149_C_CY;
  wire [0:0] CLBLM_R_X11Y149_SLICE_X15Y149_C_XOR;
  wire [0:0] CLBLM_R_X11Y149_SLICE_X15Y149_D;
  wire [0:0] CLBLM_R_X11Y149_SLICE_X15Y149_D1;
  wire [0:0] CLBLM_R_X11Y149_SLICE_X15Y149_D2;
  wire [0:0] CLBLM_R_X11Y149_SLICE_X15Y149_D3;
  wire [0:0] CLBLM_R_X11Y149_SLICE_X15Y149_D4;
  wire [0:0] CLBLM_R_X11Y149_SLICE_X15Y149_D5;
  wire [0:0] CLBLM_R_X11Y149_SLICE_X15Y149_D6;
  wire [0:0] CLBLM_R_X11Y149_SLICE_X15Y149_DO5;
  wire [0:0] CLBLM_R_X11Y149_SLICE_X15Y149_DO6;
  wire [0:0] CLBLM_R_X11Y149_SLICE_X15Y149_D_CY;
  wire [0:0] CLBLM_R_X11Y149_SLICE_X15Y149_D_XOR;
  wire [0:0] CLBLM_R_X11Y150_SLICE_X14Y150_A;
  wire [0:0] CLBLM_R_X11Y150_SLICE_X14Y150_A1;
  wire [0:0] CLBLM_R_X11Y150_SLICE_X14Y150_A2;
  wire [0:0] CLBLM_R_X11Y150_SLICE_X14Y150_A3;
  wire [0:0] CLBLM_R_X11Y150_SLICE_X14Y150_A4;
  wire [0:0] CLBLM_R_X11Y150_SLICE_X14Y150_A5;
  wire [0:0] CLBLM_R_X11Y150_SLICE_X14Y150_A6;
  wire [0:0] CLBLM_R_X11Y150_SLICE_X14Y150_AO5;
  wire [0:0] CLBLM_R_X11Y150_SLICE_X14Y150_AO6;
  wire [0:0] CLBLM_R_X11Y150_SLICE_X14Y150_AQ;
  wire [0:0] CLBLM_R_X11Y150_SLICE_X14Y150_AX;
  wire [0:0] CLBLM_R_X11Y150_SLICE_X14Y150_A_CY;
  wire [0:0] CLBLM_R_X11Y150_SLICE_X14Y150_A_XOR;
  wire [0:0] CLBLM_R_X11Y150_SLICE_X14Y150_B;
  wire [0:0] CLBLM_R_X11Y150_SLICE_X14Y150_B1;
  wire [0:0] CLBLM_R_X11Y150_SLICE_X14Y150_B2;
  wire [0:0] CLBLM_R_X11Y150_SLICE_X14Y150_B3;
  wire [0:0] CLBLM_R_X11Y150_SLICE_X14Y150_B4;
  wire [0:0] CLBLM_R_X11Y150_SLICE_X14Y150_B5;
  wire [0:0] CLBLM_R_X11Y150_SLICE_X14Y150_B6;
  wire [0:0] CLBLM_R_X11Y150_SLICE_X14Y150_BO5;
  wire [0:0] CLBLM_R_X11Y150_SLICE_X14Y150_BO6;
  wire [0:0] CLBLM_R_X11Y150_SLICE_X14Y150_B_CY;
  wire [0:0] CLBLM_R_X11Y150_SLICE_X14Y150_B_XOR;
  wire [0:0] CLBLM_R_X11Y150_SLICE_X14Y150_C;
  wire [0:0] CLBLM_R_X11Y150_SLICE_X14Y150_C1;
  wire [0:0] CLBLM_R_X11Y150_SLICE_X14Y150_C2;
  wire [0:0] CLBLM_R_X11Y150_SLICE_X14Y150_C3;
  wire [0:0] CLBLM_R_X11Y150_SLICE_X14Y150_C4;
  wire [0:0] CLBLM_R_X11Y150_SLICE_X14Y150_C5;
  wire [0:0] CLBLM_R_X11Y150_SLICE_X14Y150_C6;
  wire [0:0] CLBLM_R_X11Y150_SLICE_X14Y150_CE;
  wire [0:0] CLBLM_R_X11Y150_SLICE_X14Y150_CLK;
  wire [0:0] CLBLM_R_X11Y150_SLICE_X14Y150_CO5;
  wire [0:0] CLBLM_R_X11Y150_SLICE_X14Y150_CO6;
  wire [0:0] CLBLM_R_X11Y150_SLICE_X14Y150_C_CY;
  wire [0:0] CLBLM_R_X11Y150_SLICE_X14Y150_C_XOR;
  wire [0:0] CLBLM_R_X11Y150_SLICE_X14Y150_D;
  wire [0:0] CLBLM_R_X11Y150_SLICE_X14Y150_D1;
  wire [0:0] CLBLM_R_X11Y150_SLICE_X14Y150_D2;
  wire [0:0] CLBLM_R_X11Y150_SLICE_X14Y150_D3;
  wire [0:0] CLBLM_R_X11Y150_SLICE_X14Y150_D4;
  wire [0:0] CLBLM_R_X11Y150_SLICE_X14Y150_D5;
  wire [0:0] CLBLM_R_X11Y150_SLICE_X14Y150_D6;
  wire [0:0] CLBLM_R_X11Y150_SLICE_X14Y150_DO5;
  wire [0:0] CLBLM_R_X11Y150_SLICE_X14Y150_DO6;
  wire [0:0] CLBLM_R_X11Y150_SLICE_X14Y150_D_CY;
  wire [0:0] CLBLM_R_X11Y150_SLICE_X14Y150_D_XOR;
  wire [0:0] CLBLM_R_X11Y150_SLICE_X15Y150_A;
  wire [0:0] CLBLM_R_X11Y150_SLICE_X15Y150_A1;
  wire [0:0] CLBLM_R_X11Y150_SLICE_X15Y150_A2;
  wire [0:0] CLBLM_R_X11Y150_SLICE_X15Y150_A3;
  wire [0:0] CLBLM_R_X11Y150_SLICE_X15Y150_A4;
  wire [0:0] CLBLM_R_X11Y150_SLICE_X15Y150_A5;
  wire [0:0] CLBLM_R_X11Y150_SLICE_X15Y150_A6;
  wire [0:0] CLBLM_R_X11Y150_SLICE_X15Y150_AO5;
  wire [0:0] CLBLM_R_X11Y150_SLICE_X15Y150_AO6;
  wire [0:0] CLBLM_R_X11Y150_SLICE_X15Y150_A_CY;
  wire [0:0] CLBLM_R_X11Y150_SLICE_X15Y150_A_XOR;
  wire [0:0] CLBLM_R_X11Y150_SLICE_X15Y150_B;
  wire [0:0] CLBLM_R_X11Y150_SLICE_X15Y150_B1;
  wire [0:0] CLBLM_R_X11Y150_SLICE_X15Y150_B2;
  wire [0:0] CLBLM_R_X11Y150_SLICE_X15Y150_B3;
  wire [0:0] CLBLM_R_X11Y150_SLICE_X15Y150_B4;
  wire [0:0] CLBLM_R_X11Y150_SLICE_X15Y150_B5;
  wire [0:0] CLBLM_R_X11Y150_SLICE_X15Y150_B6;
  wire [0:0] CLBLM_R_X11Y150_SLICE_X15Y150_BO5;
  wire [0:0] CLBLM_R_X11Y150_SLICE_X15Y150_BO6;
  wire [0:0] CLBLM_R_X11Y150_SLICE_X15Y150_B_CY;
  wire [0:0] CLBLM_R_X11Y150_SLICE_X15Y150_B_XOR;
  wire [0:0] CLBLM_R_X11Y150_SLICE_X15Y150_C;
  wire [0:0] CLBLM_R_X11Y150_SLICE_X15Y150_C1;
  wire [0:0] CLBLM_R_X11Y150_SLICE_X15Y150_C2;
  wire [0:0] CLBLM_R_X11Y150_SLICE_X15Y150_C3;
  wire [0:0] CLBLM_R_X11Y150_SLICE_X15Y150_C4;
  wire [0:0] CLBLM_R_X11Y150_SLICE_X15Y150_C5;
  wire [0:0] CLBLM_R_X11Y150_SLICE_X15Y150_C6;
  wire [0:0] CLBLM_R_X11Y150_SLICE_X15Y150_CO5;
  wire [0:0] CLBLM_R_X11Y150_SLICE_X15Y150_CO6;
  wire [0:0] CLBLM_R_X11Y150_SLICE_X15Y150_C_CY;
  wire [0:0] CLBLM_R_X11Y150_SLICE_X15Y150_C_XOR;
  wire [0:0] CLBLM_R_X11Y150_SLICE_X15Y150_D;
  wire [0:0] CLBLM_R_X11Y150_SLICE_X15Y150_D1;
  wire [0:0] CLBLM_R_X11Y150_SLICE_X15Y150_D2;
  wire [0:0] CLBLM_R_X11Y150_SLICE_X15Y150_D3;
  wire [0:0] CLBLM_R_X11Y150_SLICE_X15Y150_D4;
  wire [0:0] CLBLM_R_X11Y150_SLICE_X15Y150_D5;
  wire [0:0] CLBLM_R_X11Y150_SLICE_X15Y150_D6;
  wire [0:0] CLBLM_R_X11Y150_SLICE_X15Y150_DO5;
  wire [0:0] CLBLM_R_X11Y150_SLICE_X15Y150_DO6;
  wire [0:0] CLBLM_R_X11Y150_SLICE_X15Y150_D_CY;
  wire [0:0] CLBLM_R_X11Y150_SLICE_X15Y150_D_XOR;
  wire [0:0] CLBLM_R_X11Y151_SLICE_X14Y151_A;
  wire [0:0] CLBLM_R_X11Y151_SLICE_X14Y151_A1;
  wire [0:0] CLBLM_R_X11Y151_SLICE_X14Y151_A2;
  wire [0:0] CLBLM_R_X11Y151_SLICE_X14Y151_A3;
  wire [0:0] CLBLM_R_X11Y151_SLICE_X14Y151_A4;
  wire [0:0] CLBLM_R_X11Y151_SLICE_X14Y151_A5;
  wire [0:0] CLBLM_R_X11Y151_SLICE_X14Y151_A6;
  wire [0:0] CLBLM_R_X11Y151_SLICE_X14Y151_AO5;
  wire [0:0] CLBLM_R_X11Y151_SLICE_X14Y151_AO6;
  wire [0:0] CLBLM_R_X11Y151_SLICE_X14Y151_AQ;
  wire [0:0] CLBLM_R_X11Y151_SLICE_X14Y151_A_CY;
  wire [0:0] CLBLM_R_X11Y151_SLICE_X14Y151_A_XOR;
  wire [0:0] CLBLM_R_X11Y151_SLICE_X14Y151_B;
  wire [0:0] CLBLM_R_X11Y151_SLICE_X14Y151_B1;
  wire [0:0] CLBLM_R_X11Y151_SLICE_X14Y151_B2;
  wire [0:0] CLBLM_R_X11Y151_SLICE_X14Y151_B3;
  wire [0:0] CLBLM_R_X11Y151_SLICE_X14Y151_B4;
  wire [0:0] CLBLM_R_X11Y151_SLICE_X14Y151_B5;
  wire [0:0] CLBLM_R_X11Y151_SLICE_X14Y151_B6;
  wire [0:0] CLBLM_R_X11Y151_SLICE_X14Y151_BO5;
  wire [0:0] CLBLM_R_X11Y151_SLICE_X14Y151_BO6;
  wire [0:0] CLBLM_R_X11Y151_SLICE_X14Y151_B_CY;
  wire [0:0] CLBLM_R_X11Y151_SLICE_X14Y151_B_XOR;
  wire [0:0] CLBLM_R_X11Y151_SLICE_X14Y151_C;
  wire [0:0] CLBLM_R_X11Y151_SLICE_X14Y151_C1;
  wire [0:0] CLBLM_R_X11Y151_SLICE_X14Y151_C2;
  wire [0:0] CLBLM_R_X11Y151_SLICE_X14Y151_C3;
  wire [0:0] CLBLM_R_X11Y151_SLICE_X14Y151_C4;
  wire [0:0] CLBLM_R_X11Y151_SLICE_X14Y151_C5;
  wire [0:0] CLBLM_R_X11Y151_SLICE_X14Y151_C6;
  wire [0:0] CLBLM_R_X11Y151_SLICE_X14Y151_CLK;
  wire [0:0] CLBLM_R_X11Y151_SLICE_X14Y151_CO5;
  wire [0:0] CLBLM_R_X11Y151_SLICE_X14Y151_CO6;
  wire [0:0] CLBLM_R_X11Y151_SLICE_X14Y151_C_CY;
  wire [0:0] CLBLM_R_X11Y151_SLICE_X14Y151_C_XOR;
  wire [0:0] CLBLM_R_X11Y151_SLICE_X14Y151_D;
  wire [0:0] CLBLM_R_X11Y151_SLICE_X14Y151_D1;
  wire [0:0] CLBLM_R_X11Y151_SLICE_X14Y151_D2;
  wire [0:0] CLBLM_R_X11Y151_SLICE_X14Y151_D3;
  wire [0:0] CLBLM_R_X11Y151_SLICE_X14Y151_D4;
  wire [0:0] CLBLM_R_X11Y151_SLICE_X14Y151_D5;
  wire [0:0] CLBLM_R_X11Y151_SLICE_X14Y151_D6;
  wire [0:0] CLBLM_R_X11Y151_SLICE_X14Y151_DO5;
  wire [0:0] CLBLM_R_X11Y151_SLICE_X14Y151_DO6;
  wire [0:0] CLBLM_R_X11Y151_SLICE_X14Y151_D_CY;
  wire [0:0] CLBLM_R_X11Y151_SLICE_X14Y151_D_XOR;
  wire [0:0] CLBLM_R_X11Y151_SLICE_X15Y151_A;
  wire [0:0] CLBLM_R_X11Y151_SLICE_X15Y151_A1;
  wire [0:0] CLBLM_R_X11Y151_SLICE_X15Y151_A2;
  wire [0:0] CLBLM_R_X11Y151_SLICE_X15Y151_A3;
  wire [0:0] CLBLM_R_X11Y151_SLICE_X15Y151_A4;
  wire [0:0] CLBLM_R_X11Y151_SLICE_X15Y151_A5;
  wire [0:0] CLBLM_R_X11Y151_SLICE_X15Y151_A5Q;
  wire [0:0] CLBLM_R_X11Y151_SLICE_X15Y151_A6;
  wire [0:0] CLBLM_R_X11Y151_SLICE_X15Y151_AMUX;
  wire [0:0] CLBLM_R_X11Y151_SLICE_X15Y151_AO5;
  wire [0:0] CLBLM_R_X11Y151_SLICE_X15Y151_AO6;
  wire [0:0] CLBLM_R_X11Y151_SLICE_X15Y151_AQ;
  wire [0:0] CLBLM_R_X11Y151_SLICE_X15Y151_A_CY;
  wire [0:0] CLBLM_R_X11Y151_SLICE_X15Y151_A_XOR;
  wire [0:0] CLBLM_R_X11Y151_SLICE_X15Y151_B;
  wire [0:0] CLBLM_R_X11Y151_SLICE_X15Y151_B1;
  wire [0:0] CLBLM_R_X11Y151_SLICE_X15Y151_B2;
  wire [0:0] CLBLM_R_X11Y151_SLICE_X15Y151_B3;
  wire [0:0] CLBLM_R_X11Y151_SLICE_X15Y151_B4;
  wire [0:0] CLBLM_R_X11Y151_SLICE_X15Y151_B5;
  wire [0:0] CLBLM_R_X11Y151_SLICE_X15Y151_B6;
  wire [0:0] CLBLM_R_X11Y151_SLICE_X15Y151_BO5;
  wire [0:0] CLBLM_R_X11Y151_SLICE_X15Y151_BO6;
  wire [0:0] CLBLM_R_X11Y151_SLICE_X15Y151_B_CY;
  wire [0:0] CLBLM_R_X11Y151_SLICE_X15Y151_B_XOR;
  wire [0:0] CLBLM_R_X11Y151_SLICE_X15Y151_C;
  wire [0:0] CLBLM_R_X11Y151_SLICE_X15Y151_C1;
  wire [0:0] CLBLM_R_X11Y151_SLICE_X15Y151_C2;
  wire [0:0] CLBLM_R_X11Y151_SLICE_X15Y151_C3;
  wire [0:0] CLBLM_R_X11Y151_SLICE_X15Y151_C4;
  wire [0:0] CLBLM_R_X11Y151_SLICE_X15Y151_C5;
  wire [0:0] CLBLM_R_X11Y151_SLICE_X15Y151_C6;
  wire [0:0] CLBLM_R_X11Y151_SLICE_X15Y151_CLK;
  wire [0:0] CLBLM_R_X11Y151_SLICE_X15Y151_CO5;
  wire [0:0] CLBLM_R_X11Y151_SLICE_X15Y151_CO6;
  wire [0:0] CLBLM_R_X11Y151_SLICE_X15Y151_C_CY;
  wire [0:0] CLBLM_R_X11Y151_SLICE_X15Y151_C_XOR;
  wire [0:0] CLBLM_R_X11Y151_SLICE_X15Y151_D;
  wire [0:0] CLBLM_R_X11Y151_SLICE_X15Y151_D1;
  wire [0:0] CLBLM_R_X11Y151_SLICE_X15Y151_D2;
  wire [0:0] CLBLM_R_X11Y151_SLICE_X15Y151_D3;
  wire [0:0] CLBLM_R_X11Y151_SLICE_X15Y151_D4;
  wire [0:0] CLBLM_R_X11Y151_SLICE_X15Y151_D5;
  wire [0:0] CLBLM_R_X11Y151_SLICE_X15Y151_D6;
  wire [0:0] CLBLM_R_X11Y151_SLICE_X15Y151_DO5;
  wire [0:0] CLBLM_R_X11Y151_SLICE_X15Y151_DO6;
  wire [0:0] CLBLM_R_X11Y151_SLICE_X15Y151_D_CY;
  wire [0:0] CLBLM_R_X11Y151_SLICE_X15Y151_D_XOR;
  wire [0:0] CLBLM_R_X11Y152_SLICE_X14Y152_A;
  wire [0:0] CLBLM_R_X11Y152_SLICE_X14Y152_A1;
  wire [0:0] CLBLM_R_X11Y152_SLICE_X14Y152_A2;
  wire [0:0] CLBLM_R_X11Y152_SLICE_X14Y152_A3;
  wire [0:0] CLBLM_R_X11Y152_SLICE_X14Y152_A4;
  wire [0:0] CLBLM_R_X11Y152_SLICE_X14Y152_A5;
  wire [0:0] CLBLM_R_X11Y152_SLICE_X14Y152_A6;
  wire [0:0] CLBLM_R_X11Y152_SLICE_X14Y152_AO5;
  wire [0:0] CLBLM_R_X11Y152_SLICE_X14Y152_AO6;
  wire [0:0] CLBLM_R_X11Y152_SLICE_X14Y152_A_CY;
  wire [0:0] CLBLM_R_X11Y152_SLICE_X14Y152_A_XOR;
  wire [0:0] CLBLM_R_X11Y152_SLICE_X14Y152_B;
  wire [0:0] CLBLM_R_X11Y152_SLICE_X14Y152_B1;
  wire [0:0] CLBLM_R_X11Y152_SLICE_X14Y152_B2;
  wire [0:0] CLBLM_R_X11Y152_SLICE_X14Y152_B3;
  wire [0:0] CLBLM_R_X11Y152_SLICE_X14Y152_B4;
  wire [0:0] CLBLM_R_X11Y152_SLICE_X14Y152_B5;
  wire [0:0] CLBLM_R_X11Y152_SLICE_X14Y152_B6;
  wire [0:0] CLBLM_R_X11Y152_SLICE_X14Y152_BO5;
  wire [0:0] CLBLM_R_X11Y152_SLICE_X14Y152_BO6;
  wire [0:0] CLBLM_R_X11Y152_SLICE_X14Y152_B_CY;
  wire [0:0] CLBLM_R_X11Y152_SLICE_X14Y152_B_XOR;
  wire [0:0] CLBLM_R_X11Y152_SLICE_X14Y152_C;
  wire [0:0] CLBLM_R_X11Y152_SLICE_X14Y152_C1;
  wire [0:0] CLBLM_R_X11Y152_SLICE_X14Y152_C2;
  wire [0:0] CLBLM_R_X11Y152_SLICE_X14Y152_C3;
  wire [0:0] CLBLM_R_X11Y152_SLICE_X14Y152_C4;
  wire [0:0] CLBLM_R_X11Y152_SLICE_X14Y152_C5;
  wire [0:0] CLBLM_R_X11Y152_SLICE_X14Y152_C6;
  wire [0:0] CLBLM_R_X11Y152_SLICE_X14Y152_CO5;
  wire [0:0] CLBLM_R_X11Y152_SLICE_X14Y152_CO6;
  wire [0:0] CLBLM_R_X11Y152_SLICE_X14Y152_C_CY;
  wire [0:0] CLBLM_R_X11Y152_SLICE_X14Y152_C_XOR;
  wire [0:0] CLBLM_R_X11Y152_SLICE_X14Y152_D;
  wire [0:0] CLBLM_R_X11Y152_SLICE_X14Y152_D1;
  wire [0:0] CLBLM_R_X11Y152_SLICE_X14Y152_D2;
  wire [0:0] CLBLM_R_X11Y152_SLICE_X14Y152_D3;
  wire [0:0] CLBLM_R_X11Y152_SLICE_X14Y152_D4;
  wire [0:0] CLBLM_R_X11Y152_SLICE_X14Y152_D5;
  wire [0:0] CLBLM_R_X11Y152_SLICE_X14Y152_D6;
  wire [0:0] CLBLM_R_X11Y152_SLICE_X14Y152_DO5;
  wire [0:0] CLBLM_R_X11Y152_SLICE_X14Y152_DO6;
  wire [0:0] CLBLM_R_X11Y152_SLICE_X14Y152_D_CY;
  wire [0:0] CLBLM_R_X11Y152_SLICE_X14Y152_D_XOR;
  wire [0:0] CLBLM_R_X11Y152_SLICE_X15Y152_A;
  wire [0:0] CLBLM_R_X11Y152_SLICE_X15Y152_A1;
  wire [0:0] CLBLM_R_X11Y152_SLICE_X15Y152_A2;
  wire [0:0] CLBLM_R_X11Y152_SLICE_X15Y152_A3;
  wire [0:0] CLBLM_R_X11Y152_SLICE_X15Y152_A4;
  wire [0:0] CLBLM_R_X11Y152_SLICE_X15Y152_A5;
  wire [0:0] CLBLM_R_X11Y152_SLICE_X15Y152_A5Q;
  wire [0:0] CLBLM_R_X11Y152_SLICE_X15Y152_A6;
  wire [0:0] CLBLM_R_X11Y152_SLICE_X15Y152_AMUX;
  wire [0:0] CLBLM_R_X11Y152_SLICE_X15Y152_AO5;
  wire [0:0] CLBLM_R_X11Y152_SLICE_X15Y152_AO6;
  wire [0:0] CLBLM_R_X11Y152_SLICE_X15Y152_AQ;
  wire [0:0] CLBLM_R_X11Y152_SLICE_X15Y152_A_CY;
  wire [0:0] CLBLM_R_X11Y152_SLICE_X15Y152_A_XOR;
  wire [0:0] CLBLM_R_X11Y152_SLICE_X15Y152_B;
  wire [0:0] CLBLM_R_X11Y152_SLICE_X15Y152_B1;
  wire [0:0] CLBLM_R_X11Y152_SLICE_X15Y152_B2;
  wire [0:0] CLBLM_R_X11Y152_SLICE_X15Y152_B3;
  wire [0:0] CLBLM_R_X11Y152_SLICE_X15Y152_B4;
  wire [0:0] CLBLM_R_X11Y152_SLICE_X15Y152_B5;
  wire [0:0] CLBLM_R_X11Y152_SLICE_X15Y152_B5Q;
  wire [0:0] CLBLM_R_X11Y152_SLICE_X15Y152_B6;
  wire [0:0] CLBLM_R_X11Y152_SLICE_X15Y152_BMUX;
  wire [0:0] CLBLM_R_X11Y152_SLICE_X15Y152_BO5;
  wire [0:0] CLBLM_R_X11Y152_SLICE_X15Y152_BO6;
  wire [0:0] CLBLM_R_X11Y152_SLICE_X15Y152_BQ;
  wire [0:0] CLBLM_R_X11Y152_SLICE_X15Y152_B_CY;
  wire [0:0] CLBLM_R_X11Y152_SLICE_X15Y152_B_XOR;
  wire [0:0] CLBLM_R_X11Y152_SLICE_X15Y152_C;
  wire [0:0] CLBLM_R_X11Y152_SLICE_X15Y152_C1;
  wire [0:0] CLBLM_R_X11Y152_SLICE_X15Y152_C2;
  wire [0:0] CLBLM_R_X11Y152_SLICE_X15Y152_C3;
  wire [0:0] CLBLM_R_X11Y152_SLICE_X15Y152_C4;
  wire [0:0] CLBLM_R_X11Y152_SLICE_X15Y152_C5;
  wire [0:0] CLBLM_R_X11Y152_SLICE_X15Y152_C6;
  wire [0:0] CLBLM_R_X11Y152_SLICE_X15Y152_CLK;
  wire [0:0] CLBLM_R_X11Y152_SLICE_X15Y152_CO5;
  wire [0:0] CLBLM_R_X11Y152_SLICE_X15Y152_CO6;
  wire [0:0] CLBLM_R_X11Y152_SLICE_X15Y152_CQ;
  wire [0:0] CLBLM_R_X11Y152_SLICE_X15Y152_C_CY;
  wire [0:0] CLBLM_R_X11Y152_SLICE_X15Y152_C_XOR;
  wire [0:0] CLBLM_R_X11Y152_SLICE_X15Y152_D;
  wire [0:0] CLBLM_R_X11Y152_SLICE_X15Y152_D1;
  wire [0:0] CLBLM_R_X11Y152_SLICE_X15Y152_D2;
  wire [0:0] CLBLM_R_X11Y152_SLICE_X15Y152_D3;
  wire [0:0] CLBLM_R_X11Y152_SLICE_X15Y152_D4;
  wire [0:0] CLBLM_R_X11Y152_SLICE_X15Y152_D5;
  wire [0:0] CLBLM_R_X11Y152_SLICE_X15Y152_D6;
  wire [0:0] CLBLM_R_X11Y152_SLICE_X15Y152_DO5;
  wire [0:0] CLBLM_R_X11Y152_SLICE_X15Y152_DO6;
  wire [0:0] CLBLM_R_X11Y152_SLICE_X15Y152_D_CY;
  wire [0:0] CLBLM_R_X11Y152_SLICE_X15Y152_D_XOR;
  wire [0:0] CLBLM_R_X11Y153_SLICE_X14Y153_A;
  wire [0:0] CLBLM_R_X11Y153_SLICE_X14Y153_A1;
  wire [0:0] CLBLM_R_X11Y153_SLICE_X14Y153_A2;
  wire [0:0] CLBLM_R_X11Y153_SLICE_X14Y153_A3;
  wire [0:0] CLBLM_R_X11Y153_SLICE_X14Y153_A4;
  wire [0:0] CLBLM_R_X11Y153_SLICE_X14Y153_A5;
  wire [0:0] CLBLM_R_X11Y153_SLICE_X14Y153_A5Q;
  wire [0:0] CLBLM_R_X11Y153_SLICE_X14Y153_A6;
  wire [0:0] CLBLM_R_X11Y153_SLICE_X14Y153_AMUX;
  wire [0:0] CLBLM_R_X11Y153_SLICE_X14Y153_AO5;
  wire [0:0] CLBLM_R_X11Y153_SLICE_X14Y153_AO6;
  wire [0:0] CLBLM_R_X11Y153_SLICE_X14Y153_AQ;
  wire [0:0] CLBLM_R_X11Y153_SLICE_X14Y153_A_CY;
  wire [0:0] CLBLM_R_X11Y153_SLICE_X14Y153_A_XOR;
  wire [0:0] CLBLM_R_X11Y153_SLICE_X14Y153_B;
  wire [0:0] CLBLM_R_X11Y153_SLICE_X14Y153_B1;
  wire [0:0] CLBLM_R_X11Y153_SLICE_X14Y153_B2;
  wire [0:0] CLBLM_R_X11Y153_SLICE_X14Y153_B3;
  wire [0:0] CLBLM_R_X11Y153_SLICE_X14Y153_B4;
  wire [0:0] CLBLM_R_X11Y153_SLICE_X14Y153_B5;
  wire [0:0] CLBLM_R_X11Y153_SLICE_X14Y153_B6;
  wire [0:0] CLBLM_R_X11Y153_SLICE_X14Y153_BO5;
  wire [0:0] CLBLM_R_X11Y153_SLICE_X14Y153_BO6;
  wire [0:0] CLBLM_R_X11Y153_SLICE_X14Y153_B_CY;
  wire [0:0] CLBLM_R_X11Y153_SLICE_X14Y153_B_XOR;
  wire [0:0] CLBLM_R_X11Y153_SLICE_X14Y153_C;
  wire [0:0] CLBLM_R_X11Y153_SLICE_X14Y153_C1;
  wire [0:0] CLBLM_R_X11Y153_SLICE_X14Y153_C2;
  wire [0:0] CLBLM_R_X11Y153_SLICE_X14Y153_C3;
  wire [0:0] CLBLM_R_X11Y153_SLICE_X14Y153_C4;
  wire [0:0] CLBLM_R_X11Y153_SLICE_X14Y153_C5;
  wire [0:0] CLBLM_R_X11Y153_SLICE_X14Y153_C6;
  wire [0:0] CLBLM_R_X11Y153_SLICE_X14Y153_CLK;
  wire [0:0] CLBLM_R_X11Y153_SLICE_X14Y153_CMUX;
  wire [0:0] CLBLM_R_X11Y153_SLICE_X14Y153_CO5;
  wire [0:0] CLBLM_R_X11Y153_SLICE_X14Y153_CO6;
  wire [0:0] CLBLM_R_X11Y153_SLICE_X14Y153_C_CY;
  wire [0:0] CLBLM_R_X11Y153_SLICE_X14Y153_C_XOR;
  wire [0:0] CLBLM_R_X11Y153_SLICE_X14Y153_D;
  wire [0:0] CLBLM_R_X11Y153_SLICE_X14Y153_D1;
  wire [0:0] CLBLM_R_X11Y153_SLICE_X14Y153_D2;
  wire [0:0] CLBLM_R_X11Y153_SLICE_X14Y153_D3;
  wire [0:0] CLBLM_R_X11Y153_SLICE_X14Y153_D4;
  wire [0:0] CLBLM_R_X11Y153_SLICE_X14Y153_D5;
  wire [0:0] CLBLM_R_X11Y153_SLICE_X14Y153_D6;
  wire [0:0] CLBLM_R_X11Y153_SLICE_X14Y153_DMUX;
  wire [0:0] CLBLM_R_X11Y153_SLICE_X14Y153_DO5;
  wire [0:0] CLBLM_R_X11Y153_SLICE_X14Y153_DO6;
  wire [0:0] CLBLM_R_X11Y153_SLICE_X14Y153_D_CY;
  wire [0:0] CLBLM_R_X11Y153_SLICE_X14Y153_D_XOR;
  wire [0:0] CLBLM_R_X11Y153_SLICE_X15Y153_A;
  wire [0:0] CLBLM_R_X11Y153_SLICE_X15Y153_A1;
  wire [0:0] CLBLM_R_X11Y153_SLICE_X15Y153_A2;
  wire [0:0] CLBLM_R_X11Y153_SLICE_X15Y153_A3;
  wire [0:0] CLBLM_R_X11Y153_SLICE_X15Y153_A4;
  wire [0:0] CLBLM_R_X11Y153_SLICE_X15Y153_A5;
  wire [0:0] CLBLM_R_X11Y153_SLICE_X15Y153_A6;
  wire [0:0] CLBLM_R_X11Y153_SLICE_X15Y153_AO5;
  wire [0:0] CLBLM_R_X11Y153_SLICE_X15Y153_AO6;
  wire [0:0] CLBLM_R_X11Y153_SLICE_X15Y153_AQ;
  wire [0:0] CLBLM_R_X11Y153_SLICE_X15Y153_A_CY;
  wire [0:0] CLBLM_R_X11Y153_SLICE_X15Y153_A_XOR;
  wire [0:0] CLBLM_R_X11Y153_SLICE_X15Y153_B;
  wire [0:0] CLBLM_R_X11Y153_SLICE_X15Y153_B1;
  wire [0:0] CLBLM_R_X11Y153_SLICE_X15Y153_B2;
  wire [0:0] CLBLM_R_X11Y153_SLICE_X15Y153_B3;
  wire [0:0] CLBLM_R_X11Y153_SLICE_X15Y153_B4;
  wire [0:0] CLBLM_R_X11Y153_SLICE_X15Y153_B5;
  wire [0:0] CLBLM_R_X11Y153_SLICE_X15Y153_B6;
  wire [0:0] CLBLM_R_X11Y153_SLICE_X15Y153_BMUX;
  wire [0:0] CLBLM_R_X11Y153_SLICE_X15Y153_BO5;
  wire [0:0] CLBLM_R_X11Y153_SLICE_X15Y153_BO6;
  wire [0:0] CLBLM_R_X11Y153_SLICE_X15Y153_B_CY;
  wire [0:0] CLBLM_R_X11Y153_SLICE_X15Y153_B_XOR;
  wire [0:0] CLBLM_R_X11Y153_SLICE_X15Y153_C;
  wire [0:0] CLBLM_R_X11Y153_SLICE_X15Y153_C1;
  wire [0:0] CLBLM_R_X11Y153_SLICE_X15Y153_C2;
  wire [0:0] CLBLM_R_X11Y153_SLICE_X15Y153_C3;
  wire [0:0] CLBLM_R_X11Y153_SLICE_X15Y153_C4;
  wire [0:0] CLBLM_R_X11Y153_SLICE_X15Y153_C5;
  wire [0:0] CLBLM_R_X11Y153_SLICE_X15Y153_C6;
  wire [0:0] CLBLM_R_X11Y153_SLICE_X15Y153_CLK;
  wire [0:0] CLBLM_R_X11Y153_SLICE_X15Y153_CO5;
  wire [0:0] CLBLM_R_X11Y153_SLICE_X15Y153_CO6;
  wire [0:0] CLBLM_R_X11Y153_SLICE_X15Y153_C_CY;
  wire [0:0] CLBLM_R_X11Y153_SLICE_X15Y153_C_XOR;
  wire [0:0] CLBLM_R_X11Y153_SLICE_X15Y153_D;
  wire [0:0] CLBLM_R_X11Y153_SLICE_X15Y153_D1;
  wire [0:0] CLBLM_R_X11Y153_SLICE_X15Y153_D2;
  wire [0:0] CLBLM_R_X11Y153_SLICE_X15Y153_D3;
  wire [0:0] CLBLM_R_X11Y153_SLICE_X15Y153_D4;
  wire [0:0] CLBLM_R_X11Y153_SLICE_X15Y153_D5;
  wire [0:0] CLBLM_R_X11Y153_SLICE_X15Y153_D6;
  wire [0:0] CLBLM_R_X11Y153_SLICE_X15Y153_DO5;
  wire [0:0] CLBLM_R_X11Y153_SLICE_X15Y153_DO6;
  wire [0:0] CLBLM_R_X11Y153_SLICE_X15Y153_D_CY;
  wire [0:0] CLBLM_R_X11Y153_SLICE_X15Y153_D_XOR;
  wire [0:0] CLBLM_R_X13Y146_SLICE_X18Y146_A;
  wire [0:0] CLBLM_R_X13Y146_SLICE_X18Y146_A1;
  wire [0:0] CLBLM_R_X13Y146_SLICE_X18Y146_A2;
  wire [0:0] CLBLM_R_X13Y146_SLICE_X18Y146_A3;
  wire [0:0] CLBLM_R_X13Y146_SLICE_X18Y146_A4;
  wire [0:0] CLBLM_R_X13Y146_SLICE_X18Y146_A5;
  wire [0:0] CLBLM_R_X13Y146_SLICE_X18Y146_A6;
  wire [0:0] CLBLM_R_X13Y146_SLICE_X18Y146_AMUX;
  wire [0:0] CLBLM_R_X13Y146_SLICE_X18Y146_AO5;
  wire [0:0] CLBLM_R_X13Y146_SLICE_X18Y146_AO6;
  wire [0:0] CLBLM_R_X13Y146_SLICE_X18Y146_A_CY;
  wire [0:0] CLBLM_R_X13Y146_SLICE_X18Y146_A_XOR;
  wire [0:0] CLBLM_R_X13Y146_SLICE_X18Y146_B;
  wire [0:0] CLBLM_R_X13Y146_SLICE_X18Y146_B1;
  wire [0:0] CLBLM_R_X13Y146_SLICE_X18Y146_B2;
  wire [0:0] CLBLM_R_X13Y146_SLICE_X18Y146_B3;
  wire [0:0] CLBLM_R_X13Y146_SLICE_X18Y146_B4;
  wire [0:0] CLBLM_R_X13Y146_SLICE_X18Y146_B5;
  wire [0:0] CLBLM_R_X13Y146_SLICE_X18Y146_B6;
  wire [0:0] CLBLM_R_X13Y146_SLICE_X18Y146_BO5;
  wire [0:0] CLBLM_R_X13Y146_SLICE_X18Y146_BO6;
  wire [0:0] CLBLM_R_X13Y146_SLICE_X18Y146_B_CY;
  wire [0:0] CLBLM_R_X13Y146_SLICE_X18Y146_B_XOR;
  wire [0:0] CLBLM_R_X13Y146_SLICE_X18Y146_C;
  wire [0:0] CLBLM_R_X13Y146_SLICE_X18Y146_C1;
  wire [0:0] CLBLM_R_X13Y146_SLICE_X18Y146_C2;
  wire [0:0] CLBLM_R_X13Y146_SLICE_X18Y146_C3;
  wire [0:0] CLBLM_R_X13Y146_SLICE_X18Y146_C4;
  wire [0:0] CLBLM_R_X13Y146_SLICE_X18Y146_C5;
  wire [0:0] CLBLM_R_X13Y146_SLICE_X18Y146_C6;
  wire [0:0] CLBLM_R_X13Y146_SLICE_X18Y146_CO5;
  wire [0:0] CLBLM_R_X13Y146_SLICE_X18Y146_CO6;
  wire [0:0] CLBLM_R_X13Y146_SLICE_X18Y146_C_CY;
  wire [0:0] CLBLM_R_X13Y146_SLICE_X18Y146_C_XOR;
  wire [0:0] CLBLM_R_X13Y146_SLICE_X18Y146_D;
  wire [0:0] CLBLM_R_X13Y146_SLICE_X18Y146_D1;
  wire [0:0] CLBLM_R_X13Y146_SLICE_X18Y146_D2;
  wire [0:0] CLBLM_R_X13Y146_SLICE_X18Y146_D3;
  wire [0:0] CLBLM_R_X13Y146_SLICE_X18Y146_D4;
  wire [0:0] CLBLM_R_X13Y146_SLICE_X18Y146_D5;
  wire [0:0] CLBLM_R_X13Y146_SLICE_X18Y146_D6;
  wire [0:0] CLBLM_R_X13Y146_SLICE_X18Y146_DO5;
  wire [0:0] CLBLM_R_X13Y146_SLICE_X18Y146_DO6;
  wire [0:0] CLBLM_R_X13Y146_SLICE_X18Y146_D_CY;
  wire [0:0] CLBLM_R_X13Y146_SLICE_X18Y146_D_XOR;
  wire [0:0] CLBLM_R_X13Y146_SLICE_X19Y146_A;
  wire [0:0] CLBLM_R_X13Y146_SLICE_X19Y146_A1;
  wire [0:0] CLBLM_R_X13Y146_SLICE_X19Y146_A2;
  wire [0:0] CLBLM_R_X13Y146_SLICE_X19Y146_A3;
  wire [0:0] CLBLM_R_X13Y146_SLICE_X19Y146_A4;
  wire [0:0] CLBLM_R_X13Y146_SLICE_X19Y146_A5;
  wire [0:0] CLBLM_R_X13Y146_SLICE_X19Y146_A6;
  wire [0:0] CLBLM_R_X13Y146_SLICE_X19Y146_AO5;
  wire [0:0] CLBLM_R_X13Y146_SLICE_X19Y146_AO6;
  wire [0:0] CLBLM_R_X13Y146_SLICE_X19Y146_A_CY;
  wire [0:0] CLBLM_R_X13Y146_SLICE_X19Y146_A_XOR;
  wire [0:0] CLBLM_R_X13Y146_SLICE_X19Y146_B;
  wire [0:0] CLBLM_R_X13Y146_SLICE_X19Y146_B1;
  wire [0:0] CLBLM_R_X13Y146_SLICE_X19Y146_B2;
  wire [0:0] CLBLM_R_X13Y146_SLICE_X19Y146_B3;
  wire [0:0] CLBLM_R_X13Y146_SLICE_X19Y146_B4;
  wire [0:0] CLBLM_R_X13Y146_SLICE_X19Y146_B5;
  wire [0:0] CLBLM_R_X13Y146_SLICE_X19Y146_B6;
  wire [0:0] CLBLM_R_X13Y146_SLICE_X19Y146_BO5;
  wire [0:0] CLBLM_R_X13Y146_SLICE_X19Y146_BO6;
  wire [0:0] CLBLM_R_X13Y146_SLICE_X19Y146_B_CY;
  wire [0:0] CLBLM_R_X13Y146_SLICE_X19Y146_B_XOR;
  wire [0:0] CLBLM_R_X13Y146_SLICE_X19Y146_C;
  wire [0:0] CLBLM_R_X13Y146_SLICE_X19Y146_C1;
  wire [0:0] CLBLM_R_X13Y146_SLICE_X19Y146_C2;
  wire [0:0] CLBLM_R_X13Y146_SLICE_X19Y146_C3;
  wire [0:0] CLBLM_R_X13Y146_SLICE_X19Y146_C4;
  wire [0:0] CLBLM_R_X13Y146_SLICE_X19Y146_C5;
  wire [0:0] CLBLM_R_X13Y146_SLICE_X19Y146_C6;
  wire [0:0] CLBLM_R_X13Y146_SLICE_X19Y146_CO5;
  wire [0:0] CLBLM_R_X13Y146_SLICE_X19Y146_CO6;
  wire [0:0] CLBLM_R_X13Y146_SLICE_X19Y146_C_CY;
  wire [0:0] CLBLM_R_X13Y146_SLICE_X19Y146_C_XOR;
  wire [0:0] CLBLM_R_X13Y146_SLICE_X19Y146_D;
  wire [0:0] CLBLM_R_X13Y146_SLICE_X19Y146_D1;
  wire [0:0] CLBLM_R_X13Y146_SLICE_X19Y146_D2;
  wire [0:0] CLBLM_R_X13Y146_SLICE_X19Y146_D3;
  wire [0:0] CLBLM_R_X13Y146_SLICE_X19Y146_D4;
  wire [0:0] CLBLM_R_X13Y146_SLICE_X19Y146_D5;
  wire [0:0] CLBLM_R_X13Y146_SLICE_X19Y146_D6;
  wire [0:0] CLBLM_R_X13Y146_SLICE_X19Y146_DO5;
  wire [0:0] CLBLM_R_X13Y146_SLICE_X19Y146_DO6;
  wire [0:0] CLBLM_R_X13Y146_SLICE_X19Y146_D_CY;
  wire [0:0] CLBLM_R_X13Y146_SLICE_X19Y146_D_XOR;
  wire [0:0] CLBLM_R_X13Y149_SLICE_X18Y149_A;
  wire [0:0] CLBLM_R_X13Y149_SLICE_X18Y149_A1;
  wire [0:0] CLBLM_R_X13Y149_SLICE_X18Y149_A2;
  wire [0:0] CLBLM_R_X13Y149_SLICE_X18Y149_A3;
  wire [0:0] CLBLM_R_X13Y149_SLICE_X18Y149_A4;
  wire [0:0] CLBLM_R_X13Y149_SLICE_X18Y149_A5;
  wire [0:0] CLBLM_R_X13Y149_SLICE_X18Y149_A6;
  wire [0:0] CLBLM_R_X13Y149_SLICE_X18Y149_AO5;
  wire [0:0] CLBLM_R_X13Y149_SLICE_X18Y149_AO6;
  wire [0:0] CLBLM_R_X13Y149_SLICE_X18Y149_A_CY;
  wire [0:0] CLBLM_R_X13Y149_SLICE_X18Y149_A_XOR;
  wire [0:0] CLBLM_R_X13Y149_SLICE_X18Y149_B;
  wire [0:0] CLBLM_R_X13Y149_SLICE_X18Y149_B1;
  wire [0:0] CLBLM_R_X13Y149_SLICE_X18Y149_B2;
  wire [0:0] CLBLM_R_X13Y149_SLICE_X18Y149_B3;
  wire [0:0] CLBLM_R_X13Y149_SLICE_X18Y149_B4;
  wire [0:0] CLBLM_R_X13Y149_SLICE_X18Y149_B5;
  wire [0:0] CLBLM_R_X13Y149_SLICE_X18Y149_B6;
  wire [0:0] CLBLM_R_X13Y149_SLICE_X18Y149_BO5;
  wire [0:0] CLBLM_R_X13Y149_SLICE_X18Y149_BO6;
  wire [0:0] CLBLM_R_X13Y149_SLICE_X18Y149_B_CY;
  wire [0:0] CLBLM_R_X13Y149_SLICE_X18Y149_B_XOR;
  wire [0:0] CLBLM_R_X13Y149_SLICE_X18Y149_C;
  wire [0:0] CLBLM_R_X13Y149_SLICE_X18Y149_C1;
  wire [0:0] CLBLM_R_X13Y149_SLICE_X18Y149_C2;
  wire [0:0] CLBLM_R_X13Y149_SLICE_X18Y149_C3;
  wire [0:0] CLBLM_R_X13Y149_SLICE_X18Y149_C4;
  wire [0:0] CLBLM_R_X13Y149_SLICE_X18Y149_C5;
  wire [0:0] CLBLM_R_X13Y149_SLICE_X18Y149_C6;
  wire [0:0] CLBLM_R_X13Y149_SLICE_X18Y149_CO5;
  wire [0:0] CLBLM_R_X13Y149_SLICE_X18Y149_CO6;
  wire [0:0] CLBLM_R_X13Y149_SLICE_X18Y149_C_CY;
  wire [0:0] CLBLM_R_X13Y149_SLICE_X18Y149_C_XOR;
  wire [0:0] CLBLM_R_X13Y149_SLICE_X18Y149_D;
  wire [0:0] CLBLM_R_X13Y149_SLICE_X18Y149_D1;
  wire [0:0] CLBLM_R_X13Y149_SLICE_X18Y149_D2;
  wire [0:0] CLBLM_R_X13Y149_SLICE_X18Y149_D3;
  wire [0:0] CLBLM_R_X13Y149_SLICE_X18Y149_D4;
  wire [0:0] CLBLM_R_X13Y149_SLICE_X18Y149_D5;
  wire [0:0] CLBLM_R_X13Y149_SLICE_X18Y149_D6;
  wire [0:0] CLBLM_R_X13Y149_SLICE_X18Y149_DO5;
  wire [0:0] CLBLM_R_X13Y149_SLICE_X18Y149_DO6;
  wire [0:0] CLBLM_R_X13Y149_SLICE_X18Y149_D_CY;
  wire [0:0] CLBLM_R_X13Y149_SLICE_X18Y149_D_XOR;
  wire [0:0] CLBLM_R_X13Y149_SLICE_X19Y149_A;
  wire [0:0] CLBLM_R_X13Y149_SLICE_X19Y149_A1;
  wire [0:0] CLBLM_R_X13Y149_SLICE_X19Y149_A2;
  wire [0:0] CLBLM_R_X13Y149_SLICE_X19Y149_A3;
  wire [0:0] CLBLM_R_X13Y149_SLICE_X19Y149_A4;
  wire [0:0] CLBLM_R_X13Y149_SLICE_X19Y149_A5;
  wire [0:0] CLBLM_R_X13Y149_SLICE_X19Y149_A6;
  wire [0:0] CLBLM_R_X13Y149_SLICE_X19Y149_AO5;
  wire [0:0] CLBLM_R_X13Y149_SLICE_X19Y149_AO6;
  wire [0:0] CLBLM_R_X13Y149_SLICE_X19Y149_A_CY;
  wire [0:0] CLBLM_R_X13Y149_SLICE_X19Y149_A_XOR;
  wire [0:0] CLBLM_R_X13Y149_SLICE_X19Y149_B;
  wire [0:0] CLBLM_R_X13Y149_SLICE_X19Y149_B1;
  wire [0:0] CLBLM_R_X13Y149_SLICE_X19Y149_B2;
  wire [0:0] CLBLM_R_X13Y149_SLICE_X19Y149_B3;
  wire [0:0] CLBLM_R_X13Y149_SLICE_X19Y149_B4;
  wire [0:0] CLBLM_R_X13Y149_SLICE_X19Y149_B5;
  wire [0:0] CLBLM_R_X13Y149_SLICE_X19Y149_B6;
  wire [0:0] CLBLM_R_X13Y149_SLICE_X19Y149_BO5;
  wire [0:0] CLBLM_R_X13Y149_SLICE_X19Y149_BO6;
  wire [0:0] CLBLM_R_X13Y149_SLICE_X19Y149_B_CY;
  wire [0:0] CLBLM_R_X13Y149_SLICE_X19Y149_B_XOR;
  wire [0:0] CLBLM_R_X13Y149_SLICE_X19Y149_C;
  wire [0:0] CLBLM_R_X13Y149_SLICE_X19Y149_C1;
  wire [0:0] CLBLM_R_X13Y149_SLICE_X19Y149_C2;
  wire [0:0] CLBLM_R_X13Y149_SLICE_X19Y149_C3;
  wire [0:0] CLBLM_R_X13Y149_SLICE_X19Y149_C4;
  wire [0:0] CLBLM_R_X13Y149_SLICE_X19Y149_C5;
  wire [0:0] CLBLM_R_X13Y149_SLICE_X19Y149_C6;
  wire [0:0] CLBLM_R_X13Y149_SLICE_X19Y149_CO5;
  wire [0:0] CLBLM_R_X13Y149_SLICE_X19Y149_CO6;
  wire [0:0] CLBLM_R_X13Y149_SLICE_X19Y149_C_CY;
  wire [0:0] CLBLM_R_X13Y149_SLICE_X19Y149_C_XOR;
  wire [0:0] CLBLM_R_X13Y149_SLICE_X19Y149_D;
  wire [0:0] CLBLM_R_X13Y149_SLICE_X19Y149_D1;
  wire [0:0] CLBLM_R_X13Y149_SLICE_X19Y149_D2;
  wire [0:0] CLBLM_R_X13Y149_SLICE_X19Y149_D3;
  wire [0:0] CLBLM_R_X13Y149_SLICE_X19Y149_D4;
  wire [0:0] CLBLM_R_X13Y149_SLICE_X19Y149_D5;
  wire [0:0] CLBLM_R_X13Y149_SLICE_X19Y149_D6;
  wire [0:0] CLBLM_R_X13Y149_SLICE_X19Y149_DO5;
  wire [0:0] CLBLM_R_X13Y149_SLICE_X19Y149_DO6;
  wire [0:0] CLBLM_R_X13Y149_SLICE_X19Y149_D_CY;
  wire [0:0] CLBLM_R_X13Y149_SLICE_X19Y149_D_XOR;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X2Y142_A;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X2Y142_A1;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X2Y142_A2;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X2Y142_A3;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X2Y142_A4;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X2Y142_A5;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X2Y142_A6;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X2Y142_AO5;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X2Y142_AO6;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X2Y142_AQ;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X2Y142_A_CY;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X2Y142_A_XOR;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X2Y142_B;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X2Y142_B1;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X2Y142_B2;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X2Y142_B3;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X2Y142_B4;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X2Y142_B5;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X2Y142_B6;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X2Y142_BMUX;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X2Y142_BO5;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X2Y142_BO6;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X2Y142_B_CY;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X2Y142_B_XOR;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X2Y142_C;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X2Y142_C1;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X2Y142_C2;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X2Y142_C3;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X2Y142_C4;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X2Y142_C5;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X2Y142_C6;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X2Y142_CLK;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X2Y142_CO5;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X2Y142_CO6;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X2Y142_C_CY;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X2Y142_C_XOR;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X2Y142_D;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X2Y142_D1;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X2Y142_D2;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X2Y142_D3;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X2Y142_D4;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X2Y142_D5;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X2Y142_D6;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X2Y142_DO5;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X2Y142_DO6;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X2Y142_D_CY;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X2Y142_D_XOR;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X3Y142_A;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X3Y142_A1;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X3Y142_A2;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X3Y142_A3;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X3Y142_A4;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X3Y142_A5;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X3Y142_A6;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X3Y142_AO5;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X3Y142_AO6;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X3Y142_AQ;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X3Y142_A_CY;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X3Y142_A_XOR;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X3Y142_B;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X3Y142_B1;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X3Y142_B2;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X3Y142_B3;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X3Y142_B4;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X3Y142_B5;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X3Y142_B6;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X3Y142_BO5;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X3Y142_BO6;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X3Y142_B_CY;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X3Y142_B_XOR;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X3Y142_C;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X3Y142_C1;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X3Y142_C2;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X3Y142_C3;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X3Y142_C4;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X3Y142_C5;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X3Y142_C6;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X3Y142_CLK;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X3Y142_CO5;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X3Y142_CO6;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X3Y142_C_CY;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X3Y142_C_XOR;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X3Y142_D;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X3Y142_D1;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X3Y142_D2;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X3Y142_D3;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X3Y142_D4;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X3Y142_D5;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X3Y142_D6;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X3Y142_DO5;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X3Y142_DO6;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X3Y142_D_CY;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X3Y142_D_XOR;
  wire [0:0] CLBLM_R_X3Y143_SLICE_X2Y143_A;
  wire [0:0] CLBLM_R_X3Y143_SLICE_X2Y143_A1;
  wire [0:0] CLBLM_R_X3Y143_SLICE_X2Y143_A2;
  wire [0:0] CLBLM_R_X3Y143_SLICE_X2Y143_A3;
  wire [0:0] CLBLM_R_X3Y143_SLICE_X2Y143_A4;
  wire [0:0] CLBLM_R_X3Y143_SLICE_X2Y143_A5;
  wire [0:0] CLBLM_R_X3Y143_SLICE_X2Y143_A5Q;
  wire [0:0] CLBLM_R_X3Y143_SLICE_X2Y143_A6;
  wire [0:0] CLBLM_R_X3Y143_SLICE_X2Y143_AMUX;
  wire [0:0] CLBLM_R_X3Y143_SLICE_X2Y143_AO5;
  wire [0:0] CLBLM_R_X3Y143_SLICE_X2Y143_AO6;
  wire [0:0] CLBLM_R_X3Y143_SLICE_X2Y143_AQ;
  wire [0:0] CLBLM_R_X3Y143_SLICE_X2Y143_AX;
  wire [0:0] CLBLM_R_X3Y143_SLICE_X2Y143_A_CY;
  wire [0:0] CLBLM_R_X3Y143_SLICE_X2Y143_A_XOR;
  wire [0:0] CLBLM_R_X3Y143_SLICE_X2Y143_B;
  wire [0:0] CLBLM_R_X3Y143_SLICE_X2Y143_B1;
  wire [0:0] CLBLM_R_X3Y143_SLICE_X2Y143_B2;
  wire [0:0] CLBLM_R_X3Y143_SLICE_X2Y143_B3;
  wire [0:0] CLBLM_R_X3Y143_SLICE_X2Y143_B4;
  wire [0:0] CLBLM_R_X3Y143_SLICE_X2Y143_B5;
  wire [0:0] CLBLM_R_X3Y143_SLICE_X2Y143_B6;
  wire [0:0] CLBLM_R_X3Y143_SLICE_X2Y143_BMUX;
  wire [0:0] CLBLM_R_X3Y143_SLICE_X2Y143_BO5;
  wire [0:0] CLBLM_R_X3Y143_SLICE_X2Y143_BO6;
  wire [0:0] CLBLM_R_X3Y143_SLICE_X2Y143_B_CY;
  wire [0:0] CLBLM_R_X3Y143_SLICE_X2Y143_B_XOR;
  wire [0:0] CLBLM_R_X3Y143_SLICE_X2Y143_C;
  wire [0:0] CLBLM_R_X3Y143_SLICE_X2Y143_C1;
  wire [0:0] CLBLM_R_X3Y143_SLICE_X2Y143_C2;
  wire [0:0] CLBLM_R_X3Y143_SLICE_X2Y143_C3;
  wire [0:0] CLBLM_R_X3Y143_SLICE_X2Y143_C4;
  wire [0:0] CLBLM_R_X3Y143_SLICE_X2Y143_C5;
  wire [0:0] CLBLM_R_X3Y143_SLICE_X2Y143_C6;
  wire [0:0] CLBLM_R_X3Y143_SLICE_X2Y143_CLK;
  wire [0:0] CLBLM_R_X3Y143_SLICE_X2Y143_CMUX;
  wire [0:0] CLBLM_R_X3Y143_SLICE_X2Y143_CO5;
  wire [0:0] CLBLM_R_X3Y143_SLICE_X2Y143_CO6;
  wire [0:0] CLBLM_R_X3Y143_SLICE_X2Y143_C_CY;
  wire [0:0] CLBLM_R_X3Y143_SLICE_X2Y143_C_XOR;
  wire [0:0] CLBLM_R_X3Y143_SLICE_X2Y143_D;
  wire [0:0] CLBLM_R_X3Y143_SLICE_X2Y143_D1;
  wire [0:0] CLBLM_R_X3Y143_SLICE_X2Y143_D2;
  wire [0:0] CLBLM_R_X3Y143_SLICE_X2Y143_D3;
  wire [0:0] CLBLM_R_X3Y143_SLICE_X2Y143_D4;
  wire [0:0] CLBLM_R_X3Y143_SLICE_X2Y143_D5;
  wire [0:0] CLBLM_R_X3Y143_SLICE_X2Y143_D6;
  wire [0:0] CLBLM_R_X3Y143_SLICE_X2Y143_DO5;
  wire [0:0] CLBLM_R_X3Y143_SLICE_X2Y143_DO6;
  wire [0:0] CLBLM_R_X3Y143_SLICE_X2Y143_D_CY;
  wire [0:0] CLBLM_R_X3Y143_SLICE_X2Y143_D_XOR;
  wire [0:0] CLBLM_R_X3Y143_SLICE_X3Y143_A;
  wire [0:0] CLBLM_R_X3Y143_SLICE_X3Y143_A1;
  wire [0:0] CLBLM_R_X3Y143_SLICE_X3Y143_A2;
  wire [0:0] CLBLM_R_X3Y143_SLICE_X3Y143_A3;
  wire [0:0] CLBLM_R_X3Y143_SLICE_X3Y143_A4;
  wire [0:0] CLBLM_R_X3Y143_SLICE_X3Y143_A5;
  wire [0:0] CLBLM_R_X3Y143_SLICE_X3Y143_A6;
  wire [0:0] CLBLM_R_X3Y143_SLICE_X3Y143_AO5;
  wire [0:0] CLBLM_R_X3Y143_SLICE_X3Y143_AO6;
  wire [0:0] CLBLM_R_X3Y143_SLICE_X3Y143_AQ;
  wire [0:0] CLBLM_R_X3Y143_SLICE_X3Y143_A_CY;
  wire [0:0] CLBLM_R_X3Y143_SLICE_X3Y143_A_XOR;
  wire [0:0] CLBLM_R_X3Y143_SLICE_X3Y143_B;
  wire [0:0] CLBLM_R_X3Y143_SLICE_X3Y143_B1;
  wire [0:0] CLBLM_R_X3Y143_SLICE_X3Y143_B2;
  wire [0:0] CLBLM_R_X3Y143_SLICE_X3Y143_B3;
  wire [0:0] CLBLM_R_X3Y143_SLICE_X3Y143_B4;
  wire [0:0] CLBLM_R_X3Y143_SLICE_X3Y143_B5;
  wire [0:0] CLBLM_R_X3Y143_SLICE_X3Y143_B6;
  wire [0:0] CLBLM_R_X3Y143_SLICE_X3Y143_BO5;
  wire [0:0] CLBLM_R_X3Y143_SLICE_X3Y143_BO6;
  wire [0:0] CLBLM_R_X3Y143_SLICE_X3Y143_BQ;
  wire [0:0] CLBLM_R_X3Y143_SLICE_X3Y143_B_CY;
  wire [0:0] CLBLM_R_X3Y143_SLICE_X3Y143_B_XOR;
  wire [0:0] CLBLM_R_X3Y143_SLICE_X3Y143_C;
  wire [0:0] CLBLM_R_X3Y143_SLICE_X3Y143_C1;
  wire [0:0] CLBLM_R_X3Y143_SLICE_X3Y143_C2;
  wire [0:0] CLBLM_R_X3Y143_SLICE_X3Y143_C3;
  wire [0:0] CLBLM_R_X3Y143_SLICE_X3Y143_C4;
  wire [0:0] CLBLM_R_X3Y143_SLICE_X3Y143_C5;
  wire [0:0] CLBLM_R_X3Y143_SLICE_X3Y143_C5Q;
  wire [0:0] CLBLM_R_X3Y143_SLICE_X3Y143_C6;
  wire [0:0] CLBLM_R_X3Y143_SLICE_X3Y143_CLK;
  wire [0:0] CLBLM_R_X3Y143_SLICE_X3Y143_CMUX;
  wire [0:0] CLBLM_R_X3Y143_SLICE_X3Y143_CO5;
  wire [0:0] CLBLM_R_X3Y143_SLICE_X3Y143_CO6;
  wire [0:0] CLBLM_R_X3Y143_SLICE_X3Y143_CQ;
  wire [0:0] CLBLM_R_X3Y143_SLICE_X3Y143_C_CY;
  wire [0:0] CLBLM_R_X3Y143_SLICE_X3Y143_C_XOR;
  wire [0:0] CLBLM_R_X3Y143_SLICE_X3Y143_D;
  wire [0:0] CLBLM_R_X3Y143_SLICE_X3Y143_D1;
  wire [0:0] CLBLM_R_X3Y143_SLICE_X3Y143_D2;
  wire [0:0] CLBLM_R_X3Y143_SLICE_X3Y143_D3;
  wire [0:0] CLBLM_R_X3Y143_SLICE_X3Y143_D4;
  wire [0:0] CLBLM_R_X3Y143_SLICE_X3Y143_D5;
  wire [0:0] CLBLM_R_X3Y143_SLICE_X3Y143_D6;
  wire [0:0] CLBLM_R_X3Y143_SLICE_X3Y143_DO5;
  wire [0:0] CLBLM_R_X3Y143_SLICE_X3Y143_DO6;
  wire [0:0] CLBLM_R_X3Y143_SLICE_X3Y143_D_CY;
  wire [0:0] CLBLM_R_X3Y143_SLICE_X3Y143_D_XOR;
  wire [0:0] CLBLM_R_X3Y144_SLICE_X2Y144_A;
  wire [0:0] CLBLM_R_X3Y144_SLICE_X2Y144_A1;
  wire [0:0] CLBLM_R_X3Y144_SLICE_X2Y144_A2;
  wire [0:0] CLBLM_R_X3Y144_SLICE_X2Y144_A3;
  wire [0:0] CLBLM_R_X3Y144_SLICE_X2Y144_A4;
  wire [0:0] CLBLM_R_X3Y144_SLICE_X2Y144_A5;
  wire [0:0] CLBLM_R_X3Y144_SLICE_X2Y144_A6;
  wire [0:0] CLBLM_R_X3Y144_SLICE_X2Y144_AMUX;
  wire [0:0] CLBLM_R_X3Y144_SLICE_X2Y144_AO5;
  wire [0:0] CLBLM_R_X3Y144_SLICE_X2Y144_AO6;
  wire [0:0] CLBLM_R_X3Y144_SLICE_X2Y144_AQ;
  wire [0:0] CLBLM_R_X3Y144_SLICE_X2Y144_AX;
  wire [0:0] CLBLM_R_X3Y144_SLICE_X2Y144_A_CY;
  wire [0:0] CLBLM_R_X3Y144_SLICE_X2Y144_A_XOR;
  wire [0:0] CLBLM_R_X3Y144_SLICE_X2Y144_B;
  wire [0:0] CLBLM_R_X3Y144_SLICE_X2Y144_B1;
  wire [0:0] CLBLM_R_X3Y144_SLICE_X2Y144_B2;
  wire [0:0] CLBLM_R_X3Y144_SLICE_X2Y144_B3;
  wire [0:0] CLBLM_R_X3Y144_SLICE_X2Y144_B4;
  wire [0:0] CLBLM_R_X3Y144_SLICE_X2Y144_B5;
  wire [0:0] CLBLM_R_X3Y144_SLICE_X2Y144_B6;
  wire [0:0] CLBLM_R_X3Y144_SLICE_X2Y144_BMUX;
  wire [0:0] CLBLM_R_X3Y144_SLICE_X2Y144_BO5;
  wire [0:0] CLBLM_R_X3Y144_SLICE_X2Y144_BO6;
  wire [0:0] CLBLM_R_X3Y144_SLICE_X2Y144_B_CY;
  wire [0:0] CLBLM_R_X3Y144_SLICE_X2Y144_B_XOR;
  wire [0:0] CLBLM_R_X3Y144_SLICE_X2Y144_C;
  wire [0:0] CLBLM_R_X3Y144_SLICE_X2Y144_C1;
  wire [0:0] CLBLM_R_X3Y144_SLICE_X2Y144_C2;
  wire [0:0] CLBLM_R_X3Y144_SLICE_X2Y144_C3;
  wire [0:0] CLBLM_R_X3Y144_SLICE_X2Y144_C4;
  wire [0:0] CLBLM_R_X3Y144_SLICE_X2Y144_C5;
  wire [0:0] CLBLM_R_X3Y144_SLICE_X2Y144_C6;
  wire [0:0] CLBLM_R_X3Y144_SLICE_X2Y144_CLK;
  wire [0:0] CLBLM_R_X3Y144_SLICE_X2Y144_CO5;
  wire [0:0] CLBLM_R_X3Y144_SLICE_X2Y144_CO6;
  wire [0:0] CLBLM_R_X3Y144_SLICE_X2Y144_C_CY;
  wire [0:0] CLBLM_R_X3Y144_SLICE_X2Y144_C_XOR;
  wire [0:0] CLBLM_R_X3Y144_SLICE_X2Y144_D;
  wire [0:0] CLBLM_R_X3Y144_SLICE_X2Y144_D1;
  wire [0:0] CLBLM_R_X3Y144_SLICE_X2Y144_D2;
  wire [0:0] CLBLM_R_X3Y144_SLICE_X2Y144_D3;
  wire [0:0] CLBLM_R_X3Y144_SLICE_X2Y144_D4;
  wire [0:0] CLBLM_R_X3Y144_SLICE_X2Y144_D5;
  wire [0:0] CLBLM_R_X3Y144_SLICE_X2Y144_D6;
  wire [0:0] CLBLM_R_X3Y144_SLICE_X2Y144_DO5;
  wire [0:0] CLBLM_R_X3Y144_SLICE_X2Y144_DO6;
  wire [0:0] CLBLM_R_X3Y144_SLICE_X2Y144_D_CY;
  wire [0:0] CLBLM_R_X3Y144_SLICE_X2Y144_D_XOR;
  wire [0:0] CLBLM_R_X3Y144_SLICE_X3Y144_A;
  wire [0:0] CLBLM_R_X3Y144_SLICE_X3Y144_A1;
  wire [0:0] CLBLM_R_X3Y144_SLICE_X3Y144_A2;
  wire [0:0] CLBLM_R_X3Y144_SLICE_X3Y144_A3;
  wire [0:0] CLBLM_R_X3Y144_SLICE_X3Y144_A4;
  wire [0:0] CLBLM_R_X3Y144_SLICE_X3Y144_A5;
  wire [0:0] CLBLM_R_X3Y144_SLICE_X3Y144_A6;
  wire [0:0] CLBLM_R_X3Y144_SLICE_X3Y144_AO5;
  wire [0:0] CLBLM_R_X3Y144_SLICE_X3Y144_AO6;
  wire [0:0] CLBLM_R_X3Y144_SLICE_X3Y144_AQ;
  wire [0:0] CLBLM_R_X3Y144_SLICE_X3Y144_A_CY;
  wire [0:0] CLBLM_R_X3Y144_SLICE_X3Y144_A_XOR;
  wire [0:0] CLBLM_R_X3Y144_SLICE_X3Y144_B;
  wire [0:0] CLBLM_R_X3Y144_SLICE_X3Y144_B1;
  wire [0:0] CLBLM_R_X3Y144_SLICE_X3Y144_B2;
  wire [0:0] CLBLM_R_X3Y144_SLICE_X3Y144_B3;
  wire [0:0] CLBLM_R_X3Y144_SLICE_X3Y144_B4;
  wire [0:0] CLBLM_R_X3Y144_SLICE_X3Y144_B5;
  wire [0:0] CLBLM_R_X3Y144_SLICE_X3Y144_B6;
  wire [0:0] CLBLM_R_X3Y144_SLICE_X3Y144_BO5;
  wire [0:0] CLBLM_R_X3Y144_SLICE_X3Y144_BO6;
  wire [0:0] CLBLM_R_X3Y144_SLICE_X3Y144_B_CY;
  wire [0:0] CLBLM_R_X3Y144_SLICE_X3Y144_B_XOR;
  wire [0:0] CLBLM_R_X3Y144_SLICE_X3Y144_C;
  wire [0:0] CLBLM_R_X3Y144_SLICE_X3Y144_C1;
  wire [0:0] CLBLM_R_X3Y144_SLICE_X3Y144_C2;
  wire [0:0] CLBLM_R_X3Y144_SLICE_X3Y144_C3;
  wire [0:0] CLBLM_R_X3Y144_SLICE_X3Y144_C4;
  wire [0:0] CLBLM_R_X3Y144_SLICE_X3Y144_C5;
  wire [0:0] CLBLM_R_X3Y144_SLICE_X3Y144_C6;
  wire [0:0] CLBLM_R_X3Y144_SLICE_X3Y144_CLK;
  wire [0:0] CLBLM_R_X3Y144_SLICE_X3Y144_CO5;
  wire [0:0] CLBLM_R_X3Y144_SLICE_X3Y144_CO6;
  wire [0:0] CLBLM_R_X3Y144_SLICE_X3Y144_C_CY;
  wire [0:0] CLBLM_R_X3Y144_SLICE_X3Y144_C_XOR;
  wire [0:0] CLBLM_R_X3Y144_SLICE_X3Y144_D;
  wire [0:0] CLBLM_R_X3Y144_SLICE_X3Y144_D1;
  wire [0:0] CLBLM_R_X3Y144_SLICE_X3Y144_D2;
  wire [0:0] CLBLM_R_X3Y144_SLICE_X3Y144_D3;
  wire [0:0] CLBLM_R_X3Y144_SLICE_X3Y144_D4;
  wire [0:0] CLBLM_R_X3Y144_SLICE_X3Y144_D5;
  wire [0:0] CLBLM_R_X3Y144_SLICE_X3Y144_D6;
  wire [0:0] CLBLM_R_X3Y144_SLICE_X3Y144_DO5;
  wire [0:0] CLBLM_R_X3Y144_SLICE_X3Y144_DO6;
  wire [0:0] CLBLM_R_X3Y144_SLICE_X3Y144_D_CY;
  wire [0:0] CLBLM_R_X3Y144_SLICE_X3Y144_D_XOR;
  wire [0:0] CLBLM_R_X3Y145_SLICE_X2Y145_A;
  wire [0:0] CLBLM_R_X3Y145_SLICE_X2Y145_A1;
  wire [0:0] CLBLM_R_X3Y145_SLICE_X2Y145_A2;
  wire [0:0] CLBLM_R_X3Y145_SLICE_X2Y145_A3;
  wire [0:0] CLBLM_R_X3Y145_SLICE_X2Y145_A4;
  wire [0:0] CLBLM_R_X3Y145_SLICE_X2Y145_A5;
  wire [0:0] CLBLM_R_X3Y145_SLICE_X2Y145_A6;
  wire [0:0] CLBLM_R_X3Y145_SLICE_X2Y145_AO5;
  wire [0:0] CLBLM_R_X3Y145_SLICE_X2Y145_AO6;
  wire [0:0] CLBLM_R_X3Y145_SLICE_X2Y145_AQ;
  wire [0:0] CLBLM_R_X3Y145_SLICE_X2Y145_A_CY;
  wire [0:0] CLBLM_R_X3Y145_SLICE_X2Y145_A_XOR;
  wire [0:0] CLBLM_R_X3Y145_SLICE_X2Y145_B;
  wire [0:0] CLBLM_R_X3Y145_SLICE_X2Y145_B1;
  wire [0:0] CLBLM_R_X3Y145_SLICE_X2Y145_B2;
  wire [0:0] CLBLM_R_X3Y145_SLICE_X2Y145_B3;
  wire [0:0] CLBLM_R_X3Y145_SLICE_X2Y145_B4;
  wire [0:0] CLBLM_R_X3Y145_SLICE_X2Y145_B5;
  wire [0:0] CLBLM_R_X3Y145_SLICE_X2Y145_B5Q;
  wire [0:0] CLBLM_R_X3Y145_SLICE_X2Y145_B6;
  wire [0:0] CLBLM_R_X3Y145_SLICE_X2Y145_BMUX;
  wire [0:0] CLBLM_R_X3Y145_SLICE_X2Y145_BO5;
  wire [0:0] CLBLM_R_X3Y145_SLICE_X2Y145_BO6;
  wire [0:0] CLBLM_R_X3Y145_SLICE_X2Y145_BQ;
  wire [0:0] CLBLM_R_X3Y145_SLICE_X2Y145_B_CY;
  wire [0:0] CLBLM_R_X3Y145_SLICE_X2Y145_B_XOR;
  wire [0:0] CLBLM_R_X3Y145_SLICE_X2Y145_C;
  wire [0:0] CLBLM_R_X3Y145_SLICE_X2Y145_C1;
  wire [0:0] CLBLM_R_X3Y145_SLICE_X2Y145_C2;
  wire [0:0] CLBLM_R_X3Y145_SLICE_X2Y145_C3;
  wire [0:0] CLBLM_R_X3Y145_SLICE_X2Y145_C4;
  wire [0:0] CLBLM_R_X3Y145_SLICE_X2Y145_C5;
  wire [0:0] CLBLM_R_X3Y145_SLICE_X2Y145_C5Q;
  wire [0:0] CLBLM_R_X3Y145_SLICE_X2Y145_C6;
  wire [0:0] CLBLM_R_X3Y145_SLICE_X2Y145_CLK;
  wire [0:0] CLBLM_R_X3Y145_SLICE_X2Y145_CMUX;
  wire [0:0] CLBLM_R_X3Y145_SLICE_X2Y145_CO5;
  wire [0:0] CLBLM_R_X3Y145_SLICE_X2Y145_CO6;
  wire [0:0] CLBLM_R_X3Y145_SLICE_X2Y145_CQ;
  wire [0:0] CLBLM_R_X3Y145_SLICE_X2Y145_C_CY;
  wire [0:0] CLBLM_R_X3Y145_SLICE_X2Y145_C_XOR;
  wire [0:0] CLBLM_R_X3Y145_SLICE_X2Y145_D;
  wire [0:0] CLBLM_R_X3Y145_SLICE_X2Y145_D1;
  wire [0:0] CLBLM_R_X3Y145_SLICE_X2Y145_D2;
  wire [0:0] CLBLM_R_X3Y145_SLICE_X2Y145_D3;
  wire [0:0] CLBLM_R_X3Y145_SLICE_X2Y145_D4;
  wire [0:0] CLBLM_R_X3Y145_SLICE_X2Y145_D5;
  wire [0:0] CLBLM_R_X3Y145_SLICE_X2Y145_D6;
  wire [0:0] CLBLM_R_X3Y145_SLICE_X2Y145_DO5;
  wire [0:0] CLBLM_R_X3Y145_SLICE_X2Y145_DO6;
  wire [0:0] CLBLM_R_X3Y145_SLICE_X2Y145_D_CY;
  wire [0:0] CLBLM_R_X3Y145_SLICE_X2Y145_D_XOR;
  wire [0:0] CLBLM_R_X3Y145_SLICE_X3Y145_A;
  wire [0:0] CLBLM_R_X3Y145_SLICE_X3Y145_A1;
  wire [0:0] CLBLM_R_X3Y145_SLICE_X3Y145_A2;
  wire [0:0] CLBLM_R_X3Y145_SLICE_X3Y145_A3;
  wire [0:0] CLBLM_R_X3Y145_SLICE_X3Y145_A4;
  wire [0:0] CLBLM_R_X3Y145_SLICE_X3Y145_A5;
  wire [0:0] CLBLM_R_X3Y145_SLICE_X3Y145_A6;
  wire [0:0] CLBLM_R_X3Y145_SLICE_X3Y145_AO5;
  wire [0:0] CLBLM_R_X3Y145_SLICE_X3Y145_AO6;
  wire [0:0] CLBLM_R_X3Y145_SLICE_X3Y145_AQ;
  wire [0:0] CLBLM_R_X3Y145_SLICE_X3Y145_A_CY;
  wire [0:0] CLBLM_R_X3Y145_SLICE_X3Y145_A_XOR;
  wire [0:0] CLBLM_R_X3Y145_SLICE_X3Y145_B;
  wire [0:0] CLBLM_R_X3Y145_SLICE_X3Y145_B1;
  wire [0:0] CLBLM_R_X3Y145_SLICE_X3Y145_B2;
  wire [0:0] CLBLM_R_X3Y145_SLICE_X3Y145_B3;
  wire [0:0] CLBLM_R_X3Y145_SLICE_X3Y145_B4;
  wire [0:0] CLBLM_R_X3Y145_SLICE_X3Y145_B5;
  wire [0:0] CLBLM_R_X3Y145_SLICE_X3Y145_B6;
  wire [0:0] CLBLM_R_X3Y145_SLICE_X3Y145_BO5;
  wire [0:0] CLBLM_R_X3Y145_SLICE_X3Y145_BO6;
  wire [0:0] CLBLM_R_X3Y145_SLICE_X3Y145_BQ;
  wire [0:0] CLBLM_R_X3Y145_SLICE_X3Y145_B_CY;
  wire [0:0] CLBLM_R_X3Y145_SLICE_X3Y145_B_XOR;
  wire [0:0] CLBLM_R_X3Y145_SLICE_X3Y145_C;
  wire [0:0] CLBLM_R_X3Y145_SLICE_X3Y145_C1;
  wire [0:0] CLBLM_R_X3Y145_SLICE_X3Y145_C2;
  wire [0:0] CLBLM_R_X3Y145_SLICE_X3Y145_C3;
  wire [0:0] CLBLM_R_X3Y145_SLICE_X3Y145_C4;
  wire [0:0] CLBLM_R_X3Y145_SLICE_X3Y145_C5;
  wire [0:0] CLBLM_R_X3Y145_SLICE_X3Y145_C5Q;
  wire [0:0] CLBLM_R_X3Y145_SLICE_X3Y145_C6;
  wire [0:0] CLBLM_R_X3Y145_SLICE_X3Y145_CLK;
  wire [0:0] CLBLM_R_X3Y145_SLICE_X3Y145_CMUX;
  wire [0:0] CLBLM_R_X3Y145_SLICE_X3Y145_CO5;
  wire [0:0] CLBLM_R_X3Y145_SLICE_X3Y145_CO6;
  wire [0:0] CLBLM_R_X3Y145_SLICE_X3Y145_CQ;
  wire [0:0] CLBLM_R_X3Y145_SLICE_X3Y145_C_CY;
  wire [0:0] CLBLM_R_X3Y145_SLICE_X3Y145_C_XOR;
  wire [0:0] CLBLM_R_X3Y145_SLICE_X3Y145_D;
  wire [0:0] CLBLM_R_X3Y145_SLICE_X3Y145_D1;
  wire [0:0] CLBLM_R_X3Y145_SLICE_X3Y145_D2;
  wire [0:0] CLBLM_R_X3Y145_SLICE_X3Y145_D3;
  wire [0:0] CLBLM_R_X3Y145_SLICE_X3Y145_D4;
  wire [0:0] CLBLM_R_X3Y145_SLICE_X3Y145_D5;
  wire [0:0] CLBLM_R_X3Y145_SLICE_X3Y145_D5Q;
  wire [0:0] CLBLM_R_X3Y145_SLICE_X3Y145_D6;
  wire [0:0] CLBLM_R_X3Y145_SLICE_X3Y145_DMUX;
  wire [0:0] CLBLM_R_X3Y145_SLICE_X3Y145_DO5;
  wire [0:0] CLBLM_R_X3Y145_SLICE_X3Y145_DO6;
  wire [0:0] CLBLM_R_X3Y145_SLICE_X3Y145_DQ;
  wire [0:0] CLBLM_R_X3Y145_SLICE_X3Y145_D_CY;
  wire [0:0] CLBLM_R_X3Y145_SLICE_X3Y145_D_XOR;
  wire [0:0] CLBLM_R_X3Y146_SLICE_X2Y146_A;
  wire [0:0] CLBLM_R_X3Y146_SLICE_X2Y146_A1;
  wire [0:0] CLBLM_R_X3Y146_SLICE_X2Y146_A2;
  wire [0:0] CLBLM_R_X3Y146_SLICE_X2Y146_A3;
  wire [0:0] CLBLM_R_X3Y146_SLICE_X2Y146_A4;
  wire [0:0] CLBLM_R_X3Y146_SLICE_X2Y146_A5;
  wire [0:0] CLBLM_R_X3Y146_SLICE_X2Y146_A6;
  wire [0:0] CLBLM_R_X3Y146_SLICE_X2Y146_AO5;
  wire [0:0] CLBLM_R_X3Y146_SLICE_X2Y146_AO6;
  wire [0:0] CLBLM_R_X3Y146_SLICE_X2Y146_AQ;
  wire [0:0] CLBLM_R_X3Y146_SLICE_X2Y146_A_CY;
  wire [0:0] CLBLM_R_X3Y146_SLICE_X2Y146_A_XOR;
  wire [0:0] CLBLM_R_X3Y146_SLICE_X2Y146_B;
  wire [0:0] CLBLM_R_X3Y146_SLICE_X2Y146_B1;
  wire [0:0] CLBLM_R_X3Y146_SLICE_X2Y146_B2;
  wire [0:0] CLBLM_R_X3Y146_SLICE_X2Y146_B3;
  wire [0:0] CLBLM_R_X3Y146_SLICE_X2Y146_B4;
  wire [0:0] CLBLM_R_X3Y146_SLICE_X2Y146_B5;
  wire [0:0] CLBLM_R_X3Y146_SLICE_X2Y146_B6;
  wire [0:0] CLBLM_R_X3Y146_SLICE_X2Y146_BO5;
  wire [0:0] CLBLM_R_X3Y146_SLICE_X2Y146_BO6;
  wire [0:0] CLBLM_R_X3Y146_SLICE_X2Y146_BQ;
  wire [0:0] CLBLM_R_X3Y146_SLICE_X2Y146_B_CY;
  wire [0:0] CLBLM_R_X3Y146_SLICE_X2Y146_B_XOR;
  wire [0:0] CLBLM_R_X3Y146_SLICE_X2Y146_C;
  wire [0:0] CLBLM_R_X3Y146_SLICE_X2Y146_C1;
  wire [0:0] CLBLM_R_X3Y146_SLICE_X2Y146_C2;
  wire [0:0] CLBLM_R_X3Y146_SLICE_X2Y146_C3;
  wire [0:0] CLBLM_R_X3Y146_SLICE_X2Y146_C4;
  wire [0:0] CLBLM_R_X3Y146_SLICE_X2Y146_C5;
  wire [0:0] CLBLM_R_X3Y146_SLICE_X2Y146_C5Q;
  wire [0:0] CLBLM_R_X3Y146_SLICE_X2Y146_C6;
  wire [0:0] CLBLM_R_X3Y146_SLICE_X2Y146_CLK;
  wire [0:0] CLBLM_R_X3Y146_SLICE_X2Y146_CMUX;
  wire [0:0] CLBLM_R_X3Y146_SLICE_X2Y146_CO5;
  wire [0:0] CLBLM_R_X3Y146_SLICE_X2Y146_CO6;
  wire [0:0] CLBLM_R_X3Y146_SLICE_X2Y146_CQ;
  wire [0:0] CLBLM_R_X3Y146_SLICE_X2Y146_C_CY;
  wire [0:0] CLBLM_R_X3Y146_SLICE_X2Y146_C_XOR;
  wire [0:0] CLBLM_R_X3Y146_SLICE_X2Y146_D;
  wire [0:0] CLBLM_R_X3Y146_SLICE_X2Y146_D1;
  wire [0:0] CLBLM_R_X3Y146_SLICE_X2Y146_D2;
  wire [0:0] CLBLM_R_X3Y146_SLICE_X2Y146_D3;
  wire [0:0] CLBLM_R_X3Y146_SLICE_X2Y146_D4;
  wire [0:0] CLBLM_R_X3Y146_SLICE_X2Y146_D5;
  wire [0:0] CLBLM_R_X3Y146_SLICE_X2Y146_D5Q;
  wire [0:0] CLBLM_R_X3Y146_SLICE_X2Y146_D6;
  wire [0:0] CLBLM_R_X3Y146_SLICE_X2Y146_DMUX;
  wire [0:0] CLBLM_R_X3Y146_SLICE_X2Y146_DO5;
  wire [0:0] CLBLM_R_X3Y146_SLICE_X2Y146_DO6;
  wire [0:0] CLBLM_R_X3Y146_SLICE_X2Y146_DQ;
  wire [0:0] CLBLM_R_X3Y146_SLICE_X2Y146_D_CY;
  wire [0:0] CLBLM_R_X3Y146_SLICE_X2Y146_D_XOR;
  wire [0:0] CLBLM_R_X3Y146_SLICE_X3Y146_A;
  wire [0:0] CLBLM_R_X3Y146_SLICE_X3Y146_A1;
  wire [0:0] CLBLM_R_X3Y146_SLICE_X3Y146_A2;
  wire [0:0] CLBLM_R_X3Y146_SLICE_X3Y146_A3;
  wire [0:0] CLBLM_R_X3Y146_SLICE_X3Y146_A4;
  wire [0:0] CLBLM_R_X3Y146_SLICE_X3Y146_A5;
  wire [0:0] CLBLM_R_X3Y146_SLICE_X3Y146_A6;
  wire [0:0] CLBLM_R_X3Y146_SLICE_X3Y146_AO5;
  wire [0:0] CLBLM_R_X3Y146_SLICE_X3Y146_AO6;
  wire [0:0] CLBLM_R_X3Y146_SLICE_X3Y146_AQ;
  wire [0:0] CLBLM_R_X3Y146_SLICE_X3Y146_A_CY;
  wire [0:0] CLBLM_R_X3Y146_SLICE_X3Y146_A_XOR;
  wire [0:0] CLBLM_R_X3Y146_SLICE_X3Y146_B;
  wire [0:0] CLBLM_R_X3Y146_SLICE_X3Y146_B1;
  wire [0:0] CLBLM_R_X3Y146_SLICE_X3Y146_B2;
  wire [0:0] CLBLM_R_X3Y146_SLICE_X3Y146_B3;
  wire [0:0] CLBLM_R_X3Y146_SLICE_X3Y146_B4;
  wire [0:0] CLBLM_R_X3Y146_SLICE_X3Y146_B5;
  wire [0:0] CLBLM_R_X3Y146_SLICE_X3Y146_B6;
  wire [0:0] CLBLM_R_X3Y146_SLICE_X3Y146_BO5;
  wire [0:0] CLBLM_R_X3Y146_SLICE_X3Y146_BO6;
  wire [0:0] CLBLM_R_X3Y146_SLICE_X3Y146_BQ;
  wire [0:0] CLBLM_R_X3Y146_SLICE_X3Y146_B_CY;
  wire [0:0] CLBLM_R_X3Y146_SLICE_X3Y146_B_XOR;
  wire [0:0] CLBLM_R_X3Y146_SLICE_X3Y146_C;
  wire [0:0] CLBLM_R_X3Y146_SLICE_X3Y146_C1;
  wire [0:0] CLBLM_R_X3Y146_SLICE_X3Y146_C2;
  wire [0:0] CLBLM_R_X3Y146_SLICE_X3Y146_C3;
  wire [0:0] CLBLM_R_X3Y146_SLICE_X3Y146_C4;
  wire [0:0] CLBLM_R_X3Y146_SLICE_X3Y146_C5;
  wire [0:0] CLBLM_R_X3Y146_SLICE_X3Y146_C6;
  wire [0:0] CLBLM_R_X3Y146_SLICE_X3Y146_CLK;
  wire [0:0] CLBLM_R_X3Y146_SLICE_X3Y146_CO5;
  wire [0:0] CLBLM_R_X3Y146_SLICE_X3Y146_CO6;
  wire [0:0] CLBLM_R_X3Y146_SLICE_X3Y146_C_CY;
  wire [0:0] CLBLM_R_X3Y146_SLICE_X3Y146_C_XOR;
  wire [0:0] CLBLM_R_X3Y146_SLICE_X3Y146_D;
  wire [0:0] CLBLM_R_X3Y146_SLICE_X3Y146_D1;
  wire [0:0] CLBLM_R_X3Y146_SLICE_X3Y146_D2;
  wire [0:0] CLBLM_R_X3Y146_SLICE_X3Y146_D3;
  wire [0:0] CLBLM_R_X3Y146_SLICE_X3Y146_D4;
  wire [0:0] CLBLM_R_X3Y146_SLICE_X3Y146_D5;
  wire [0:0] CLBLM_R_X3Y146_SLICE_X3Y146_D6;
  wire [0:0] CLBLM_R_X3Y146_SLICE_X3Y146_DO5;
  wire [0:0] CLBLM_R_X3Y146_SLICE_X3Y146_DO6;
  wire [0:0] CLBLM_R_X3Y146_SLICE_X3Y146_D_CY;
  wire [0:0] CLBLM_R_X3Y146_SLICE_X3Y146_D_XOR;
  wire [0:0] CLBLM_R_X3Y147_SLICE_X2Y147_A;
  wire [0:0] CLBLM_R_X3Y147_SLICE_X2Y147_A1;
  wire [0:0] CLBLM_R_X3Y147_SLICE_X2Y147_A2;
  wire [0:0] CLBLM_R_X3Y147_SLICE_X2Y147_A3;
  wire [0:0] CLBLM_R_X3Y147_SLICE_X2Y147_A4;
  wire [0:0] CLBLM_R_X3Y147_SLICE_X2Y147_A5;
  wire [0:0] CLBLM_R_X3Y147_SLICE_X2Y147_A6;
  wire [0:0] CLBLM_R_X3Y147_SLICE_X2Y147_AO5;
  wire [0:0] CLBLM_R_X3Y147_SLICE_X2Y147_AO6;
  wire [0:0] CLBLM_R_X3Y147_SLICE_X2Y147_AQ;
  wire [0:0] CLBLM_R_X3Y147_SLICE_X2Y147_A_CY;
  wire [0:0] CLBLM_R_X3Y147_SLICE_X2Y147_A_XOR;
  wire [0:0] CLBLM_R_X3Y147_SLICE_X2Y147_B;
  wire [0:0] CLBLM_R_X3Y147_SLICE_X2Y147_B1;
  wire [0:0] CLBLM_R_X3Y147_SLICE_X2Y147_B2;
  wire [0:0] CLBLM_R_X3Y147_SLICE_X2Y147_B3;
  wire [0:0] CLBLM_R_X3Y147_SLICE_X2Y147_B4;
  wire [0:0] CLBLM_R_X3Y147_SLICE_X2Y147_B5;
  wire [0:0] CLBLM_R_X3Y147_SLICE_X2Y147_B6;
  wire [0:0] CLBLM_R_X3Y147_SLICE_X2Y147_BO5;
  wire [0:0] CLBLM_R_X3Y147_SLICE_X2Y147_BO6;
  wire [0:0] CLBLM_R_X3Y147_SLICE_X2Y147_BQ;
  wire [0:0] CLBLM_R_X3Y147_SLICE_X2Y147_B_CY;
  wire [0:0] CLBLM_R_X3Y147_SLICE_X2Y147_B_XOR;
  wire [0:0] CLBLM_R_X3Y147_SLICE_X2Y147_C;
  wire [0:0] CLBLM_R_X3Y147_SLICE_X2Y147_C1;
  wire [0:0] CLBLM_R_X3Y147_SLICE_X2Y147_C2;
  wire [0:0] CLBLM_R_X3Y147_SLICE_X2Y147_C3;
  wire [0:0] CLBLM_R_X3Y147_SLICE_X2Y147_C4;
  wire [0:0] CLBLM_R_X3Y147_SLICE_X2Y147_C5;
  wire [0:0] CLBLM_R_X3Y147_SLICE_X2Y147_C6;
  wire [0:0] CLBLM_R_X3Y147_SLICE_X2Y147_CLK;
  wire [0:0] CLBLM_R_X3Y147_SLICE_X2Y147_CO5;
  wire [0:0] CLBLM_R_X3Y147_SLICE_X2Y147_CO6;
  wire [0:0] CLBLM_R_X3Y147_SLICE_X2Y147_CQ;
  wire [0:0] CLBLM_R_X3Y147_SLICE_X2Y147_C_CY;
  wire [0:0] CLBLM_R_X3Y147_SLICE_X2Y147_C_XOR;
  wire [0:0] CLBLM_R_X3Y147_SLICE_X2Y147_D;
  wire [0:0] CLBLM_R_X3Y147_SLICE_X2Y147_D1;
  wire [0:0] CLBLM_R_X3Y147_SLICE_X2Y147_D2;
  wire [0:0] CLBLM_R_X3Y147_SLICE_X2Y147_D3;
  wire [0:0] CLBLM_R_X3Y147_SLICE_X2Y147_D4;
  wire [0:0] CLBLM_R_X3Y147_SLICE_X2Y147_D5;
  wire [0:0] CLBLM_R_X3Y147_SLICE_X2Y147_D5Q;
  wire [0:0] CLBLM_R_X3Y147_SLICE_X2Y147_D6;
  wire [0:0] CLBLM_R_X3Y147_SLICE_X2Y147_DMUX;
  wire [0:0] CLBLM_R_X3Y147_SLICE_X2Y147_DO5;
  wire [0:0] CLBLM_R_X3Y147_SLICE_X2Y147_DO6;
  wire [0:0] CLBLM_R_X3Y147_SLICE_X2Y147_DQ;
  wire [0:0] CLBLM_R_X3Y147_SLICE_X2Y147_D_CY;
  wire [0:0] CLBLM_R_X3Y147_SLICE_X2Y147_D_XOR;
  wire [0:0] CLBLM_R_X3Y147_SLICE_X3Y147_A;
  wire [0:0] CLBLM_R_X3Y147_SLICE_X3Y147_A1;
  wire [0:0] CLBLM_R_X3Y147_SLICE_X3Y147_A2;
  wire [0:0] CLBLM_R_X3Y147_SLICE_X3Y147_A3;
  wire [0:0] CLBLM_R_X3Y147_SLICE_X3Y147_A4;
  wire [0:0] CLBLM_R_X3Y147_SLICE_X3Y147_A5;
  wire [0:0] CLBLM_R_X3Y147_SLICE_X3Y147_A6;
  wire [0:0] CLBLM_R_X3Y147_SLICE_X3Y147_AO5;
  wire [0:0] CLBLM_R_X3Y147_SLICE_X3Y147_AO6;
  wire [0:0] CLBLM_R_X3Y147_SLICE_X3Y147_AQ;
  wire [0:0] CLBLM_R_X3Y147_SLICE_X3Y147_A_CY;
  wire [0:0] CLBLM_R_X3Y147_SLICE_X3Y147_A_XOR;
  wire [0:0] CLBLM_R_X3Y147_SLICE_X3Y147_B;
  wire [0:0] CLBLM_R_X3Y147_SLICE_X3Y147_B1;
  wire [0:0] CLBLM_R_X3Y147_SLICE_X3Y147_B2;
  wire [0:0] CLBLM_R_X3Y147_SLICE_X3Y147_B3;
  wire [0:0] CLBLM_R_X3Y147_SLICE_X3Y147_B4;
  wire [0:0] CLBLM_R_X3Y147_SLICE_X3Y147_B5;
  wire [0:0] CLBLM_R_X3Y147_SLICE_X3Y147_B5Q;
  wire [0:0] CLBLM_R_X3Y147_SLICE_X3Y147_B6;
  wire [0:0] CLBLM_R_X3Y147_SLICE_X3Y147_BMUX;
  wire [0:0] CLBLM_R_X3Y147_SLICE_X3Y147_BO5;
  wire [0:0] CLBLM_R_X3Y147_SLICE_X3Y147_BO6;
  wire [0:0] CLBLM_R_X3Y147_SLICE_X3Y147_BQ;
  wire [0:0] CLBLM_R_X3Y147_SLICE_X3Y147_B_CY;
  wire [0:0] CLBLM_R_X3Y147_SLICE_X3Y147_B_XOR;
  wire [0:0] CLBLM_R_X3Y147_SLICE_X3Y147_C;
  wire [0:0] CLBLM_R_X3Y147_SLICE_X3Y147_C1;
  wire [0:0] CLBLM_R_X3Y147_SLICE_X3Y147_C2;
  wire [0:0] CLBLM_R_X3Y147_SLICE_X3Y147_C3;
  wire [0:0] CLBLM_R_X3Y147_SLICE_X3Y147_C4;
  wire [0:0] CLBLM_R_X3Y147_SLICE_X3Y147_C5;
  wire [0:0] CLBLM_R_X3Y147_SLICE_X3Y147_C5Q;
  wire [0:0] CLBLM_R_X3Y147_SLICE_X3Y147_C6;
  wire [0:0] CLBLM_R_X3Y147_SLICE_X3Y147_CLK;
  wire [0:0] CLBLM_R_X3Y147_SLICE_X3Y147_CMUX;
  wire [0:0] CLBLM_R_X3Y147_SLICE_X3Y147_CO5;
  wire [0:0] CLBLM_R_X3Y147_SLICE_X3Y147_CO6;
  wire [0:0] CLBLM_R_X3Y147_SLICE_X3Y147_CQ;
  wire [0:0] CLBLM_R_X3Y147_SLICE_X3Y147_C_CY;
  wire [0:0] CLBLM_R_X3Y147_SLICE_X3Y147_C_XOR;
  wire [0:0] CLBLM_R_X3Y147_SLICE_X3Y147_D;
  wire [0:0] CLBLM_R_X3Y147_SLICE_X3Y147_D1;
  wire [0:0] CLBLM_R_X3Y147_SLICE_X3Y147_D2;
  wire [0:0] CLBLM_R_X3Y147_SLICE_X3Y147_D3;
  wire [0:0] CLBLM_R_X3Y147_SLICE_X3Y147_D4;
  wire [0:0] CLBLM_R_X3Y147_SLICE_X3Y147_D5;
  wire [0:0] CLBLM_R_X3Y147_SLICE_X3Y147_D6;
  wire [0:0] CLBLM_R_X3Y147_SLICE_X3Y147_DO5;
  wire [0:0] CLBLM_R_X3Y147_SLICE_X3Y147_DO6;
  wire [0:0] CLBLM_R_X3Y147_SLICE_X3Y147_D_CY;
  wire [0:0] CLBLM_R_X3Y147_SLICE_X3Y147_D_XOR;
  wire [0:0] CLBLM_R_X3Y148_SLICE_X2Y148_A;
  wire [0:0] CLBLM_R_X3Y148_SLICE_X2Y148_A1;
  wire [0:0] CLBLM_R_X3Y148_SLICE_X2Y148_A2;
  wire [0:0] CLBLM_R_X3Y148_SLICE_X2Y148_A3;
  wire [0:0] CLBLM_R_X3Y148_SLICE_X2Y148_A4;
  wire [0:0] CLBLM_R_X3Y148_SLICE_X2Y148_A5;
  wire [0:0] CLBLM_R_X3Y148_SLICE_X2Y148_A5Q;
  wire [0:0] CLBLM_R_X3Y148_SLICE_X2Y148_A6;
  wire [0:0] CLBLM_R_X3Y148_SLICE_X2Y148_AMUX;
  wire [0:0] CLBLM_R_X3Y148_SLICE_X2Y148_AO5;
  wire [0:0] CLBLM_R_X3Y148_SLICE_X2Y148_AO6;
  wire [0:0] CLBLM_R_X3Y148_SLICE_X2Y148_AQ;
  wire [0:0] CLBLM_R_X3Y148_SLICE_X2Y148_A_CY;
  wire [0:0] CLBLM_R_X3Y148_SLICE_X2Y148_A_XOR;
  wire [0:0] CLBLM_R_X3Y148_SLICE_X2Y148_B;
  wire [0:0] CLBLM_R_X3Y148_SLICE_X2Y148_B1;
  wire [0:0] CLBLM_R_X3Y148_SLICE_X2Y148_B2;
  wire [0:0] CLBLM_R_X3Y148_SLICE_X2Y148_B3;
  wire [0:0] CLBLM_R_X3Y148_SLICE_X2Y148_B4;
  wire [0:0] CLBLM_R_X3Y148_SLICE_X2Y148_B5;
  wire [0:0] CLBLM_R_X3Y148_SLICE_X2Y148_B5Q;
  wire [0:0] CLBLM_R_X3Y148_SLICE_X2Y148_B6;
  wire [0:0] CLBLM_R_X3Y148_SLICE_X2Y148_BMUX;
  wire [0:0] CLBLM_R_X3Y148_SLICE_X2Y148_BO5;
  wire [0:0] CLBLM_R_X3Y148_SLICE_X2Y148_BO6;
  wire [0:0] CLBLM_R_X3Y148_SLICE_X2Y148_BQ;
  wire [0:0] CLBLM_R_X3Y148_SLICE_X2Y148_B_CY;
  wire [0:0] CLBLM_R_X3Y148_SLICE_X2Y148_B_XOR;
  wire [0:0] CLBLM_R_X3Y148_SLICE_X2Y148_C;
  wire [0:0] CLBLM_R_X3Y148_SLICE_X2Y148_C1;
  wire [0:0] CLBLM_R_X3Y148_SLICE_X2Y148_C2;
  wire [0:0] CLBLM_R_X3Y148_SLICE_X2Y148_C3;
  wire [0:0] CLBLM_R_X3Y148_SLICE_X2Y148_C4;
  wire [0:0] CLBLM_R_X3Y148_SLICE_X2Y148_C5;
  wire [0:0] CLBLM_R_X3Y148_SLICE_X2Y148_C6;
  wire [0:0] CLBLM_R_X3Y148_SLICE_X2Y148_CLK;
  wire [0:0] CLBLM_R_X3Y148_SLICE_X2Y148_CMUX;
  wire [0:0] CLBLM_R_X3Y148_SLICE_X2Y148_CO5;
  wire [0:0] CLBLM_R_X3Y148_SLICE_X2Y148_CO6;
  wire [0:0] CLBLM_R_X3Y148_SLICE_X2Y148_C_CY;
  wire [0:0] CLBLM_R_X3Y148_SLICE_X2Y148_C_XOR;
  wire [0:0] CLBLM_R_X3Y148_SLICE_X2Y148_D;
  wire [0:0] CLBLM_R_X3Y148_SLICE_X2Y148_D1;
  wire [0:0] CLBLM_R_X3Y148_SLICE_X2Y148_D2;
  wire [0:0] CLBLM_R_X3Y148_SLICE_X2Y148_D3;
  wire [0:0] CLBLM_R_X3Y148_SLICE_X2Y148_D4;
  wire [0:0] CLBLM_R_X3Y148_SLICE_X2Y148_D5;
  wire [0:0] CLBLM_R_X3Y148_SLICE_X2Y148_D6;
  wire [0:0] CLBLM_R_X3Y148_SLICE_X2Y148_DO5;
  wire [0:0] CLBLM_R_X3Y148_SLICE_X2Y148_DO6;
  wire [0:0] CLBLM_R_X3Y148_SLICE_X2Y148_D_CY;
  wire [0:0] CLBLM_R_X3Y148_SLICE_X2Y148_D_XOR;
  wire [0:0] CLBLM_R_X3Y148_SLICE_X3Y148_A;
  wire [0:0] CLBLM_R_X3Y148_SLICE_X3Y148_A1;
  wire [0:0] CLBLM_R_X3Y148_SLICE_X3Y148_A2;
  wire [0:0] CLBLM_R_X3Y148_SLICE_X3Y148_A3;
  wire [0:0] CLBLM_R_X3Y148_SLICE_X3Y148_A4;
  wire [0:0] CLBLM_R_X3Y148_SLICE_X3Y148_A5;
  wire [0:0] CLBLM_R_X3Y148_SLICE_X3Y148_A6;
  wire [0:0] CLBLM_R_X3Y148_SLICE_X3Y148_AO5;
  wire [0:0] CLBLM_R_X3Y148_SLICE_X3Y148_AO6;
  wire [0:0] CLBLM_R_X3Y148_SLICE_X3Y148_AQ;
  wire [0:0] CLBLM_R_X3Y148_SLICE_X3Y148_A_CY;
  wire [0:0] CLBLM_R_X3Y148_SLICE_X3Y148_A_XOR;
  wire [0:0] CLBLM_R_X3Y148_SLICE_X3Y148_B;
  wire [0:0] CLBLM_R_X3Y148_SLICE_X3Y148_B1;
  wire [0:0] CLBLM_R_X3Y148_SLICE_X3Y148_B2;
  wire [0:0] CLBLM_R_X3Y148_SLICE_X3Y148_B3;
  wire [0:0] CLBLM_R_X3Y148_SLICE_X3Y148_B4;
  wire [0:0] CLBLM_R_X3Y148_SLICE_X3Y148_B5;
  wire [0:0] CLBLM_R_X3Y148_SLICE_X3Y148_B5Q;
  wire [0:0] CLBLM_R_X3Y148_SLICE_X3Y148_B6;
  wire [0:0] CLBLM_R_X3Y148_SLICE_X3Y148_BMUX;
  wire [0:0] CLBLM_R_X3Y148_SLICE_X3Y148_BO5;
  wire [0:0] CLBLM_R_X3Y148_SLICE_X3Y148_BO6;
  wire [0:0] CLBLM_R_X3Y148_SLICE_X3Y148_BQ;
  wire [0:0] CLBLM_R_X3Y148_SLICE_X3Y148_B_CY;
  wire [0:0] CLBLM_R_X3Y148_SLICE_X3Y148_B_XOR;
  wire [0:0] CLBLM_R_X3Y148_SLICE_X3Y148_C;
  wire [0:0] CLBLM_R_X3Y148_SLICE_X3Y148_C1;
  wire [0:0] CLBLM_R_X3Y148_SLICE_X3Y148_C2;
  wire [0:0] CLBLM_R_X3Y148_SLICE_X3Y148_C3;
  wire [0:0] CLBLM_R_X3Y148_SLICE_X3Y148_C4;
  wire [0:0] CLBLM_R_X3Y148_SLICE_X3Y148_C5;
  wire [0:0] CLBLM_R_X3Y148_SLICE_X3Y148_C5Q;
  wire [0:0] CLBLM_R_X3Y148_SLICE_X3Y148_C6;
  wire [0:0] CLBLM_R_X3Y148_SLICE_X3Y148_CLK;
  wire [0:0] CLBLM_R_X3Y148_SLICE_X3Y148_CMUX;
  wire [0:0] CLBLM_R_X3Y148_SLICE_X3Y148_CO5;
  wire [0:0] CLBLM_R_X3Y148_SLICE_X3Y148_CO6;
  wire [0:0] CLBLM_R_X3Y148_SLICE_X3Y148_CQ;
  wire [0:0] CLBLM_R_X3Y148_SLICE_X3Y148_C_CY;
  wire [0:0] CLBLM_R_X3Y148_SLICE_X3Y148_C_XOR;
  wire [0:0] CLBLM_R_X3Y148_SLICE_X3Y148_D;
  wire [0:0] CLBLM_R_X3Y148_SLICE_X3Y148_D1;
  wire [0:0] CLBLM_R_X3Y148_SLICE_X3Y148_D2;
  wire [0:0] CLBLM_R_X3Y148_SLICE_X3Y148_D3;
  wire [0:0] CLBLM_R_X3Y148_SLICE_X3Y148_D4;
  wire [0:0] CLBLM_R_X3Y148_SLICE_X3Y148_D5;
  wire [0:0] CLBLM_R_X3Y148_SLICE_X3Y148_D6;
  wire [0:0] CLBLM_R_X3Y148_SLICE_X3Y148_DMUX;
  wire [0:0] CLBLM_R_X3Y148_SLICE_X3Y148_DO5;
  wire [0:0] CLBLM_R_X3Y148_SLICE_X3Y148_DO6;
  wire [0:0] CLBLM_R_X3Y148_SLICE_X3Y148_D_CY;
  wire [0:0] CLBLM_R_X3Y148_SLICE_X3Y148_D_XOR;
  wire [0:0] CLBLM_R_X3Y149_SLICE_X2Y149_A;
  wire [0:0] CLBLM_R_X3Y149_SLICE_X2Y149_A1;
  wire [0:0] CLBLM_R_X3Y149_SLICE_X2Y149_A2;
  wire [0:0] CLBLM_R_X3Y149_SLICE_X2Y149_A3;
  wire [0:0] CLBLM_R_X3Y149_SLICE_X2Y149_A4;
  wire [0:0] CLBLM_R_X3Y149_SLICE_X2Y149_A5;
  wire [0:0] CLBLM_R_X3Y149_SLICE_X2Y149_A6;
  wire [0:0] CLBLM_R_X3Y149_SLICE_X2Y149_AO5;
  wire [0:0] CLBLM_R_X3Y149_SLICE_X2Y149_AO6;
  wire [0:0] CLBLM_R_X3Y149_SLICE_X2Y149_AQ;
  wire [0:0] CLBLM_R_X3Y149_SLICE_X2Y149_A_CY;
  wire [0:0] CLBLM_R_X3Y149_SLICE_X2Y149_A_XOR;
  wire [0:0] CLBLM_R_X3Y149_SLICE_X2Y149_B;
  wire [0:0] CLBLM_R_X3Y149_SLICE_X2Y149_B1;
  wire [0:0] CLBLM_R_X3Y149_SLICE_X2Y149_B2;
  wire [0:0] CLBLM_R_X3Y149_SLICE_X2Y149_B3;
  wire [0:0] CLBLM_R_X3Y149_SLICE_X2Y149_B4;
  wire [0:0] CLBLM_R_X3Y149_SLICE_X2Y149_B5;
  wire [0:0] CLBLM_R_X3Y149_SLICE_X2Y149_B6;
  wire [0:0] CLBLM_R_X3Y149_SLICE_X2Y149_BO5;
  wire [0:0] CLBLM_R_X3Y149_SLICE_X2Y149_BO6;
  wire [0:0] CLBLM_R_X3Y149_SLICE_X2Y149_BQ;
  wire [0:0] CLBLM_R_X3Y149_SLICE_X2Y149_B_CY;
  wire [0:0] CLBLM_R_X3Y149_SLICE_X2Y149_B_XOR;
  wire [0:0] CLBLM_R_X3Y149_SLICE_X2Y149_C;
  wire [0:0] CLBLM_R_X3Y149_SLICE_X2Y149_C1;
  wire [0:0] CLBLM_R_X3Y149_SLICE_X2Y149_C2;
  wire [0:0] CLBLM_R_X3Y149_SLICE_X2Y149_C3;
  wire [0:0] CLBLM_R_X3Y149_SLICE_X2Y149_C4;
  wire [0:0] CLBLM_R_X3Y149_SLICE_X2Y149_C5;
  wire [0:0] CLBLM_R_X3Y149_SLICE_X2Y149_C5Q;
  wire [0:0] CLBLM_R_X3Y149_SLICE_X2Y149_C6;
  wire [0:0] CLBLM_R_X3Y149_SLICE_X2Y149_CLK;
  wire [0:0] CLBLM_R_X3Y149_SLICE_X2Y149_CMUX;
  wire [0:0] CLBLM_R_X3Y149_SLICE_X2Y149_CO5;
  wire [0:0] CLBLM_R_X3Y149_SLICE_X2Y149_CO6;
  wire [0:0] CLBLM_R_X3Y149_SLICE_X2Y149_CQ;
  wire [0:0] CLBLM_R_X3Y149_SLICE_X2Y149_C_CY;
  wire [0:0] CLBLM_R_X3Y149_SLICE_X2Y149_C_XOR;
  wire [0:0] CLBLM_R_X3Y149_SLICE_X2Y149_D;
  wire [0:0] CLBLM_R_X3Y149_SLICE_X2Y149_D1;
  wire [0:0] CLBLM_R_X3Y149_SLICE_X2Y149_D2;
  wire [0:0] CLBLM_R_X3Y149_SLICE_X2Y149_D3;
  wire [0:0] CLBLM_R_X3Y149_SLICE_X2Y149_D4;
  wire [0:0] CLBLM_R_X3Y149_SLICE_X2Y149_D5;
  wire [0:0] CLBLM_R_X3Y149_SLICE_X2Y149_D6;
  wire [0:0] CLBLM_R_X3Y149_SLICE_X2Y149_DO5;
  wire [0:0] CLBLM_R_X3Y149_SLICE_X2Y149_DO6;
  wire [0:0] CLBLM_R_X3Y149_SLICE_X2Y149_DQ;
  wire [0:0] CLBLM_R_X3Y149_SLICE_X2Y149_D_CY;
  wire [0:0] CLBLM_R_X3Y149_SLICE_X2Y149_D_XOR;
  wire [0:0] CLBLM_R_X3Y149_SLICE_X3Y149_A;
  wire [0:0] CLBLM_R_X3Y149_SLICE_X3Y149_A1;
  wire [0:0] CLBLM_R_X3Y149_SLICE_X3Y149_A2;
  wire [0:0] CLBLM_R_X3Y149_SLICE_X3Y149_A3;
  wire [0:0] CLBLM_R_X3Y149_SLICE_X3Y149_A4;
  wire [0:0] CLBLM_R_X3Y149_SLICE_X3Y149_A5;
  wire [0:0] CLBLM_R_X3Y149_SLICE_X3Y149_A6;
  wire [0:0] CLBLM_R_X3Y149_SLICE_X3Y149_AO5;
  wire [0:0] CLBLM_R_X3Y149_SLICE_X3Y149_AO6;
  wire [0:0] CLBLM_R_X3Y149_SLICE_X3Y149_AQ;
  wire [0:0] CLBLM_R_X3Y149_SLICE_X3Y149_A_CY;
  wire [0:0] CLBLM_R_X3Y149_SLICE_X3Y149_A_XOR;
  wire [0:0] CLBLM_R_X3Y149_SLICE_X3Y149_B;
  wire [0:0] CLBLM_R_X3Y149_SLICE_X3Y149_B1;
  wire [0:0] CLBLM_R_X3Y149_SLICE_X3Y149_B2;
  wire [0:0] CLBLM_R_X3Y149_SLICE_X3Y149_B3;
  wire [0:0] CLBLM_R_X3Y149_SLICE_X3Y149_B4;
  wire [0:0] CLBLM_R_X3Y149_SLICE_X3Y149_B5;
  wire [0:0] CLBLM_R_X3Y149_SLICE_X3Y149_B6;
  wire [0:0] CLBLM_R_X3Y149_SLICE_X3Y149_BO5;
  wire [0:0] CLBLM_R_X3Y149_SLICE_X3Y149_BO6;
  wire [0:0] CLBLM_R_X3Y149_SLICE_X3Y149_BQ;
  wire [0:0] CLBLM_R_X3Y149_SLICE_X3Y149_B_CY;
  wire [0:0] CLBLM_R_X3Y149_SLICE_X3Y149_B_XOR;
  wire [0:0] CLBLM_R_X3Y149_SLICE_X3Y149_C;
  wire [0:0] CLBLM_R_X3Y149_SLICE_X3Y149_C1;
  wire [0:0] CLBLM_R_X3Y149_SLICE_X3Y149_C2;
  wire [0:0] CLBLM_R_X3Y149_SLICE_X3Y149_C3;
  wire [0:0] CLBLM_R_X3Y149_SLICE_X3Y149_C4;
  wire [0:0] CLBLM_R_X3Y149_SLICE_X3Y149_C5;
  wire [0:0] CLBLM_R_X3Y149_SLICE_X3Y149_C6;
  wire [0:0] CLBLM_R_X3Y149_SLICE_X3Y149_CLK;
  wire [0:0] CLBLM_R_X3Y149_SLICE_X3Y149_CO5;
  wire [0:0] CLBLM_R_X3Y149_SLICE_X3Y149_CO6;
  wire [0:0] CLBLM_R_X3Y149_SLICE_X3Y149_CQ;
  wire [0:0] CLBLM_R_X3Y149_SLICE_X3Y149_C_CY;
  wire [0:0] CLBLM_R_X3Y149_SLICE_X3Y149_C_XOR;
  wire [0:0] CLBLM_R_X3Y149_SLICE_X3Y149_D;
  wire [0:0] CLBLM_R_X3Y149_SLICE_X3Y149_D1;
  wire [0:0] CLBLM_R_X3Y149_SLICE_X3Y149_D2;
  wire [0:0] CLBLM_R_X3Y149_SLICE_X3Y149_D3;
  wire [0:0] CLBLM_R_X3Y149_SLICE_X3Y149_D4;
  wire [0:0] CLBLM_R_X3Y149_SLICE_X3Y149_D5;
  wire [0:0] CLBLM_R_X3Y149_SLICE_X3Y149_D5Q;
  wire [0:0] CLBLM_R_X3Y149_SLICE_X3Y149_D6;
  wire [0:0] CLBLM_R_X3Y149_SLICE_X3Y149_DMUX;
  wire [0:0] CLBLM_R_X3Y149_SLICE_X3Y149_DO5;
  wire [0:0] CLBLM_R_X3Y149_SLICE_X3Y149_DO6;
  wire [0:0] CLBLM_R_X3Y149_SLICE_X3Y149_DQ;
  wire [0:0] CLBLM_R_X3Y149_SLICE_X3Y149_D_CY;
  wire [0:0] CLBLM_R_X3Y149_SLICE_X3Y149_D_XOR;
  wire [0:0] CLBLM_R_X3Y150_SLICE_X2Y150_A;
  wire [0:0] CLBLM_R_X3Y150_SLICE_X2Y150_A1;
  wire [0:0] CLBLM_R_X3Y150_SLICE_X2Y150_A2;
  wire [0:0] CLBLM_R_X3Y150_SLICE_X2Y150_A3;
  wire [0:0] CLBLM_R_X3Y150_SLICE_X2Y150_A4;
  wire [0:0] CLBLM_R_X3Y150_SLICE_X2Y150_A5;
  wire [0:0] CLBLM_R_X3Y150_SLICE_X2Y150_A6;
  wire [0:0] CLBLM_R_X3Y150_SLICE_X2Y150_AO5;
  wire [0:0] CLBLM_R_X3Y150_SLICE_X2Y150_AO6;
  wire [0:0] CLBLM_R_X3Y150_SLICE_X2Y150_AQ;
  wire [0:0] CLBLM_R_X3Y150_SLICE_X2Y150_A_CY;
  wire [0:0] CLBLM_R_X3Y150_SLICE_X2Y150_A_XOR;
  wire [0:0] CLBLM_R_X3Y150_SLICE_X2Y150_B;
  wire [0:0] CLBLM_R_X3Y150_SLICE_X2Y150_B1;
  wire [0:0] CLBLM_R_X3Y150_SLICE_X2Y150_B2;
  wire [0:0] CLBLM_R_X3Y150_SLICE_X2Y150_B3;
  wire [0:0] CLBLM_R_X3Y150_SLICE_X2Y150_B4;
  wire [0:0] CLBLM_R_X3Y150_SLICE_X2Y150_B5;
  wire [0:0] CLBLM_R_X3Y150_SLICE_X2Y150_B6;
  wire [0:0] CLBLM_R_X3Y150_SLICE_X2Y150_BO5;
  wire [0:0] CLBLM_R_X3Y150_SLICE_X2Y150_BO6;
  wire [0:0] CLBLM_R_X3Y150_SLICE_X2Y150_BQ;
  wire [0:0] CLBLM_R_X3Y150_SLICE_X2Y150_B_CY;
  wire [0:0] CLBLM_R_X3Y150_SLICE_X2Y150_B_XOR;
  wire [0:0] CLBLM_R_X3Y150_SLICE_X2Y150_C;
  wire [0:0] CLBLM_R_X3Y150_SLICE_X2Y150_C1;
  wire [0:0] CLBLM_R_X3Y150_SLICE_X2Y150_C2;
  wire [0:0] CLBLM_R_X3Y150_SLICE_X2Y150_C3;
  wire [0:0] CLBLM_R_X3Y150_SLICE_X2Y150_C4;
  wire [0:0] CLBLM_R_X3Y150_SLICE_X2Y150_C5;
  wire [0:0] CLBLM_R_X3Y150_SLICE_X2Y150_C6;
  wire [0:0] CLBLM_R_X3Y150_SLICE_X2Y150_CLK;
  wire [0:0] CLBLM_R_X3Y150_SLICE_X2Y150_CO5;
  wire [0:0] CLBLM_R_X3Y150_SLICE_X2Y150_CO6;
  wire [0:0] CLBLM_R_X3Y150_SLICE_X2Y150_CQ;
  wire [0:0] CLBLM_R_X3Y150_SLICE_X2Y150_C_CY;
  wire [0:0] CLBLM_R_X3Y150_SLICE_X2Y150_C_XOR;
  wire [0:0] CLBLM_R_X3Y150_SLICE_X2Y150_D;
  wire [0:0] CLBLM_R_X3Y150_SLICE_X2Y150_D1;
  wire [0:0] CLBLM_R_X3Y150_SLICE_X2Y150_D2;
  wire [0:0] CLBLM_R_X3Y150_SLICE_X2Y150_D3;
  wire [0:0] CLBLM_R_X3Y150_SLICE_X2Y150_D4;
  wire [0:0] CLBLM_R_X3Y150_SLICE_X2Y150_D5;
  wire [0:0] CLBLM_R_X3Y150_SLICE_X2Y150_D5Q;
  wire [0:0] CLBLM_R_X3Y150_SLICE_X2Y150_D6;
  wire [0:0] CLBLM_R_X3Y150_SLICE_X2Y150_DMUX;
  wire [0:0] CLBLM_R_X3Y150_SLICE_X2Y150_DO5;
  wire [0:0] CLBLM_R_X3Y150_SLICE_X2Y150_DO6;
  wire [0:0] CLBLM_R_X3Y150_SLICE_X2Y150_DQ;
  wire [0:0] CLBLM_R_X3Y150_SLICE_X2Y150_D_CY;
  wire [0:0] CLBLM_R_X3Y150_SLICE_X2Y150_D_XOR;
  wire [0:0] CLBLM_R_X3Y150_SLICE_X3Y150_A;
  wire [0:0] CLBLM_R_X3Y150_SLICE_X3Y150_A1;
  wire [0:0] CLBLM_R_X3Y150_SLICE_X3Y150_A2;
  wire [0:0] CLBLM_R_X3Y150_SLICE_X3Y150_A3;
  wire [0:0] CLBLM_R_X3Y150_SLICE_X3Y150_A4;
  wire [0:0] CLBLM_R_X3Y150_SLICE_X3Y150_A5;
  wire [0:0] CLBLM_R_X3Y150_SLICE_X3Y150_A5Q;
  wire [0:0] CLBLM_R_X3Y150_SLICE_X3Y150_A6;
  wire [0:0] CLBLM_R_X3Y150_SLICE_X3Y150_AMUX;
  wire [0:0] CLBLM_R_X3Y150_SLICE_X3Y150_AO5;
  wire [0:0] CLBLM_R_X3Y150_SLICE_X3Y150_AO6;
  wire [0:0] CLBLM_R_X3Y150_SLICE_X3Y150_AQ;
  wire [0:0] CLBLM_R_X3Y150_SLICE_X3Y150_A_CY;
  wire [0:0] CLBLM_R_X3Y150_SLICE_X3Y150_A_XOR;
  wire [0:0] CLBLM_R_X3Y150_SLICE_X3Y150_B;
  wire [0:0] CLBLM_R_X3Y150_SLICE_X3Y150_B1;
  wire [0:0] CLBLM_R_X3Y150_SLICE_X3Y150_B2;
  wire [0:0] CLBLM_R_X3Y150_SLICE_X3Y150_B3;
  wire [0:0] CLBLM_R_X3Y150_SLICE_X3Y150_B4;
  wire [0:0] CLBLM_R_X3Y150_SLICE_X3Y150_B5;
  wire [0:0] CLBLM_R_X3Y150_SLICE_X3Y150_B5Q;
  wire [0:0] CLBLM_R_X3Y150_SLICE_X3Y150_B6;
  wire [0:0] CLBLM_R_X3Y150_SLICE_X3Y150_BMUX;
  wire [0:0] CLBLM_R_X3Y150_SLICE_X3Y150_BO5;
  wire [0:0] CLBLM_R_X3Y150_SLICE_X3Y150_BO6;
  wire [0:0] CLBLM_R_X3Y150_SLICE_X3Y150_BQ;
  wire [0:0] CLBLM_R_X3Y150_SLICE_X3Y150_B_CY;
  wire [0:0] CLBLM_R_X3Y150_SLICE_X3Y150_B_XOR;
  wire [0:0] CLBLM_R_X3Y150_SLICE_X3Y150_C;
  wire [0:0] CLBLM_R_X3Y150_SLICE_X3Y150_C1;
  wire [0:0] CLBLM_R_X3Y150_SLICE_X3Y150_C2;
  wire [0:0] CLBLM_R_X3Y150_SLICE_X3Y150_C3;
  wire [0:0] CLBLM_R_X3Y150_SLICE_X3Y150_C4;
  wire [0:0] CLBLM_R_X3Y150_SLICE_X3Y150_C5;
  wire [0:0] CLBLM_R_X3Y150_SLICE_X3Y150_C6;
  wire [0:0] CLBLM_R_X3Y150_SLICE_X3Y150_CLK;
  wire [0:0] CLBLM_R_X3Y150_SLICE_X3Y150_CO5;
  wire [0:0] CLBLM_R_X3Y150_SLICE_X3Y150_CO6;
  wire [0:0] CLBLM_R_X3Y150_SLICE_X3Y150_CQ;
  wire [0:0] CLBLM_R_X3Y150_SLICE_X3Y150_C_CY;
  wire [0:0] CLBLM_R_X3Y150_SLICE_X3Y150_C_XOR;
  wire [0:0] CLBLM_R_X3Y150_SLICE_X3Y150_D;
  wire [0:0] CLBLM_R_X3Y150_SLICE_X3Y150_D1;
  wire [0:0] CLBLM_R_X3Y150_SLICE_X3Y150_D2;
  wire [0:0] CLBLM_R_X3Y150_SLICE_X3Y150_D3;
  wire [0:0] CLBLM_R_X3Y150_SLICE_X3Y150_D4;
  wire [0:0] CLBLM_R_X3Y150_SLICE_X3Y150_D5;
  wire [0:0] CLBLM_R_X3Y150_SLICE_X3Y150_D5Q;
  wire [0:0] CLBLM_R_X3Y150_SLICE_X3Y150_D6;
  wire [0:0] CLBLM_R_X3Y150_SLICE_X3Y150_DMUX;
  wire [0:0] CLBLM_R_X3Y150_SLICE_X3Y150_DO5;
  wire [0:0] CLBLM_R_X3Y150_SLICE_X3Y150_DO6;
  wire [0:0] CLBLM_R_X3Y150_SLICE_X3Y150_DQ;
  wire [0:0] CLBLM_R_X3Y150_SLICE_X3Y150_D_CY;
  wire [0:0] CLBLM_R_X3Y150_SLICE_X3Y150_D_XOR;
  wire [0:0] CLBLM_R_X3Y151_SLICE_X2Y151_A;
  wire [0:0] CLBLM_R_X3Y151_SLICE_X2Y151_A1;
  wire [0:0] CLBLM_R_X3Y151_SLICE_X2Y151_A2;
  wire [0:0] CLBLM_R_X3Y151_SLICE_X2Y151_A3;
  wire [0:0] CLBLM_R_X3Y151_SLICE_X2Y151_A4;
  wire [0:0] CLBLM_R_X3Y151_SLICE_X2Y151_A5;
  wire [0:0] CLBLM_R_X3Y151_SLICE_X2Y151_A6;
  wire [0:0] CLBLM_R_X3Y151_SLICE_X2Y151_AMUX;
  wire [0:0] CLBLM_R_X3Y151_SLICE_X2Y151_AO5;
  wire [0:0] CLBLM_R_X3Y151_SLICE_X2Y151_AO6;
  wire [0:0] CLBLM_R_X3Y151_SLICE_X2Y151_AQ;
  wire [0:0] CLBLM_R_X3Y151_SLICE_X2Y151_AX;
  wire [0:0] CLBLM_R_X3Y151_SLICE_X2Y151_A_CY;
  wire [0:0] CLBLM_R_X3Y151_SLICE_X2Y151_A_XOR;
  wire [0:0] CLBLM_R_X3Y151_SLICE_X2Y151_B;
  wire [0:0] CLBLM_R_X3Y151_SLICE_X2Y151_B1;
  wire [0:0] CLBLM_R_X3Y151_SLICE_X2Y151_B2;
  wire [0:0] CLBLM_R_X3Y151_SLICE_X2Y151_B3;
  wire [0:0] CLBLM_R_X3Y151_SLICE_X2Y151_B4;
  wire [0:0] CLBLM_R_X3Y151_SLICE_X2Y151_B5;
  wire [0:0] CLBLM_R_X3Y151_SLICE_X2Y151_B6;
  wire [0:0] CLBLM_R_X3Y151_SLICE_X2Y151_BMUX;
  wire [0:0] CLBLM_R_X3Y151_SLICE_X2Y151_BO5;
  wire [0:0] CLBLM_R_X3Y151_SLICE_X2Y151_BO6;
  wire [0:0] CLBLM_R_X3Y151_SLICE_X2Y151_B_CY;
  wire [0:0] CLBLM_R_X3Y151_SLICE_X2Y151_B_XOR;
  wire [0:0] CLBLM_R_X3Y151_SLICE_X2Y151_C;
  wire [0:0] CLBLM_R_X3Y151_SLICE_X2Y151_C1;
  wire [0:0] CLBLM_R_X3Y151_SLICE_X2Y151_C2;
  wire [0:0] CLBLM_R_X3Y151_SLICE_X2Y151_C3;
  wire [0:0] CLBLM_R_X3Y151_SLICE_X2Y151_C4;
  wire [0:0] CLBLM_R_X3Y151_SLICE_X2Y151_C5;
  wire [0:0] CLBLM_R_X3Y151_SLICE_X2Y151_C6;
  wire [0:0] CLBLM_R_X3Y151_SLICE_X2Y151_CE;
  wire [0:0] CLBLM_R_X3Y151_SLICE_X2Y151_CLK;
  wire [0:0] CLBLM_R_X3Y151_SLICE_X2Y151_CO5;
  wire [0:0] CLBLM_R_X3Y151_SLICE_X2Y151_CO6;
  wire [0:0] CLBLM_R_X3Y151_SLICE_X2Y151_C_CY;
  wire [0:0] CLBLM_R_X3Y151_SLICE_X2Y151_C_XOR;
  wire [0:0] CLBLM_R_X3Y151_SLICE_X2Y151_D;
  wire [0:0] CLBLM_R_X3Y151_SLICE_X2Y151_D1;
  wire [0:0] CLBLM_R_X3Y151_SLICE_X2Y151_D2;
  wire [0:0] CLBLM_R_X3Y151_SLICE_X2Y151_D3;
  wire [0:0] CLBLM_R_X3Y151_SLICE_X2Y151_D4;
  wire [0:0] CLBLM_R_X3Y151_SLICE_X2Y151_D5;
  wire [0:0] CLBLM_R_X3Y151_SLICE_X2Y151_D6;
  wire [0:0] CLBLM_R_X3Y151_SLICE_X2Y151_DO5;
  wire [0:0] CLBLM_R_X3Y151_SLICE_X2Y151_DO6;
  wire [0:0] CLBLM_R_X3Y151_SLICE_X2Y151_D_CY;
  wire [0:0] CLBLM_R_X3Y151_SLICE_X2Y151_D_XOR;
  wire [0:0] CLBLM_R_X3Y151_SLICE_X3Y151_A;
  wire [0:0] CLBLM_R_X3Y151_SLICE_X3Y151_A1;
  wire [0:0] CLBLM_R_X3Y151_SLICE_X3Y151_A2;
  wire [0:0] CLBLM_R_X3Y151_SLICE_X3Y151_A3;
  wire [0:0] CLBLM_R_X3Y151_SLICE_X3Y151_A4;
  wire [0:0] CLBLM_R_X3Y151_SLICE_X3Y151_A5;
  wire [0:0] CLBLM_R_X3Y151_SLICE_X3Y151_A5Q;
  wire [0:0] CLBLM_R_X3Y151_SLICE_X3Y151_A6;
  wire [0:0] CLBLM_R_X3Y151_SLICE_X3Y151_AMUX;
  wire [0:0] CLBLM_R_X3Y151_SLICE_X3Y151_AO5;
  wire [0:0] CLBLM_R_X3Y151_SLICE_X3Y151_AO6;
  wire [0:0] CLBLM_R_X3Y151_SLICE_X3Y151_AQ;
  wire [0:0] CLBLM_R_X3Y151_SLICE_X3Y151_AX;
  wire [0:0] CLBLM_R_X3Y151_SLICE_X3Y151_A_CY;
  wire [0:0] CLBLM_R_X3Y151_SLICE_X3Y151_A_XOR;
  wire [0:0] CLBLM_R_X3Y151_SLICE_X3Y151_B;
  wire [0:0] CLBLM_R_X3Y151_SLICE_X3Y151_B1;
  wire [0:0] CLBLM_R_X3Y151_SLICE_X3Y151_B2;
  wire [0:0] CLBLM_R_X3Y151_SLICE_X3Y151_B3;
  wire [0:0] CLBLM_R_X3Y151_SLICE_X3Y151_B4;
  wire [0:0] CLBLM_R_X3Y151_SLICE_X3Y151_B5;
  wire [0:0] CLBLM_R_X3Y151_SLICE_X3Y151_B6;
  wire [0:0] CLBLM_R_X3Y151_SLICE_X3Y151_BO5;
  wire [0:0] CLBLM_R_X3Y151_SLICE_X3Y151_BO6;
  wire [0:0] CLBLM_R_X3Y151_SLICE_X3Y151_BQ;
  wire [0:0] CLBLM_R_X3Y151_SLICE_X3Y151_B_CY;
  wire [0:0] CLBLM_R_X3Y151_SLICE_X3Y151_B_XOR;
  wire [0:0] CLBLM_R_X3Y151_SLICE_X3Y151_C;
  wire [0:0] CLBLM_R_X3Y151_SLICE_X3Y151_C1;
  wire [0:0] CLBLM_R_X3Y151_SLICE_X3Y151_C2;
  wire [0:0] CLBLM_R_X3Y151_SLICE_X3Y151_C3;
  wire [0:0] CLBLM_R_X3Y151_SLICE_X3Y151_C4;
  wire [0:0] CLBLM_R_X3Y151_SLICE_X3Y151_C5;
  wire [0:0] CLBLM_R_X3Y151_SLICE_X3Y151_C6;
  wire [0:0] CLBLM_R_X3Y151_SLICE_X3Y151_CLK;
  wire [0:0] CLBLM_R_X3Y151_SLICE_X3Y151_CO5;
  wire [0:0] CLBLM_R_X3Y151_SLICE_X3Y151_CO6;
  wire [0:0] CLBLM_R_X3Y151_SLICE_X3Y151_CQ;
  wire [0:0] CLBLM_R_X3Y151_SLICE_X3Y151_C_CY;
  wire [0:0] CLBLM_R_X3Y151_SLICE_X3Y151_C_XOR;
  wire [0:0] CLBLM_R_X3Y151_SLICE_X3Y151_D;
  wire [0:0] CLBLM_R_X3Y151_SLICE_X3Y151_D1;
  wire [0:0] CLBLM_R_X3Y151_SLICE_X3Y151_D2;
  wire [0:0] CLBLM_R_X3Y151_SLICE_X3Y151_D3;
  wire [0:0] CLBLM_R_X3Y151_SLICE_X3Y151_D4;
  wire [0:0] CLBLM_R_X3Y151_SLICE_X3Y151_D5;
  wire [0:0] CLBLM_R_X3Y151_SLICE_X3Y151_D6;
  wire [0:0] CLBLM_R_X3Y151_SLICE_X3Y151_DMUX;
  wire [0:0] CLBLM_R_X3Y151_SLICE_X3Y151_DO5;
  wire [0:0] CLBLM_R_X3Y151_SLICE_X3Y151_DO6;
  wire [0:0] CLBLM_R_X3Y151_SLICE_X3Y151_D_CY;
  wire [0:0] CLBLM_R_X3Y151_SLICE_X3Y151_D_XOR;
  wire [0:0] CLBLM_R_X3Y152_SLICE_X2Y152_A;
  wire [0:0] CLBLM_R_X3Y152_SLICE_X2Y152_A1;
  wire [0:0] CLBLM_R_X3Y152_SLICE_X2Y152_A2;
  wire [0:0] CLBLM_R_X3Y152_SLICE_X2Y152_A3;
  wire [0:0] CLBLM_R_X3Y152_SLICE_X2Y152_A4;
  wire [0:0] CLBLM_R_X3Y152_SLICE_X2Y152_A5;
  wire [0:0] CLBLM_R_X3Y152_SLICE_X2Y152_A6;
  wire [0:0] CLBLM_R_X3Y152_SLICE_X2Y152_AO5;
  wire [0:0] CLBLM_R_X3Y152_SLICE_X2Y152_AO6;
  wire [0:0] CLBLM_R_X3Y152_SLICE_X2Y152_A_CY;
  wire [0:0] CLBLM_R_X3Y152_SLICE_X2Y152_A_XOR;
  wire [0:0] CLBLM_R_X3Y152_SLICE_X2Y152_B;
  wire [0:0] CLBLM_R_X3Y152_SLICE_X2Y152_B1;
  wire [0:0] CLBLM_R_X3Y152_SLICE_X2Y152_B2;
  wire [0:0] CLBLM_R_X3Y152_SLICE_X2Y152_B3;
  wire [0:0] CLBLM_R_X3Y152_SLICE_X2Y152_B4;
  wire [0:0] CLBLM_R_X3Y152_SLICE_X2Y152_B5;
  wire [0:0] CLBLM_R_X3Y152_SLICE_X2Y152_B6;
  wire [0:0] CLBLM_R_X3Y152_SLICE_X2Y152_BO5;
  wire [0:0] CLBLM_R_X3Y152_SLICE_X2Y152_BO6;
  wire [0:0] CLBLM_R_X3Y152_SLICE_X2Y152_B_CY;
  wire [0:0] CLBLM_R_X3Y152_SLICE_X2Y152_B_XOR;
  wire [0:0] CLBLM_R_X3Y152_SLICE_X2Y152_C;
  wire [0:0] CLBLM_R_X3Y152_SLICE_X2Y152_C1;
  wire [0:0] CLBLM_R_X3Y152_SLICE_X2Y152_C2;
  wire [0:0] CLBLM_R_X3Y152_SLICE_X2Y152_C3;
  wire [0:0] CLBLM_R_X3Y152_SLICE_X2Y152_C4;
  wire [0:0] CLBLM_R_X3Y152_SLICE_X2Y152_C5;
  wire [0:0] CLBLM_R_X3Y152_SLICE_X2Y152_C6;
  wire [0:0] CLBLM_R_X3Y152_SLICE_X2Y152_CO5;
  wire [0:0] CLBLM_R_X3Y152_SLICE_X2Y152_CO6;
  wire [0:0] CLBLM_R_X3Y152_SLICE_X2Y152_C_CY;
  wire [0:0] CLBLM_R_X3Y152_SLICE_X2Y152_C_XOR;
  wire [0:0] CLBLM_R_X3Y152_SLICE_X2Y152_D;
  wire [0:0] CLBLM_R_X3Y152_SLICE_X2Y152_D1;
  wire [0:0] CLBLM_R_X3Y152_SLICE_X2Y152_D2;
  wire [0:0] CLBLM_R_X3Y152_SLICE_X2Y152_D3;
  wire [0:0] CLBLM_R_X3Y152_SLICE_X2Y152_D4;
  wire [0:0] CLBLM_R_X3Y152_SLICE_X2Y152_D5;
  wire [0:0] CLBLM_R_X3Y152_SLICE_X2Y152_D6;
  wire [0:0] CLBLM_R_X3Y152_SLICE_X2Y152_DO5;
  wire [0:0] CLBLM_R_X3Y152_SLICE_X2Y152_DO6;
  wire [0:0] CLBLM_R_X3Y152_SLICE_X2Y152_D_CY;
  wire [0:0] CLBLM_R_X3Y152_SLICE_X2Y152_D_XOR;
  wire [0:0] CLBLM_R_X3Y152_SLICE_X3Y152_A;
  wire [0:0] CLBLM_R_X3Y152_SLICE_X3Y152_A1;
  wire [0:0] CLBLM_R_X3Y152_SLICE_X3Y152_A2;
  wire [0:0] CLBLM_R_X3Y152_SLICE_X3Y152_A3;
  wire [0:0] CLBLM_R_X3Y152_SLICE_X3Y152_A4;
  wire [0:0] CLBLM_R_X3Y152_SLICE_X3Y152_A5;
  wire [0:0] CLBLM_R_X3Y152_SLICE_X3Y152_A6;
  wire [0:0] CLBLM_R_X3Y152_SLICE_X3Y152_AO5;
  wire [0:0] CLBLM_R_X3Y152_SLICE_X3Y152_AO6;
  wire [0:0] CLBLM_R_X3Y152_SLICE_X3Y152_AQ;
  wire [0:0] CLBLM_R_X3Y152_SLICE_X3Y152_A_CY;
  wire [0:0] CLBLM_R_X3Y152_SLICE_X3Y152_A_XOR;
  wire [0:0] CLBLM_R_X3Y152_SLICE_X3Y152_B;
  wire [0:0] CLBLM_R_X3Y152_SLICE_X3Y152_B1;
  wire [0:0] CLBLM_R_X3Y152_SLICE_X3Y152_B2;
  wire [0:0] CLBLM_R_X3Y152_SLICE_X3Y152_B3;
  wire [0:0] CLBLM_R_X3Y152_SLICE_X3Y152_B4;
  wire [0:0] CLBLM_R_X3Y152_SLICE_X3Y152_B5;
  wire [0:0] CLBLM_R_X3Y152_SLICE_X3Y152_B6;
  wire [0:0] CLBLM_R_X3Y152_SLICE_X3Y152_BO5;
  wire [0:0] CLBLM_R_X3Y152_SLICE_X3Y152_BO6;
  wire [0:0] CLBLM_R_X3Y152_SLICE_X3Y152_BQ;
  wire [0:0] CLBLM_R_X3Y152_SLICE_X3Y152_B_CY;
  wire [0:0] CLBLM_R_X3Y152_SLICE_X3Y152_B_XOR;
  wire [0:0] CLBLM_R_X3Y152_SLICE_X3Y152_C;
  wire [0:0] CLBLM_R_X3Y152_SLICE_X3Y152_C1;
  wire [0:0] CLBLM_R_X3Y152_SLICE_X3Y152_C2;
  wire [0:0] CLBLM_R_X3Y152_SLICE_X3Y152_C3;
  wire [0:0] CLBLM_R_X3Y152_SLICE_X3Y152_C4;
  wire [0:0] CLBLM_R_X3Y152_SLICE_X3Y152_C5;
  wire [0:0] CLBLM_R_X3Y152_SLICE_X3Y152_C6;
  wire [0:0] CLBLM_R_X3Y152_SLICE_X3Y152_CLK;
  wire [0:0] CLBLM_R_X3Y152_SLICE_X3Y152_CO5;
  wire [0:0] CLBLM_R_X3Y152_SLICE_X3Y152_CO6;
  wire [0:0] CLBLM_R_X3Y152_SLICE_X3Y152_CQ;
  wire [0:0] CLBLM_R_X3Y152_SLICE_X3Y152_C_CY;
  wire [0:0] CLBLM_R_X3Y152_SLICE_X3Y152_C_XOR;
  wire [0:0] CLBLM_R_X3Y152_SLICE_X3Y152_D;
  wire [0:0] CLBLM_R_X3Y152_SLICE_X3Y152_D1;
  wire [0:0] CLBLM_R_X3Y152_SLICE_X3Y152_D2;
  wire [0:0] CLBLM_R_X3Y152_SLICE_X3Y152_D3;
  wire [0:0] CLBLM_R_X3Y152_SLICE_X3Y152_D4;
  wire [0:0] CLBLM_R_X3Y152_SLICE_X3Y152_D5;
  wire [0:0] CLBLM_R_X3Y152_SLICE_X3Y152_D6;
  wire [0:0] CLBLM_R_X3Y152_SLICE_X3Y152_DO5;
  wire [0:0] CLBLM_R_X3Y152_SLICE_X3Y152_DO6;
  wire [0:0] CLBLM_R_X3Y152_SLICE_X3Y152_D_CY;
  wire [0:0] CLBLM_R_X3Y152_SLICE_X3Y152_D_XOR;
  wire [0:0] CLBLM_R_X3Y153_SLICE_X2Y153_A;
  wire [0:0] CLBLM_R_X3Y153_SLICE_X2Y153_A1;
  wire [0:0] CLBLM_R_X3Y153_SLICE_X2Y153_A2;
  wire [0:0] CLBLM_R_X3Y153_SLICE_X2Y153_A3;
  wire [0:0] CLBLM_R_X3Y153_SLICE_X2Y153_A4;
  wire [0:0] CLBLM_R_X3Y153_SLICE_X2Y153_A5;
  wire [0:0] CLBLM_R_X3Y153_SLICE_X2Y153_A6;
  wire [0:0] CLBLM_R_X3Y153_SLICE_X2Y153_AO5;
  wire [0:0] CLBLM_R_X3Y153_SLICE_X2Y153_AO6;
  wire [0:0] CLBLM_R_X3Y153_SLICE_X2Y153_AQ;
  wire [0:0] CLBLM_R_X3Y153_SLICE_X2Y153_AX;
  wire [0:0] CLBLM_R_X3Y153_SLICE_X2Y153_A_CY;
  wire [0:0] CLBLM_R_X3Y153_SLICE_X2Y153_A_XOR;
  wire [0:0] CLBLM_R_X3Y153_SLICE_X2Y153_B;
  wire [0:0] CLBLM_R_X3Y153_SLICE_X2Y153_B1;
  wire [0:0] CLBLM_R_X3Y153_SLICE_X2Y153_B2;
  wire [0:0] CLBLM_R_X3Y153_SLICE_X2Y153_B3;
  wire [0:0] CLBLM_R_X3Y153_SLICE_X2Y153_B4;
  wire [0:0] CLBLM_R_X3Y153_SLICE_X2Y153_B5;
  wire [0:0] CLBLM_R_X3Y153_SLICE_X2Y153_B6;
  wire [0:0] CLBLM_R_X3Y153_SLICE_X2Y153_BO5;
  wire [0:0] CLBLM_R_X3Y153_SLICE_X2Y153_BO6;
  wire [0:0] CLBLM_R_X3Y153_SLICE_X2Y153_B_CY;
  wire [0:0] CLBLM_R_X3Y153_SLICE_X2Y153_B_XOR;
  wire [0:0] CLBLM_R_X3Y153_SLICE_X2Y153_C;
  wire [0:0] CLBLM_R_X3Y153_SLICE_X2Y153_C1;
  wire [0:0] CLBLM_R_X3Y153_SLICE_X2Y153_C2;
  wire [0:0] CLBLM_R_X3Y153_SLICE_X2Y153_C3;
  wire [0:0] CLBLM_R_X3Y153_SLICE_X2Y153_C4;
  wire [0:0] CLBLM_R_X3Y153_SLICE_X2Y153_C5;
  wire [0:0] CLBLM_R_X3Y153_SLICE_X2Y153_C6;
  wire [0:0] CLBLM_R_X3Y153_SLICE_X2Y153_CLK;
  wire [0:0] CLBLM_R_X3Y153_SLICE_X2Y153_CO5;
  wire [0:0] CLBLM_R_X3Y153_SLICE_X2Y153_CO6;
  wire [0:0] CLBLM_R_X3Y153_SLICE_X2Y153_C_CY;
  wire [0:0] CLBLM_R_X3Y153_SLICE_X2Y153_C_XOR;
  wire [0:0] CLBLM_R_X3Y153_SLICE_X2Y153_D;
  wire [0:0] CLBLM_R_X3Y153_SLICE_X2Y153_D1;
  wire [0:0] CLBLM_R_X3Y153_SLICE_X2Y153_D2;
  wire [0:0] CLBLM_R_X3Y153_SLICE_X2Y153_D3;
  wire [0:0] CLBLM_R_X3Y153_SLICE_X2Y153_D4;
  wire [0:0] CLBLM_R_X3Y153_SLICE_X2Y153_D5;
  wire [0:0] CLBLM_R_X3Y153_SLICE_X2Y153_D6;
  wire [0:0] CLBLM_R_X3Y153_SLICE_X2Y153_DO5;
  wire [0:0] CLBLM_R_X3Y153_SLICE_X2Y153_DO6;
  wire [0:0] CLBLM_R_X3Y153_SLICE_X2Y153_D_CY;
  wire [0:0] CLBLM_R_X3Y153_SLICE_X2Y153_D_XOR;
  wire [0:0] CLBLM_R_X3Y153_SLICE_X3Y153_A;
  wire [0:0] CLBLM_R_X3Y153_SLICE_X3Y153_A1;
  wire [0:0] CLBLM_R_X3Y153_SLICE_X3Y153_A2;
  wire [0:0] CLBLM_R_X3Y153_SLICE_X3Y153_A3;
  wire [0:0] CLBLM_R_X3Y153_SLICE_X3Y153_A4;
  wire [0:0] CLBLM_R_X3Y153_SLICE_X3Y153_A5;
  wire [0:0] CLBLM_R_X3Y153_SLICE_X3Y153_A6;
  wire [0:0] CLBLM_R_X3Y153_SLICE_X3Y153_AO5;
  wire [0:0] CLBLM_R_X3Y153_SLICE_X3Y153_AO6;
  wire [0:0] CLBLM_R_X3Y153_SLICE_X3Y153_A_CY;
  wire [0:0] CLBLM_R_X3Y153_SLICE_X3Y153_A_XOR;
  wire [0:0] CLBLM_R_X3Y153_SLICE_X3Y153_B;
  wire [0:0] CLBLM_R_X3Y153_SLICE_X3Y153_B1;
  wire [0:0] CLBLM_R_X3Y153_SLICE_X3Y153_B2;
  wire [0:0] CLBLM_R_X3Y153_SLICE_X3Y153_B3;
  wire [0:0] CLBLM_R_X3Y153_SLICE_X3Y153_B4;
  wire [0:0] CLBLM_R_X3Y153_SLICE_X3Y153_B5;
  wire [0:0] CLBLM_R_X3Y153_SLICE_X3Y153_B6;
  wire [0:0] CLBLM_R_X3Y153_SLICE_X3Y153_BO5;
  wire [0:0] CLBLM_R_X3Y153_SLICE_X3Y153_BO6;
  wire [0:0] CLBLM_R_X3Y153_SLICE_X3Y153_B_CY;
  wire [0:0] CLBLM_R_X3Y153_SLICE_X3Y153_B_XOR;
  wire [0:0] CLBLM_R_X3Y153_SLICE_X3Y153_C;
  wire [0:0] CLBLM_R_X3Y153_SLICE_X3Y153_C1;
  wire [0:0] CLBLM_R_X3Y153_SLICE_X3Y153_C2;
  wire [0:0] CLBLM_R_X3Y153_SLICE_X3Y153_C3;
  wire [0:0] CLBLM_R_X3Y153_SLICE_X3Y153_C4;
  wire [0:0] CLBLM_R_X3Y153_SLICE_X3Y153_C5;
  wire [0:0] CLBLM_R_X3Y153_SLICE_X3Y153_C6;
  wire [0:0] CLBLM_R_X3Y153_SLICE_X3Y153_CO5;
  wire [0:0] CLBLM_R_X3Y153_SLICE_X3Y153_CO6;
  wire [0:0] CLBLM_R_X3Y153_SLICE_X3Y153_C_CY;
  wire [0:0] CLBLM_R_X3Y153_SLICE_X3Y153_C_XOR;
  wire [0:0] CLBLM_R_X3Y153_SLICE_X3Y153_D;
  wire [0:0] CLBLM_R_X3Y153_SLICE_X3Y153_D1;
  wire [0:0] CLBLM_R_X3Y153_SLICE_X3Y153_D2;
  wire [0:0] CLBLM_R_X3Y153_SLICE_X3Y153_D3;
  wire [0:0] CLBLM_R_X3Y153_SLICE_X3Y153_D4;
  wire [0:0] CLBLM_R_X3Y153_SLICE_X3Y153_D5;
  wire [0:0] CLBLM_R_X3Y153_SLICE_X3Y153_D6;
  wire [0:0] CLBLM_R_X3Y153_SLICE_X3Y153_DO5;
  wire [0:0] CLBLM_R_X3Y153_SLICE_X3Y153_DO6;
  wire [0:0] CLBLM_R_X3Y153_SLICE_X3Y153_D_CY;
  wire [0:0] CLBLM_R_X3Y153_SLICE_X3Y153_D_XOR;
  wire [0:0] CLBLM_R_X5Y140_SLICE_X6Y140_A;
  wire [0:0] CLBLM_R_X5Y140_SLICE_X6Y140_A1;
  wire [0:0] CLBLM_R_X5Y140_SLICE_X6Y140_A2;
  wire [0:0] CLBLM_R_X5Y140_SLICE_X6Y140_A3;
  wire [0:0] CLBLM_R_X5Y140_SLICE_X6Y140_A4;
  wire [0:0] CLBLM_R_X5Y140_SLICE_X6Y140_A5;
  wire [0:0] CLBLM_R_X5Y140_SLICE_X6Y140_A5Q;
  wire [0:0] CLBLM_R_X5Y140_SLICE_X6Y140_A6;
  wire [0:0] CLBLM_R_X5Y140_SLICE_X6Y140_AMUX;
  wire [0:0] CLBLM_R_X5Y140_SLICE_X6Y140_AO5;
  wire [0:0] CLBLM_R_X5Y140_SLICE_X6Y140_AO6;
  wire [0:0] CLBLM_R_X5Y140_SLICE_X6Y140_AQ;
  wire [0:0] CLBLM_R_X5Y140_SLICE_X6Y140_AX;
  wire [0:0] CLBLM_R_X5Y140_SLICE_X6Y140_A_CY;
  wire [0:0] CLBLM_R_X5Y140_SLICE_X6Y140_A_XOR;
  wire [0:0] CLBLM_R_X5Y140_SLICE_X6Y140_B;
  wire [0:0] CLBLM_R_X5Y140_SLICE_X6Y140_B1;
  wire [0:0] CLBLM_R_X5Y140_SLICE_X6Y140_B2;
  wire [0:0] CLBLM_R_X5Y140_SLICE_X6Y140_B3;
  wire [0:0] CLBLM_R_X5Y140_SLICE_X6Y140_B4;
  wire [0:0] CLBLM_R_X5Y140_SLICE_X6Y140_B5;
  wire [0:0] CLBLM_R_X5Y140_SLICE_X6Y140_B6;
  wire [0:0] CLBLM_R_X5Y140_SLICE_X6Y140_BO5;
  wire [0:0] CLBLM_R_X5Y140_SLICE_X6Y140_BO6;
  wire [0:0] CLBLM_R_X5Y140_SLICE_X6Y140_BQ;
  wire [0:0] CLBLM_R_X5Y140_SLICE_X6Y140_B_CY;
  wire [0:0] CLBLM_R_X5Y140_SLICE_X6Y140_B_XOR;
  wire [0:0] CLBLM_R_X5Y140_SLICE_X6Y140_C;
  wire [0:0] CLBLM_R_X5Y140_SLICE_X6Y140_C1;
  wire [0:0] CLBLM_R_X5Y140_SLICE_X6Y140_C2;
  wire [0:0] CLBLM_R_X5Y140_SLICE_X6Y140_C3;
  wire [0:0] CLBLM_R_X5Y140_SLICE_X6Y140_C4;
  wire [0:0] CLBLM_R_X5Y140_SLICE_X6Y140_C5;
  wire [0:0] CLBLM_R_X5Y140_SLICE_X6Y140_C6;
  wire [0:0] CLBLM_R_X5Y140_SLICE_X6Y140_CLK;
  wire [0:0] CLBLM_R_X5Y140_SLICE_X6Y140_CO5;
  wire [0:0] CLBLM_R_X5Y140_SLICE_X6Y140_CO6;
  wire [0:0] CLBLM_R_X5Y140_SLICE_X6Y140_CQ;
  wire [0:0] CLBLM_R_X5Y140_SLICE_X6Y140_C_CY;
  wire [0:0] CLBLM_R_X5Y140_SLICE_X6Y140_C_XOR;
  wire [0:0] CLBLM_R_X5Y140_SLICE_X6Y140_D;
  wire [0:0] CLBLM_R_X5Y140_SLICE_X6Y140_D1;
  wire [0:0] CLBLM_R_X5Y140_SLICE_X6Y140_D2;
  wire [0:0] CLBLM_R_X5Y140_SLICE_X6Y140_D3;
  wire [0:0] CLBLM_R_X5Y140_SLICE_X6Y140_D4;
  wire [0:0] CLBLM_R_X5Y140_SLICE_X6Y140_D5;
  wire [0:0] CLBLM_R_X5Y140_SLICE_X6Y140_D6;
  wire [0:0] CLBLM_R_X5Y140_SLICE_X6Y140_DMUX;
  wire [0:0] CLBLM_R_X5Y140_SLICE_X6Y140_DO5;
  wire [0:0] CLBLM_R_X5Y140_SLICE_X6Y140_DO6;
  wire [0:0] CLBLM_R_X5Y140_SLICE_X6Y140_D_CY;
  wire [0:0] CLBLM_R_X5Y140_SLICE_X6Y140_D_XOR;
  wire [0:0] CLBLM_R_X5Y140_SLICE_X7Y140_A;
  wire [0:0] CLBLM_R_X5Y140_SLICE_X7Y140_A1;
  wire [0:0] CLBLM_R_X5Y140_SLICE_X7Y140_A2;
  wire [0:0] CLBLM_R_X5Y140_SLICE_X7Y140_A3;
  wire [0:0] CLBLM_R_X5Y140_SLICE_X7Y140_A4;
  wire [0:0] CLBLM_R_X5Y140_SLICE_X7Y140_A5;
  wire [0:0] CLBLM_R_X5Y140_SLICE_X7Y140_A6;
  wire [0:0] CLBLM_R_X5Y140_SLICE_X7Y140_AO5;
  wire [0:0] CLBLM_R_X5Y140_SLICE_X7Y140_AO6;
  wire [0:0] CLBLM_R_X5Y140_SLICE_X7Y140_A_CY;
  wire [0:0] CLBLM_R_X5Y140_SLICE_X7Y140_A_XOR;
  wire [0:0] CLBLM_R_X5Y140_SLICE_X7Y140_B;
  wire [0:0] CLBLM_R_X5Y140_SLICE_X7Y140_B1;
  wire [0:0] CLBLM_R_X5Y140_SLICE_X7Y140_B2;
  wire [0:0] CLBLM_R_X5Y140_SLICE_X7Y140_B3;
  wire [0:0] CLBLM_R_X5Y140_SLICE_X7Y140_B4;
  wire [0:0] CLBLM_R_X5Y140_SLICE_X7Y140_B5;
  wire [0:0] CLBLM_R_X5Y140_SLICE_X7Y140_B6;
  wire [0:0] CLBLM_R_X5Y140_SLICE_X7Y140_BO5;
  wire [0:0] CLBLM_R_X5Y140_SLICE_X7Y140_BO6;
  wire [0:0] CLBLM_R_X5Y140_SLICE_X7Y140_B_CY;
  wire [0:0] CLBLM_R_X5Y140_SLICE_X7Y140_B_XOR;
  wire [0:0] CLBLM_R_X5Y140_SLICE_X7Y140_C;
  wire [0:0] CLBLM_R_X5Y140_SLICE_X7Y140_C1;
  wire [0:0] CLBLM_R_X5Y140_SLICE_X7Y140_C2;
  wire [0:0] CLBLM_R_X5Y140_SLICE_X7Y140_C3;
  wire [0:0] CLBLM_R_X5Y140_SLICE_X7Y140_C4;
  wire [0:0] CLBLM_R_X5Y140_SLICE_X7Y140_C5;
  wire [0:0] CLBLM_R_X5Y140_SLICE_X7Y140_C6;
  wire [0:0] CLBLM_R_X5Y140_SLICE_X7Y140_CO5;
  wire [0:0] CLBLM_R_X5Y140_SLICE_X7Y140_CO6;
  wire [0:0] CLBLM_R_X5Y140_SLICE_X7Y140_C_CY;
  wire [0:0] CLBLM_R_X5Y140_SLICE_X7Y140_C_XOR;
  wire [0:0] CLBLM_R_X5Y140_SLICE_X7Y140_D;
  wire [0:0] CLBLM_R_X5Y140_SLICE_X7Y140_D1;
  wire [0:0] CLBLM_R_X5Y140_SLICE_X7Y140_D2;
  wire [0:0] CLBLM_R_X5Y140_SLICE_X7Y140_D3;
  wire [0:0] CLBLM_R_X5Y140_SLICE_X7Y140_D4;
  wire [0:0] CLBLM_R_X5Y140_SLICE_X7Y140_D5;
  wire [0:0] CLBLM_R_X5Y140_SLICE_X7Y140_D6;
  wire [0:0] CLBLM_R_X5Y140_SLICE_X7Y140_DO5;
  wire [0:0] CLBLM_R_X5Y140_SLICE_X7Y140_DO6;
  wire [0:0] CLBLM_R_X5Y140_SLICE_X7Y140_D_CY;
  wire [0:0] CLBLM_R_X5Y140_SLICE_X7Y140_D_XOR;
  wire [0:0] CLBLM_R_X5Y141_SLICE_X6Y141_A;
  wire [0:0] CLBLM_R_X5Y141_SLICE_X6Y141_A1;
  wire [0:0] CLBLM_R_X5Y141_SLICE_X6Y141_A2;
  wire [0:0] CLBLM_R_X5Y141_SLICE_X6Y141_A3;
  wire [0:0] CLBLM_R_X5Y141_SLICE_X6Y141_A4;
  wire [0:0] CLBLM_R_X5Y141_SLICE_X6Y141_A5;
  wire [0:0] CLBLM_R_X5Y141_SLICE_X6Y141_A6;
  wire [0:0] CLBLM_R_X5Y141_SLICE_X6Y141_AO5;
  wire [0:0] CLBLM_R_X5Y141_SLICE_X6Y141_AO6;
  wire [0:0] CLBLM_R_X5Y141_SLICE_X6Y141_AQ;
  wire [0:0] CLBLM_R_X5Y141_SLICE_X6Y141_A_CY;
  wire [0:0] CLBLM_R_X5Y141_SLICE_X6Y141_A_XOR;
  wire [0:0] CLBLM_R_X5Y141_SLICE_X6Y141_B;
  wire [0:0] CLBLM_R_X5Y141_SLICE_X6Y141_B1;
  wire [0:0] CLBLM_R_X5Y141_SLICE_X6Y141_B2;
  wire [0:0] CLBLM_R_X5Y141_SLICE_X6Y141_B3;
  wire [0:0] CLBLM_R_X5Y141_SLICE_X6Y141_B4;
  wire [0:0] CLBLM_R_X5Y141_SLICE_X6Y141_B5;
  wire [0:0] CLBLM_R_X5Y141_SLICE_X6Y141_B5Q;
  wire [0:0] CLBLM_R_X5Y141_SLICE_X6Y141_B6;
  wire [0:0] CLBLM_R_X5Y141_SLICE_X6Y141_BMUX;
  wire [0:0] CLBLM_R_X5Y141_SLICE_X6Y141_BO5;
  wire [0:0] CLBLM_R_X5Y141_SLICE_X6Y141_BO6;
  wire [0:0] CLBLM_R_X5Y141_SLICE_X6Y141_BQ;
  wire [0:0] CLBLM_R_X5Y141_SLICE_X6Y141_B_CY;
  wire [0:0] CLBLM_R_X5Y141_SLICE_X6Y141_B_XOR;
  wire [0:0] CLBLM_R_X5Y141_SLICE_X6Y141_C;
  wire [0:0] CLBLM_R_X5Y141_SLICE_X6Y141_C1;
  wire [0:0] CLBLM_R_X5Y141_SLICE_X6Y141_C2;
  wire [0:0] CLBLM_R_X5Y141_SLICE_X6Y141_C3;
  wire [0:0] CLBLM_R_X5Y141_SLICE_X6Y141_C4;
  wire [0:0] CLBLM_R_X5Y141_SLICE_X6Y141_C5;
  wire [0:0] CLBLM_R_X5Y141_SLICE_X6Y141_C6;
  wire [0:0] CLBLM_R_X5Y141_SLICE_X6Y141_CLK;
  wire [0:0] CLBLM_R_X5Y141_SLICE_X6Y141_CMUX;
  wire [0:0] CLBLM_R_X5Y141_SLICE_X6Y141_CO5;
  wire [0:0] CLBLM_R_X5Y141_SLICE_X6Y141_CO6;
  wire [0:0] CLBLM_R_X5Y141_SLICE_X6Y141_C_CY;
  wire [0:0] CLBLM_R_X5Y141_SLICE_X6Y141_C_XOR;
  wire [0:0] CLBLM_R_X5Y141_SLICE_X6Y141_D;
  wire [0:0] CLBLM_R_X5Y141_SLICE_X6Y141_D1;
  wire [0:0] CLBLM_R_X5Y141_SLICE_X6Y141_D2;
  wire [0:0] CLBLM_R_X5Y141_SLICE_X6Y141_D3;
  wire [0:0] CLBLM_R_X5Y141_SLICE_X6Y141_D4;
  wire [0:0] CLBLM_R_X5Y141_SLICE_X6Y141_D5;
  wire [0:0] CLBLM_R_X5Y141_SLICE_X6Y141_D5Q;
  wire [0:0] CLBLM_R_X5Y141_SLICE_X6Y141_D6;
  wire [0:0] CLBLM_R_X5Y141_SLICE_X6Y141_DMUX;
  wire [0:0] CLBLM_R_X5Y141_SLICE_X6Y141_DO5;
  wire [0:0] CLBLM_R_X5Y141_SLICE_X6Y141_DO6;
  wire [0:0] CLBLM_R_X5Y141_SLICE_X6Y141_DQ;
  wire [0:0] CLBLM_R_X5Y141_SLICE_X6Y141_D_CY;
  wire [0:0] CLBLM_R_X5Y141_SLICE_X6Y141_D_XOR;
  wire [0:0] CLBLM_R_X5Y141_SLICE_X7Y141_A;
  wire [0:0] CLBLM_R_X5Y141_SLICE_X7Y141_A1;
  wire [0:0] CLBLM_R_X5Y141_SLICE_X7Y141_A2;
  wire [0:0] CLBLM_R_X5Y141_SLICE_X7Y141_A3;
  wire [0:0] CLBLM_R_X5Y141_SLICE_X7Y141_A4;
  wire [0:0] CLBLM_R_X5Y141_SLICE_X7Y141_A5;
  wire [0:0] CLBLM_R_X5Y141_SLICE_X7Y141_A6;
  wire [0:0] CLBLM_R_X5Y141_SLICE_X7Y141_AO5;
  wire [0:0] CLBLM_R_X5Y141_SLICE_X7Y141_AO6;
  wire [0:0] CLBLM_R_X5Y141_SLICE_X7Y141_A_CY;
  wire [0:0] CLBLM_R_X5Y141_SLICE_X7Y141_A_XOR;
  wire [0:0] CLBLM_R_X5Y141_SLICE_X7Y141_B;
  wire [0:0] CLBLM_R_X5Y141_SLICE_X7Y141_B1;
  wire [0:0] CLBLM_R_X5Y141_SLICE_X7Y141_B2;
  wire [0:0] CLBLM_R_X5Y141_SLICE_X7Y141_B3;
  wire [0:0] CLBLM_R_X5Y141_SLICE_X7Y141_B4;
  wire [0:0] CLBLM_R_X5Y141_SLICE_X7Y141_B5;
  wire [0:0] CLBLM_R_X5Y141_SLICE_X7Y141_B6;
  wire [0:0] CLBLM_R_X5Y141_SLICE_X7Y141_BO5;
  wire [0:0] CLBLM_R_X5Y141_SLICE_X7Y141_BO6;
  wire [0:0] CLBLM_R_X5Y141_SLICE_X7Y141_B_CY;
  wire [0:0] CLBLM_R_X5Y141_SLICE_X7Y141_B_XOR;
  wire [0:0] CLBLM_R_X5Y141_SLICE_X7Y141_C;
  wire [0:0] CLBLM_R_X5Y141_SLICE_X7Y141_C1;
  wire [0:0] CLBLM_R_X5Y141_SLICE_X7Y141_C2;
  wire [0:0] CLBLM_R_X5Y141_SLICE_X7Y141_C3;
  wire [0:0] CLBLM_R_X5Y141_SLICE_X7Y141_C4;
  wire [0:0] CLBLM_R_X5Y141_SLICE_X7Y141_C5;
  wire [0:0] CLBLM_R_X5Y141_SLICE_X7Y141_C6;
  wire [0:0] CLBLM_R_X5Y141_SLICE_X7Y141_CO5;
  wire [0:0] CLBLM_R_X5Y141_SLICE_X7Y141_CO6;
  wire [0:0] CLBLM_R_X5Y141_SLICE_X7Y141_C_CY;
  wire [0:0] CLBLM_R_X5Y141_SLICE_X7Y141_C_XOR;
  wire [0:0] CLBLM_R_X5Y141_SLICE_X7Y141_D;
  wire [0:0] CLBLM_R_X5Y141_SLICE_X7Y141_D1;
  wire [0:0] CLBLM_R_X5Y141_SLICE_X7Y141_D2;
  wire [0:0] CLBLM_R_X5Y141_SLICE_X7Y141_D3;
  wire [0:0] CLBLM_R_X5Y141_SLICE_X7Y141_D4;
  wire [0:0] CLBLM_R_X5Y141_SLICE_X7Y141_D5;
  wire [0:0] CLBLM_R_X5Y141_SLICE_X7Y141_D6;
  wire [0:0] CLBLM_R_X5Y141_SLICE_X7Y141_DO5;
  wire [0:0] CLBLM_R_X5Y141_SLICE_X7Y141_DO6;
  wire [0:0] CLBLM_R_X5Y141_SLICE_X7Y141_D_CY;
  wire [0:0] CLBLM_R_X5Y141_SLICE_X7Y141_D_XOR;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X6Y142_A;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X6Y142_A1;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X6Y142_A2;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X6Y142_A3;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X6Y142_A4;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X6Y142_A5;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X6Y142_A6;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X6Y142_AO5;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X6Y142_AO6;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X6Y142_AQ;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X6Y142_A_CY;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X6Y142_A_XOR;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X6Y142_B;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X6Y142_B1;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X6Y142_B2;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X6Y142_B3;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X6Y142_B4;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X6Y142_B5;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X6Y142_B6;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X6Y142_BO5;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X6Y142_BO6;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X6Y142_BQ;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X6Y142_B_CY;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X6Y142_B_XOR;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X6Y142_C;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X6Y142_C1;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X6Y142_C2;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X6Y142_C3;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X6Y142_C4;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X6Y142_C5;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X6Y142_C6;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X6Y142_CLK;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X6Y142_CO5;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X6Y142_CO6;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X6Y142_CQ;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X6Y142_C_CY;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X6Y142_C_XOR;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X6Y142_D;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X6Y142_D1;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X6Y142_D2;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X6Y142_D3;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X6Y142_D4;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X6Y142_D5;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X6Y142_D5Q;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X6Y142_D6;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X6Y142_DMUX;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X6Y142_DO5;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X6Y142_DO6;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X6Y142_DQ;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X6Y142_D_CY;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X6Y142_D_XOR;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X7Y142_A;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X7Y142_A1;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X7Y142_A2;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X7Y142_A3;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X7Y142_A4;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X7Y142_A5;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X7Y142_A5Q;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X7Y142_A6;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X7Y142_AMUX;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X7Y142_AO5;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X7Y142_AO6;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X7Y142_AQ;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X7Y142_A_CY;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X7Y142_A_XOR;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X7Y142_B;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X7Y142_B1;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X7Y142_B2;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X7Y142_B3;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X7Y142_B4;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X7Y142_B5;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X7Y142_B6;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X7Y142_BO5;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X7Y142_BO6;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X7Y142_BQ;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X7Y142_BX;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X7Y142_B_CY;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X7Y142_B_XOR;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X7Y142_C;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X7Y142_C1;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X7Y142_C2;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X7Y142_C3;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X7Y142_C4;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X7Y142_C5;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X7Y142_C6;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X7Y142_CLK;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X7Y142_CO5;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X7Y142_CO6;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X7Y142_C_CY;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X7Y142_C_XOR;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X7Y142_D;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X7Y142_D1;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X7Y142_D2;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X7Y142_D3;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X7Y142_D4;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X7Y142_D5;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X7Y142_D6;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X7Y142_DO5;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X7Y142_DO6;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X7Y142_D_CY;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X7Y142_D_XOR;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X6Y143_A;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X6Y143_A1;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X6Y143_A2;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X6Y143_A3;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X6Y143_A4;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X6Y143_A5;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X6Y143_A6;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X6Y143_AO5;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X6Y143_AO6;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X6Y143_AQ;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X6Y143_A_CY;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X6Y143_A_XOR;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X6Y143_B;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X6Y143_B1;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X6Y143_B2;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X6Y143_B3;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X6Y143_B4;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X6Y143_B5;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X6Y143_B6;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X6Y143_BO5;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X6Y143_BO6;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X6Y143_BQ;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X6Y143_B_CY;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X6Y143_B_XOR;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X6Y143_C;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X6Y143_C1;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X6Y143_C2;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X6Y143_C3;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X6Y143_C4;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X6Y143_C5;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X6Y143_C5Q;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X6Y143_C6;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X6Y143_CLK;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X6Y143_CMUX;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X6Y143_CO5;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X6Y143_CO6;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X6Y143_CQ;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X6Y143_C_CY;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X6Y143_C_XOR;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X6Y143_D;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X6Y143_D1;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X6Y143_D2;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X6Y143_D3;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X6Y143_D4;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X6Y143_D5;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X6Y143_D5Q;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X6Y143_D6;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X6Y143_DMUX;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X6Y143_DO5;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X6Y143_DO6;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X6Y143_DQ;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X6Y143_D_CY;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X6Y143_D_XOR;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X7Y143_A;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X7Y143_A1;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X7Y143_A2;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X7Y143_A3;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X7Y143_A4;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X7Y143_A5;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X7Y143_A6;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X7Y143_AO5;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X7Y143_AO6;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X7Y143_AQ;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X7Y143_A_CY;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X7Y143_A_XOR;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X7Y143_B;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X7Y143_B1;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X7Y143_B2;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X7Y143_B3;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X7Y143_B4;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X7Y143_B5;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X7Y143_B6;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X7Y143_BO5;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X7Y143_BO6;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X7Y143_BQ;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X7Y143_B_CY;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X7Y143_B_XOR;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X7Y143_C;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X7Y143_C1;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X7Y143_C2;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X7Y143_C3;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X7Y143_C4;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X7Y143_C5;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X7Y143_C5Q;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X7Y143_C6;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X7Y143_CLK;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X7Y143_CMUX;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X7Y143_CO5;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X7Y143_CO6;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X7Y143_CQ;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X7Y143_C_CY;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X7Y143_C_XOR;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X7Y143_D;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X7Y143_D1;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X7Y143_D2;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X7Y143_D3;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X7Y143_D4;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X7Y143_D5;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X7Y143_D6;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X7Y143_DMUX;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X7Y143_DO5;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X7Y143_DO6;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X7Y143_D_CY;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X7Y143_D_XOR;
  wire [0:0] CLBLM_R_X5Y144_SLICE_X6Y144_A;
  wire [0:0] CLBLM_R_X5Y144_SLICE_X6Y144_A1;
  wire [0:0] CLBLM_R_X5Y144_SLICE_X6Y144_A2;
  wire [0:0] CLBLM_R_X5Y144_SLICE_X6Y144_A3;
  wire [0:0] CLBLM_R_X5Y144_SLICE_X6Y144_A4;
  wire [0:0] CLBLM_R_X5Y144_SLICE_X6Y144_A5;
  wire [0:0] CLBLM_R_X5Y144_SLICE_X6Y144_A6;
  wire [0:0] CLBLM_R_X5Y144_SLICE_X6Y144_AO5;
  wire [0:0] CLBLM_R_X5Y144_SLICE_X6Y144_AO6;
  wire [0:0] CLBLM_R_X5Y144_SLICE_X6Y144_AQ;
  wire [0:0] CLBLM_R_X5Y144_SLICE_X6Y144_A_CY;
  wire [0:0] CLBLM_R_X5Y144_SLICE_X6Y144_A_XOR;
  wire [0:0] CLBLM_R_X5Y144_SLICE_X6Y144_B;
  wire [0:0] CLBLM_R_X5Y144_SLICE_X6Y144_B1;
  wire [0:0] CLBLM_R_X5Y144_SLICE_X6Y144_B2;
  wire [0:0] CLBLM_R_X5Y144_SLICE_X6Y144_B3;
  wire [0:0] CLBLM_R_X5Y144_SLICE_X6Y144_B4;
  wire [0:0] CLBLM_R_X5Y144_SLICE_X6Y144_B5;
  wire [0:0] CLBLM_R_X5Y144_SLICE_X6Y144_B6;
  wire [0:0] CLBLM_R_X5Y144_SLICE_X6Y144_BO5;
  wire [0:0] CLBLM_R_X5Y144_SLICE_X6Y144_BO6;
  wire [0:0] CLBLM_R_X5Y144_SLICE_X6Y144_BQ;
  wire [0:0] CLBLM_R_X5Y144_SLICE_X6Y144_B_CY;
  wire [0:0] CLBLM_R_X5Y144_SLICE_X6Y144_B_XOR;
  wire [0:0] CLBLM_R_X5Y144_SLICE_X6Y144_C;
  wire [0:0] CLBLM_R_X5Y144_SLICE_X6Y144_C1;
  wire [0:0] CLBLM_R_X5Y144_SLICE_X6Y144_C2;
  wire [0:0] CLBLM_R_X5Y144_SLICE_X6Y144_C3;
  wire [0:0] CLBLM_R_X5Y144_SLICE_X6Y144_C4;
  wire [0:0] CLBLM_R_X5Y144_SLICE_X6Y144_C5;
  wire [0:0] CLBLM_R_X5Y144_SLICE_X6Y144_C6;
  wire [0:0] CLBLM_R_X5Y144_SLICE_X6Y144_CLK;
  wire [0:0] CLBLM_R_X5Y144_SLICE_X6Y144_CO5;
  wire [0:0] CLBLM_R_X5Y144_SLICE_X6Y144_CO6;
  wire [0:0] CLBLM_R_X5Y144_SLICE_X6Y144_CQ;
  wire [0:0] CLBLM_R_X5Y144_SLICE_X6Y144_C_CY;
  wire [0:0] CLBLM_R_X5Y144_SLICE_X6Y144_C_XOR;
  wire [0:0] CLBLM_R_X5Y144_SLICE_X6Y144_D;
  wire [0:0] CLBLM_R_X5Y144_SLICE_X6Y144_D1;
  wire [0:0] CLBLM_R_X5Y144_SLICE_X6Y144_D2;
  wire [0:0] CLBLM_R_X5Y144_SLICE_X6Y144_D3;
  wire [0:0] CLBLM_R_X5Y144_SLICE_X6Y144_D4;
  wire [0:0] CLBLM_R_X5Y144_SLICE_X6Y144_D5;
  wire [0:0] CLBLM_R_X5Y144_SLICE_X6Y144_D5Q;
  wire [0:0] CLBLM_R_X5Y144_SLICE_X6Y144_D6;
  wire [0:0] CLBLM_R_X5Y144_SLICE_X6Y144_DMUX;
  wire [0:0] CLBLM_R_X5Y144_SLICE_X6Y144_DO5;
  wire [0:0] CLBLM_R_X5Y144_SLICE_X6Y144_DO6;
  wire [0:0] CLBLM_R_X5Y144_SLICE_X6Y144_DQ;
  wire [0:0] CLBLM_R_X5Y144_SLICE_X6Y144_D_CY;
  wire [0:0] CLBLM_R_X5Y144_SLICE_X6Y144_D_XOR;
  wire [0:0] CLBLM_R_X5Y144_SLICE_X7Y144_A;
  wire [0:0] CLBLM_R_X5Y144_SLICE_X7Y144_A1;
  wire [0:0] CLBLM_R_X5Y144_SLICE_X7Y144_A2;
  wire [0:0] CLBLM_R_X5Y144_SLICE_X7Y144_A3;
  wire [0:0] CLBLM_R_X5Y144_SLICE_X7Y144_A4;
  wire [0:0] CLBLM_R_X5Y144_SLICE_X7Y144_A5;
  wire [0:0] CLBLM_R_X5Y144_SLICE_X7Y144_A6;
  wire [0:0] CLBLM_R_X5Y144_SLICE_X7Y144_AO5;
  wire [0:0] CLBLM_R_X5Y144_SLICE_X7Y144_AO6;
  wire [0:0] CLBLM_R_X5Y144_SLICE_X7Y144_AQ;
  wire [0:0] CLBLM_R_X5Y144_SLICE_X7Y144_A_CY;
  wire [0:0] CLBLM_R_X5Y144_SLICE_X7Y144_A_XOR;
  wire [0:0] CLBLM_R_X5Y144_SLICE_X7Y144_B;
  wire [0:0] CLBLM_R_X5Y144_SLICE_X7Y144_B1;
  wire [0:0] CLBLM_R_X5Y144_SLICE_X7Y144_B2;
  wire [0:0] CLBLM_R_X5Y144_SLICE_X7Y144_B3;
  wire [0:0] CLBLM_R_X5Y144_SLICE_X7Y144_B4;
  wire [0:0] CLBLM_R_X5Y144_SLICE_X7Y144_B5;
  wire [0:0] CLBLM_R_X5Y144_SLICE_X7Y144_B5Q;
  wire [0:0] CLBLM_R_X5Y144_SLICE_X7Y144_B6;
  wire [0:0] CLBLM_R_X5Y144_SLICE_X7Y144_BMUX;
  wire [0:0] CLBLM_R_X5Y144_SLICE_X7Y144_BO5;
  wire [0:0] CLBLM_R_X5Y144_SLICE_X7Y144_BO6;
  wire [0:0] CLBLM_R_X5Y144_SLICE_X7Y144_BQ;
  wire [0:0] CLBLM_R_X5Y144_SLICE_X7Y144_B_CY;
  wire [0:0] CLBLM_R_X5Y144_SLICE_X7Y144_B_XOR;
  wire [0:0] CLBLM_R_X5Y144_SLICE_X7Y144_C;
  wire [0:0] CLBLM_R_X5Y144_SLICE_X7Y144_C1;
  wire [0:0] CLBLM_R_X5Y144_SLICE_X7Y144_C2;
  wire [0:0] CLBLM_R_X5Y144_SLICE_X7Y144_C3;
  wire [0:0] CLBLM_R_X5Y144_SLICE_X7Y144_C4;
  wire [0:0] CLBLM_R_X5Y144_SLICE_X7Y144_C5;
  wire [0:0] CLBLM_R_X5Y144_SLICE_X7Y144_C5Q;
  wire [0:0] CLBLM_R_X5Y144_SLICE_X7Y144_C6;
  wire [0:0] CLBLM_R_X5Y144_SLICE_X7Y144_CLK;
  wire [0:0] CLBLM_R_X5Y144_SLICE_X7Y144_CMUX;
  wire [0:0] CLBLM_R_X5Y144_SLICE_X7Y144_CO5;
  wire [0:0] CLBLM_R_X5Y144_SLICE_X7Y144_CO6;
  wire [0:0] CLBLM_R_X5Y144_SLICE_X7Y144_CQ;
  wire [0:0] CLBLM_R_X5Y144_SLICE_X7Y144_C_CY;
  wire [0:0] CLBLM_R_X5Y144_SLICE_X7Y144_C_XOR;
  wire [0:0] CLBLM_R_X5Y144_SLICE_X7Y144_D;
  wire [0:0] CLBLM_R_X5Y144_SLICE_X7Y144_D1;
  wire [0:0] CLBLM_R_X5Y144_SLICE_X7Y144_D2;
  wire [0:0] CLBLM_R_X5Y144_SLICE_X7Y144_D3;
  wire [0:0] CLBLM_R_X5Y144_SLICE_X7Y144_D4;
  wire [0:0] CLBLM_R_X5Y144_SLICE_X7Y144_D5;
  wire [0:0] CLBLM_R_X5Y144_SLICE_X7Y144_D6;
  wire [0:0] CLBLM_R_X5Y144_SLICE_X7Y144_DMUX;
  wire [0:0] CLBLM_R_X5Y144_SLICE_X7Y144_DO5;
  wire [0:0] CLBLM_R_X5Y144_SLICE_X7Y144_DO6;
  wire [0:0] CLBLM_R_X5Y144_SLICE_X7Y144_D_CY;
  wire [0:0] CLBLM_R_X5Y144_SLICE_X7Y144_D_XOR;
  wire [0:0] CLBLM_R_X5Y145_SLICE_X6Y145_A;
  wire [0:0] CLBLM_R_X5Y145_SLICE_X6Y145_A1;
  wire [0:0] CLBLM_R_X5Y145_SLICE_X6Y145_A2;
  wire [0:0] CLBLM_R_X5Y145_SLICE_X6Y145_A3;
  wire [0:0] CLBLM_R_X5Y145_SLICE_X6Y145_A4;
  wire [0:0] CLBLM_R_X5Y145_SLICE_X6Y145_A5;
  wire [0:0] CLBLM_R_X5Y145_SLICE_X6Y145_A6;
  wire [0:0] CLBLM_R_X5Y145_SLICE_X6Y145_AO5;
  wire [0:0] CLBLM_R_X5Y145_SLICE_X6Y145_AO6;
  wire [0:0] CLBLM_R_X5Y145_SLICE_X6Y145_AQ;
  wire [0:0] CLBLM_R_X5Y145_SLICE_X6Y145_A_CY;
  wire [0:0] CLBLM_R_X5Y145_SLICE_X6Y145_A_XOR;
  wire [0:0] CLBLM_R_X5Y145_SLICE_X6Y145_B;
  wire [0:0] CLBLM_R_X5Y145_SLICE_X6Y145_B1;
  wire [0:0] CLBLM_R_X5Y145_SLICE_X6Y145_B2;
  wire [0:0] CLBLM_R_X5Y145_SLICE_X6Y145_B3;
  wire [0:0] CLBLM_R_X5Y145_SLICE_X6Y145_B4;
  wire [0:0] CLBLM_R_X5Y145_SLICE_X6Y145_B5;
  wire [0:0] CLBLM_R_X5Y145_SLICE_X6Y145_B5Q;
  wire [0:0] CLBLM_R_X5Y145_SLICE_X6Y145_B6;
  wire [0:0] CLBLM_R_X5Y145_SLICE_X6Y145_BMUX;
  wire [0:0] CLBLM_R_X5Y145_SLICE_X6Y145_BO5;
  wire [0:0] CLBLM_R_X5Y145_SLICE_X6Y145_BO6;
  wire [0:0] CLBLM_R_X5Y145_SLICE_X6Y145_BQ;
  wire [0:0] CLBLM_R_X5Y145_SLICE_X6Y145_B_CY;
  wire [0:0] CLBLM_R_X5Y145_SLICE_X6Y145_B_XOR;
  wire [0:0] CLBLM_R_X5Y145_SLICE_X6Y145_C;
  wire [0:0] CLBLM_R_X5Y145_SLICE_X6Y145_C1;
  wire [0:0] CLBLM_R_X5Y145_SLICE_X6Y145_C2;
  wire [0:0] CLBLM_R_X5Y145_SLICE_X6Y145_C3;
  wire [0:0] CLBLM_R_X5Y145_SLICE_X6Y145_C4;
  wire [0:0] CLBLM_R_X5Y145_SLICE_X6Y145_C5;
  wire [0:0] CLBLM_R_X5Y145_SLICE_X6Y145_C5Q;
  wire [0:0] CLBLM_R_X5Y145_SLICE_X6Y145_C6;
  wire [0:0] CLBLM_R_X5Y145_SLICE_X6Y145_CLK;
  wire [0:0] CLBLM_R_X5Y145_SLICE_X6Y145_CMUX;
  wire [0:0] CLBLM_R_X5Y145_SLICE_X6Y145_CO5;
  wire [0:0] CLBLM_R_X5Y145_SLICE_X6Y145_CO6;
  wire [0:0] CLBLM_R_X5Y145_SLICE_X6Y145_CQ;
  wire [0:0] CLBLM_R_X5Y145_SLICE_X6Y145_C_CY;
  wire [0:0] CLBLM_R_X5Y145_SLICE_X6Y145_C_XOR;
  wire [0:0] CLBLM_R_X5Y145_SLICE_X6Y145_D;
  wire [0:0] CLBLM_R_X5Y145_SLICE_X6Y145_D1;
  wire [0:0] CLBLM_R_X5Y145_SLICE_X6Y145_D2;
  wire [0:0] CLBLM_R_X5Y145_SLICE_X6Y145_D3;
  wire [0:0] CLBLM_R_X5Y145_SLICE_X6Y145_D4;
  wire [0:0] CLBLM_R_X5Y145_SLICE_X6Y145_D5;
  wire [0:0] CLBLM_R_X5Y145_SLICE_X6Y145_D5Q;
  wire [0:0] CLBLM_R_X5Y145_SLICE_X6Y145_D6;
  wire [0:0] CLBLM_R_X5Y145_SLICE_X6Y145_DMUX;
  wire [0:0] CLBLM_R_X5Y145_SLICE_X6Y145_DO5;
  wire [0:0] CLBLM_R_X5Y145_SLICE_X6Y145_DO6;
  wire [0:0] CLBLM_R_X5Y145_SLICE_X6Y145_DQ;
  wire [0:0] CLBLM_R_X5Y145_SLICE_X6Y145_D_CY;
  wire [0:0] CLBLM_R_X5Y145_SLICE_X6Y145_D_XOR;
  wire [0:0] CLBLM_R_X5Y145_SLICE_X7Y145_A;
  wire [0:0] CLBLM_R_X5Y145_SLICE_X7Y145_A1;
  wire [0:0] CLBLM_R_X5Y145_SLICE_X7Y145_A2;
  wire [0:0] CLBLM_R_X5Y145_SLICE_X7Y145_A3;
  wire [0:0] CLBLM_R_X5Y145_SLICE_X7Y145_A4;
  wire [0:0] CLBLM_R_X5Y145_SLICE_X7Y145_A5;
  wire [0:0] CLBLM_R_X5Y145_SLICE_X7Y145_A5Q;
  wire [0:0] CLBLM_R_X5Y145_SLICE_X7Y145_A6;
  wire [0:0] CLBLM_R_X5Y145_SLICE_X7Y145_AMUX;
  wire [0:0] CLBLM_R_X5Y145_SLICE_X7Y145_AO5;
  wire [0:0] CLBLM_R_X5Y145_SLICE_X7Y145_AO6;
  wire [0:0] CLBLM_R_X5Y145_SLICE_X7Y145_AQ;
  wire [0:0] CLBLM_R_X5Y145_SLICE_X7Y145_A_CY;
  wire [0:0] CLBLM_R_X5Y145_SLICE_X7Y145_A_XOR;
  wire [0:0] CLBLM_R_X5Y145_SLICE_X7Y145_B;
  wire [0:0] CLBLM_R_X5Y145_SLICE_X7Y145_B1;
  wire [0:0] CLBLM_R_X5Y145_SLICE_X7Y145_B2;
  wire [0:0] CLBLM_R_X5Y145_SLICE_X7Y145_B3;
  wire [0:0] CLBLM_R_X5Y145_SLICE_X7Y145_B4;
  wire [0:0] CLBLM_R_X5Y145_SLICE_X7Y145_B5;
  wire [0:0] CLBLM_R_X5Y145_SLICE_X7Y145_B5Q;
  wire [0:0] CLBLM_R_X5Y145_SLICE_X7Y145_B6;
  wire [0:0] CLBLM_R_X5Y145_SLICE_X7Y145_BMUX;
  wire [0:0] CLBLM_R_X5Y145_SLICE_X7Y145_BO5;
  wire [0:0] CLBLM_R_X5Y145_SLICE_X7Y145_BO6;
  wire [0:0] CLBLM_R_X5Y145_SLICE_X7Y145_BQ;
  wire [0:0] CLBLM_R_X5Y145_SLICE_X7Y145_B_CY;
  wire [0:0] CLBLM_R_X5Y145_SLICE_X7Y145_B_XOR;
  wire [0:0] CLBLM_R_X5Y145_SLICE_X7Y145_C;
  wire [0:0] CLBLM_R_X5Y145_SLICE_X7Y145_C1;
  wire [0:0] CLBLM_R_X5Y145_SLICE_X7Y145_C2;
  wire [0:0] CLBLM_R_X5Y145_SLICE_X7Y145_C3;
  wire [0:0] CLBLM_R_X5Y145_SLICE_X7Y145_C4;
  wire [0:0] CLBLM_R_X5Y145_SLICE_X7Y145_C5;
  wire [0:0] CLBLM_R_X5Y145_SLICE_X7Y145_C6;
  wire [0:0] CLBLM_R_X5Y145_SLICE_X7Y145_CLK;
  wire [0:0] CLBLM_R_X5Y145_SLICE_X7Y145_CO5;
  wire [0:0] CLBLM_R_X5Y145_SLICE_X7Y145_CO6;
  wire [0:0] CLBLM_R_X5Y145_SLICE_X7Y145_C_CY;
  wire [0:0] CLBLM_R_X5Y145_SLICE_X7Y145_C_XOR;
  wire [0:0] CLBLM_R_X5Y145_SLICE_X7Y145_D;
  wire [0:0] CLBLM_R_X5Y145_SLICE_X7Y145_D1;
  wire [0:0] CLBLM_R_X5Y145_SLICE_X7Y145_D2;
  wire [0:0] CLBLM_R_X5Y145_SLICE_X7Y145_D3;
  wire [0:0] CLBLM_R_X5Y145_SLICE_X7Y145_D4;
  wire [0:0] CLBLM_R_X5Y145_SLICE_X7Y145_D5;
  wire [0:0] CLBLM_R_X5Y145_SLICE_X7Y145_D6;
  wire [0:0] CLBLM_R_X5Y145_SLICE_X7Y145_DO5;
  wire [0:0] CLBLM_R_X5Y145_SLICE_X7Y145_DO6;
  wire [0:0] CLBLM_R_X5Y145_SLICE_X7Y145_D_CY;
  wire [0:0] CLBLM_R_X5Y145_SLICE_X7Y145_D_XOR;
  wire [0:0] CLBLM_R_X5Y146_SLICE_X6Y146_A;
  wire [0:0] CLBLM_R_X5Y146_SLICE_X6Y146_A1;
  wire [0:0] CLBLM_R_X5Y146_SLICE_X6Y146_A2;
  wire [0:0] CLBLM_R_X5Y146_SLICE_X6Y146_A3;
  wire [0:0] CLBLM_R_X5Y146_SLICE_X6Y146_A4;
  wire [0:0] CLBLM_R_X5Y146_SLICE_X6Y146_A5;
  wire [0:0] CLBLM_R_X5Y146_SLICE_X6Y146_A6;
  wire [0:0] CLBLM_R_X5Y146_SLICE_X6Y146_AO5;
  wire [0:0] CLBLM_R_X5Y146_SLICE_X6Y146_AO6;
  wire [0:0] CLBLM_R_X5Y146_SLICE_X6Y146_AQ;
  wire [0:0] CLBLM_R_X5Y146_SLICE_X6Y146_A_CY;
  wire [0:0] CLBLM_R_X5Y146_SLICE_X6Y146_A_XOR;
  wire [0:0] CLBLM_R_X5Y146_SLICE_X6Y146_B;
  wire [0:0] CLBLM_R_X5Y146_SLICE_X6Y146_B1;
  wire [0:0] CLBLM_R_X5Y146_SLICE_X6Y146_B2;
  wire [0:0] CLBLM_R_X5Y146_SLICE_X6Y146_B3;
  wire [0:0] CLBLM_R_X5Y146_SLICE_X6Y146_B4;
  wire [0:0] CLBLM_R_X5Y146_SLICE_X6Y146_B5;
  wire [0:0] CLBLM_R_X5Y146_SLICE_X6Y146_B5Q;
  wire [0:0] CLBLM_R_X5Y146_SLICE_X6Y146_B6;
  wire [0:0] CLBLM_R_X5Y146_SLICE_X6Y146_BMUX;
  wire [0:0] CLBLM_R_X5Y146_SLICE_X6Y146_BO5;
  wire [0:0] CLBLM_R_X5Y146_SLICE_X6Y146_BO6;
  wire [0:0] CLBLM_R_X5Y146_SLICE_X6Y146_BQ;
  wire [0:0] CLBLM_R_X5Y146_SLICE_X6Y146_B_CY;
  wire [0:0] CLBLM_R_X5Y146_SLICE_X6Y146_B_XOR;
  wire [0:0] CLBLM_R_X5Y146_SLICE_X6Y146_C;
  wire [0:0] CLBLM_R_X5Y146_SLICE_X6Y146_C1;
  wire [0:0] CLBLM_R_X5Y146_SLICE_X6Y146_C2;
  wire [0:0] CLBLM_R_X5Y146_SLICE_X6Y146_C3;
  wire [0:0] CLBLM_R_X5Y146_SLICE_X6Y146_C4;
  wire [0:0] CLBLM_R_X5Y146_SLICE_X6Y146_C5;
  wire [0:0] CLBLM_R_X5Y146_SLICE_X6Y146_C6;
  wire [0:0] CLBLM_R_X5Y146_SLICE_X6Y146_CLK;
  wire [0:0] CLBLM_R_X5Y146_SLICE_X6Y146_CO5;
  wire [0:0] CLBLM_R_X5Y146_SLICE_X6Y146_CO6;
  wire [0:0] CLBLM_R_X5Y146_SLICE_X6Y146_C_CY;
  wire [0:0] CLBLM_R_X5Y146_SLICE_X6Y146_C_XOR;
  wire [0:0] CLBLM_R_X5Y146_SLICE_X6Y146_D;
  wire [0:0] CLBLM_R_X5Y146_SLICE_X6Y146_D1;
  wire [0:0] CLBLM_R_X5Y146_SLICE_X6Y146_D2;
  wire [0:0] CLBLM_R_X5Y146_SLICE_X6Y146_D3;
  wire [0:0] CLBLM_R_X5Y146_SLICE_X6Y146_D4;
  wire [0:0] CLBLM_R_X5Y146_SLICE_X6Y146_D5;
  wire [0:0] CLBLM_R_X5Y146_SLICE_X6Y146_D6;
  wire [0:0] CLBLM_R_X5Y146_SLICE_X6Y146_DO5;
  wire [0:0] CLBLM_R_X5Y146_SLICE_X6Y146_DO6;
  wire [0:0] CLBLM_R_X5Y146_SLICE_X6Y146_D_CY;
  wire [0:0] CLBLM_R_X5Y146_SLICE_X6Y146_D_XOR;
  wire [0:0] CLBLM_R_X5Y146_SLICE_X7Y146_A;
  wire [0:0] CLBLM_R_X5Y146_SLICE_X7Y146_A1;
  wire [0:0] CLBLM_R_X5Y146_SLICE_X7Y146_A2;
  wire [0:0] CLBLM_R_X5Y146_SLICE_X7Y146_A3;
  wire [0:0] CLBLM_R_X5Y146_SLICE_X7Y146_A4;
  wire [0:0] CLBLM_R_X5Y146_SLICE_X7Y146_A5;
  wire [0:0] CLBLM_R_X5Y146_SLICE_X7Y146_A6;
  wire [0:0] CLBLM_R_X5Y146_SLICE_X7Y146_AO5;
  wire [0:0] CLBLM_R_X5Y146_SLICE_X7Y146_AO6;
  wire [0:0] CLBLM_R_X5Y146_SLICE_X7Y146_AQ;
  wire [0:0] CLBLM_R_X5Y146_SLICE_X7Y146_A_CY;
  wire [0:0] CLBLM_R_X5Y146_SLICE_X7Y146_A_XOR;
  wire [0:0] CLBLM_R_X5Y146_SLICE_X7Y146_B;
  wire [0:0] CLBLM_R_X5Y146_SLICE_X7Y146_B1;
  wire [0:0] CLBLM_R_X5Y146_SLICE_X7Y146_B2;
  wire [0:0] CLBLM_R_X5Y146_SLICE_X7Y146_B3;
  wire [0:0] CLBLM_R_X5Y146_SLICE_X7Y146_B4;
  wire [0:0] CLBLM_R_X5Y146_SLICE_X7Y146_B5;
  wire [0:0] CLBLM_R_X5Y146_SLICE_X7Y146_B6;
  wire [0:0] CLBLM_R_X5Y146_SLICE_X7Y146_BO5;
  wire [0:0] CLBLM_R_X5Y146_SLICE_X7Y146_BO6;
  wire [0:0] CLBLM_R_X5Y146_SLICE_X7Y146_BQ;
  wire [0:0] CLBLM_R_X5Y146_SLICE_X7Y146_B_CY;
  wire [0:0] CLBLM_R_X5Y146_SLICE_X7Y146_B_XOR;
  wire [0:0] CLBLM_R_X5Y146_SLICE_X7Y146_C;
  wire [0:0] CLBLM_R_X5Y146_SLICE_X7Y146_C1;
  wire [0:0] CLBLM_R_X5Y146_SLICE_X7Y146_C2;
  wire [0:0] CLBLM_R_X5Y146_SLICE_X7Y146_C3;
  wire [0:0] CLBLM_R_X5Y146_SLICE_X7Y146_C4;
  wire [0:0] CLBLM_R_X5Y146_SLICE_X7Y146_C5;
  wire [0:0] CLBLM_R_X5Y146_SLICE_X7Y146_C5Q;
  wire [0:0] CLBLM_R_X5Y146_SLICE_X7Y146_C6;
  wire [0:0] CLBLM_R_X5Y146_SLICE_X7Y146_CLK;
  wire [0:0] CLBLM_R_X5Y146_SLICE_X7Y146_CMUX;
  wire [0:0] CLBLM_R_X5Y146_SLICE_X7Y146_CO5;
  wire [0:0] CLBLM_R_X5Y146_SLICE_X7Y146_CO6;
  wire [0:0] CLBLM_R_X5Y146_SLICE_X7Y146_CQ;
  wire [0:0] CLBLM_R_X5Y146_SLICE_X7Y146_C_CY;
  wire [0:0] CLBLM_R_X5Y146_SLICE_X7Y146_C_XOR;
  wire [0:0] CLBLM_R_X5Y146_SLICE_X7Y146_D;
  wire [0:0] CLBLM_R_X5Y146_SLICE_X7Y146_D1;
  wire [0:0] CLBLM_R_X5Y146_SLICE_X7Y146_D2;
  wire [0:0] CLBLM_R_X5Y146_SLICE_X7Y146_D3;
  wire [0:0] CLBLM_R_X5Y146_SLICE_X7Y146_D4;
  wire [0:0] CLBLM_R_X5Y146_SLICE_X7Y146_D5;
  wire [0:0] CLBLM_R_X5Y146_SLICE_X7Y146_D5Q;
  wire [0:0] CLBLM_R_X5Y146_SLICE_X7Y146_D6;
  wire [0:0] CLBLM_R_X5Y146_SLICE_X7Y146_DMUX;
  wire [0:0] CLBLM_R_X5Y146_SLICE_X7Y146_DO5;
  wire [0:0] CLBLM_R_X5Y146_SLICE_X7Y146_DO6;
  wire [0:0] CLBLM_R_X5Y146_SLICE_X7Y146_DQ;
  wire [0:0] CLBLM_R_X5Y146_SLICE_X7Y146_D_CY;
  wire [0:0] CLBLM_R_X5Y146_SLICE_X7Y146_D_XOR;
  wire [0:0] CLBLM_R_X5Y147_SLICE_X6Y147_A;
  wire [0:0] CLBLM_R_X5Y147_SLICE_X6Y147_A1;
  wire [0:0] CLBLM_R_X5Y147_SLICE_X6Y147_A2;
  wire [0:0] CLBLM_R_X5Y147_SLICE_X6Y147_A3;
  wire [0:0] CLBLM_R_X5Y147_SLICE_X6Y147_A4;
  wire [0:0] CLBLM_R_X5Y147_SLICE_X6Y147_A5;
  wire [0:0] CLBLM_R_X5Y147_SLICE_X6Y147_A6;
  wire [0:0] CLBLM_R_X5Y147_SLICE_X6Y147_AO5;
  wire [0:0] CLBLM_R_X5Y147_SLICE_X6Y147_AO6;
  wire [0:0] CLBLM_R_X5Y147_SLICE_X6Y147_AQ;
  wire [0:0] CLBLM_R_X5Y147_SLICE_X6Y147_A_CY;
  wire [0:0] CLBLM_R_X5Y147_SLICE_X6Y147_A_XOR;
  wire [0:0] CLBLM_R_X5Y147_SLICE_X6Y147_B;
  wire [0:0] CLBLM_R_X5Y147_SLICE_X6Y147_B1;
  wire [0:0] CLBLM_R_X5Y147_SLICE_X6Y147_B2;
  wire [0:0] CLBLM_R_X5Y147_SLICE_X6Y147_B3;
  wire [0:0] CLBLM_R_X5Y147_SLICE_X6Y147_B4;
  wire [0:0] CLBLM_R_X5Y147_SLICE_X6Y147_B5;
  wire [0:0] CLBLM_R_X5Y147_SLICE_X6Y147_B5Q;
  wire [0:0] CLBLM_R_X5Y147_SLICE_X6Y147_B6;
  wire [0:0] CLBLM_R_X5Y147_SLICE_X6Y147_BMUX;
  wire [0:0] CLBLM_R_X5Y147_SLICE_X6Y147_BO5;
  wire [0:0] CLBLM_R_X5Y147_SLICE_X6Y147_BO6;
  wire [0:0] CLBLM_R_X5Y147_SLICE_X6Y147_BQ;
  wire [0:0] CLBLM_R_X5Y147_SLICE_X6Y147_B_CY;
  wire [0:0] CLBLM_R_X5Y147_SLICE_X6Y147_B_XOR;
  wire [0:0] CLBLM_R_X5Y147_SLICE_X6Y147_C;
  wire [0:0] CLBLM_R_X5Y147_SLICE_X6Y147_C1;
  wire [0:0] CLBLM_R_X5Y147_SLICE_X6Y147_C2;
  wire [0:0] CLBLM_R_X5Y147_SLICE_X6Y147_C3;
  wire [0:0] CLBLM_R_X5Y147_SLICE_X6Y147_C4;
  wire [0:0] CLBLM_R_X5Y147_SLICE_X6Y147_C5;
  wire [0:0] CLBLM_R_X5Y147_SLICE_X6Y147_C5Q;
  wire [0:0] CLBLM_R_X5Y147_SLICE_X6Y147_C6;
  wire [0:0] CLBLM_R_X5Y147_SLICE_X6Y147_CLK;
  wire [0:0] CLBLM_R_X5Y147_SLICE_X6Y147_CMUX;
  wire [0:0] CLBLM_R_X5Y147_SLICE_X6Y147_CO5;
  wire [0:0] CLBLM_R_X5Y147_SLICE_X6Y147_CO6;
  wire [0:0] CLBLM_R_X5Y147_SLICE_X6Y147_CQ;
  wire [0:0] CLBLM_R_X5Y147_SLICE_X6Y147_C_CY;
  wire [0:0] CLBLM_R_X5Y147_SLICE_X6Y147_C_XOR;
  wire [0:0] CLBLM_R_X5Y147_SLICE_X6Y147_D;
  wire [0:0] CLBLM_R_X5Y147_SLICE_X6Y147_D1;
  wire [0:0] CLBLM_R_X5Y147_SLICE_X6Y147_D2;
  wire [0:0] CLBLM_R_X5Y147_SLICE_X6Y147_D3;
  wire [0:0] CLBLM_R_X5Y147_SLICE_X6Y147_D4;
  wire [0:0] CLBLM_R_X5Y147_SLICE_X6Y147_D5;
  wire [0:0] CLBLM_R_X5Y147_SLICE_X6Y147_D6;
  wire [0:0] CLBLM_R_X5Y147_SLICE_X6Y147_DO5;
  wire [0:0] CLBLM_R_X5Y147_SLICE_X6Y147_DO6;
  wire [0:0] CLBLM_R_X5Y147_SLICE_X6Y147_D_CY;
  wire [0:0] CLBLM_R_X5Y147_SLICE_X6Y147_D_XOR;
  wire [0:0] CLBLM_R_X5Y147_SLICE_X7Y147_A;
  wire [0:0] CLBLM_R_X5Y147_SLICE_X7Y147_A1;
  wire [0:0] CLBLM_R_X5Y147_SLICE_X7Y147_A2;
  wire [0:0] CLBLM_R_X5Y147_SLICE_X7Y147_A3;
  wire [0:0] CLBLM_R_X5Y147_SLICE_X7Y147_A4;
  wire [0:0] CLBLM_R_X5Y147_SLICE_X7Y147_A5;
  wire [0:0] CLBLM_R_X5Y147_SLICE_X7Y147_A6;
  wire [0:0] CLBLM_R_X5Y147_SLICE_X7Y147_AO5;
  wire [0:0] CLBLM_R_X5Y147_SLICE_X7Y147_AO6;
  wire [0:0] CLBLM_R_X5Y147_SLICE_X7Y147_AQ;
  wire [0:0] CLBLM_R_X5Y147_SLICE_X7Y147_A_CY;
  wire [0:0] CLBLM_R_X5Y147_SLICE_X7Y147_A_XOR;
  wire [0:0] CLBLM_R_X5Y147_SLICE_X7Y147_B;
  wire [0:0] CLBLM_R_X5Y147_SLICE_X7Y147_B1;
  wire [0:0] CLBLM_R_X5Y147_SLICE_X7Y147_B2;
  wire [0:0] CLBLM_R_X5Y147_SLICE_X7Y147_B3;
  wire [0:0] CLBLM_R_X5Y147_SLICE_X7Y147_B4;
  wire [0:0] CLBLM_R_X5Y147_SLICE_X7Y147_B5;
  wire [0:0] CLBLM_R_X5Y147_SLICE_X7Y147_B5Q;
  wire [0:0] CLBLM_R_X5Y147_SLICE_X7Y147_B6;
  wire [0:0] CLBLM_R_X5Y147_SLICE_X7Y147_BMUX;
  wire [0:0] CLBLM_R_X5Y147_SLICE_X7Y147_BO5;
  wire [0:0] CLBLM_R_X5Y147_SLICE_X7Y147_BO6;
  wire [0:0] CLBLM_R_X5Y147_SLICE_X7Y147_BQ;
  wire [0:0] CLBLM_R_X5Y147_SLICE_X7Y147_B_CY;
  wire [0:0] CLBLM_R_X5Y147_SLICE_X7Y147_B_XOR;
  wire [0:0] CLBLM_R_X5Y147_SLICE_X7Y147_C;
  wire [0:0] CLBLM_R_X5Y147_SLICE_X7Y147_C1;
  wire [0:0] CLBLM_R_X5Y147_SLICE_X7Y147_C2;
  wire [0:0] CLBLM_R_X5Y147_SLICE_X7Y147_C3;
  wire [0:0] CLBLM_R_X5Y147_SLICE_X7Y147_C4;
  wire [0:0] CLBLM_R_X5Y147_SLICE_X7Y147_C5;
  wire [0:0] CLBLM_R_X5Y147_SLICE_X7Y147_C5Q;
  wire [0:0] CLBLM_R_X5Y147_SLICE_X7Y147_C6;
  wire [0:0] CLBLM_R_X5Y147_SLICE_X7Y147_CLK;
  wire [0:0] CLBLM_R_X5Y147_SLICE_X7Y147_CMUX;
  wire [0:0] CLBLM_R_X5Y147_SLICE_X7Y147_CO5;
  wire [0:0] CLBLM_R_X5Y147_SLICE_X7Y147_CO6;
  wire [0:0] CLBLM_R_X5Y147_SLICE_X7Y147_CQ;
  wire [0:0] CLBLM_R_X5Y147_SLICE_X7Y147_C_CY;
  wire [0:0] CLBLM_R_X5Y147_SLICE_X7Y147_C_XOR;
  wire [0:0] CLBLM_R_X5Y147_SLICE_X7Y147_D;
  wire [0:0] CLBLM_R_X5Y147_SLICE_X7Y147_D1;
  wire [0:0] CLBLM_R_X5Y147_SLICE_X7Y147_D2;
  wire [0:0] CLBLM_R_X5Y147_SLICE_X7Y147_D3;
  wire [0:0] CLBLM_R_X5Y147_SLICE_X7Y147_D4;
  wire [0:0] CLBLM_R_X5Y147_SLICE_X7Y147_D5;
  wire [0:0] CLBLM_R_X5Y147_SLICE_X7Y147_D6;
  wire [0:0] CLBLM_R_X5Y147_SLICE_X7Y147_DO5;
  wire [0:0] CLBLM_R_X5Y147_SLICE_X7Y147_DO6;
  wire [0:0] CLBLM_R_X5Y147_SLICE_X7Y147_D_CY;
  wire [0:0] CLBLM_R_X5Y147_SLICE_X7Y147_D_XOR;
  wire [0:0] CLBLM_R_X5Y148_SLICE_X6Y148_A;
  wire [0:0] CLBLM_R_X5Y148_SLICE_X6Y148_A1;
  wire [0:0] CLBLM_R_X5Y148_SLICE_X6Y148_A2;
  wire [0:0] CLBLM_R_X5Y148_SLICE_X6Y148_A3;
  wire [0:0] CLBLM_R_X5Y148_SLICE_X6Y148_A4;
  wire [0:0] CLBLM_R_X5Y148_SLICE_X6Y148_A5;
  wire [0:0] CLBLM_R_X5Y148_SLICE_X6Y148_A6;
  wire [0:0] CLBLM_R_X5Y148_SLICE_X6Y148_AMUX;
  wire [0:0] CLBLM_R_X5Y148_SLICE_X6Y148_AO5;
  wire [0:0] CLBLM_R_X5Y148_SLICE_X6Y148_AO6;
  wire [0:0] CLBLM_R_X5Y148_SLICE_X6Y148_AQ;
  wire [0:0] CLBLM_R_X5Y148_SLICE_X6Y148_AX;
  wire [0:0] CLBLM_R_X5Y148_SLICE_X6Y148_A_CY;
  wire [0:0] CLBLM_R_X5Y148_SLICE_X6Y148_A_XOR;
  wire [0:0] CLBLM_R_X5Y148_SLICE_X6Y148_B;
  wire [0:0] CLBLM_R_X5Y148_SLICE_X6Y148_B1;
  wire [0:0] CLBLM_R_X5Y148_SLICE_X6Y148_B2;
  wire [0:0] CLBLM_R_X5Y148_SLICE_X6Y148_B3;
  wire [0:0] CLBLM_R_X5Y148_SLICE_X6Y148_B4;
  wire [0:0] CLBLM_R_X5Y148_SLICE_X6Y148_B5;
  wire [0:0] CLBLM_R_X5Y148_SLICE_X6Y148_B6;
  wire [0:0] CLBLM_R_X5Y148_SLICE_X6Y148_BO5;
  wire [0:0] CLBLM_R_X5Y148_SLICE_X6Y148_BO6;
  wire [0:0] CLBLM_R_X5Y148_SLICE_X6Y148_BQ;
  wire [0:0] CLBLM_R_X5Y148_SLICE_X6Y148_BX;
  wire [0:0] CLBLM_R_X5Y148_SLICE_X6Y148_B_CY;
  wire [0:0] CLBLM_R_X5Y148_SLICE_X6Y148_B_XOR;
  wire [0:0] CLBLM_R_X5Y148_SLICE_X6Y148_C;
  wire [0:0] CLBLM_R_X5Y148_SLICE_X6Y148_C1;
  wire [0:0] CLBLM_R_X5Y148_SLICE_X6Y148_C2;
  wire [0:0] CLBLM_R_X5Y148_SLICE_X6Y148_C3;
  wire [0:0] CLBLM_R_X5Y148_SLICE_X6Y148_C4;
  wire [0:0] CLBLM_R_X5Y148_SLICE_X6Y148_C5;
  wire [0:0] CLBLM_R_X5Y148_SLICE_X6Y148_C6;
  wire [0:0] CLBLM_R_X5Y148_SLICE_X6Y148_CE;
  wire [0:0] CLBLM_R_X5Y148_SLICE_X6Y148_CLK;
  wire [0:0] CLBLM_R_X5Y148_SLICE_X6Y148_CO5;
  wire [0:0] CLBLM_R_X5Y148_SLICE_X6Y148_CO6;
  wire [0:0] CLBLM_R_X5Y148_SLICE_X6Y148_CQ;
  wire [0:0] CLBLM_R_X5Y148_SLICE_X6Y148_CX;
  wire [0:0] CLBLM_R_X5Y148_SLICE_X6Y148_C_CY;
  wire [0:0] CLBLM_R_X5Y148_SLICE_X6Y148_C_XOR;
  wire [0:0] CLBLM_R_X5Y148_SLICE_X6Y148_D;
  wire [0:0] CLBLM_R_X5Y148_SLICE_X6Y148_D1;
  wire [0:0] CLBLM_R_X5Y148_SLICE_X6Y148_D2;
  wire [0:0] CLBLM_R_X5Y148_SLICE_X6Y148_D3;
  wire [0:0] CLBLM_R_X5Y148_SLICE_X6Y148_D4;
  wire [0:0] CLBLM_R_X5Y148_SLICE_X6Y148_D5;
  wire [0:0] CLBLM_R_X5Y148_SLICE_X6Y148_D6;
  wire [0:0] CLBLM_R_X5Y148_SLICE_X6Y148_DO5;
  wire [0:0] CLBLM_R_X5Y148_SLICE_X6Y148_DO6;
  wire [0:0] CLBLM_R_X5Y148_SLICE_X6Y148_D_CY;
  wire [0:0] CLBLM_R_X5Y148_SLICE_X6Y148_D_XOR;
  wire [0:0] CLBLM_R_X5Y148_SLICE_X7Y148_A;
  wire [0:0] CLBLM_R_X5Y148_SLICE_X7Y148_A1;
  wire [0:0] CLBLM_R_X5Y148_SLICE_X7Y148_A2;
  wire [0:0] CLBLM_R_X5Y148_SLICE_X7Y148_A3;
  wire [0:0] CLBLM_R_X5Y148_SLICE_X7Y148_A4;
  wire [0:0] CLBLM_R_X5Y148_SLICE_X7Y148_A5;
  wire [0:0] CLBLM_R_X5Y148_SLICE_X7Y148_A6;
  wire [0:0] CLBLM_R_X5Y148_SLICE_X7Y148_AO5;
  wire [0:0] CLBLM_R_X5Y148_SLICE_X7Y148_AO6;
  wire [0:0] CLBLM_R_X5Y148_SLICE_X7Y148_AQ;
  wire [0:0] CLBLM_R_X5Y148_SLICE_X7Y148_A_CY;
  wire [0:0] CLBLM_R_X5Y148_SLICE_X7Y148_A_XOR;
  wire [0:0] CLBLM_R_X5Y148_SLICE_X7Y148_B;
  wire [0:0] CLBLM_R_X5Y148_SLICE_X7Y148_B1;
  wire [0:0] CLBLM_R_X5Y148_SLICE_X7Y148_B2;
  wire [0:0] CLBLM_R_X5Y148_SLICE_X7Y148_B3;
  wire [0:0] CLBLM_R_X5Y148_SLICE_X7Y148_B4;
  wire [0:0] CLBLM_R_X5Y148_SLICE_X7Y148_B5;
  wire [0:0] CLBLM_R_X5Y148_SLICE_X7Y148_B6;
  wire [0:0] CLBLM_R_X5Y148_SLICE_X7Y148_BO5;
  wire [0:0] CLBLM_R_X5Y148_SLICE_X7Y148_BO6;
  wire [0:0] CLBLM_R_X5Y148_SLICE_X7Y148_BQ;
  wire [0:0] CLBLM_R_X5Y148_SLICE_X7Y148_B_CY;
  wire [0:0] CLBLM_R_X5Y148_SLICE_X7Y148_B_XOR;
  wire [0:0] CLBLM_R_X5Y148_SLICE_X7Y148_C;
  wire [0:0] CLBLM_R_X5Y148_SLICE_X7Y148_C1;
  wire [0:0] CLBLM_R_X5Y148_SLICE_X7Y148_C2;
  wire [0:0] CLBLM_R_X5Y148_SLICE_X7Y148_C3;
  wire [0:0] CLBLM_R_X5Y148_SLICE_X7Y148_C4;
  wire [0:0] CLBLM_R_X5Y148_SLICE_X7Y148_C5;
  wire [0:0] CLBLM_R_X5Y148_SLICE_X7Y148_C5Q;
  wire [0:0] CLBLM_R_X5Y148_SLICE_X7Y148_C6;
  wire [0:0] CLBLM_R_X5Y148_SLICE_X7Y148_CLK;
  wire [0:0] CLBLM_R_X5Y148_SLICE_X7Y148_CMUX;
  wire [0:0] CLBLM_R_X5Y148_SLICE_X7Y148_CO5;
  wire [0:0] CLBLM_R_X5Y148_SLICE_X7Y148_CO6;
  wire [0:0] CLBLM_R_X5Y148_SLICE_X7Y148_CQ;
  wire [0:0] CLBLM_R_X5Y148_SLICE_X7Y148_C_CY;
  wire [0:0] CLBLM_R_X5Y148_SLICE_X7Y148_C_XOR;
  wire [0:0] CLBLM_R_X5Y148_SLICE_X7Y148_D;
  wire [0:0] CLBLM_R_X5Y148_SLICE_X7Y148_D1;
  wire [0:0] CLBLM_R_X5Y148_SLICE_X7Y148_D2;
  wire [0:0] CLBLM_R_X5Y148_SLICE_X7Y148_D3;
  wire [0:0] CLBLM_R_X5Y148_SLICE_X7Y148_D4;
  wire [0:0] CLBLM_R_X5Y148_SLICE_X7Y148_D5;
  wire [0:0] CLBLM_R_X5Y148_SLICE_X7Y148_D6;
  wire [0:0] CLBLM_R_X5Y148_SLICE_X7Y148_DMUX;
  wire [0:0] CLBLM_R_X5Y148_SLICE_X7Y148_DO5;
  wire [0:0] CLBLM_R_X5Y148_SLICE_X7Y148_DO6;
  wire [0:0] CLBLM_R_X5Y148_SLICE_X7Y148_D_CY;
  wire [0:0] CLBLM_R_X5Y148_SLICE_X7Y148_D_XOR;
  wire [0:0] CLBLM_R_X5Y149_SLICE_X6Y149_A;
  wire [0:0] CLBLM_R_X5Y149_SLICE_X6Y149_A1;
  wire [0:0] CLBLM_R_X5Y149_SLICE_X6Y149_A2;
  wire [0:0] CLBLM_R_X5Y149_SLICE_X6Y149_A3;
  wire [0:0] CLBLM_R_X5Y149_SLICE_X6Y149_A4;
  wire [0:0] CLBLM_R_X5Y149_SLICE_X6Y149_A5;
  wire [0:0] CLBLM_R_X5Y149_SLICE_X6Y149_A6;
  wire [0:0] CLBLM_R_X5Y149_SLICE_X6Y149_AO5;
  wire [0:0] CLBLM_R_X5Y149_SLICE_X6Y149_AO6;
  wire [0:0] CLBLM_R_X5Y149_SLICE_X6Y149_AQ;
  wire [0:0] CLBLM_R_X5Y149_SLICE_X6Y149_A_CY;
  wire [0:0] CLBLM_R_X5Y149_SLICE_X6Y149_A_XOR;
  wire [0:0] CLBLM_R_X5Y149_SLICE_X6Y149_B;
  wire [0:0] CLBLM_R_X5Y149_SLICE_X6Y149_B1;
  wire [0:0] CLBLM_R_X5Y149_SLICE_X6Y149_B2;
  wire [0:0] CLBLM_R_X5Y149_SLICE_X6Y149_B3;
  wire [0:0] CLBLM_R_X5Y149_SLICE_X6Y149_B4;
  wire [0:0] CLBLM_R_X5Y149_SLICE_X6Y149_B5;
  wire [0:0] CLBLM_R_X5Y149_SLICE_X6Y149_B5Q;
  wire [0:0] CLBLM_R_X5Y149_SLICE_X6Y149_B6;
  wire [0:0] CLBLM_R_X5Y149_SLICE_X6Y149_BMUX;
  wire [0:0] CLBLM_R_X5Y149_SLICE_X6Y149_BO5;
  wire [0:0] CLBLM_R_X5Y149_SLICE_X6Y149_BO6;
  wire [0:0] CLBLM_R_X5Y149_SLICE_X6Y149_BQ;
  wire [0:0] CLBLM_R_X5Y149_SLICE_X6Y149_B_CY;
  wire [0:0] CLBLM_R_X5Y149_SLICE_X6Y149_B_XOR;
  wire [0:0] CLBLM_R_X5Y149_SLICE_X6Y149_C;
  wire [0:0] CLBLM_R_X5Y149_SLICE_X6Y149_C1;
  wire [0:0] CLBLM_R_X5Y149_SLICE_X6Y149_C2;
  wire [0:0] CLBLM_R_X5Y149_SLICE_X6Y149_C3;
  wire [0:0] CLBLM_R_X5Y149_SLICE_X6Y149_C4;
  wire [0:0] CLBLM_R_X5Y149_SLICE_X6Y149_C5;
  wire [0:0] CLBLM_R_X5Y149_SLICE_X6Y149_C5Q;
  wire [0:0] CLBLM_R_X5Y149_SLICE_X6Y149_C6;
  wire [0:0] CLBLM_R_X5Y149_SLICE_X6Y149_CLK;
  wire [0:0] CLBLM_R_X5Y149_SLICE_X6Y149_CMUX;
  wire [0:0] CLBLM_R_X5Y149_SLICE_X6Y149_CO5;
  wire [0:0] CLBLM_R_X5Y149_SLICE_X6Y149_CO6;
  wire [0:0] CLBLM_R_X5Y149_SLICE_X6Y149_CQ;
  wire [0:0] CLBLM_R_X5Y149_SLICE_X6Y149_C_CY;
  wire [0:0] CLBLM_R_X5Y149_SLICE_X6Y149_C_XOR;
  wire [0:0] CLBLM_R_X5Y149_SLICE_X6Y149_D;
  wire [0:0] CLBLM_R_X5Y149_SLICE_X6Y149_D1;
  wire [0:0] CLBLM_R_X5Y149_SLICE_X6Y149_D2;
  wire [0:0] CLBLM_R_X5Y149_SLICE_X6Y149_D3;
  wire [0:0] CLBLM_R_X5Y149_SLICE_X6Y149_D4;
  wire [0:0] CLBLM_R_X5Y149_SLICE_X6Y149_D5;
  wire [0:0] CLBLM_R_X5Y149_SLICE_X6Y149_D6;
  wire [0:0] CLBLM_R_X5Y149_SLICE_X6Y149_DO5;
  wire [0:0] CLBLM_R_X5Y149_SLICE_X6Y149_DO6;
  wire [0:0] CLBLM_R_X5Y149_SLICE_X6Y149_D_CY;
  wire [0:0] CLBLM_R_X5Y149_SLICE_X6Y149_D_XOR;
  wire [0:0] CLBLM_R_X5Y149_SLICE_X7Y149_A;
  wire [0:0] CLBLM_R_X5Y149_SLICE_X7Y149_A1;
  wire [0:0] CLBLM_R_X5Y149_SLICE_X7Y149_A2;
  wire [0:0] CLBLM_R_X5Y149_SLICE_X7Y149_A3;
  wire [0:0] CLBLM_R_X5Y149_SLICE_X7Y149_A4;
  wire [0:0] CLBLM_R_X5Y149_SLICE_X7Y149_A5;
  wire [0:0] CLBLM_R_X5Y149_SLICE_X7Y149_A6;
  wire [0:0] CLBLM_R_X5Y149_SLICE_X7Y149_AO5;
  wire [0:0] CLBLM_R_X5Y149_SLICE_X7Y149_AO6;
  wire [0:0] CLBLM_R_X5Y149_SLICE_X7Y149_AQ;
  wire [0:0] CLBLM_R_X5Y149_SLICE_X7Y149_A_CY;
  wire [0:0] CLBLM_R_X5Y149_SLICE_X7Y149_A_XOR;
  wire [0:0] CLBLM_R_X5Y149_SLICE_X7Y149_B;
  wire [0:0] CLBLM_R_X5Y149_SLICE_X7Y149_B1;
  wire [0:0] CLBLM_R_X5Y149_SLICE_X7Y149_B2;
  wire [0:0] CLBLM_R_X5Y149_SLICE_X7Y149_B3;
  wire [0:0] CLBLM_R_X5Y149_SLICE_X7Y149_B4;
  wire [0:0] CLBLM_R_X5Y149_SLICE_X7Y149_B5;
  wire [0:0] CLBLM_R_X5Y149_SLICE_X7Y149_B6;
  wire [0:0] CLBLM_R_X5Y149_SLICE_X7Y149_BO5;
  wire [0:0] CLBLM_R_X5Y149_SLICE_X7Y149_BO6;
  wire [0:0] CLBLM_R_X5Y149_SLICE_X7Y149_BQ;
  wire [0:0] CLBLM_R_X5Y149_SLICE_X7Y149_B_CY;
  wire [0:0] CLBLM_R_X5Y149_SLICE_X7Y149_B_XOR;
  wire [0:0] CLBLM_R_X5Y149_SLICE_X7Y149_C;
  wire [0:0] CLBLM_R_X5Y149_SLICE_X7Y149_C1;
  wire [0:0] CLBLM_R_X5Y149_SLICE_X7Y149_C2;
  wire [0:0] CLBLM_R_X5Y149_SLICE_X7Y149_C3;
  wire [0:0] CLBLM_R_X5Y149_SLICE_X7Y149_C4;
  wire [0:0] CLBLM_R_X5Y149_SLICE_X7Y149_C5;
  wire [0:0] CLBLM_R_X5Y149_SLICE_X7Y149_C5Q;
  wire [0:0] CLBLM_R_X5Y149_SLICE_X7Y149_C6;
  wire [0:0] CLBLM_R_X5Y149_SLICE_X7Y149_CLK;
  wire [0:0] CLBLM_R_X5Y149_SLICE_X7Y149_CMUX;
  wire [0:0] CLBLM_R_X5Y149_SLICE_X7Y149_CO5;
  wire [0:0] CLBLM_R_X5Y149_SLICE_X7Y149_CO6;
  wire [0:0] CLBLM_R_X5Y149_SLICE_X7Y149_CQ;
  wire [0:0] CLBLM_R_X5Y149_SLICE_X7Y149_C_CY;
  wire [0:0] CLBLM_R_X5Y149_SLICE_X7Y149_C_XOR;
  wire [0:0] CLBLM_R_X5Y149_SLICE_X7Y149_D;
  wire [0:0] CLBLM_R_X5Y149_SLICE_X7Y149_D1;
  wire [0:0] CLBLM_R_X5Y149_SLICE_X7Y149_D2;
  wire [0:0] CLBLM_R_X5Y149_SLICE_X7Y149_D3;
  wire [0:0] CLBLM_R_X5Y149_SLICE_X7Y149_D4;
  wire [0:0] CLBLM_R_X5Y149_SLICE_X7Y149_D5;
  wire [0:0] CLBLM_R_X5Y149_SLICE_X7Y149_D5Q;
  wire [0:0] CLBLM_R_X5Y149_SLICE_X7Y149_D6;
  wire [0:0] CLBLM_R_X5Y149_SLICE_X7Y149_DMUX;
  wire [0:0] CLBLM_R_X5Y149_SLICE_X7Y149_DO5;
  wire [0:0] CLBLM_R_X5Y149_SLICE_X7Y149_DO6;
  wire [0:0] CLBLM_R_X5Y149_SLICE_X7Y149_DQ;
  wire [0:0] CLBLM_R_X5Y149_SLICE_X7Y149_D_CY;
  wire [0:0] CLBLM_R_X5Y149_SLICE_X7Y149_D_XOR;
  wire [0:0] CLBLM_R_X5Y150_SLICE_X6Y150_A;
  wire [0:0] CLBLM_R_X5Y150_SLICE_X6Y150_A1;
  wire [0:0] CLBLM_R_X5Y150_SLICE_X6Y150_A2;
  wire [0:0] CLBLM_R_X5Y150_SLICE_X6Y150_A3;
  wire [0:0] CLBLM_R_X5Y150_SLICE_X6Y150_A4;
  wire [0:0] CLBLM_R_X5Y150_SLICE_X6Y150_A5;
  wire [0:0] CLBLM_R_X5Y150_SLICE_X6Y150_A5Q;
  wire [0:0] CLBLM_R_X5Y150_SLICE_X6Y150_A6;
  wire [0:0] CLBLM_R_X5Y150_SLICE_X6Y150_AMUX;
  wire [0:0] CLBLM_R_X5Y150_SLICE_X6Y150_AO5;
  wire [0:0] CLBLM_R_X5Y150_SLICE_X6Y150_AO6;
  wire [0:0] CLBLM_R_X5Y150_SLICE_X6Y150_AQ;
  wire [0:0] CLBLM_R_X5Y150_SLICE_X6Y150_A_CY;
  wire [0:0] CLBLM_R_X5Y150_SLICE_X6Y150_A_XOR;
  wire [0:0] CLBLM_R_X5Y150_SLICE_X6Y150_B;
  wire [0:0] CLBLM_R_X5Y150_SLICE_X6Y150_B1;
  wire [0:0] CLBLM_R_X5Y150_SLICE_X6Y150_B2;
  wire [0:0] CLBLM_R_X5Y150_SLICE_X6Y150_B3;
  wire [0:0] CLBLM_R_X5Y150_SLICE_X6Y150_B4;
  wire [0:0] CLBLM_R_X5Y150_SLICE_X6Y150_B5;
  wire [0:0] CLBLM_R_X5Y150_SLICE_X6Y150_B5Q;
  wire [0:0] CLBLM_R_X5Y150_SLICE_X6Y150_B6;
  wire [0:0] CLBLM_R_X5Y150_SLICE_X6Y150_BMUX;
  wire [0:0] CLBLM_R_X5Y150_SLICE_X6Y150_BO5;
  wire [0:0] CLBLM_R_X5Y150_SLICE_X6Y150_BO6;
  wire [0:0] CLBLM_R_X5Y150_SLICE_X6Y150_BQ;
  wire [0:0] CLBLM_R_X5Y150_SLICE_X6Y150_B_CY;
  wire [0:0] CLBLM_R_X5Y150_SLICE_X6Y150_B_XOR;
  wire [0:0] CLBLM_R_X5Y150_SLICE_X6Y150_C;
  wire [0:0] CLBLM_R_X5Y150_SLICE_X6Y150_C1;
  wire [0:0] CLBLM_R_X5Y150_SLICE_X6Y150_C2;
  wire [0:0] CLBLM_R_X5Y150_SLICE_X6Y150_C3;
  wire [0:0] CLBLM_R_X5Y150_SLICE_X6Y150_C4;
  wire [0:0] CLBLM_R_X5Y150_SLICE_X6Y150_C5;
  wire [0:0] CLBLM_R_X5Y150_SLICE_X6Y150_C5Q;
  wire [0:0] CLBLM_R_X5Y150_SLICE_X6Y150_C6;
  wire [0:0] CLBLM_R_X5Y150_SLICE_X6Y150_CLK;
  wire [0:0] CLBLM_R_X5Y150_SLICE_X6Y150_CMUX;
  wire [0:0] CLBLM_R_X5Y150_SLICE_X6Y150_CO5;
  wire [0:0] CLBLM_R_X5Y150_SLICE_X6Y150_CO6;
  wire [0:0] CLBLM_R_X5Y150_SLICE_X6Y150_CQ;
  wire [0:0] CLBLM_R_X5Y150_SLICE_X6Y150_C_CY;
  wire [0:0] CLBLM_R_X5Y150_SLICE_X6Y150_C_XOR;
  wire [0:0] CLBLM_R_X5Y150_SLICE_X6Y150_D;
  wire [0:0] CLBLM_R_X5Y150_SLICE_X6Y150_D1;
  wire [0:0] CLBLM_R_X5Y150_SLICE_X6Y150_D2;
  wire [0:0] CLBLM_R_X5Y150_SLICE_X6Y150_D3;
  wire [0:0] CLBLM_R_X5Y150_SLICE_X6Y150_D4;
  wire [0:0] CLBLM_R_X5Y150_SLICE_X6Y150_D5;
  wire [0:0] CLBLM_R_X5Y150_SLICE_X6Y150_D6;
  wire [0:0] CLBLM_R_X5Y150_SLICE_X6Y150_DO5;
  wire [0:0] CLBLM_R_X5Y150_SLICE_X6Y150_DO6;
  wire [0:0] CLBLM_R_X5Y150_SLICE_X6Y150_D_CY;
  wire [0:0] CLBLM_R_X5Y150_SLICE_X6Y150_D_XOR;
  wire [0:0] CLBLM_R_X5Y150_SLICE_X7Y150_A;
  wire [0:0] CLBLM_R_X5Y150_SLICE_X7Y150_A1;
  wire [0:0] CLBLM_R_X5Y150_SLICE_X7Y150_A2;
  wire [0:0] CLBLM_R_X5Y150_SLICE_X7Y150_A3;
  wire [0:0] CLBLM_R_X5Y150_SLICE_X7Y150_A4;
  wire [0:0] CLBLM_R_X5Y150_SLICE_X7Y150_A5;
  wire [0:0] CLBLM_R_X5Y150_SLICE_X7Y150_A5Q;
  wire [0:0] CLBLM_R_X5Y150_SLICE_X7Y150_A6;
  wire [0:0] CLBLM_R_X5Y150_SLICE_X7Y150_AMUX;
  wire [0:0] CLBLM_R_X5Y150_SLICE_X7Y150_AO5;
  wire [0:0] CLBLM_R_X5Y150_SLICE_X7Y150_AO6;
  wire [0:0] CLBLM_R_X5Y150_SLICE_X7Y150_AQ;
  wire [0:0] CLBLM_R_X5Y150_SLICE_X7Y150_A_CY;
  wire [0:0] CLBLM_R_X5Y150_SLICE_X7Y150_A_XOR;
  wire [0:0] CLBLM_R_X5Y150_SLICE_X7Y150_B;
  wire [0:0] CLBLM_R_X5Y150_SLICE_X7Y150_B1;
  wire [0:0] CLBLM_R_X5Y150_SLICE_X7Y150_B2;
  wire [0:0] CLBLM_R_X5Y150_SLICE_X7Y150_B3;
  wire [0:0] CLBLM_R_X5Y150_SLICE_X7Y150_B4;
  wire [0:0] CLBLM_R_X5Y150_SLICE_X7Y150_B5;
  wire [0:0] CLBLM_R_X5Y150_SLICE_X7Y150_B6;
  wire [0:0] CLBLM_R_X5Y150_SLICE_X7Y150_BO5;
  wire [0:0] CLBLM_R_X5Y150_SLICE_X7Y150_BO6;
  wire [0:0] CLBLM_R_X5Y150_SLICE_X7Y150_B_CY;
  wire [0:0] CLBLM_R_X5Y150_SLICE_X7Y150_B_XOR;
  wire [0:0] CLBLM_R_X5Y150_SLICE_X7Y150_C;
  wire [0:0] CLBLM_R_X5Y150_SLICE_X7Y150_C1;
  wire [0:0] CLBLM_R_X5Y150_SLICE_X7Y150_C2;
  wire [0:0] CLBLM_R_X5Y150_SLICE_X7Y150_C3;
  wire [0:0] CLBLM_R_X5Y150_SLICE_X7Y150_C4;
  wire [0:0] CLBLM_R_X5Y150_SLICE_X7Y150_C5;
  wire [0:0] CLBLM_R_X5Y150_SLICE_X7Y150_C6;
  wire [0:0] CLBLM_R_X5Y150_SLICE_X7Y150_CLK;
  wire [0:0] CLBLM_R_X5Y150_SLICE_X7Y150_CO5;
  wire [0:0] CLBLM_R_X5Y150_SLICE_X7Y150_CO6;
  wire [0:0] CLBLM_R_X5Y150_SLICE_X7Y150_C_CY;
  wire [0:0] CLBLM_R_X5Y150_SLICE_X7Y150_C_XOR;
  wire [0:0] CLBLM_R_X5Y150_SLICE_X7Y150_D;
  wire [0:0] CLBLM_R_X5Y150_SLICE_X7Y150_D1;
  wire [0:0] CLBLM_R_X5Y150_SLICE_X7Y150_D2;
  wire [0:0] CLBLM_R_X5Y150_SLICE_X7Y150_D3;
  wire [0:0] CLBLM_R_X5Y150_SLICE_X7Y150_D4;
  wire [0:0] CLBLM_R_X5Y150_SLICE_X7Y150_D5;
  wire [0:0] CLBLM_R_X5Y150_SLICE_X7Y150_D6;
  wire [0:0] CLBLM_R_X5Y150_SLICE_X7Y150_DMUX;
  wire [0:0] CLBLM_R_X5Y150_SLICE_X7Y150_DO5;
  wire [0:0] CLBLM_R_X5Y150_SLICE_X7Y150_DO6;
  wire [0:0] CLBLM_R_X5Y150_SLICE_X7Y150_D_CY;
  wire [0:0] CLBLM_R_X5Y150_SLICE_X7Y150_D_XOR;
  wire [0:0] CLBLM_R_X5Y151_SLICE_X6Y151_A;
  wire [0:0] CLBLM_R_X5Y151_SLICE_X6Y151_A1;
  wire [0:0] CLBLM_R_X5Y151_SLICE_X6Y151_A2;
  wire [0:0] CLBLM_R_X5Y151_SLICE_X6Y151_A3;
  wire [0:0] CLBLM_R_X5Y151_SLICE_X6Y151_A4;
  wire [0:0] CLBLM_R_X5Y151_SLICE_X6Y151_A5;
  wire [0:0] CLBLM_R_X5Y151_SLICE_X6Y151_A6;
  wire [0:0] CLBLM_R_X5Y151_SLICE_X6Y151_AO5;
  wire [0:0] CLBLM_R_X5Y151_SLICE_X6Y151_AO6;
  wire [0:0] CLBLM_R_X5Y151_SLICE_X6Y151_AQ;
  wire [0:0] CLBLM_R_X5Y151_SLICE_X6Y151_A_CY;
  wire [0:0] CLBLM_R_X5Y151_SLICE_X6Y151_A_XOR;
  wire [0:0] CLBLM_R_X5Y151_SLICE_X6Y151_B;
  wire [0:0] CLBLM_R_X5Y151_SLICE_X6Y151_B1;
  wire [0:0] CLBLM_R_X5Y151_SLICE_X6Y151_B2;
  wire [0:0] CLBLM_R_X5Y151_SLICE_X6Y151_B3;
  wire [0:0] CLBLM_R_X5Y151_SLICE_X6Y151_B4;
  wire [0:0] CLBLM_R_X5Y151_SLICE_X6Y151_B5;
  wire [0:0] CLBLM_R_X5Y151_SLICE_X6Y151_B6;
  wire [0:0] CLBLM_R_X5Y151_SLICE_X6Y151_BO5;
  wire [0:0] CLBLM_R_X5Y151_SLICE_X6Y151_BO6;
  wire [0:0] CLBLM_R_X5Y151_SLICE_X6Y151_BQ;
  wire [0:0] CLBLM_R_X5Y151_SLICE_X6Y151_B_CY;
  wire [0:0] CLBLM_R_X5Y151_SLICE_X6Y151_B_XOR;
  wire [0:0] CLBLM_R_X5Y151_SLICE_X6Y151_C;
  wire [0:0] CLBLM_R_X5Y151_SLICE_X6Y151_C1;
  wire [0:0] CLBLM_R_X5Y151_SLICE_X6Y151_C2;
  wire [0:0] CLBLM_R_X5Y151_SLICE_X6Y151_C3;
  wire [0:0] CLBLM_R_X5Y151_SLICE_X6Y151_C4;
  wire [0:0] CLBLM_R_X5Y151_SLICE_X6Y151_C5;
  wire [0:0] CLBLM_R_X5Y151_SLICE_X6Y151_C5Q;
  wire [0:0] CLBLM_R_X5Y151_SLICE_X6Y151_C6;
  wire [0:0] CLBLM_R_X5Y151_SLICE_X6Y151_CLK;
  wire [0:0] CLBLM_R_X5Y151_SLICE_X6Y151_CMUX;
  wire [0:0] CLBLM_R_X5Y151_SLICE_X6Y151_CO5;
  wire [0:0] CLBLM_R_X5Y151_SLICE_X6Y151_CO6;
  wire [0:0] CLBLM_R_X5Y151_SLICE_X6Y151_CQ;
  wire [0:0] CLBLM_R_X5Y151_SLICE_X6Y151_C_CY;
  wire [0:0] CLBLM_R_X5Y151_SLICE_X6Y151_C_XOR;
  wire [0:0] CLBLM_R_X5Y151_SLICE_X6Y151_D;
  wire [0:0] CLBLM_R_X5Y151_SLICE_X6Y151_D1;
  wire [0:0] CLBLM_R_X5Y151_SLICE_X6Y151_D2;
  wire [0:0] CLBLM_R_X5Y151_SLICE_X6Y151_D3;
  wire [0:0] CLBLM_R_X5Y151_SLICE_X6Y151_D4;
  wire [0:0] CLBLM_R_X5Y151_SLICE_X6Y151_D5;
  wire [0:0] CLBLM_R_X5Y151_SLICE_X6Y151_D6;
  wire [0:0] CLBLM_R_X5Y151_SLICE_X6Y151_DO5;
  wire [0:0] CLBLM_R_X5Y151_SLICE_X6Y151_DO6;
  wire [0:0] CLBLM_R_X5Y151_SLICE_X6Y151_D_CY;
  wire [0:0] CLBLM_R_X5Y151_SLICE_X6Y151_D_XOR;
  wire [0:0] CLBLM_R_X5Y151_SLICE_X7Y151_A;
  wire [0:0] CLBLM_R_X5Y151_SLICE_X7Y151_A1;
  wire [0:0] CLBLM_R_X5Y151_SLICE_X7Y151_A2;
  wire [0:0] CLBLM_R_X5Y151_SLICE_X7Y151_A3;
  wire [0:0] CLBLM_R_X5Y151_SLICE_X7Y151_A4;
  wire [0:0] CLBLM_R_X5Y151_SLICE_X7Y151_A5;
  wire [0:0] CLBLM_R_X5Y151_SLICE_X7Y151_A6;
  wire [0:0] CLBLM_R_X5Y151_SLICE_X7Y151_AO5;
  wire [0:0] CLBLM_R_X5Y151_SLICE_X7Y151_AO6;
  wire [0:0] CLBLM_R_X5Y151_SLICE_X7Y151_AQ;
  wire [0:0] CLBLM_R_X5Y151_SLICE_X7Y151_A_CY;
  wire [0:0] CLBLM_R_X5Y151_SLICE_X7Y151_A_XOR;
  wire [0:0] CLBLM_R_X5Y151_SLICE_X7Y151_B;
  wire [0:0] CLBLM_R_X5Y151_SLICE_X7Y151_B1;
  wire [0:0] CLBLM_R_X5Y151_SLICE_X7Y151_B2;
  wire [0:0] CLBLM_R_X5Y151_SLICE_X7Y151_B3;
  wire [0:0] CLBLM_R_X5Y151_SLICE_X7Y151_B4;
  wire [0:0] CLBLM_R_X5Y151_SLICE_X7Y151_B5;
  wire [0:0] CLBLM_R_X5Y151_SLICE_X7Y151_B5Q;
  wire [0:0] CLBLM_R_X5Y151_SLICE_X7Y151_B6;
  wire [0:0] CLBLM_R_X5Y151_SLICE_X7Y151_BMUX;
  wire [0:0] CLBLM_R_X5Y151_SLICE_X7Y151_BO5;
  wire [0:0] CLBLM_R_X5Y151_SLICE_X7Y151_BO6;
  wire [0:0] CLBLM_R_X5Y151_SLICE_X7Y151_BQ;
  wire [0:0] CLBLM_R_X5Y151_SLICE_X7Y151_B_CY;
  wire [0:0] CLBLM_R_X5Y151_SLICE_X7Y151_B_XOR;
  wire [0:0] CLBLM_R_X5Y151_SLICE_X7Y151_C;
  wire [0:0] CLBLM_R_X5Y151_SLICE_X7Y151_C1;
  wire [0:0] CLBLM_R_X5Y151_SLICE_X7Y151_C2;
  wire [0:0] CLBLM_R_X5Y151_SLICE_X7Y151_C3;
  wire [0:0] CLBLM_R_X5Y151_SLICE_X7Y151_C4;
  wire [0:0] CLBLM_R_X5Y151_SLICE_X7Y151_C5;
  wire [0:0] CLBLM_R_X5Y151_SLICE_X7Y151_C6;
  wire [0:0] CLBLM_R_X5Y151_SLICE_X7Y151_CLK;
  wire [0:0] CLBLM_R_X5Y151_SLICE_X7Y151_CO5;
  wire [0:0] CLBLM_R_X5Y151_SLICE_X7Y151_CO6;
  wire [0:0] CLBLM_R_X5Y151_SLICE_X7Y151_C_CY;
  wire [0:0] CLBLM_R_X5Y151_SLICE_X7Y151_C_XOR;
  wire [0:0] CLBLM_R_X5Y151_SLICE_X7Y151_D;
  wire [0:0] CLBLM_R_X5Y151_SLICE_X7Y151_D1;
  wire [0:0] CLBLM_R_X5Y151_SLICE_X7Y151_D2;
  wire [0:0] CLBLM_R_X5Y151_SLICE_X7Y151_D3;
  wire [0:0] CLBLM_R_X5Y151_SLICE_X7Y151_D4;
  wire [0:0] CLBLM_R_X5Y151_SLICE_X7Y151_D5;
  wire [0:0] CLBLM_R_X5Y151_SLICE_X7Y151_D6;
  wire [0:0] CLBLM_R_X5Y151_SLICE_X7Y151_DMUX;
  wire [0:0] CLBLM_R_X5Y151_SLICE_X7Y151_DO5;
  wire [0:0] CLBLM_R_X5Y151_SLICE_X7Y151_DO6;
  wire [0:0] CLBLM_R_X5Y151_SLICE_X7Y151_D_CY;
  wire [0:0] CLBLM_R_X5Y151_SLICE_X7Y151_D_XOR;
  wire [0:0] CLBLM_R_X5Y152_SLICE_X6Y152_A;
  wire [0:0] CLBLM_R_X5Y152_SLICE_X6Y152_A1;
  wire [0:0] CLBLM_R_X5Y152_SLICE_X6Y152_A2;
  wire [0:0] CLBLM_R_X5Y152_SLICE_X6Y152_A3;
  wire [0:0] CLBLM_R_X5Y152_SLICE_X6Y152_A4;
  wire [0:0] CLBLM_R_X5Y152_SLICE_X6Y152_A5;
  wire [0:0] CLBLM_R_X5Y152_SLICE_X6Y152_A6;
  wire [0:0] CLBLM_R_X5Y152_SLICE_X6Y152_AO5;
  wire [0:0] CLBLM_R_X5Y152_SLICE_X6Y152_AO6;
  wire [0:0] CLBLM_R_X5Y152_SLICE_X6Y152_AQ;
  wire [0:0] CLBLM_R_X5Y152_SLICE_X6Y152_A_CY;
  wire [0:0] CLBLM_R_X5Y152_SLICE_X6Y152_A_XOR;
  wire [0:0] CLBLM_R_X5Y152_SLICE_X6Y152_B;
  wire [0:0] CLBLM_R_X5Y152_SLICE_X6Y152_B1;
  wire [0:0] CLBLM_R_X5Y152_SLICE_X6Y152_B2;
  wire [0:0] CLBLM_R_X5Y152_SLICE_X6Y152_B3;
  wire [0:0] CLBLM_R_X5Y152_SLICE_X6Y152_B4;
  wire [0:0] CLBLM_R_X5Y152_SLICE_X6Y152_B5;
  wire [0:0] CLBLM_R_X5Y152_SLICE_X6Y152_B5Q;
  wire [0:0] CLBLM_R_X5Y152_SLICE_X6Y152_B6;
  wire [0:0] CLBLM_R_X5Y152_SLICE_X6Y152_BMUX;
  wire [0:0] CLBLM_R_X5Y152_SLICE_X6Y152_BO5;
  wire [0:0] CLBLM_R_X5Y152_SLICE_X6Y152_BO6;
  wire [0:0] CLBLM_R_X5Y152_SLICE_X6Y152_BQ;
  wire [0:0] CLBLM_R_X5Y152_SLICE_X6Y152_B_CY;
  wire [0:0] CLBLM_R_X5Y152_SLICE_X6Y152_B_XOR;
  wire [0:0] CLBLM_R_X5Y152_SLICE_X6Y152_C;
  wire [0:0] CLBLM_R_X5Y152_SLICE_X6Y152_C1;
  wire [0:0] CLBLM_R_X5Y152_SLICE_X6Y152_C2;
  wire [0:0] CLBLM_R_X5Y152_SLICE_X6Y152_C3;
  wire [0:0] CLBLM_R_X5Y152_SLICE_X6Y152_C4;
  wire [0:0] CLBLM_R_X5Y152_SLICE_X6Y152_C5;
  wire [0:0] CLBLM_R_X5Y152_SLICE_X6Y152_C6;
  wire [0:0] CLBLM_R_X5Y152_SLICE_X6Y152_CLK;
  wire [0:0] CLBLM_R_X5Y152_SLICE_X6Y152_CO5;
  wire [0:0] CLBLM_R_X5Y152_SLICE_X6Y152_CO6;
  wire [0:0] CLBLM_R_X5Y152_SLICE_X6Y152_CQ;
  wire [0:0] CLBLM_R_X5Y152_SLICE_X6Y152_C_CY;
  wire [0:0] CLBLM_R_X5Y152_SLICE_X6Y152_C_XOR;
  wire [0:0] CLBLM_R_X5Y152_SLICE_X6Y152_D;
  wire [0:0] CLBLM_R_X5Y152_SLICE_X6Y152_D1;
  wire [0:0] CLBLM_R_X5Y152_SLICE_X6Y152_D2;
  wire [0:0] CLBLM_R_X5Y152_SLICE_X6Y152_D3;
  wire [0:0] CLBLM_R_X5Y152_SLICE_X6Y152_D4;
  wire [0:0] CLBLM_R_X5Y152_SLICE_X6Y152_D5;
  wire [0:0] CLBLM_R_X5Y152_SLICE_X6Y152_D6;
  wire [0:0] CLBLM_R_X5Y152_SLICE_X6Y152_DO5;
  wire [0:0] CLBLM_R_X5Y152_SLICE_X6Y152_DO6;
  wire [0:0] CLBLM_R_X5Y152_SLICE_X6Y152_DQ;
  wire [0:0] CLBLM_R_X5Y152_SLICE_X6Y152_D_CY;
  wire [0:0] CLBLM_R_X5Y152_SLICE_X6Y152_D_XOR;
  wire [0:0] CLBLM_R_X5Y152_SLICE_X7Y152_A;
  wire [0:0] CLBLM_R_X5Y152_SLICE_X7Y152_A1;
  wire [0:0] CLBLM_R_X5Y152_SLICE_X7Y152_A2;
  wire [0:0] CLBLM_R_X5Y152_SLICE_X7Y152_A3;
  wire [0:0] CLBLM_R_X5Y152_SLICE_X7Y152_A4;
  wire [0:0] CLBLM_R_X5Y152_SLICE_X7Y152_A5;
  wire [0:0] CLBLM_R_X5Y152_SLICE_X7Y152_A5Q;
  wire [0:0] CLBLM_R_X5Y152_SLICE_X7Y152_A6;
  wire [0:0] CLBLM_R_X5Y152_SLICE_X7Y152_AMUX;
  wire [0:0] CLBLM_R_X5Y152_SLICE_X7Y152_AO5;
  wire [0:0] CLBLM_R_X5Y152_SLICE_X7Y152_AO6;
  wire [0:0] CLBLM_R_X5Y152_SLICE_X7Y152_AQ;
  wire [0:0] CLBLM_R_X5Y152_SLICE_X7Y152_A_CY;
  wire [0:0] CLBLM_R_X5Y152_SLICE_X7Y152_A_XOR;
  wire [0:0] CLBLM_R_X5Y152_SLICE_X7Y152_B;
  wire [0:0] CLBLM_R_X5Y152_SLICE_X7Y152_B1;
  wire [0:0] CLBLM_R_X5Y152_SLICE_X7Y152_B2;
  wire [0:0] CLBLM_R_X5Y152_SLICE_X7Y152_B3;
  wire [0:0] CLBLM_R_X5Y152_SLICE_X7Y152_B4;
  wire [0:0] CLBLM_R_X5Y152_SLICE_X7Y152_B5;
  wire [0:0] CLBLM_R_X5Y152_SLICE_X7Y152_B5Q;
  wire [0:0] CLBLM_R_X5Y152_SLICE_X7Y152_B6;
  wire [0:0] CLBLM_R_X5Y152_SLICE_X7Y152_BMUX;
  wire [0:0] CLBLM_R_X5Y152_SLICE_X7Y152_BO5;
  wire [0:0] CLBLM_R_X5Y152_SLICE_X7Y152_BO6;
  wire [0:0] CLBLM_R_X5Y152_SLICE_X7Y152_BQ;
  wire [0:0] CLBLM_R_X5Y152_SLICE_X7Y152_B_CY;
  wire [0:0] CLBLM_R_X5Y152_SLICE_X7Y152_B_XOR;
  wire [0:0] CLBLM_R_X5Y152_SLICE_X7Y152_C;
  wire [0:0] CLBLM_R_X5Y152_SLICE_X7Y152_C1;
  wire [0:0] CLBLM_R_X5Y152_SLICE_X7Y152_C2;
  wire [0:0] CLBLM_R_X5Y152_SLICE_X7Y152_C3;
  wire [0:0] CLBLM_R_X5Y152_SLICE_X7Y152_C4;
  wire [0:0] CLBLM_R_X5Y152_SLICE_X7Y152_C5;
  wire [0:0] CLBLM_R_X5Y152_SLICE_X7Y152_C5Q;
  wire [0:0] CLBLM_R_X5Y152_SLICE_X7Y152_C6;
  wire [0:0] CLBLM_R_X5Y152_SLICE_X7Y152_CLK;
  wire [0:0] CLBLM_R_X5Y152_SLICE_X7Y152_CMUX;
  wire [0:0] CLBLM_R_X5Y152_SLICE_X7Y152_CO5;
  wire [0:0] CLBLM_R_X5Y152_SLICE_X7Y152_CO6;
  wire [0:0] CLBLM_R_X5Y152_SLICE_X7Y152_CQ;
  wire [0:0] CLBLM_R_X5Y152_SLICE_X7Y152_C_CY;
  wire [0:0] CLBLM_R_X5Y152_SLICE_X7Y152_C_XOR;
  wire [0:0] CLBLM_R_X5Y152_SLICE_X7Y152_D;
  wire [0:0] CLBLM_R_X5Y152_SLICE_X7Y152_D1;
  wire [0:0] CLBLM_R_X5Y152_SLICE_X7Y152_D2;
  wire [0:0] CLBLM_R_X5Y152_SLICE_X7Y152_D3;
  wire [0:0] CLBLM_R_X5Y152_SLICE_X7Y152_D4;
  wire [0:0] CLBLM_R_X5Y152_SLICE_X7Y152_D5;
  wire [0:0] CLBLM_R_X5Y152_SLICE_X7Y152_D6;
  wire [0:0] CLBLM_R_X5Y152_SLICE_X7Y152_DO5;
  wire [0:0] CLBLM_R_X5Y152_SLICE_X7Y152_DO6;
  wire [0:0] CLBLM_R_X5Y152_SLICE_X7Y152_DQ;
  wire [0:0] CLBLM_R_X5Y152_SLICE_X7Y152_D_CY;
  wire [0:0] CLBLM_R_X5Y152_SLICE_X7Y152_D_XOR;
  wire [0:0] CLBLM_R_X5Y153_SLICE_X6Y153_A;
  wire [0:0] CLBLM_R_X5Y153_SLICE_X6Y153_A1;
  wire [0:0] CLBLM_R_X5Y153_SLICE_X6Y153_A2;
  wire [0:0] CLBLM_R_X5Y153_SLICE_X6Y153_A3;
  wire [0:0] CLBLM_R_X5Y153_SLICE_X6Y153_A4;
  wire [0:0] CLBLM_R_X5Y153_SLICE_X6Y153_A5;
  wire [0:0] CLBLM_R_X5Y153_SLICE_X6Y153_A5Q;
  wire [0:0] CLBLM_R_X5Y153_SLICE_X6Y153_A6;
  wire [0:0] CLBLM_R_X5Y153_SLICE_X6Y153_AMUX;
  wire [0:0] CLBLM_R_X5Y153_SLICE_X6Y153_AO5;
  wire [0:0] CLBLM_R_X5Y153_SLICE_X6Y153_AO6;
  wire [0:0] CLBLM_R_X5Y153_SLICE_X6Y153_AQ;
  wire [0:0] CLBLM_R_X5Y153_SLICE_X6Y153_A_CY;
  wire [0:0] CLBLM_R_X5Y153_SLICE_X6Y153_A_XOR;
  wire [0:0] CLBLM_R_X5Y153_SLICE_X6Y153_B;
  wire [0:0] CLBLM_R_X5Y153_SLICE_X6Y153_B1;
  wire [0:0] CLBLM_R_X5Y153_SLICE_X6Y153_B2;
  wire [0:0] CLBLM_R_X5Y153_SLICE_X6Y153_B3;
  wire [0:0] CLBLM_R_X5Y153_SLICE_X6Y153_B4;
  wire [0:0] CLBLM_R_X5Y153_SLICE_X6Y153_B5;
  wire [0:0] CLBLM_R_X5Y153_SLICE_X6Y153_B5Q;
  wire [0:0] CLBLM_R_X5Y153_SLICE_X6Y153_B6;
  wire [0:0] CLBLM_R_X5Y153_SLICE_X6Y153_BMUX;
  wire [0:0] CLBLM_R_X5Y153_SLICE_X6Y153_BO5;
  wire [0:0] CLBLM_R_X5Y153_SLICE_X6Y153_BO6;
  wire [0:0] CLBLM_R_X5Y153_SLICE_X6Y153_BQ;
  wire [0:0] CLBLM_R_X5Y153_SLICE_X6Y153_B_CY;
  wire [0:0] CLBLM_R_X5Y153_SLICE_X6Y153_B_XOR;
  wire [0:0] CLBLM_R_X5Y153_SLICE_X6Y153_C;
  wire [0:0] CLBLM_R_X5Y153_SLICE_X6Y153_C1;
  wire [0:0] CLBLM_R_X5Y153_SLICE_X6Y153_C2;
  wire [0:0] CLBLM_R_X5Y153_SLICE_X6Y153_C3;
  wire [0:0] CLBLM_R_X5Y153_SLICE_X6Y153_C4;
  wire [0:0] CLBLM_R_X5Y153_SLICE_X6Y153_C5;
  wire [0:0] CLBLM_R_X5Y153_SLICE_X6Y153_C6;
  wire [0:0] CLBLM_R_X5Y153_SLICE_X6Y153_CLK;
  wire [0:0] CLBLM_R_X5Y153_SLICE_X6Y153_CO5;
  wire [0:0] CLBLM_R_X5Y153_SLICE_X6Y153_CO6;
  wire [0:0] CLBLM_R_X5Y153_SLICE_X6Y153_CQ;
  wire [0:0] CLBLM_R_X5Y153_SLICE_X6Y153_C_CY;
  wire [0:0] CLBLM_R_X5Y153_SLICE_X6Y153_C_XOR;
  wire [0:0] CLBLM_R_X5Y153_SLICE_X6Y153_D;
  wire [0:0] CLBLM_R_X5Y153_SLICE_X6Y153_D1;
  wire [0:0] CLBLM_R_X5Y153_SLICE_X6Y153_D2;
  wire [0:0] CLBLM_R_X5Y153_SLICE_X6Y153_D3;
  wire [0:0] CLBLM_R_X5Y153_SLICE_X6Y153_D4;
  wire [0:0] CLBLM_R_X5Y153_SLICE_X6Y153_D5;
  wire [0:0] CLBLM_R_X5Y153_SLICE_X6Y153_D5Q;
  wire [0:0] CLBLM_R_X5Y153_SLICE_X6Y153_D6;
  wire [0:0] CLBLM_R_X5Y153_SLICE_X6Y153_DMUX;
  wire [0:0] CLBLM_R_X5Y153_SLICE_X6Y153_DO5;
  wire [0:0] CLBLM_R_X5Y153_SLICE_X6Y153_DO6;
  wire [0:0] CLBLM_R_X5Y153_SLICE_X6Y153_DQ;
  wire [0:0] CLBLM_R_X5Y153_SLICE_X6Y153_D_CY;
  wire [0:0] CLBLM_R_X5Y153_SLICE_X6Y153_D_XOR;
  wire [0:0] CLBLM_R_X5Y153_SLICE_X7Y153_A;
  wire [0:0] CLBLM_R_X5Y153_SLICE_X7Y153_A1;
  wire [0:0] CLBLM_R_X5Y153_SLICE_X7Y153_A2;
  wire [0:0] CLBLM_R_X5Y153_SLICE_X7Y153_A3;
  wire [0:0] CLBLM_R_X5Y153_SLICE_X7Y153_A4;
  wire [0:0] CLBLM_R_X5Y153_SLICE_X7Y153_A5;
  wire [0:0] CLBLM_R_X5Y153_SLICE_X7Y153_A6;
  wire [0:0] CLBLM_R_X5Y153_SLICE_X7Y153_AO5;
  wire [0:0] CLBLM_R_X5Y153_SLICE_X7Y153_AO6;
  wire [0:0] CLBLM_R_X5Y153_SLICE_X7Y153_AQ;
  wire [0:0] CLBLM_R_X5Y153_SLICE_X7Y153_A_CY;
  wire [0:0] CLBLM_R_X5Y153_SLICE_X7Y153_A_XOR;
  wire [0:0] CLBLM_R_X5Y153_SLICE_X7Y153_B;
  wire [0:0] CLBLM_R_X5Y153_SLICE_X7Y153_B1;
  wire [0:0] CLBLM_R_X5Y153_SLICE_X7Y153_B2;
  wire [0:0] CLBLM_R_X5Y153_SLICE_X7Y153_B3;
  wire [0:0] CLBLM_R_X5Y153_SLICE_X7Y153_B4;
  wire [0:0] CLBLM_R_X5Y153_SLICE_X7Y153_B5;
  wire [0:0] CLBLM_R_X5Y153_SLICE_X7Y153_B6;
  wire [0:0] CLBLM_R_X5Y153_SLICE_X7Y153_BO5;
  wire [0:0] CLBLM_R_X5Y153_SLICE_X7Y153_BO6;
  wire [0:0] CLBLM_R_X5Y153_SLICE_X7Y153_BQ;
  wire [0:0] CLBLM_R_X5Y153_SLICE_X7Y153_B_CY;
  wire [0:0] CLBLM_R_X5Y153_SLICE_X7Y153_B_XOR;
  wire [0:0] CLBLM_R_X5Y153_SLICE_X7Y153_C;
  wire [0:0] CLBLM_R_X5Y153_SLICE_X7Y153_C1;
  wire [0:0] CLBLM_R_X5Y153_SLICE_X7Y153_C2;
  wire [0:0] CLBLM_R_X5Y153_SLICE_X7Y153_C3;
  wire [0:0] CLBLM_R_X5Y153_SLICE_X7Y153_C4;
  wire [0:0] CLBLM_R_X5Y153_SLICE_X7Y153_C5;
  wire [0:0] CLBLM_R_X5Y153_SLICE_X7Y153_C6;
  wire [0:0] CLBLM_R_X5Y153_SLICE_X7Y153_CLK;
  wire [0:0] CLBLM_R_X5Y153_SLICE_X7Y153_CO5;
  wire [0:0] CLBLM_R_X5Y153_SLICE_X7Y153_CO6;
  wire [0:0] CLBLM_R_X5Y153_SLICE_X7Y153_CQ;
  wire [0:0] CLBLM_R_X5Y153_SLICE_X7Y153_C_CY;
  wire [0:0] CLBLM_R_X5Y153_SLICE_X7Y153_C_XOR;
  wire [0:0] CLBLM_R_X5Y153_SLICE_X7Y153_D;
  wire [0:0] CLBLM_R_X5Y153_SLICE_X7Y153_D1;
  wire [0:0] CLBLM_R_X5Y153_SLICE_X7Y153_D2;
  wire [0:0] CLBLM_R_X5Y153_SLICE_X7Y153_D3;
  wire [0:0] CLBLM_R_X5Y153_SLICE_X7Y153_D4;
  wire [0:0] CLBLM_R_X5Y153_SLICE_X7Y153_D5;
  wire [0:0] CLBLM_R_X5Y153_SLICE_X7Y153_D6;
  wire [0:0] CLBLM_R_X5Y153_SLICE_X7Y153_DMUX;
  wire [0:0] CLBLM_R_X5Y153_SLICE_X7Y153_DO5;
  wire [0:0] CLBLM_R_X5Y153_SLICE_X7Y153_DO6;
  wire [0:0] CLBLM_R_X5Y153_SLICE_X7Y153_D_CY;
  wire [0:0] CLBLM_R_X5Y153_SLICE_X7Y153_D_XOR;
  wire [0:0] CLBLM_R_X5Y154_SLICE_X6Y154_A;
  wire [0:0] CLBLM_R_X5Y154_SLICE_X6Y154_A1;
  wire [0:0] CLBLM_R_X5Y154_SLICE_X6Y154_A2;
  wire [0:0] CLBLM_R_X5Y154_SLICE_X6Y154_A3;
  wire [0:0] CLBLM_R_X5Y154_SLICE_X6Y154_A4;
  wire [0:0] CLBLM_R_X5Y154_SLICE_X6Y154_A5;
  wire [0:0] CLBLM_R_X5Y154_SLICE_X6Y154_A6;
  wire [0:0] CLBLM_R_X5Y154_SLICE_X6Y154_AO5;
  wire [0:0] CLBLM_R_X5Y154_SLICE_X6Y154_AO6;
  wire [0:0] CLBLM_R_X5Y154_SLICE_X6Y154_AQ;
  wire [0:0] CLBLM_R_X5Y154_SLICE_X6Y154_A_CY;
  wire [0:0] CLBLM_R_X5Y154_SLICE_X6Y154_A_XOR;
  wire [0:0] CLBLM_R_X5Y154_SLICE_X6Y154_B;
  wire [0:0] CLBLM_R_X5Y154_SLICE_X6Y154_B1;
  wire [0:0] CLBLM_R_X5Y154_SLICE_X6Y154_B2;
  wire [0:0] CLBLM_R_X5Y154_SLICE_X6Y154_B3;
  wire [0:0] CLBLM_R_X5Y154_SLICE_X6Y154_B4;
  wire [0:0] CLBLM_R_X5Y154_SLICE_X6Y154_B5;
  wire [0:0] CLBLM_R_X5Y154_SLICE_X6Y154_B6;
  wire [0:0] CLBLM_R_X5Y154_SLICE_X6Y154_BO5;
  wire [0:0] CLBLM_R_X5Y154_SLICE_X6Y154_BO6;
  wire [0:0] CLBLM_R_X5Y154_SLICE_X6Y154_BQ;
  wire [0:0] CLBLM_R_X5Y154_SLICE_X6Y154_B_CY;
  wire [0:0] CLBLM_R_X5Y154_SLICE_X6Y154_B_XOR;
  wire [0:0] CLBLM_R_X5Y154_SLICE_X6Y154_C;
  wire [0:0] CLBLM_R_X5Y154_SLICE_X6Y154_C1;
  wire [0:0] CLBLM_R_X5Y154_SLICE_X6Y154_C2;
  wire [0:0] CLBLM_R_X5Y154_SLICE_X6Y154_C3;
  wire [0:0] CLBLM_R_X5Y154_SLICE_X6Y154_C4;
  wire [0:0] CLBLM_R_X5Y154_SLICE_X6Y154_C5;
  wire [0:0] CLBLM_R_X5Y154_SLICE_X6Y154_C6;
  wire [0:0] CLBLM_R_X5Y154_SLICE_X6Y154_CLK;
  wire [0:0] CLBLM_R_X5Y154_SLICE_X6Y154_CO5;
  wire [0:0] CLBLM_R_X5Y154_SLICE_X6Y154_CO6;
  wire [0:0] CLBLM_R_X5Y154_SLICE_X6Y154_C_CY;
  wire [0:0] CLBLM_R_X5Y154_SLICE_X6Y154_C_XOR;
  wire [0:0] CLBLM_R_X5Y154_SLICE_X6Y154_D;
  wire [0:0] CLBLM_R_X5Y154_SLICE_X6Y154_D1;
  wire [0:0] CLBLM_R_X5Y154_SLICE_X6Y154_D2;
  wire [0:0] CLBLM_R_X5Y154_SLICE_X6Y154_D3;
  wire [0:0] CLBLM_R_X5Y154_SLICE_X6Y154_D4;
  wire [0:0] CLBLM_R_X5Y154_SLICE_X6Y154_D5;
  wire [0:0] CLBLM_R_X5Y154_SLICE_X6Y154_D6;
  wire [0:0] CLBLM_R_X5Y154_SLICE_X6Y154_DO5;
  wire [0:0] CLBLM_R_X5Y154_SLICE_X6Y154_DO6;
  wire [0:0] CLBLM_R_X5Y154_SLICE_X6Y154_D_CY;
  wire [0:0] CLBLM_R_X5Y154_SLICE_X6Y154_D_XOR;
  wire [0:0] CLBLM_R_X5Y154_SLICE_X7Y154_A;
  wire [0:0] CLBLM_R_X5Y154_SLICE_X7Y154_A1;
  wire [0:0] CLBLM_R_X5Y154_SLICE_X7Y154_A2;
  wire [0:0] CLBLM_R_X5Y154_SLICE_X7Y154_A3;
  wire [0:0] CLBLM_R_X5Y154_SLICE_X7Y154_A4;
  wire [0:0] CLBLM_R_X5Y154_SLICE_X7Y154_A5;
  wire [0:0] CLBLM_R_X5Y154_SLICE_X7Y154_A6;
  wire [0:0] CLBLM_R_X5Y154_SLICE_X7Y154_AO5;
  wire [0:0] CLBLM_R_X5Y154_SLICE_X7Y154_AO6;
  wire [0:0] CLBLM_R_X5Y154_SLICE_X7Y154_AQ;
  wire [0:0] CLBLM_R_X5Y154_SLICE_X7Y154_A_CY;
  wire [0:0] CLBLM_R_X5Y154_SLICE_X7Y154_A_XOR;
  wire [0:0] CLBLM_R_X5Y154_SLICE_X7Y154_B;
  wire [0:0] CLBLM_R_X5Y154_SLICE_X7Y154_B1;
  wire [0:0] CLBLM_R_X5Y154_SLICE_X7Y154_B2;
  wire [0:0] CLBLM_R_X5Y154_SLICE_X7Y154_B3;
  wire [0:0] CLBLM_R_X5Y154_SLICE_X7Y154_B4;
  wire [0:0] CLBLM_R_X5Y154_SLICE_X7Y154_B5;
  wire [0:0] CLBLM_R_X5Y154_SLICE_X7Y154_B6;
  wire [0:0] CLBLM_R_X5Y154_SLICE_X7Y154_BO5;
  wire [0:0] CLBLM_R_X5Y154_SLICE_X7Y154_BO6;
  wire [0:0] CLBLM_R_X5Y154_SLICE_X7Y154_B_CY;
  wire [0:0] CLBLM_R_X5Y154_SLICE_X7Y154_B_XOR;
  wire [0:0] CLBLM_R_X5Y154_SLICE_X7Y154_C;
  wire [0:0] CLBLM_R_X5Y154_SLICE_X7Y154_C1;
  wire [0:0] CLBLM_R_X5Y154_SLICE_X7Y154_C2;
  wire [0:0] CLBLM_R_X5Y154_SLICE_X7Y154_C3;
  wire [0:0] CLBLM_R_X5Y154_SLICE_X7Y154_C4;
  wire [0:0] CLBLM_R_X5Y154_SLICE_X7Y154_C5;
  wire [0:0] CLBLM_R_X5Y154_SLICE_X7Y154_C6;
  wire [0:0] CLBLM_R_X5Y154_SLICE_X7Y154_CLK;
  wire [0:0] CLBLM_R_X5Y154_SLICE_X7Y154_CO5;
  wire [0:0] CLBLM_R_X5Y154_SLICE_X7Y154_CO6;
  wire [0:0] CLBLM_R_X5Y154_SLICE_X7Y154_C_CY;
  wire [0:0] CLBLM_R_X5Y154_SLICE_X7Y154_C_XOR;
  wire [0:0] CLBLM_R_X5Y154_SLICE_X7Y154_D;
  wire [0:0] CLBLM_R_X5Y154_SLICE_X7Y154_D1;
  wire [0:0] CLBLM_R_X5Y154_SLICE_X7Y154_D2;
  wire [0:0] CLBLM_R_X5Y154_SLICE_X7Y154_D3;
  wire [0:0] CLBLM_R_X5Y154_SLICE_X7Y154_D4;
  wire [0:0] CLBLM_R_X5Y154_SLICE_X7Y154_D5;
  wire [0:0] CLBLM_R_X5Y154_SLICE_X7Y154_D6;
  wire [0:0] CLBLM_R_X5Y154_SLICE_X7Y154_DO5;
  wire [0:0] CLBLM_R_X5Y154_SLICE_X7Y154_DO6;
  wire [0:0] CLBLM_R_X5Y154_SLICE_X7Y154_D_CY;
  wire [0:0] CLBLM_R_X5Y154_SLICE_X7Y154_D_XOR;
  wire [0:0] CLBLM_R_X7Y141_SLICE_X8Y141_A;
  wire [0:0] CLBLM_R_X7Y141_SLICE_X8Y141_A1;
  wire [0:0] CLBLM_R_X7Y141_SLICE_X8Y141_A2;
  wire [0:0] CLBLM_R_X7Y141_SLICE_X8Y141_A3;
  wire [0:0] CLBLM_R_X7Y141_SLICE_X8Y141_A4;
  wire [0:0] CLBLM_R_X7Y141_SLICE_X8Y141_A5;
  wire [0:0] CLBLM_R_X7Y141_SLICE_X8Y141_A6;
  wire [0:0] CLBLM_R_X7Y141_SLICE_X8Y141_AMUX;
  wire [0:0] CLBLM_R_X7Y141_SLICE_X8Y141_AO5;
  wire [0:0] CLBLM_R_X7Y141_SLICE_X8Y141_AO6;
  wire [0:0] CLBLM_R_X7Y141_SLICE_X8Y141_A_CY;
  wire [0:0] CLBLM_R_X7Y141_SLICE_X8Y141_A_XOR;
  wire [0:0] CLBLM_R_X7Y141_SLICE_X8Y141_B;
  wire [0:0] CLBLM_R_X7Y141_SLICE_X8Y141_B1;
  wire [0:0] CLBLM_R_X7Y141_SLICE_X8Y141_B2;
  wire [0:0] CLBLM_R_X7Y141_SLICE_X8Y141_B3;
  wire [0:0] CLBLM_R_X7Y141_SLICE_X8Y141_B4;
  wire [0:0] CLBLM_R_X7Y141_SLICE_X8Y141_B5;
  wire [0:0] CLBLM_R_X7Y141_SLICE_X8Y141_B6;
  wire [0:0] CLBLM_R_X7Y141_SLICE_X8Y141_BO5;
  wire [0:0] CLBLM_R_X7Y141_SLICE_X8Y141_BO6;
  wire [0:0] CLBLM_R_X7Y141_SLICE_X8Y141_B_CY;
  wire [0:0] CLBLM_R_X7Y141_SLICE_X8Y141_B_XOR;
  wire [0:0] CLBLM_R_X7Y141_SLICE_X8Y141_C;
  wire [0:0] CLBLM_R_X7Y141_SLICE_X8Y141_C1;
  wire [0:0] CLBLM_R_X7Y141_SLICE_X8Y141_C2;
  wire [0:0] CLBLM_R_X7Y141_SLICE_X8Y141_C3;
  wire [0:0] CLBLM_R_X7Y141_SLICE_X8Y141_C4;
  wire [0:0] CLBLM_R_X7Y141_SLICE_X8Y141_C5;
  wire [0:0] CLBLM_R_X7Y141_SLICE_X8Y141_C6;
  wire [0:0] CLBLM_R_X7Y141_SLICE_X8Y141_CO5;
  wire [0:0] CLBLM_R_X7Y141_SLICE_X8Y141_CO6;
  wire [0:0] CLBLM_R_X7Y141_SLICE_X8Y141_C_CY;
  wire [0:0] CLBLM_R_X7Y141_SLICE_X8Y141_C_XOR;
  wire [0:0] CLBLM_R_X7Y141_SLICE_X8Y141_D;
  wire [0:0] CLBLM_R_X7Y141_SLICE_X8Y141_D1;
  wire [0:0] CLBLM_R_X7Y141_SLICE_X8Y141_D2;
  wire [0:0] CLBLM_R_X7Y141_SLICE_X8Y141_D3;
  wire [0:0] CLBLM_R_X7Y141_SLICE_X8Y141_D4;
  wire [0:0] CLBLM_R_X7Y141_SLICE_X8Y141_D5;
  wire [0:0] CLBLM_R_X7Y141_SLICE_X8Y141_D6;
  wire [0:0] CLBLM_R_X7Y141_SLICE_X8Y141_DO5;
  wire [0:0] CLBLM_R_X7Y141_SLICE_X8Y141_DO6;
  wire [0:0] CLBLM_R_X7Y141_SLICE_X8Y141_D_CY;
  wire [0:0] CLBLM_R_X7Y141_SLICE_X8Y141_D_XOR;
  wire [0:0] CLBLM_R_X7Y141_SLICE_X9Y141_A;
  wire [0:0] CLBLM_R_X7Y141_SLICE_X9Y141_A1;
  wire [0:0] CLBLM_R_X7Y141_SLICE_X9Y141_A2;
  wire [0:0] CLBLM_R_X7Y141_SLICE_X9Y141_A3;
  wire [0:0] CLBLM_R_X7Y141_SLICE_X9Y141_A4;
  wire [0:0] CLBLM_R_X7Y141_SLICE_X9Y141_A5;
  wire [0:0] CLBLM_R_X7Y141_SLICE_X9Y141_A6;
  wire [0:0] CLBLM_R_X7Y141_SLICE_X9Y141_AO5;
  wire [0:0] CLBLM_R_X7Y141_SLICE_X9Y141_AO6;
  wire [0:0] CLBLM_R_X7Y141_SLICE_X9Y141_AQ;
  wire [0:0] CLBLM_R_X7Y141_SLICE_X9Y141_A_CY;
  wire [0:0] CLBLM_R_X7Y141_SLICE_X9Y141_A_XOR;
  wire [0:0] CLBLM_R_X7Y141_SLICE_X9Y141_B;
  wire [0:0] CLBLM_R_X7Y141_SLICE_X9Y141_B1;
  wire [0:0] CLBLM_R_X7Y141_SLICE_X9Y141_B2;
  wire [0:0] CLBLM_R_X7Y141_SLICE_X9Y141_B3;
  wire [0:0] CLBLM_R_X7Y141_SLICE_X9Y141_B4;
  wire [0:0] CLBLM_R_X7Y141_SLICE_X9Y141_B5;
  wire [0:0] CLBLM_R_X7Y141_SLICE_X9Y141_B6;
  wire [0:0] CLBLM_R_X7Y141_SLICE_X9Y141_BO5;
  wire [0:0] CLBLM_R_X7Y141_SLICE_X9Y141_BO6;
  wire [0:0] CLBLM_R_X7Y141_SLICE_X9Y141_B_CY;
  wire [0:0] CLBLM_R_X7Y141_SLICE_X9Y141_B_XOR;
  wire [0:0] CLBLM_R_X7Y141_SLICE_X9Y141_C;
  wire [0:0] CLBLM_R_X7Y141_SLICE_X9Y141_C1;
  wire [0:0] CLBLM_R_X7Y141_SLICE_X9Y141_C2;
  wire [0:0] CLBLM_R_X7Y141_SLICE_X9Y141_C3;
  wire [0:0] CLBLM_R_X7Y141_SLICE_X9Y141_C4;
  wire [0:0] CLBLM_R_X7Y141_SLICE_X9Y141_C5;
  wire [0:0] CLBLM_R_X7Y141_SLICE_X9Y141_C6;
  wire [0:0] CLBLM_R_X7Y141_SLICE_X9Y141_CLK;
  wire [0:0] CLBLM_R_X7Y141_SLICE_X9Y141_CO5;
  wire [0:0] CLBLM_R_X7Y141_SLICE_X9Y141_CO6;
  wire [0:0] CLBLM_R_X7Y141_SLICE_X9Y141_C_CY;
  wire [0:0] CLBLM_R_X7Y141_SLICE_X9Y141_C_XOR;
  wire [0:0] CLBLM_R_X7Y141_SLICE_X9Y141_D;
  wire [0:0] CLBLM_R_X7Y141_SLICE_X9Y141_D1;
  wire [0:0] CLBLM_R_X7Y141_SLICE_X9Y141_D2;
  wire [0:0] CLBLM_R_X7Y141_SLICE_X9Y141_D3;
  wire [0:0] CLBLM_R_X7Y141_SLICE_X9Y141_D4;
  wire [0:0] CLBLM_R_X7Y141_SLICE_X9Y141_D5;
  wire [0:0] CLBLM_R_X7Y141_SLICE_X9Y141_D6;
  wire [0:0] CLBLM_R_X7Y141_SLICE_X9Y141_DO5;
  wire [0:0] CLBLM_R_X7Y141_SLICE_X9Y141_DO6;
  wire [0:0] CLBLM_R_X7Y141_SLICE_X9Y141_D_CY;
  wire [0:0] CLBLM_R_X7Y141_SLICE_X9Y141_D_XOR;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X8Y142_A;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X8Y142_A1;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X8Y142_A2;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X8Y142_A3;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X8Y142_A4;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X8Y142_A5;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X8Y142_A6;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X8Y142_AO5;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X8Y142_AO6;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X8Y142_AQ;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X8Y142_A_CY;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X8Y142_A_XOR;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X8Y142_B;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X8Y142_B1;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X8Y142_B2;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X8Y142_B3;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X8Y142_B4;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X8Y142_B5;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X8Y142_B6;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X8Y142_BO5;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X8Y142_BO6;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X8Y142_BQ;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X8Y142_B_CY;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X8Y142_B_XOR;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X8Y142_C;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X8Y142_C1;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X8Y142_C2;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X8Y142_C3;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X8Y142_C4;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X8Y142_C5;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X8Y142_C5Q;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X8Y142_C6;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X8Y142_CLK;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X8Y142_CMUX;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X8Y142_CO5;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X8Y142_CO6;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X8Y142_CQ;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X8Y142_C_CY;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X8Y142_C_XOR;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X8Y142_D;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X8Y142_D1;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X8Y142_D2;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X8Y142_D3;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X8Y142_D4;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X8Y142_D5;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X8Y142_D5Q;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X8Y142_D6;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X8Y142_DMUX;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X8Y142_DO5;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X8Y142_DO6;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X8Y142_DQ;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X8Y142_D_CY;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X8Y142_D_XOR;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X9Y142_A;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X9Y142_A1;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X9Y142_A2;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X9Y142_A3;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X9Y142_A4;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X9Y142_A5;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X9Y142_A6;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X9Y142_AO5;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X9Y142_AO6;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X9Y142_AQ;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X9Y142_A_CY;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X9Y142_A_XOR;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X9Y142_B;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X9Y142_B1;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X9Y142_B2;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X9Y142_B3;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X9Y142_B4;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X9Y142_B5;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X9Y142_B6;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X9Y142_BO5;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X9Y142_BO6;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X9Y142_BQ;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X9Y142_B_CY;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X9Y142_B_XOR;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X9Y142_C;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X9Y142_C1;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X9Y142_C2;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X9Y142_C3;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X9Y142_C4;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X9Y142_C5;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X9Y142_C6;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X9Y142_CLK;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X9Y142_CO5;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X9Y142_CO6;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X9Y142_CQ;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X9Y142_C_CY;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X9Y142_C_XOR;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X9Y142_D;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X9Y142_D1;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X9Y142_D2;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X9Y142_D3;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X9Y142_D4;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X9Y142_D5;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X9Y142_D6;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X9Y142_DO5;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X9Y142_DO6;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X9Y142_D_CY;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X9Y142_D_XOR;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X8Y143_A;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X8Y143_A1;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X8Y143_A2;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X8Y143_A3;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X8Y143_A4;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X8Y143_A5;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X8Y143_A6;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X8Y143_AO5;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X8Y143_AO6;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X8Y143_AQ;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X8Y143_A_CY;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X8Y143_A_XOR;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X8Y143_B;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X8Y143_B1;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X8Y143_B2;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X8Y143_B3;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X8Y143_B4;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X8Y143_B5;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X8Y143_B6;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X8Y143_BO5;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X8Y143_BO6;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X8Y143_BQ;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X8Y143_B_CY;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X8Y143_B_XOR;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X8Y143_C;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X8Y143_C1;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X8Y143_C2;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X8Y143_C3;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X8Y143_C4;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X8Y143_C5;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X8Y143_C6;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X8Y143_CLK;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X8Y143_CMUX;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X8Y143_CO5;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X8Y143_CO6;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X8Y143_C_CY;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X8Y143_C_XOR;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X8Y143_D;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X8Y143_D1;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X8Y143_D2;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X8Y143_D3;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X8Y143_D4;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X8Y143_D5;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X8Y143_D6;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X8Y143_DO5;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X8Y143_DO6;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X8Y143_D_CY;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X8Y143_D_XOR;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X9Y143_A;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X9Y143_A1;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X9Y143_A2;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X9Y143_A3;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X9Y143_A4;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X9Y143_A5;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X9Y143_A6;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X9Y143_AO5;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X9Y143_AO6;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X9Y143_AQ;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X9Y143_A_CY;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X9Y143_A_XOR;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X9Y143_B;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X9Y143_B1;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X9Y143_B2;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X9Y143_B3;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X9Y143_B4;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X9Y143_B5;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X9Y143_B5Q;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X9Y143_B6;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X9Y143_BMUX;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X9Y143_BO5;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X9Y143_BO6;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X9Y143_BQ;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X9Y143_B_CY;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X9Y143_B_XOR;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X9Y143_C;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X9Y143_C1;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X9Y143_C2;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X9Y143_C3;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X9Y143_C4;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X9Y143_C5;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X9Y143_C6;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X9Y143_CLK;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X9Y143_CO5;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X9Y143_CO6;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X9Y143_CQ;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X9Y143_C_CY;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X9Y143_C_XOR;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X9Y143_D;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X9Y143_D1;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X9Y143_D2;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X9Y143_D3;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X9Y143_D4;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X9Y143_D5;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X9Y143_D6;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X9Y143_DO5;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X9Y143_DO6;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X9Y143_D_CY;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X9Y143_D_XOR;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X8Y144_A;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X8Y144_A1;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X8Y144_A2;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X8Y144_A3;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X8Y144_A4;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X8Y144_A5;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X8Y144_A6;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X8Y144_AO5;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X8Y144_AO6;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X8Y144_AQ;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X8Y144_A_CY;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X8Y144_A_XOR;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X8Y144_B;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X8Y144_B1;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X8Y144_B2;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X8Y144_B3;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X8Y144_B4;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X8Y144_B5;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X8Y144_B5Q;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X8Y144_B6;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X8Y144_BMUX;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X8Y144_BO5;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X8Y144_BO6;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X8Y144_BQ;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X8Y144_B_CY;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X8Y144_B_XOR;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X8Y144_C;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X8Y144_C1;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X8Y144_C2;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X8Y144_C3;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X8Y144_C4;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X8Y144_C5;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X8Y144_C5Q;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X8Y144_C6;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X8Y144_CLK;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X8Y144_CMUX;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X8Y144_CO5;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X8Y144_CO6;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X8Y144_CQ;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X8Y144_C_CY;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X8Y144_C_XOR;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X8Y144_D;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X8Y144_D1;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X8Y144_D2;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X8Y144_D3;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X8Y144_D4;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X8Y144_D5;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X8Y144_D5Q;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X8Y144_D6;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X8Y144_DMUX;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X8Y144_DO5;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X8Y144_DO6;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X8Y144_DQ;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X8Y144_D_CY;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X8Y144_D_XOR;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X9Y144_A;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X9Y144_A1;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X9Y144_A2;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X9Y144_A3;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X9Y144_A4;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X9Y144_A5;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X9Y144_A5Q;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X9Y144_A6;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X9Y144_AMUX;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X9Y144_AO5;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X9Y144_AO6;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X9Y144_AQ;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X9Y144_AX;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X9Y144_A_CY;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X9Y144_A_XOR;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X9Y144_B;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X9Y144_B1;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X9Y144_B2;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X9Y144_B3;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X9Y144_B4;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X9Y144_B5;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X9Y144_B5Q;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X9Y144_B6;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X9Y144_BMUX;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X9Y144_BO5;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X9Y144_BO6;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X9Y144_BQ;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X9Y144_B_CY;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X9Y144_B_XOR;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X9Y144_C;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X9Y144_C1;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X9Y144_C2;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X9Y144_C3;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X9Y144_C4;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X9Y144_C5;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X9Y144_C6;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X9Y144_CLK;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X9Y144_CO5;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X9Y144_CO6;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X9Y144_C_CY;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X9Y144_C_XOR;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X9Y144_D;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X9Y144_D1;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X9Y144_D2;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X9Y144_D3;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X9Y144_D4;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X9Y144_D5;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X9Y144_D6;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X9Y144_DO5;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X9Y144_DO6;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X9Y144_D_CY;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X9Y144_D_XOR;
  wire [0:0] CLBLM_R_X7Y145_SLICE_X8Y145_A;
  wire [0:0] CLBLM_R_X7Y145_SLICE_X8Y145_A1;
  wire [0:0] CLBLM_R_X7Y145_SLICE_X8Y145_A2;
  wire [0:0] CLBLM_R_X7Y145_SLICE_X8Y145_A3;
  wire [0:0] CLBLM_R_X7Y145_SLICE_X8Y145_A4;
  wire [0:0] CLBLM_R_X7Y145_SLICE_X8Y145_A5;
  wire [0:0] CLBLM_R_X7Y145_SLICE_X8Y145_A5Q;
  wire [0:0] CLBLM_R_X7Y145_SLICE_X8Y145_A6;
  wire [0:0] CLBLM_R_X7Y145_SLICE_X8Y145_AMUX;
  wire [0:0] CLBLM_R_X7Y145_SLICE_X8Y145_AO5;
  wire [0:0] CLBLM_R_X7Y145_SLICE_X8Y145_AO6;
  wire [0:0] CLBLM_R_X7Y145_SLICE_X8Y145_AQ;
  wire [0:0] CLBLM_R_X7Y145_SLICE_X8Y145_A_CY;
  wire [0:0] CLBLM_R_X7Y145_SLICE_X8Y145_A_XOR;
  wire [0:0] CLBLM_R_X7Y145_SLICE_X8Y145_B;
  wire [0:0] CLBLM_R_X7Y145_SLICE_X8Y145_B1;
  wire [0:0] CLBLM_R_X7Y145_SLICE_X8Y145_B2;
  wire [0:0] CLBLM_R_X7Y145_SLICE_X8Y145_B3;
  wire [0:0] CLBLM_R_X7Y145_SLICE_X8Y145_B4;
  wire [0:0] CLBLM_R_X7Y145_SLICE_X8Y145_B5;
  wire [0:0] CLBLM_R_X7Y145_SLICE_X8Y145_B5Q;
  wire [0:0] CLBLM_R_X7Y145_SLICE_X8Y145_B6;
  wire [0:0] CLBLM_R_X7Y145_SLICE_X8Y145_BMUX;
  wire [0:0] CLBLM_R_X7Y145_SLICE_X8Y145_BO5;
  wire [0:0] CLBLM_R_X7Y145_SLICE_X8Y145_BO6;
  wire [0:0] CLBLM_R_X7Y145_SLICE_X8Y145_BQ;
  wire [0:0] CLBLM_R_X7Y145_SLICE_X8Y145_B_CY;
  wire [0:0] CLBLM_R_X7Y145_SLICE_X8Y145_B_XOR;
  wire [0:0] CLBLM_R_X7Y145_SLICE_X8Y145_C;
  wire [0:0] CLBLM_R_X7Y145_SLICE_X8Y145_C1;
  wire [0:0] CLBLM_R_X7Y145_SLICE_X8Y145_C2;
  wire [0:0] CLBLM_R_X7Y145_SLICE_X8Y145_C3;
  wire [0:0] CLBLM_R_X7Y145_SLICE_X8Y145_C4;
  wire [0:0] CLBLM_R_X7Y145_SLICE_X8Y145_C5;
  wire [0:0] CLBLM_R_X7Y145_SLICE_X8Y145_C5Q;
  wire [0:0] CLBLM_R_X7Y145_SLICE_X8Y145_C6;
  wire [0:0] CLBLM_R_X7Y145_SLICE_X8Y145_CLK;
  wire [0:0] CLBLM_R_X7Y145_SLICE_X8Y145_CMUX;
  wire [0:0] CLBLM_R_X7Y145_SLICE_X8Y145_CO5;
  wire [0:0] CLBLM_R_X7Y145_SLICE_X8Y145_CO6;
  wire [0:0] CLBLM_R_X7Y145_SLICE_X8Y145_CQ;
  wire [0:0] CLBLM_R_X7Y145_SLICE_X8Y145_C_CY;
  wire [0:0] CLBLM_R_X7Y145_SLICE_X8Y145_C_XOR;
  wire [0:0] CLBLM_R_X7Y145_SLICE_X8Y145_D;
  wire [0:0] CLBLM_R_X7Y145_SLICE_X8Y145_D1;
  wire [0:0] CLBLM_R_X7Y145_SLICE_X8Y145_D2;
  wire [0:0] CLBLM_R_X7Y145_SLICE_X8Y145_D3;
  wire [0:0] CLBLM_R_X7Y145_SLICE_X8Y145_D4;
  wire [0:0] CLBLM_R_X7Y145_SLICE_X8Y145_D5;
  wire [0:0] CLBLM_R_X7Y145_SLICE_X8Y145_D5Q;
  wire [0:0] CLBLM_R_X7Y145_SLICE_X8Y145_D6;
  wire [0:0] CLBLM_R_X7Y145_SLICE_X8Y145_DMUX;
  wire [0:0] CLBLM_R_X7Y145_SLICE_X8Y145_DO5;
  wire [0:0] CLBLM_R_X7Y145_SLICE_X8Y145_DO6;
  wire [0:0] CLBLM_R_X7Y145_SLICE_X8Y145_DQ;
  wire [0:0] CLBLM_R_X7Y145_SLICE_X8Y145_D_CY;
  wire [0:0] CLBLM_R_X7Y145_SLICE_X8Y145_D_XOR;
  wire [0:0] CLBLM_R_X7Y145_SLICE_X9Y145_A;
  wire [0:0] CLBLM_R_X7Y145_SLICE_X9Y145_A1;
  wire [0:0] CLBLM_R_X7Y145_SLICE_X9Y145_A2;
  wire [0:0] CLBLM_R_X7Y145_SLICE_X9Y145_A3;
  wire [0:0] CLBLM_R_X7Y145_SLICE_X9Y145_A4;
  wire [0:0] CLBLM_R_X7Y145_SLICE_X9Y145_A5;
  wire [0:0] CLBLM_R_X7Y145_SLICE_X9Y145_A6;
  wire [0:0] CLBLM_R_X7Y145_SLICE_X9Y145_AO5;
  wire [0:0] CLBLM_R_X7Y145_SLICE_X9Y145_AO6;
  wire [0:0] CLBLM_R_X7Y145_SLICE_X9Y145_A_CY;
  wire [0:0] CLBLM_R_X7Y145_SLICE_X9Y145_A_XOR;
  wire [0:0] CLBLM_R_X7Y145_SLICE_X9Y145_B;
  wire [0:0] CLBLM_R_X7Y145_SLICE_X9Y145_B1;
  wire [0:0] CLBLM_R_X7Y145_SLICE_X9Y145_B2;
  wire [0:0] CLBLM_R_X7Y145_SLICE_X9Y145_B3;
  wire [0:0] CLBLM_R_X7Y145_SLICE_X9Y145_B4;
  wire [0:0] CLBLM_R_X7Y145_SLICE_X9Y145_B5;
  wire [0:0] CLBLM_R_X7Y145_SLICE_X9Y145_B6;
  wire [0:0] CLBLM_R_X7Y145_SLICE_X9Y145_BO5;
  wire [0:0] CLBLM_R_X7Y145_SLICE_X9Y145_BO6;
  wire [0:0] CLBLM_R_X7Y145_SLICE_X9Y145_B_CY;
  wire [0:0] CLBLM_R_X7Y145_SLICE_X9Y145_B_XOR;
  wire [0:0] CLBLM_R_X7Y145_SLICE_X9Y145_C;
  wire [0:0] CLBLM_R_X7Y145_SLICE_X9Y145_C1;
  wire [0:0] CLBLM_R_X7Y145_SLICE_X9Y145_C2;
  wire [0:0] CLBLM_R_X7Y145_SLICE_X9Y145_C3;
  wire [0:0] CLBLM_R_X7Y145_SLICE_X9Y145_C4;
  wire [0:0] CLBLM_R_X7Y145_SLICE_X9Y145_C5;
  wire [0:0] CLBLM_R_X7Y145_SLICE_X9Y145_C6;
  wire [0:0] CLBLM_R_X7Y145_SLICE_X9Y145_CO5;
  wire [0:0] CLBLM_R_X7Y145_SLICE_X9Y145_CO6;
  wire [0:0] CLBLM_R_X7Y145_SLICE_X9Y145_C_CY;
  wire [0:0] CLBLM_R_X7Y145_SLICE_X9Y145_C_XOR;
  wire [0:0] CLBLM_R_X7Y145_SLICE_X9Y145_D;
  wire [0:0] CLBLM_R_X7Y145_SLICE_X9Y145_D1;
  wire [0:0] CLBLM_R_X7Y145_SLICE_X9Y145_D2;
  wire [0:0] CLBLM_R_X7Y145_SLICE_X9Y145_D3;
  wire [0:0] CLBLM_R_X7Y145_SLICE_X9Y145_D4;
  wire [0:0] CLBLM_R_X7Y145_SLICE_X9Y145_D5;
  wire [0:0] CLBLM_R_X7Y145_SLICE_X9Y145_D6;
  wire [0:0] CLBLM_R_X7Y145_SLICE_X9Y145_DMUX;
  wire [0:0] CLBLM_R_X7Y145_SLICE_X9Y145_DO5;
  wire [0:0] CLBLM_R_X7Y145_SLICE_X9Y145_DO6;
  wire [0:0] CLBLM_R_X7Y145_SLICE_X9Y145_D_CY;
  wire [0:0] CLBLM_R_X7Y145_SLICE_X9Y145_D_XOR;
  wire [0:0] CLBLM_R_X7Y146_SLICE_X8Y146_A;
  wire [0:0] CLBLM_R_X7Y146_SLICE_X8Y146_A1;
  wire [0:0] CLBLM_R_X7Y146_SLICE_X8Y146_A2;
  wire [0:0] CLBLM_R_X7Y146_SLICE_X8Y146_A3;
  wire [0:0] CLBLM_R_X7Y146_SLICE_X8Y146_A4;
  wire [0:0] CLBLM_R_X7Y146_SLICE_X8Y146_A5;
  wire [0:0] CLBLM_R_X7Y146_SLICE_X8Y146_A5Q;
  wire [0:0] CLBLM_R_X7Y146_SLICE_X8Y146_A6;
  wire [0:0] CLBLM_R_X7Y146_SLICE_X8Y146_AMUX;
  wire [0:0] CLBLM_R_X7Y146_SLICE_X8Y146_AO5;
  wire [0:0] CLBLM_R_X7Y146_SLICE_X8Y146_AO6;
  wire [0:0] CLBLM_R_X7Y146_SLICE_X8Y146_AQ;
  wire [0:0] CLBLM_R_X7Y146_SLICE_X8Y146_A_CY;
  wire [0:0] CLBLM_R_X7Y146_SLICE_X8Y146_A_XOR;
  wire [0:0] CLBLM_R_X7Y146_SLICE_X8Y146_B;
  wire [0:0] CLBLM_R_X7Y146_SLICE_X8Y146_B1;
  wire [0:0] CLBLM_R_X7Y146_SLICE_X8Y146_B2;
  wire [0:0] CLBLM_R_X7Y146_SLICE_X8Y146_B3;
  wire [0:0] CLBLM_R_X7Y146_SLICE_X8Y146_B4;
  wire [0:0] CLBLM_R_X7Y146_SLICE_X8Y146_B5;
  wire [0:0] CLBLM_R_X7Y146_SLICE_X8Y146_B5Q;
  wire [0:0] CLBLM_R_X7Y146_SLICE_X8Y146_B6;
  wire [0:0] CLBLM_R_X7Y146_SLICE_X8Y146_BMUX;
  wire [0:0] CLBLM_R_X7Y146_SLICE_X8Y146_BO5;
  wire [0:0] CLBLM_R_X7Y146_SLICE_X8Y146_BO6;
  wire [0:0] CLBLM_R_X7Y146_SLICE_X8Y146_BQ;
  wire [0:0] CLBLM_R_X7Y146_SLICE_X8Y146_B_CY;
  wire [0:0] CLBLM_R_X7Y146_SLICE_X8Y146_B_XOR;
  wire [0:0] CLBLM_R_X7Y146_SLICE_X8Y146_C;
  wire [0:0] CLBLM_R_X7Y146_SLICE_X8Y146_C1;
  wire [0:0] CLBLM_R_X7Y146_SLICE_X8Y146_C2;
  wire [0:0] CLBLM_R_X7Y146_SLICE_X8Y146_C3;
  wire [0:0] CLBLM_R_X7Y146_SLICE_X8Y146_C4;
  wire [0:0] CLBLM_R_X7Y146_SLICE_X8Y146_C5;
  wire [0:0] CLBLM_R_X7Y146_SLICE_X8Y146_C5Q;
  wire [0:0] CLBLM_R_X7Y146_SLICE_X8Y146_C6;
  wire [0:0] CLBLM_R_X7Y146_SLICE_X8Y146_CLK;
  wire [0:0] CLBLM_R_X7Y146_SLICE_X8Y146_CMUX;
  wire [0:0] CLBLM_R_X7Y146_SLICE_X8Y146_CO5;
  wire [0:0] CLBLM_R_X7Y146_SLICE_X8Y146_CO6;
  wire [0:0] CLBLM_R_X7Y146_SLICE_X8Y146_CQ;
  wire [0:0] CLBLM_R_X7Y146_SLICE_X8Y146_C_CY;
  wire [0:0] CLBLM_R_X7Y146_SLICE_X8Y146_C_XOR;
  wire [0:0] CLBLM_R_X7Y146_SLICE_X8Y146_D;
  wire [0:0] CLBLM_R_X7Y146_SLICE_X8Y146_D1;
  wire [0:0] CLBLM_R_X7Y146_SLICE_X8Y146_D2;
  wire [0:0] CLBLM_R_X7Y146_SLICE_X8Y146_D3;
  wire [0:0] CLBLM_R_X7Y146_SLICE_X8Y146_D4;
  wire [0:0] CLBLM_R_X7Y146_SLICE_X8Y146_D5;
  wire [0:0] CLBLM_R_X7Y146_SLICE_X8Y146_D5Q;
  wire [0:0] CLBLM_R_X7Y146_SLICE_X8Y146_D6;
  wire [0:0] CLBLM_R_X7Y146_SLICE_X8Y146_DMUX;
  wire [0:0] CLBLM_R_X7Y146_SLICE_X8Y146_DO5;
  wire [0:0] CLBLM_R_X7Y146_SLICE_X8Y146_DO6;
  wire [0:0] CLBLM_R_X7Y146_SLICE_X8Y146_DQ;
  wire [0:0] CLBLM_R_X7Y146_SLICE_X8Y146_D_CY;
  wire [0:0] CLBLM_R_X7Y146_SLICE_X8Y146_D_XOR;
  wire [0:0] CLBLM_R_X7Y146_SLICE_X9Y146_A;
  wire [0:0] CLBLM_R_X7Y146_SLICE_X9Y146_A1;
  wire [0:0] CLBLM_R_X7Y146_SLICE_X9Y146_A2;
  wire [0:0] CLBLM_R_X7Y146_SLICE_X9Y146_A3;
  wire [0:0] CLBLM_R_X7Y146_SLICE_X9Y146_A4;
  wire [0:0] CLBLM_R_X7Y146_SLICE_X9Y146_A5;
  wire [0:0] CLBLM_R_X7Y146_SLICE_X9Y146_A6;
  wire [0:0] CLBLM_R_X7Y146_SLICE_X9Y146_AO5;
  wire [0:0] CLBLM_R_X7Y146_SLICE_X9Y146_AO6;
  wire [0:0] CLBLM_R_X7Y146_SLICE_X9Y146_AQ;
  wire [0:0] CLBLM_R_X7Y146_SLICE_X9Y146_A_CY;
  wire [0:0] CLBLM_R_X7Y146_SLICE_X9Y146_A_XOR;
  wire [0:0] CLBLM_R_X7Y146_SLICE_X9Y146_B;
  wire [0:0] CLBLM_R_X7Y146_SLICE_X9Y146_B1;
  wire [0:0] CLBLM_R_X7Y146_SLICE_X9Y146_B2;
  wire [0:0] CLBLM_R_X7Y146_SLICE_X9Y146_B3;
  wire [0:0] CLBLM_R_X7Y146_SLICE_X9Y146_B4;
  wire [0:0] CLBLM_R_X7Y146_SLICE_X9Y146_B5;
  wire [0:0] CLBLM_R_X7Y146_SLICE_X9Y146_B6;
  wire [0:0] CLBLM_R_X7Y146_SLICE_X9Y146_BO5;
  wire [0:0] CLBLM_R_X7Y146_SLICE_X9Y146_BO6;
  wire [0:0] CLBLM_R_X7Y146_SLICE_X9Y146_BQ;
  wire [0:0] CLBLM_R_X7Y146_SLICE_X9Y146_B_CY;
  wire [0:0] CLBLM_R_X7Y146_SLICE_X9Y146_B_XOR;
  wire [0:0] CLBLM_R_X7Y146_SLICE_X9Y146_C;
  wire [0:0] CLBLM_R_X7Y146_SLICE_X9Y146_C1;
  wire [0:0] CLBLM_R_X7Y146_SLICE_X9Y146_C2;
  wire [0:0] CLBLM_R_X7Y146_SLICE_X9Y146_C3;
  wire [0:0] CLBLM_R_X7Y146_SLICE_X9Y146_C4;
  wire [0:0] CLBLM_R_X7Y146_SLICE_X9Y146_C5;
  wire [0:0] CLBLM_R_X7Y146_SLICE_X9Y146_C6;
  wire [0:0] CLBLM_R_X7Y146_SLICE_X9Y146_CLK;
  wire [0:0] CLBLM_R_X7Y146_SLICE_X9Y146_CMUX;
  wire [0:0] CLBLM_R_X7Y146_SLICE_X9Y146_CO5;
  wire [0:0] CLBLM_R_X7Y146_SLICE_X9Y146_CO6;
  wire [0:0] CLBLM_R_X7Y146_SLICE_X9Y146_C_CY;
  wire [0:0] CLBLM_R_X7Y146_SLICE_X9Y146_C_XOR;
  wire [0:0] CLBLM_R_X7Y146_SLICE_X9Y146_D;
  wire [0:0] CLBLM_R_X7Y146_SLICE_X9Y146_D1;
  wire [0:0] CLBLM_R_X7Y146_SLICE_X9Y146_D2;
  wire [0:0] CLBLM_R_X7Y146_SLICE_X9Y146_D3;
  wire [0:0] CLBLM_R_X7Y146_SLICE_X9Y146_D4;
  wire [0:0] CLBLM_R_X7Y146_SLICE_X9Y146_D5;
  wire [0:0] CLBLM_R_X7Y146_SLICE_X9Y146_D6;
  wire [0:0] CLBLM_R_X7Y146_SLICE_X9Y146_DO5;
  wire [0:0] CLBLM_R_X7Y146_SLICE_X9Y146_DO6;
  wire [0:0] CLBLM_R_X7Y146_SLICE_X9Y146_D_CY;
  wire [0:0] CLBLM_R_X7Y146_SLICE_X9Y146_D_XOR;
  wire [0:0] CLBLM_R_X7Y147_SLICE_X8Y147_A;
  wire [0:0] CLBLM_R_X7Y147_SLICE_X8Y147_A1;
  wire [0:0] CLBLM_R_X7Y147_SLICE_X8Y147_A2;
  wire [0:0] CLBLM_R_X7Y147_SLICE_X8Y147_A3;
  wire [0:0] CLBLM_R_X7Y147_SLICE_X8Y147_A4;
  wire [0:0] CLBLM_R_X7Y147_SLICE_X8Y147_A5;
  wire [0:0] CLBLM_R_X7Y147_SLICE_X8Y147_A6;
  wire [0:0] CLBLM_R_X7Y147_SLICE_X8Y147_AO5;
  wire [0:0] CLBLM_R_X7Y147_SLICE_X8Y147_AO6;
  wire [0:0] CLBLM_R_X7Y147_SLICE_X8Y147_AQ;
  wire [0:0] CLBLM_R_X7Y147_SLICE_X8Y147_AX;
  wire [0:0] CLBLM_R_X7Y147_SLICE_X8Y147_A_CY;
  wire [0:0] CLBLM_R_X7Y147_SLICE_X8Y147_A_XOR;
  wire [0:0] CLBLM_R_X7Y147_SLICE_X8Y147_B;
  wire [0:0] CLBLM_R_X7Y147_SLICE_X8Y147_B1;
  wire [0:0] CLBLM_R_X7Y147_SLICE_X8Y147_B2;
  wire [0:0] CLBLM_R_X7Y147_SLICE_X8Y147_B3;
  wire [0:0] CLBLM_R_X7Y147_SLICE_X8Y147_B4;
  wire [0:0] CLBLM_R_X7Y147_SLICE_X8Y147_B5;
  wire [0:0] CLBLM_R_X7Y147_SLICE_X8Y147_B6;
  wire [0:0] CLBLM_R_X7Y147_SLICE_X8Y147_BMUX;
  wire [0:0] CLBLM_R_X7Y147_SLICE_X8Y147_BO5;
  wire [0:0] CLBLM_R_X7Y147_SLICE_X8Y147_BO6;
  wire [0:0] CLBLM_R_X7Y147_SLICE_X8Y147_B_CY;
  wire [0:0] CLBLM_R_X7Y147_SLICE_X8Y147_B_XOR;
  wire [0:0] CLBLM_R_X7Y147_SLICE_X8Y147_C;
  wire [0:0] CLBLM_R_X7Y147_SLICE_X8Y147_C1;
  wire [0:0] CLBLM_R_X7Y147_SLICE_X8Y147_C2;
  wire [0:0] CLBLM_R_X7Y147_SLICE_X8Y147_C3;
  wire [0:0] CLBLM_R_X7Y147_SLICE_X8Y147_C4;
  wire [0:0] CLBLM_R_X7Y147_SLICE_X8Y147_C5;
  wire [0:0] CLBLM_R_X7Y147_SLICE_X8Y147_C6;
  wire [0:0] CLBLM_R_X7Y147_SLICE_X8Y147_CE;
  wire [0:0] CLBLM_R_X7Y147_SLICE_X8Y147_CLK;
  wire [0:0] CLBLM_R_X7Y147_SLICE_X8Y147_CMUX;
  wire [0:0] CLBLM_R_X7Y147_SLICE_X8Y147_CO5;
  wire [0:0] CLBLM_R_X7Y147_SLICE_X8Y147_CO6;
  wire [0:0] CLBLM_R_X7Y147_SLICE_X8Y147_C_CY;
  wire [0:0] CLBLM_R_X7Y147_SLICE_X8Y147_C_XOR;
  wire [0:0] CLBLM_R_X7Y147_SLICE_X8Y147_D;
  wire [0:0] CLBLM_R_X7Y147_SLICE_X8Y147_D1;
  wire [0:0] CLBLM_R_X7Y147_SLICE_X8Y147_D2;
  wire [0:0] CLBLM_R_X7Y147_SLICE_X8Y147_D3;
  wire [0:0] CLBLM_R_X7Y147_SLICE_X8Y147_D4;
  wire [0:0] CLBLM_R_X7Y147_SLICE_X8Y147_D5;
  wire [0:0] CLBLM_R_X7Y147_SLICE_X8Y147_D6;
  wire [0:0] CLBLM_R_X7Y147_SLICE_X8Y147_DO5;
  wire [0:0] CLBLM_R_X7Y147_SLICE_X8Y147_DO6;
  wire [0:0] CLBLM_R_X7Y147_SLICE_X8Y147_D_CY;
  wire [0:0] CLBLM_R_X7Y147_SLICE_X8Y147_D_XOR;
  wire [0:0] CLBLM_R_X7Y147_SLICE_X9Y147_A;
  wire [0:0] CLBLM_R_X7Y147_SLICE_X9Y147_A1;
  wire [0:0] CLBLM_R_X7Y147_SLICE_X9Y147_A2;
  wire [0:0] CLBLM_R_X7Y147_SLICE_X9Y147_A3;
  wire [0:0] CLBLM_R_X7Y147_SLICE_X9Y147_A4;
  wire [0:0] CLBLM_R_X7Y147_SLICE_X9Y147_A5;
  wire [0:0] CLBLM_R_X7Y147_SLICE_X9Y147_A5Q;
  wire [0:0] CLBLM_R_X7Y147_SLICE_X9Y147_A6;
  wire [0:0] CLBLM_R_X7Y147_SLICE_X9Y147_AMUX;
  wire [0:0] CLBLM_R_X7Y147_SLICE_X9Y147_AO5;
  wire [0:0] CLBLM_R_X7Y147_SLICE_X9Y147_AO6;
  wire [0:0] CLBLM_R_X7Y147_SLICE_X9Y147_AQ;
  wire [0:0] CLBLM_R_X7Y147_SLICE_X9Y147_A_CY;
  wire [0:0] CLBLM_R_X7Y147_SLICE_X9Y147_A_XOR;
  wire [0:0] CLBLM_R_X7Y147_SLICE_X9Y147_B;
  wire [0:0] CLBLM_R_X7Y147_SLICE_X9Y147_B1;
  wire [0:0] CLBLM_R_X7Y147_SLICE_X9Y147_B2;
  wire [0:0] CLBLM_R_X7Y147_SLICE_X9Y147_B3;
  wire [0:0] CLBLM_R_X7Y147_SLICE_X9Y147_B4;
  wire [0:0] CLBLM_R_X7Y147_SLICE_X9Y147_B5;
  wire [0:0] CLBLM_R_X7Y147_SLICE_X9Y147_B6;
  wire [0:0] CLBLM_R_X7Y147_SLICE_X9Y147_BO5;
  wire [0:0] CLBLM_R_X7Y147_SLICE_X9Y147_BO6;
  wire [0:0] CLBLM_R_X7Y147_SLICE_X9Y147_BQ;
  wire [0:0] CLBLM_R_X7Y147_SLICE_X9Y147_B_CY;
  wire [0:0] CLBLM_R_X7Y147_SLICE_X9Y147_B_XOR;
  wire [0:0] CLBLM_R_X7Y147_SLICE_X9Y147_C;
  wire [0:0] CLBLM_R_X7Y147_SLICE_X9Y147_C1;
  wire [0:0] CLBLM_R_X7Y147_SLICE_X9Y147_C2;
  wire [0:0] CLBLM_R_X7Y147_SLICE_X9Y147_C3;
  wire [0:0] CLBLM_R_X7Y147_SLICE_X9Y147_C4;
  wire [0:0] CLBLM_R_X7Y147_SLICE_X9Y147_C5;
  wire [0:0] CLBLM_R_X7Y147_SLICE_X9Y147_C5Q;
  wire [0:0] CLBLM_R_X7Y147_SLICE_X9Y147_C6;
  wire [0:0] CLBLM_R_X7Y147_SLICE_X9Y147_CLK;
  wire [0:0] CLBLM_R_X7Y147_SLICE_X9Y147_CMUX;
  wire [0:0] CLBLM_R_X7Y147_SLICE_X9Y147_CO5;
  wire [0:0] CLBLM_R_X7Y147_SLICE_X9Y147_CO6;
  wire [0:0] CLBLM_R_X7Y147_SLICE_X9Y147_CQ;
  wire [0:0] CLBLM_R_X7Y147_SLICE_X9Y147_C_CY;
  wire [0:0] CLBLM_R_X7Y147_SLICE_X9Y147_C_XOR;
  wire [0:0] CLBLM_R_X7Y147_SLICE_X9Y147_D;
  wire [0:0] CLBLM_R_X7Y147_SLICE_X9Y147_D1;
  wire [0:0] CLBLM_R_X7Y147_SLICE_X9Y147_D2;
  wire [0:0] CLBLM_R_X7Y147_SLICE_X9Y147_D3;
  wire [0:0] CLBLM_R_X7Y147_SLICE_X9Y147_D4;
  wire [0:0] CLBLM_R_X7Y147_SLICE_X9Y147_D5;
  wire [0:0] CLBLM_R_X7Y147_SLICE_X9Y147_D5Q;
  wire [0:0] CLBLM_R_X7Y147_SLICE_X9Y147_D6;
  wire [0:0] CLBLM_R_X7Y147_SLICE_X9Y147_DMUX;
  wire [0:0] CLBLM_R_X7Y147_SLICE_X9Y147_DO5;
  wire [0:0] CLBLM_R_X7Y147_SLICE_X9Y147_DO6;
  wire [0:0] CLBLM_R_X7Y147_SLICE_X9Y147_DQ;
  wire [0:0] CLBLM_R_X7Y147_SLICE_X9Y147_D_CY;
  wire [0:0] CLBLM_R_X7Y147_SLICE_X9Y147_D_XOR;
  wire [0:0] CLBLM_R_X7Y148_SLICE_X8Y148_A;
  wire [0:0] CLBLM_R_X7Y148_SLICE_X8Y148_A1;
  wire [0:0] CLBLM_R_X7Y148_SLICE_X8Y148_A2;
  wire [0:0] CLBLM_R_X7Y148_SLICE_X8Y148_A3;
  wire [0:0] CLBLM_R_X7Y148_SLICE_X8Y148_A4;
  wire [0:0] CLBLM_R_X7Y148_SLICE_X8Y148_A5;
  wire [0:0] CLBLM_R_X7Y148_SLICE_X8Y148_A6;
  wire [0:0] CLBLM_R_X7Y148_SLICE_X8Y148_AMUX;
  wire [0:0] CLBLM_R_X7Y148_SLICE_X8Y148_AO5;
  wire [0:0] CLBLM_R_X7Y148_SLICE_X8Y148_AO6;
  wire [0:0] CLBLM_R_X7Y148_SLICE_X8Y148_AQ;
  wire [0:0] CLBLM_R_X7Y148_SLICE_X8Y148_AX;
  wire [0:0] CLBLM_R_X7Y148_SLICE_X8Y148_A_CY;
  wire [0:0] CLBLM_R_X7Y148_SLICE_X8Y148_A_XOR;
  wire [0:0] CLBLM_R_X7Y148_SLICE_X8Y148_B;
  wire [0:0] CLBLM_R_X7Y148_SLICE_X8Y148_B1;
  wire [0:0] CLBLM_R_X7Y148_SLICE_X8Y148_B2;
  wire [0:0] CLBLM_R_X7Y148_SLICE_X8Y148_B3;
  wire [0:0] CLBLM_R_X7Y148_SLICE_X8Y148_B4;
  wire [0:0] CLBLM_R_X7Y148_SLICE_X8Y148_B5;
  wire [0:0] CLBLM_R_X7Y148_SLICE_X8Y148_B6;
  wire [0:0] CLBLM_R_X7Y148_SLICE_X8Y148_BO5;
  wire [0:0] CLBLM_R_X7Y148_SLICE_X8Y148_BO6;
  wire [0:0] CLBLM_R_X7Y148_SLICE_X8Y148_B_CY;
  wire [0:0] CLBLM_R_X7Y148_SLICE_X8Y148_B_XOR;
  wire [0:0] CLBLM_R_X7Y148_SLICE_X8Y148_C;
  wire [0:0] CLBLM_R_X7Y148_SLICE_X8Y148_C1;
  wire [0:0] CLBLM_R_X7Y148_SLICE_X8Y148_C2;
  wire [0:0] CLBLM_R_X7Y148_SLICE_X8Y148_C3;
  wire [0:0] CLBLM_R_X7Y148_SLICE_X8Y148_C4;
  wire [0:0] CLBLM_R_X7Y148_SLICE_X8Y148_C5;
  wire [0:0] CLBLM_R_X7Y148_SLICE_X8Y148_C6;
  wire [0:0] CLBLM_R_X7Y148_SLICE_X8Y148_CE;
  wire [0:0] CLBLM_R_X7Y148_SLICE_X8Y148_CLK;
  wire [0:0] CLBLM_R_X7Y148_SLICE_X8Y148_CO5;
  wire [0:0] CLBLM_R_X7Y148_SLICE_X8Y148_CO6;
  wire [0:0] CLBLM_R_X7Y148_SLICE_X8Y148_C_CY;
  wire [0:0] CLBLM_R_X7Y148_SLICE_X8Y148_C_XOR;
  wire [0:0] CLBLM_R_X7Y148_SLICE_X8Y148_D;
  wire [0:0] CLBLM_R_X7Y148_SLICE_X8Y148_D1;
  wire [0:0] CLBLM_R_X7Y148_SLICE_X8Y148_D2;
  wire [0:0] CLBLM_R_X7Y148_SLICE_X8Y148_D3;
  wire [0:0] CLBLM_R_X7Y148_SLICE_X8Y148_D4;
  wire [0:0] CLBLM_R_X7Y148_SLICE_X8Y148_D5;
  wire [0:0] CLBLM_R_X7Y148_SLICE_X8Y148_D6;
  wire [0:0] CLBLM_R_X7Y148_SLICE_X8Y148_DO5;
  wire [0:0] CLBLM_R_X7Y148_SLICE_X8Y148_DO6;
  wire [0:0] CLBLM_R_X7Y148_SLICE_X8Y148_D_CY;
  wire [0:0] CLBLM_R_X7Y148_SLICE_X8Y148_D_XOR;
  wire [0:0] CLBLM_R_X7Y148_SLICE_X9Y148_A;
  wire [0:0] CLBLM_R_X7Y148_SLICE_X9Y148_A1;
  wire [0:0] CLBLM_R_X7Y148_SLICE_X9Y148_A2;
  wire [0:0] CLBLM_R_X7Y148_SLICE_X9Y148_A3;
  wire [0:0] CLBLM_R_X7Y148_SLICE_X9Y148_A4;
  wire [0:0] CLBLM_R_X7Y148_SLICE_X9Y148_A5;
  wire [0:0] CLBLM_R_X7Y148_SLICE_X9Y148_A5Q;
  wire [0:0] CLBLM_R_X7Y148_SLICE_X9Y148_A6;
  wire [0:0] CLBLM_R_X7Y148_SLICE_X9Y148_AMUX;
  wire [0:0] CLBLM_R_X7Y148_SLICE_X9Y148_AO5;
  wire [0:0] CLBLM_R_X7Y148_SLICE_X9Y148_AO6;
  wire [0:0] CLBLM_R_X7Y148_SLICE_X9Y148_AQ;
  wire [0:0] CLBLM_R_X7Y148_SLICE_X9Y148_A_CY;
  wire [0:0] CLBLM_R_X7Y148_SLICE_X9Y148_A_XOR;
  wire [0:0] CLBLM_R_X7Y148_SLICE_X9Y148_B;
  wire [0:0] CLBLM_R_X7Y148_SLICE_X9Y148_B1;
  wire [0:0] CLBLM_R_X7Y148_SLICE_X9Y148_B2;
  wire [0:0] CLBLM_R_X7Y148_SLICE_X9Y148_B3;
  wire [0:0] CLBLM_R_X7Y148_SLICE_X9Y148_B4;
  wire [0:0] CLBLM_R_X7Y148_SLICE_X9Y148_B5;
  wire [0:0] CLBLM_R_X7Y148_SLICE_X9Y148_B6;
  wire [0:0] CLBLM_R_X7Y148_SLICE_X9Y148_BO5;
  wire [0:0] CLBLM_R_X7Y148_SLICE_X9Y148_BO6;
  wire [0:0] CLBLM_R_X7Y148_SLICE_X9Y148_BQ;
  wire [0:0] CLBLM_R_X7Y148_SLICE_X9Y148_B_CY;
  wire [0:0] CLBLM_R_X7Y148_SLICE_X9Y148_B_XOR;
  wire [0:0] CLBLM_R_X7Y148_SLICE_X9Y148_C;
  wire [0:0] CLBLM_R_X7Y148_SLICE_X9Y148_C1;
  wire [0:0] CLBLM_R_X7Y148_SLICE_X9Y148_C2;
  wire [0:0] CLBLM_R_X7Y148_SLICE_X9Y148_C3;
  wire [0:0] CLBLM_R_X7Y148_SLICE_X9Y148_C4;
  wire [0:0] CLBLM_R_X7Y148_SLICE_X9Y148_C5;
  wire [0:0] CLBLM_R_X7Y148_SLICE_X9Y148_C5Q;
  wire [0:0] CLBLM_R_X7Y148_SLICE_X9Y148_C6;
  wire [0:0] CLBLM_R_X7Y148_SLICE_X9Y148_CLK;
  wire [0:0] CLBLM_R_X7Y148_SLICE_X9Y148_CMUX;
  wire [0:0] CLBLM_R_X7Y148_SLICE_X9Y148_CO5;
  wire [0:0] CLBLM_R_X7Y148_SLICE_X9Y148_CO6;
  wire [0:0] CLBLM_R_X7Y148_SLICE_X9Y148_CQ;
  wire [0:0] CLBLM_R_X7Y148_SLICE_X9Y148_C_CY;
  wire [0:0] CLBLM_R_X7Y148_SLICE_X9Y148_C_XOR;
  wire [0:0] CLBLM_R_X7Y148_SLICE_X9Y148_D;
  wire [0:0] CLBLM_R_X7Y148_SLICE_X9Y148_D1;
  wire [0:0] CLBLM_R_X7Y148_SLICE_X9Y148_D2;
  wire [0:0] CLBLM_R_X7Y148_SLICE_X9Y148_D3;
  wire [0:0] CLBLM_R_X7Y148_SLICE_X9Y148_D4;
  wire [0:0] CLBLM_R_X7Y148_SLICE_X9Y148_D5;
  wire [0:0] CLBLM_R_X7Y148_SLICE_X9Y148_D6;
  wire [0:0] CLBLM_R_X7Y148_SLICE_X9Y148_DMUX;
  wire [0:0] CLBLM_R_X7Y148_SLICE_X9Y148_DO5;
  wire [0:0] CLBLM_R_X7Y148_SLICE_X9Y148_DO6;
  wire [0:0] CLBLM_R_X7Y148_SLICE_X9Y148_D_CY;
  wire [0:0] CLBLM_R_X7Y148_SLICE_X9Y148_D_XOR;
  wire [0:0] CLBLM_R_X7Y149_SLICE_X8Y149_A;
  wire [0:0] CLBLM_R_X7Y149_SLICE_X8Y149_A1;
  wire [0:0] CLBLM_R_X7Y149_SLICE_X8Y149_A2;
  wire [0:0] CLBLM_R_X7Y149_SLICE_X8Y149_A3;
  wire [0:0] CLBLM_R_X7Y149_SLICE_X8Y149_A4;
  wire [0:0] CLBLM_R_X7Y149_SLICE_X8Y149_A5;
  wire [0:0] CLBLM_R_X7Y149_SLICE_X8Y149_A5Q;
  wire [0:0] CLBLM_R_X7Y149_SLICE_X8Y149_A6;
  wire [0:0] CLBLM_R_X7Y149_SLICE_X8Y149_AMUX;
  wire [0:0] CLBLM_R_X7Y149_SLICE_X8Y149_AO5;
  wire [0:0] CLBLM_R_X7Y149_SLICE_X8Y149_AO6;
  wire [0:0] CLBLM_R_X7Y149_SLICE_X8Y149_AQ;
  wire [0:0] CLBLM_R_X7Y149_SLICE_X8Y149_A_CY;
  wire [0:0] CLBLM_R_X7Y149_SLICE_X8Y149_A_XOR;
  wire [0:0] CLBLM_R_X7Y149_SLICE_X8Y149_B;
  wire [0:0] CLBLM_R_X7Y149_SLICE_X8Y149_B1;
  wire [0:0] CLBLM_R_X7Y149_SLICE_X8Y149_B2;
  wire [0:0] CLBLM_R_X7Y149_SLICE_X8Y149_B3;
  wire [0:0] CLBLM_R_X7Y149_SLICE_X8Y149_B4;
  wire [0:0] CLBLM_R_X7Y149_SLICE_X8Y149_B5;
  wire [0:0] CLBLM_R_X7Y149_SLICE_X8Y149_B6;
  wire [0:0] CLBLM_R_X7Y149_SLICE_X8Y149_BO5;
  wire [0:0] CLBLM_R_X7Y149_SLICE_X8Y149_BO6;
  wire [0:0] CLBLM_R_X7Y149_SLICE_X8Y149_B_CY;
  wire [0:0] CLBLM_R_X7Y149_SLICE_X8Y149_B_XOR;
  wire [0:0] CLBLM_R_X7Y149_SLICE_X8Y149_C;
  wire [0:0] CLBLM_R_X7Y149_SLICE_X8Y149_C1;
  wire [0:0] CLBLM_R_X7Y149_SLICE_X8Y149_C2;
  wire [0:0] CLBLM_R_X7Y149_SLICE_X8Y149_C3;
  wire [0:0] CLBLM_R_X7Y149_SLICE_X8Y149_C4;
  wire [0:0] CLBLM_R_X7Y149_SLICE_X8Y149_C5;
  wire [0:0] CLBLM_R_X7Y149_SLICE_X8Y149_C6;
  wire [0:0] CLBLM_R_X7Y149_SLICE_X8Y149_CLK;
  wire [0:0] CLBLM_R_X7Y149_SLICE_X8Y149_CO5;
  wire [0:0] CLBLM_R_X7Y149_SLICE_X8Y149_CO6;
  wire [0:0] CLBLM_R_X7Y149_SLICE_X8Y149_C_CY;
  wire [0:0] CLBLM_R_X7Y149_SLICE_X8Y149_C_XOR;
  wire [0:0] CLBLM_R_X7Y149_SLICE_X8Y149_D;
  wire [0:0] CLBLM_R_X7Y149_SLICE_X8Y149_D1;
  wire [0:0] CLBLM_R_X7Y149_SLICE_X8Y149_D2;
  wire [0:0] CLBLM_R_X7Y149_SLICE_X8Y149_D3;
  wire [0:0] CLBLM_R_X7Y149_SLICE_X8Y149_D4;
  wire [0:0] CLBLM_R_X7Y149_SLICE_X8Y149_D5;
  wire [0:0] CLBLM_R_X7Y149_SLICE_X8Y149_D6;
  wire [0:0] CLBLM_R_X7Y149_SLICE_X8Y149_DO5;
  wire [0:0] CLBLM_R_X7Y149_SLICE_X8Y149_DO6;
  wire [0:0] CLBLM_R_X7Y149_SLICE_X8Y149_D_CY;
  wire [0:0] CLBLM_R_X7Y149_SLICE_X8Y149_D_XOR;
  wire [0:0] CLBLM_R_X7Y149_SLICE_X9Y149_A;
  wire [0:0] CLBLM_R_X7Y149_SLICE_X9Y149_A1;
  wire [0:0] CLBLM_R_X7Y149_SLICE_X9Y149_A2;
  wire [0:0] CLBLM_R_X7Y149_SLICE_X9Y149_A3;
  wire [0:0] CLBLM_R_X7Y149_SLICE_X9Y149_A4;
  wire [0:0] CLBLM_R_X7Y149_SLICE_X9Y149_A5;
  wire [0:0] CLBLM_R_X7Y149_SLICE_X9Y149_A5Q;
  wire [0:0] CLBLM_R_X7Y149_SLICE_X9Y149_A6;
  wire [0:0] CLBLM_R_X7Y149_SLICE_X9Y149_AMUX;
  wire [0:0] CLBLM_R_X7Y149_SLICE_X9Y149_AO5;
  wire [0:0] CLBLM_R_X7Y149_SLICE_X9Y149_AO6;
  wire [0:0] CLBLM_R_X7Y149_SLICE_X9Y149_AQ;
  wire [0:0] CLBLM_R_X7Y149_SLICE_X9Y149_A_CY;
  wire [0:0] CLBLM_R_X7Y149_SLICE_X9Y149_A_XOR;
  wire [0:0] CLBLM_R_X7Y149_SLICE_X9Y149_B;
  wire [0:0] CLBLM_R_X7Y149_SLICE_X9Y149_B1;
  wire [0:0] CLBLM_R_X7Y149_SLICE_X9Y149_B2;
  wire [0:0] CLBLM_R_X7Y149_SLICE_X9Y149_B3;
  wire [0:0] CLBLM_R_X7Y149_SLICE_X9Y149_B4;
  wire [0:0] CLBLM_R_X7Y149_SLICE_X9Y149_B5;
  wire [0:0] CLBLM_R_X7Y149_SLICE_X9Y149_B5Q;
  wire [0:0] CLBLM_R_X7Y149_SLICE_X9Y149_B6;
  wire [0:0] CLBLM_R_X7Y149_SLICE_X9Y149_BMUX;
  wire [0:0] CLBLM_R_X7Y149_SLICE_X9Y149_BO5;
  wire [0:0] CLBLM_R_X7Y149_SLICE_X9Y149_BO6;
  wire [0:0] CLBLM_R_X7Y149_SLICE_X9Y149_BQ;
  wire [0:0] CLBLM_R_X7Y149_SLICE_X9Y149_B_CY;
  wire [0:0] CLBLM_R_X7Y149_SLICE_X9Y149_B_XOR;
  wire [0:0] CLBLM_R_X7Y149_SLICE_X9Y149_C;
  wire [0:0] CLBLM_R_X7Y149_SLICE_X9Y149_C1;
  wire [0:0] CLBLM_R_X7Y149_SLICE_X9Y149_C2;
  wire [0:0] CLBLM_R_X7Y149_SLICE_X9Y149_C3;
  wire [0:0] CLBLM_R_X7Y149_SLICE_X9Y149_C4;
  wire [0:0] CLBLM_R_X7Y149_SLICE_X9Y149_C5;
  wire [0:0] CLBLM_R_X7Y149_SLICE_X9Y149_C5Q;
  wire [0:0] CLBLM_R_X7Y149_SLICE_X9Y149_C6;
  wire [0:0] CLBLM_R_X7Y149_SLICE_X9Y149_CLK;
  wire [0:0] CLBLM_R_X7Y149_SLICE_X9Y149_CMUX;
  wire [0:0] CLBLM_R_X7Y149_SLICE_X9Y149_CO5;
  wire [0:0] CLBLM_R_X7Y149_SLICE_X9Y149_CO6;
  wire [0:0] CLBLM_R_X7Y149_SLICE_X9Y149_CQ;
  wire [0:0] CLBLM_R_X7Y149_SLICE_X9Y149_C_CY;
  wire [0:0] CLBLM_R_X7Y149_SLICE_X9Y149_C_XOR;
  wire [0:0] CLBLM_R_X7Y149_SLICE_X9Y149_D;
  wire [0:0] CLBLM_R_X7Y149_SLICE_X9Y149_D1;
  wire [0:0] CLBLM_R_X7Y149_SLICE_X9Y149_D2;
  wire [0:0] CLBLM_R_X7Y149_SLICE_X9Y149_D3;
  wire [0:0] CLBLM_R_X7Y149_SLICE_X9Y149_D4;
  wire [0:0] CLBLM_R_X7Y149_SLICE_X9Y149_D5;
  wire [0:0] CLBLM_R_X7Y149_SLICE_X9Y149_D6;
  wire [0:0] CLBLM_R_X7Y149_SLICE_X9Y149_DO5;
  wire [0:0] CLBLM_R_X7Y149_SLICE_X9Y149_DO6;
  wire [0:0] CLBLM_R_X7Y149_SLICE_X9Y149_D_CY;
  wire [0:0] CLBLM_R_X7Y149_SLICE_X9Y149_D_XOR;
  wire [0:0] CLBLM_R_X7Y150_SLICE_X8Y150_A;
  wire [0:0] CLBLM_R_X7Y150_SLICE_X8Y150_A1;
  wire [0:0] CLBLM_R_X7Y150_SLICE_X8Y150_A2;
  wire [0:0] CLBLM_R_X7Y150_SLICE_X8Y150_A3;
  wire [0:0] CLBLM_R_X7Y150_SLICE_X8Y150_A4;
  wire [0:0] CLBLM_R_X7Y150_SLICE_X8Y150_A5;
  wire [0:0] CLBLM_R_X7Y150_SLICE_X8Y150_A6;
  wire [0:0] CLBLM_R_X7Y150_SLICE_X8Y150_AO5;
  wire [0:0] CLBLM_R_X7Y150_SLICE_X8Y150_AO6;
  wire [0:0] CLBLM_R_X7Y150_SLICE_X8Y150_AQ;
  wire [0:0] CLBLM_R_X7Y150_SLICE_X8Y150_A_CY;
  wire [0:0] CLBLM_R_X7Y150_SLICE_X8Y150_A_XOR;
  wire [0:0] CLBLM_R_X7Y150_SLICE_X8Y150_B;
  wire [0:0] CLBLM_R_X7Y150_SLICE_X8Y150_B1;
  wire [0:0] CLBLM_R_X7Y150_SLICE_X8Y150_B2;
  wire [0:0] CLBLM_R_X7Y150_SLICE_X8Y150_B3;
  wire [0:0] CLBLM_R_X7Y150_SLICE_X8Y150_B4;
  wire [0:0] CLBLM_R_X7Y150_SLICE_X8Y150_B5;
  wire [0:0] CLBLM_R_X7Y150_SLICE_X8Y150_B6;
  wire [0:0] CLBLM_R_X7Y150_SLICE_X8Y150_BMUX;
  wire [0:0] CLBLM_R_X7Y150_SLICE_X8Y150_BO5;
  wire [0:0] CLBLM_R_X7Y150_SLICE_X8Y150_BO6;
  wire [0:0] CLBLM_R_X7Y150_SLICE_X8Y150_B_CY;
  wire [0:0] CLBLM_R_X7Y150_SLICE_X8Y150_B_XOR;
  wire [0:0] CLBLM_R_X7Y150_SLICE_X8Y150_C;
  wire [0:0] CLBLM_R_X7Y150_SLICE_X8Y150_C1;
  wire [0:0] CLBLM_R_X7Y150_SLICE_X8Y150_C2;
  wire [0:0] CLBLM_R_X7Y150_SLICE_X8Y150_C3;
  wire [0:0] CLBLM_R_X7Y150_SLICE_X8Y150_C4;
  wire [0:0] CLBLM_R_X7Y150_SLICE_X8Y150_C5;
  wire [0:0] CLBLM_R_X7Y150_SLICE_X8Y150_C6;
  wire [0:0] CLBLM_R_X7Y150_SLICE_X8Y150_CLK;
  wire [0:0] CLBLM_R_X7Y150_SLICE_X8Y150_CO5;
  wire [0:0] CLBLM_R_X7Y150_SLICE_X8Y150_CO6;
  wire [0:0] CLBLM_R_X7Y150_SLICE_X8Y150_C_CY;
  wire [0:0] CLBLM_R_X7Y150_SLICE_X8Y150_C_XOR;
  wire [0:0] CLBLM_R_X7Y150_SLICE_X8Y150_D;
  wire [0:0] CLBLM_R_X7Y150_SLICE_X8Y150_D1;
  wire [0:0] CLBLM_R_X7Y150_SLICE_X8Y150_D2;
  wire [0:0] CLBLM_R_X7Y150_SLICE_X8Y150_D3;
  wire [0:0] CLBLM_R_X7Y150_SLICE_X8Y150_D4;
  wire [0:0] CLBLM_R_X7Y150_SLICE_X8Y150_D5;
  wire [0:0] CLBLM_R_X7Y150_SLICE_X8Y150_D6;
  wire [0:0] CLBLM_R_X7Y150_SLICE_X8Y150_DO5;
  wire [0:0] CLBLM_R_X7Y150_SLICE_X8Y150_DO6;
  wire [0:0] CLBLM_R_X7Y150_SLICE_X8Y150_D_CY;
  wire [0:0] CLBLM_R_X7Y150_SLICE_X8Y150_D_XOR;
  wire [0:0] CLBLM_R_X7Y150_SLICE_X9Y150_A;
  wire [0:0] CLBLM_R_X7Y150_SLICE_X9Y150_A1;
  wire [0:0] CLBLM_R_X7Y150_SLICE_X9Y150_A2;
  wire [0:0] CLBLM_R_X7Y150_SLICE_X9Y150_A3;
  wire [0:0] CLBLM_R_X7Y150_SLICE_X9Y150_A4;
  wire [0:0] CLBLM_R_X7Y150_SLICE_X9Y150_A5;
  wire [0:0] CLBLM_R_X7Y150_SLICE_X9Y150_A6;
  wire [0:0] CLBLM_R_X7Y150_SLICE_X9Y150_AO5;
  wire [0:0] CLBLM_R_X7Y150_SLICE_X9Y150_AO6;
  wire [0:0] CLBLM_R_X7Y150_SLICE_X9Y150_A_CY;
  wire [0:0] CLBLM_R_X7Y150_SLICE_X9Y150_A_XOR;
  wire [0:0] CLBLM_R_X7Y150_SLICE_X9Y150_B;
  wire [0:0] CLBLM_R_X7Y150_SLICE_X9Y150_B1;
  wire [0:0] CLBLM_R_X7Y150_SLICE_X9Y150_B2;
  wire [0:0] CLBLM_R_X7Y150_SLICE_X9Y150_B3;
  wire [0:0] CLBLM_R_X7Y150_SLICE_X9Y150_B4;
  wire [0:0] CLBLM_R_X7Y150_SLICE_X9Y150_B5;
  wire [0:0] CLBLM_R_X7Y150_SLICE_X9Y150_B6;
  wire [0:0] CLBLM_R_X7Y150_SLICE_X9Y150_BO5;
  wire [0:0] CLBLM_R_X7Y150_SLICE_X9Y150_BO6;
  wire [0:0] CLBLM_R_X7Y150_SLICE_X9Y150_B_CY;
  wire [0:0] CLBLM_R_X7Y150_SLICE_X9Y150_B_XOR;
  wire [0:0] CLBLM_R_X7Y150_SLICE_X9Y150_C;
  wire [0:0] CLBLM_R_X7Y150_SLICE_X9Y150_C1;
  wire [0:0] CLBLM_R_X7Y150_SLICE_X9Y150_C2;
  wire [0:0] CLBLM_R_X7Y150_SLICE_X9Y150_C3;
  wire [0:0] CLBLM_R_X7Y150_SLICE_X9Y150_C4;
  wire [0:0] CLBLM_R_X7Y150_SLICE_X9Y150_C5;
  wire [0:0] CLBLM_R_X7Y150_SLICE_X9Y150_C6;
  wire [0:0] CLBLM_R_X7Y150_SLICE_X9Y150_CO5;
  wire [0:0] CLBLM_R_X7Y150_SLICE_X9Y150_CO6;
  wire [0:0] CLBLM_R_X7Y150_SLICE_X9Y150_C_CY;
  wire [0:0] CLBLM_R_X7Y150_SLICE_X9Y150_C_XOR;
  wire [0:0] CLBLM_R_X7Y150_SLICE_X9Y150_D;
  wire [0:0] CLBLM_R_X7Y150_SLICE_X9Y150_D1;
  wire [0:0] CLBLM_R_X7Y150_SLICE_X9Y150_D2;
  wire [0:0] CLBLM_R_X7Y150_SLICE_X9Y150_D3;
  wire [0:0] CLBLM_R_X7Y150_SLICE_X9Y150_D4;
  wire [0:0] CLBLM_R_X7Y150_SLICE_X9Y150_D5;
  wire [0:0] CLBLM_R_X7Y150_SLICE_X9Y150_D6;
  wire [0:0] CLBLM_R_X7Y150_SLICE_X9Y150_DO5;
  wire [0:0] CLBLM_R_X7Y150_SLICE_X9Y150_DO6;
  wire [0:0] CLBLM_R_X7Y150_SLICE_X9Y150_D_CY;
  wire [0:0] CLBLM_R_X7Y150_SLICE_X9Y150_D_XOR;
  wire [0:0] CLBLM_R_X7Y151_SLICE_X8Y151_A;
  wire [0:0] CLBLM_R_X7Y151_SLICE_X8Y151_A1;
  wire [0:0] CLBLM_R_X7Y151_SLICE_X8Y151_A2;
  wire [0:0] CLBLM_R_X7Y151_SLICE_X8Y151_A3;
  wire [0:0] CLBLM_R_X7Y151_SLICE_X8Y151_A4;
  wire [0:0] CLBLM_R_X7Y151_SLICE_X8Y151_A5;
  wire [0:0] CLBLM_R_X7Y151_SLICE_X8Y151_A6;
  wire [0:0] CLBLM_R_X7Y151_SLICE_X8Y151_AO5;
  wire [0:0] CLBLM_R_X7Y151_SLICE_X8Y151_AO6;
  wire [0:0] CLBLM_R_X7Y151_SLICE_X8Y151_AQ;
  wire [0:0] CLBLM_R_X7Y151_SLICE_X8Y151_A_CY;
  wire [0:0] CLBLM_R_X7Y151_SLICE_X8Y151_A_XOR;
  wire [0:0] CLBLM_R_X7Y151_SLICE_X8Y151_B;
  wire [0:0] CLBLM_R_X7Y151_SLICE_X8Y151_B1;
  wire [0:0] CLBLM_R_X7Y151_SLICE_X8Y151_B2;
  wire [0:0] CLBLM_R_X7Y151_SLICE_X8Y151_B3;
  wire [0:0] CLBLM_R_X7Y151_SLICE_X8Y151_B4;
  wire [0:0] CLBLM_R_X7Y151_SLICE_X8Y151_B5;
  wire [0:0] CLBLM_R_X7Y151_SLICE_X8Y151_B6;
  wire [0:0] CLBLM_R_X7Y151_SLICE_X8Y151_BO5;
  wire [0:0] CLBLM_R_X7Y151_SLICE_X8Y151_BO6;
  wire [0:0] CLBLM_R_X7Y151_SLICE_X8Y151_BQ;
  wire [0:0] CLBLM_R_X7Y151_SLICE_X8Y151_B_CY;
  wire [0:0] CLBLM_R_X7Y151_SLICE_X8Y151_B_XOR;
  wire [0:0] CLBLM_R_X7Y151_SLICE_X8Y151_C;
  wire [0:0] CLBLM_R_X7Y151_SLICE_X8Y151_C1;
  wire [0:0] CLBLM_R_X7Y151_SLICE_X8Y151_C2;
  wire [0:0] CLBLM_R_X7Y151_SLICE_X8Y151_C3;
  wire [0:0] CLBLM_R_X7Y151_SLICE_X8Y151_C4;
  wire [0:0] CLBLM_R_X7Y151_SLICE_X8Y151_C5;
  wire [0:0] CLBLM_R_X7Y151_SLICE_X8Y151_C5Q;
  wire [0:0] CLBLM_R_X7Y151_SLICE_X8Y151_C6;
  wire [0:0] CLBLM_R_X7Y151_SLICE_X8Y151_CLK;
  wire [0:0] CLBLM_R_X7Y151_SLICE_X8Y151_CMUX;
  wire [0:0] CLBLM_R_X7Y151_SLICE_X8Y151_CO5;
  wire [0:0] CLBLM_R_X7Y151_SLICE_X8Y151_CO6;
  wire [0:0] CLBLM_R_X7Y151_SLICE_X8Y151_CQ;
  wire [0:0] CLBLM_R_X7Y151_SLICE_X8Y151_C_CY;
  wire [0:0] CLBLM_R_X7Y151_SLICE_X8Y151_C_XOR;
  wire [0:0] CLBLM_R_X7Y151_SLICE_X8Y151_D;
  wire [0:0] CLBLM_R_X7Y151_SLICE_X8Y151_D1;
  wire [0:0] CLBLM_R_X7Y151_SLICE_X8Y151_D2;
  wire [0:0] CLBLM_R_X7Y151_SLICE_X8Y151_D3;
  wire [0:0] CLBLM_R_X7Y151_SLICE_X8Y151_D4;
  wire [0:0] CLBLM_R_X7Y151_SLICE_X8Y151_D5;
  wire [0:0] CLBLM_R_X7Y151_SLICE_X8Y151_D5Q;
  wire [0:0] CLBLM_R_X7Y151_SLICE_X8Y151_D6;
  wire [0:0] CLBLM_R_X7Y151_SLICE_X8Y151_DMUX;
  wire [0:0] CLBLM_R_X7Y151_SLICE_X8Y151_DO5;
  wire [0:0] CLBLM_R_X7Y151_SLICE_X8Y151_DO6;
  wire [0:0] CLBLM_R_X7Y151_SLICE_X8Y151_DQ;
  wire [0:0] CLBLM_R_X7Y151_SLICE_X8Y151_D_CY;
  wire [0:0] CLBLM_R_X7Y151_SLICE_X8Y151_D_XOR;
  wire [0:0] CLBLM_R_X7Y151_SLICE_X9Y151_A;
  wire [0:0] CLBLM_R_X7Y151_SLICE_X9Y151_A1;
  wire [0:0] CLBLM_R_X7Y151_SLICE_X9Y151_A2;
  wire [0:0] CLBLM_R_X7Y151_SLICE_X9Y151_A3;
  wire [0:0] CLBLM_R_X7Y151_SLICE_X9Y151_A4;
  wire [0:0] CLBLM_R_X7Y151_SLICE_X9Y151_A5;
  wire [0:0] CLBLM_R_X7Y151_SLICE_X9Y151_A5Q;
  wire [0:0] CLBLM_R_X7Y151_SLICE_X9Y151_A6;
  wire [0:0] CLBLM_R_X7Y151_SLICE_X9Y151_AMUX;
  wire [0:0] CLBLM_R_X7Y151_SLICE_X9Y151_AO5;
  wire [0:0] CLBLM_R_X7Y151_SLICE_X9Y151_AO6;
  wire [0:0] CLBLM_R_X7Y151_SLICE_X9Y151_AQ;
  wire [0:0] CLBLM_R_X7Y151_SLICE_X9Y151_AX;
  wire [0:0] CLBLM_R_X7Y151_SLICE_X9Y151_A_CY;
  wire [0:0] CLBLM_R_X7Y151_SLICE_X9Y151_A_XOR;
  wire [0:0] CLBLM_R_X7Y151_SLICE_X9Y151_B;
  wire [0:0] CLBLM_R_X7Y151_SLICE_X9Y151_B1;
  wire [0:0] CLBLM_R_X7Y151_SLICE_X9Y151_B2;
  wire [0:0] CLBLM_R_X7Y151_SLICE_X9Y151_B3;
  wire [0:0] CLBLM_R_X7Y151_SLICE_X9Y151_B4;
  wire [0:0] CLBLM_R_X7Y151_SLICE_X9Y151_B5;
  wire [0:0] CLBLM_R_X7Y151_SLICE_X9Y151_B6;
  wire [0:0] CLBLM_R_X7Y151_SLICE_X9Y151_BO5;
  wire [0:0] CLBLM_R_X7Y151_SLICE_X9Y151_BO6;
  wire [0:0] CLBLM_R_X7Y151_SLICE_X9Y151_BQ;
  wire [0:0] CLBLM_R_X7Y151_SLICE_X9Y151_B_CY;
  wire [0:0] CLBLM_R_X7Y151_SLICE_X9Y151_B_XOR;
  wire [0:0] CLBLM_R_X7Y151_SLICE_X9Y151_C;
  wire [0:0] CLBLM_R_X7Y151_SLICE_X9Y151_C1;
  wire [0:0] CLBLM_R_X7Y151_SLICE_X9Y151_C2;
  wire [0:0] CLBLM_R_X7Y151_SLICE_X9Y151_C3;
  wire [0:0] CLBLM_R_X7Y151_SLICE_X9Y151_C4;
  wire [0:0] CLBLM_R_X7Y151_SLICE_X9Y151_C5;
  wire [0:0] CLBLM_R_X7Y151_SLICE_X9Y151_C5Q;
  wire [0:0] CLBLM_R_X7Y151_SLICE_X9Y151_C6;
  wire [0:0] CLBLM_R_X7Y151_SLICE_X9Y151_CLK;
  wire [0:0] CLBLM_R_X7Y151_SLICE_X9Y151_CMUX;
  wire [0:0] CLBLM_R_X7Y151_SLICE_X9Y151_CO5;
  wire [0:0] CLBLM_R_X7Y151_SLICE_X9Y151_CO6;
  wire [0:0] CLBLM_R_X7Y151_SLICE_X9Y151_CQ;
  wire [0:0] CLBLM_R_X7Y151_SLICE_X9Y151_C_CY;
  wire [0:0] CLBLM_R_X7Y151_SLICE_X9Y151_C_XOR;
  wire [0:0] CLBLM_R_X7Y151_SLICE_X9Y151_D;
  wire [0:0] CLBLM_R_X7Y151_SLICE_X9Y151_D1;
  wire [0:0] CLBLM_R_X7Y151_SLICE_X9Y151_D2;
  wire [0:0] CLBLM_R_X7Y151_SLICE_X9Y151_D3;
  wire [0:0] CLBLM_R_X7Y151_SLICE_X9Y151_D4;
  wire [0:0] CLBLM_R_X7Y151_SLICE_X9Y151_D5;
  wire [0:0] CLBLM_R_X7Y151_SLICE_X9Y151_D5Q;
  wire [0:0] CLBLM_R_X7Y151_SLICE_X9Y151_D6;
  wire [0:0] CLBLM_R_X7Y151_SLICE_X9Y151_DMUX;
  wire [0:0] CLBLM_R_X7Y151_SLICE_X9Y151_DO5;
  wire [0:0] CLBLM_R_X7Y151_SLICE_X9Y151_DO6;
  wire [0:0] CLBLM_R_X7Y151_SLICE_X9Y151_DQ;
  wire [0:0] CLBLM_R_X7Y151_SLICE_X9Y151_D_CY;
  wire [0:0] CLBLM_R_X7Y151_SLICE_X9Y151_D_XOR;
  wire [0:0] CLBLM_R_X7Y152_SLICE_X8Y152_A;
  wire [0:0] CLBLM_R_X7Y152_SLICE_X8Y152_A1;
  wire [0:0] CLBLM_R_X7Y152_SLICE_X8Y152_A2;
  wire [0:0] CLBLM_R_X7Y152_SLICE_X8Y152_A3;
  wire [0:0] CLBLM_R_X7Y152_SLICE_X8Y152_A4;
  wire [0:0] CLBLM_R_X7Y152_SLICE_X8Y152_A5;
  wire [0:0] CLBLM_R_X7Y152_SLICE_X8Y152_A6;
  wire [0:0] CLBLM_R_X7Y152_SLICE_X8Y152_AO5;
  wire [0:0] CLBLM_R_X7Y152_SLICE_X8Y152_AO6;
  wire [0:0] CLBLM_R_X7Y152_SLICE_X8Y152_AQ;
  wire [0:0] CLBLM_R_X7Y152_SLICE_X8Y152_A_CY;
  wire [0:0] CLBLM_R_X7Y152_SLICE_X8Y152_A_XOR;
  wire [0:0] CLBLM_R_X7Y152_SLICE_X8Y152_B;
  wire [0:0] CLBLM_R_X7Y152_SLICE_X8Y152_B1;
  wire [0:0] CLBLM_R_X7Y152_SLICE_X8Y152_B2;
  wire [0:0] CLBLM_R_X7Y152_SLICE_X8Y152_B3;
  wire [0:0] CLBLM_R_X7Y152_SLICE_X8Y152_B4;
  wire [0:0] CLBLM_R_X7Y152_SLICE_X8Y152_B5;
  wire [0:0] CLBLM_R_X7Y152_SLICE_X8Y152_B5Q;
  wire [0:0] CLBLM_R_X7Y152_SLICE_X8Y152_B6;
  wire [0:0] CLBLM_R_X7Y152_SLICE_X8Y152_BMUX;
  wire [0:0] CLBLM_R_X7Y152_SLICE_X8Y152_BO5;
  wire [0:0] CLBLM_R_X7Y152_SLICE_X8Y152_BO6;
  wire [0:0] CLBLM_R_X7Y152_SLICE_X8Y152_BQ;
  wire [0:0] CLBLM_R_X7Y152_SLICE_X8Y152_B_CY;
  wire [0:0] CLBLM_R_X7Y152_SLICE_X8Y152_B_XOR;
  wire [0:0] CLBLM_R_X7Y152_SLICE_X8Y152_C;
  wire [0:0] CLBLM_R_X7Y152_SLICE_X8Y152_C1;
  wire [0:0] CLBLM_R_X7Y152_SLICE_X8Y152_C2;
  wire [0:0] CLBLM_R_X7Y152_SLICE_X8Y152_C3;
  wire [0:0] CLBLM_R_X7Y152_SLICE_X8Y152_C4;
  wire [0:0] CLBLM_R_X7Y152_SLICE_X8Y152_C5;
  wire [0:0] CLBLM_R_X7Y152_SLICE_X8Y152_C6;
  wire [0:0] CLBLM_R_X7Y152_SLICE_X8Y152_CLK;
  wire [0:0] CLBLM_R_X7Y152_SLICE_X8Y152_CO5;
  wire [0:0] CLBLM_R_X7Y152_SLICE_X8Y152_CO6;
  wire [0:0] CLBLM_R_X7Y152_SLICE_X8Y152_CQ;
  wire [0:0] CLBLM_R_X7Y152_SLICE_X8Y152_C_CY;
  wire [0:0] CLBLM_R_X7Y152_SLICE_X8Y152_C_XOR;
  wire [0:0] CLBLM_R_X7Y152_SLICE_X8Y152_D;
  wire [0:0] CLBLM_R_X7Y152_SLICE_X8Y152_D1;
  wire [0:0] CLBLM_R_X7Y152_SLICE_X8Y152_D2;
  wire [0:0] CLBLM_R_X7Y152_SLICE_X8Y152_D3;
  wire [0:0] CLBLM_R_X7Y152_SLICE_X8Y152_D4;
  wire [0:0] CLBLM_R_X7Y152_SLICE_X8Y152_D5;
  wire [0:0] CLBLM_R_X7Y152_SLICE_X8Y152_D5Q;
  wire [0:0] CLBLM_R_X7Y152_SLICE_X8Y152_D6;
  wire [0:0] CLBLM_R_X7Y152_SLICE_X8Y152_DMUX;
  wire [0:0] CLBLM_R_X7Y152_SLICE_X8Y152_DO5;
  wire [0:0] CLBLM_R_X7Y152_SLICE_X8Y152_DO6;
  wire [0:0] CLBLM_R_X7Y152_SLICE_X8Y152_DQ;
  wire [0:0] CLBLM_R_X7Y152_SLICE_X8Y152_D_CY;
  wire [0:0] CLBLM_R_X7Y152_SLICE_X8Y152_D_XOR;
  wire [0:0] CLBLM_R_X7Y152_SLICE_X9Y152_A;
  wire [0:0] CLBLM_R_X7Y152_SLICE_X9Y152_A1;
  wire [0:0] CLBLM_R_X7Y152_SLICE_X9Y152_A2;
  wire [0:0] CLBLM_R_X7Y152_SLICE_X9Y152_A3;
  wire [0:0] CLBLM_R_X7Y152_SLICE_X9Y152_A4;
  wire [0:0] CLBLM_R_X7Y152_SLICE_X9Y152_A5;
  wire [0:0] CLBLM_R_X7Y152_SLICE_X9Y152_A6;
  wire [0:0] CLBLM_R_X7Y152_SLICE_X9Y152_AO5;
  wire [0:0] CLBLM_R_X7Y152_SLICE_X9Y152_AO6;
  wire [0:0] CLBLM_R_X7Y152_SLICE_X9Y152_AQ;
  wire [0:0] CLBLM_R_X7Y152_SLICE_X9Y152_A_CY;
  wire [0:0] CLBLM_R_X7Y152_SLICE_X9Y152_A_XOR;
  wire [0:0] CLBLM_R_X7Y152_SLICE_X9Y152_B;
  wire [0:0] CLBLM_R_X7Y152_SLICE_X9Y152_B1;
  wire [0:0] CLBLM_R_X7Y152_SLICE_X9Y152_B2;
  wire [0:0] CLBLM_R_X7Y152_SLICE_X9Y152_B3;
  wire [0:0] CLBLM_R_X7Y152_SLICE_X9Y152_B4;
  wire [0:0] CLBLM_R_X7Y152_SLICE_X9Y152_B5;
  wire [0:0] CLBLM_R_X7Y152_SLICE_X9Y152_B5Q;
  wire [0:0] CLBLM_R_X7Y152_SLICE_X9Y152_B6;
  wire [0:0] CLBLM_R_X7Y152_SLICE_X9Y152_BMUX;
  wire [0:0] CLBLM_R_X7Y152_SLICE_X9Y152_BO5;
  wire [0:0] CLBLM_R_X7Y152_SLICE_X9Y152_BO6;
  wire [0:0] CLBLM_R_X7Y152_SLICE_X9Y152_BQ;
  wire [0:0] CLBLM_R_X7Y152_SLICE_X9Y152_B_CY;
  wire [0:0] CLBLM_R_X7Y152_SLICE_X9Y152_B_XOR;
  wire [0:0] CLBLM_R_X7Y152_SLICE_X9Y152_C;
  wire [0:0] CLBLM_R_X7Y152_SLICE_X9Y152_C1;
  wire [0:0] CLBLM_R_X7Y152_SLICE_X9Y152_C2;
  wire [0:0] CLBLM_R_X7Y152_SLICE_X9Y152_C3;
  wire [0:0] CLBLM_R_X7Y152_SLICE_X9Y152_C4;
  wire [0:0] CLBLM_R_X7Y152_SLICE_X9Y152_C5;
  wire [0:0] CLBLM_R_X7Y152_SLICE_X9Y152_C5Q;
  wire [0:0] CLBLM_R_X7Y152_SLICE_X9Y152_C6;
  wire [0:0] CLBLM_R_X7Y152_SLICE_X9Y152_CLK;
  wire [0:0] CLBLM_R_X7Y152_SLICE_X9Y152_CMUX;
  wire [0:0] CLBLM_R_X7Y152_SLICE_X9Y152_CO5;
  wire [0:0] CLBLM_R_X7Y152_SLICE_X9Y152_CO6;
  wire [0:0] CLBLM_R_X7Y152_SLICE_X9Y152_CQ;
  wire [0:0] CLBLM_R_X7Y152_SLICE_X9Y152_C_CY;
  wire [0:0] CLBLM_R_X7Y152_SLICE_X9Y152_C_XOR;
  wire [0:0] CLBLM_R_X7Y152_SLICE_X9Y152_D;
  wire [0:0] CLBLM_R_X7Y152_SLICE_X9Y152_D1;
  wire [0:0] CLBLM_R_X7Y152_SLICE_X9Y152_D2;
  wire [0:0] CLBLM_R_X7Y152_SLICE_X9Y152_D3;
  wire [0:0] CLBLM_R_X7Y152_SLICE_X9Y152_D4;
  wire [0:0] CLBLM_R_X7Y152_SLICE_X9Y152_D5;
  wire [0:0] CLBLM_R_X7Y152_SLICE_X9Y152_D6;
  wire [0:0] CLBLM_R_X7Y152_SLICE_X9Y152_DMUX;
  wire [0:0] CLBLM_R_X7Y152_SLICE_X9Y152_DO5;
  wire [0:0] CLBLM_R_X7Y152_SLICE_X9Y152_DO6;
  wire [0:0] CLBLM_R_X7Y152_SLICE_X9Y152_D_CY;
  wire [0:0] CLBLM_R_X7Y152_SLICE_X9Y152_D_XOR;
  wire [0:0] CLBLM_R_X7Y153_SLICE_X8Y153_A;
  wire [0:0] CLBLM_R_X7Y153_SLICE_X8Y153_A1;
  wire [0:0] CLBLM_R_X7Y153_SLICE_X8Y153_A2;
  wire [0:0] CLBLM_R_X7Y153_SLICE_X8Y153_A3;
  wire [0:0] CLBLM_R_X7Y153_SLICE_X8Y153_A4;
  wire [0:0] CLBLM_R_X7Y153_SLICE_X8Y153_A5;
  wire [0:0] CLBLM_R_X7Y153_SLICE_X8Y153_A5Q;
  wire [0:0] CLBLM_R_X7Y153_SLICE_X8Y153_A6;
  wire [0:0] CLBLM_R_X7Y153_SLICE_X8Y153_AMUX;
  wire [0:0] CLBLM_R_X7Y153_SLICE_X8Y153_AO5;
  wire [0:0] CLBLM_R_X7Y153_SLICE_X8Y153_AO6;
  wire [0:0] CLBLM_R_X7Y153_SLICE_X8Y153_AQ;
  wire [0:0] CLBLM_R_X7Y153_SLICE_X8Y153_A_CY;
  wire [0:0] CLBLM_R_X7Y153_SLICE_X8Y153_A_XOR;
  wire [0:0] CLBLM_R_X7Y153_SLICE_X8Y153_B;
  wire [0:0] CLBLM_R_X7Y153_SLICE_X8Y153_B1;
  wire [0:0] CLBLM_R_X7Y153_SLICE_X8Y153_B2;
  wire [0:0] CLBLM_R_X7Y153_SLICE_X8Y153_B3;
  wire [0:0] CLBLM_R_X7Y153_SLICE_X8Y153_B4;
  wire [0:0] CLBLM_R_X7Y153_SLICE_X8Y153_B5;
  wire [0:0] CLBLM_R_X7Y153_SLICE_X8Y153_B6;
  wire [0:0] CLBLM_R_X7Y153_SLICE_X8Y153_BO5;
  wire [0:0] CLBLM_R_X7Y153_SLICE_X8Y153_BO6;
  wire [0:0] CLBLM_R_X7Y153_SLICE_X8Y153_BQ;
  wire [0:0] CLBLM_R_X7Y153_SLICE_X8Y153_B_CY;
  wire [0:0] CLBLM_R_X7Y153_SLICE_X8Y153_B_XOR;
  wire [0:0] CLBLM_R_X7Y153_SLICE_X8Y153_C;
  wire [0:0] CLBLM_R_X7Y153_SLICE_X8Y153_C1;
  wire [0:0] CLBLM_R_X7Y153_SLICE_X8Y153_C2;
  wire [0:0] CLBLM_R_X7Y153_SLICE_X8Y153_C3;
  wire [0:0] CLBLM_R_X7Y153_SLICE_X8Y153_C4;
  wire [0:0] CLBLM_R_X7Y153_SLICE_X8Y153_C5;
  wire [0:0] CLBLM_R_X7Y153_SLICE_X8Y153_C6;
  wire [0:0] CLBLM_R_X7Y153_SLICE_X8Y153_CLK;
  wire [0:0] CLBLM_R_X7Y153_SLICE_X8Y153_CO5;
  wire [0:0] CLBLM_R_X7Y153_SLICE_X8Y153_CO6;
  wire [0:0] CLBLM_R_X7Y153_SLICE_X8Y153_CQ;
  wire [0:0] CLBLM_R_X7Y153_SLICE_X8Y153_C_CY;
  wire [0:0] CLBLM_R_X7Y153_SLICE_X8Y153_C_XOR;
  wire [0:0] CLBLM_R_X7Y153_SLICE_X8Y153_D;
  wire [0:0] CLBLM_R_X7Y153_SLICE_X8Y153_D1;
  wire [0:0] CLBLM_R_X7Y153_SLICE_X8Y153_D2;
  wire [0:0] CLBLM_R_X7Y153_SLICE_X8Y153_D3;
  wire [0:0] CLBLM_R_X7Y153_SLICE_X8Y153_D4;
  wire [0:0] CLBLM_R_X7Y153_SLICE_X8Y153_D5;
  wire [0:0] CLBLM_R_X7Y153_SLICE_X8Y153_D6;
  wire [0:0] CLBLM_R_X7Y153_SLICE_X8Y153_DO5;
  wire [0:0] CLBLM_R_X7Y153_SLICE_X8Y153_DO6;
  wire [0:0] CLBLM_R_X7Y153_SLICE_X8Y153_DQ;
  wire [0:0] CLBLM_R_X7Y153_SLICE_X8Y153_D_CY;
  wire [0:0] CLBLM_R_X7Y153_SLICE_X8Y153_D_XOR;
  wire [0:0] CLBLM_R_X7Y153_SLICE_X9Y153_A;
  wire [0:0] CLBLM_R_X7Y153_SLICE_X9Y153_A1;
  wire [0:0] CLBLM_R_X7Y153_SLICE_X9Y153_A2;
  wire [0:0] CLBLM_R_X7Y153_SLICE_X9Y153_A3;
  wire [0:0] CLBLM_R_X7Y153_SLICE_X9Y153_A4;
  wire [0:0] CLBLM_R_X7Y153_SLICE_X9Y153_A5;
  wire [0:0] CLBLM_R_X7Y153_SLICE_X9Y153_A5Q;
  wire [0:0] CLBLM_R_X7Y153_SLICE_X9Y153_A6;
  wire [0:0] CLBLM_R_X7Y153_SLICE_X9Y153_AMUX;
  wire [0:0] CLBLM_R_X7Y153_SLICE_X9Y153_AO5;
  wire [0:0] CLBLM_R_X7Y153_SLICE_X9Y153_AO6;
  wire [0:0] CLBLM_R_X7Y153_SLICE_X9Y153_AQ;
  wire [0:0] CLBLM_R_X7Y153_SLICE_X9Y153_A_CY;
  wire [0:0] CLBLM_R_X7Y153_SLICE_X9Y153_A_XOR;
  wire [0:0] CLBLM_R_X7Y153_SLICE_X9Y153_B;
  wire [0:0] CLBLM_R_X7Y153_SLICE_X9Y153_B1;
  wire [0:0] CLBLM_R_X7Y153_SLICE_X9Y153_B2;
  wire [0:0] CLBLM_R_X7Y153_SLICE_X9Y153_B3;
  wire [0:0] CLBLM_R_X7Y153_SLICE_X9Y153_B4;
  wire [0:0] CLBLM_R_X7Y153_SLICE_X9Y153_B5;
  wire [0:0] CLBLM_R_X7Y153_SLICE_X9Y153_B6;
  wire [0:0] CLBLM_R_X7Y153_SLICE_X9Y153_BO5;
  wire [0:0] CLBLM_R_X7Y153_SLICE_X9Y153_BO6;
  wire [0:0] CLBLM_R_X7Y153_SLICE_X9Y153_BQ;
  wire [0:0] CLBLM_R_X7Y153_SLICE_X9Y153_B_CY;
  wire [0:0] CLBLM_R_X7Y153_SLICE_X9Y153_B_XOR;
  wire [0:0] CLBLM_R_X7Y153_SLICE_X9Y153_C;
  wire [0:0] CLBLM_R_X7Y153_SLICE_X9Y153_C1;
  wire [0:0] CLBLM_R_X7Y153_SLICE_X9Y153_C2;
  wire [0:0] CLBLM_R_X7Y153_SLICE_X9Y153_C3;
  wire [0:0] CLBLM_R_X7Y153_SLICE_X9Y153_C4;
  wire [0:0] CLBLM_R_X7Y153_SLICE_X9Y153_C5;
  wire [0:0] CLBLM_R_X7Y153_SLICE_X9Y153_C5Q;
  wire [0:0] CLBLM_R_X7Y153_SLICE_X9Y153_C6;
  wire [0:0] CLBLM_R_X7Y153_SLICE_X9Y153_CLK;
  wire [0:0] CLBLM_R_X7Y153_SLICE_X9Y153_CMUX;
  wire [0:0] CLBLM_R_X7Y153_SLICE_X9Y153_CO5;
  wire [0:0] CLBLM_R_X7Y153_SLICE_X9Y153_CO6;
  wire [0:0] CLBLM_R_X7Y153_SLICE_X9Y153_CQ;
  wire [0:0] CLBLM_R_X7Y153_SLICE_X9Y153_C_CY;
  wire [0:0] CLBLM_R_X7Y153_SLICE_X9Y153_C_XOR;
  wire [0:0] CLBLM_R_X7Y153_SLICE_X9Y153_D;
  wire [0:0] CLBLM_R_X7Y153_SLICE_X9Y153_D1;
  wire [0:0] CLBLM_R_X7Y153_SLICE_X9Y153_D2;
  wire [0:0] CLBLM_R_X7Y153_SLICE_X9Y153_D3;
  wire [0:0] CLBLM_R_X7Y153_SLICE_X9Y153_D4;
  wire [0:0] CLBLM_R_X7Y153_SLICE_X9Y153_D5;
  wire [0:0] CLBLM_R_X7Y153_SLICE_X9Y153_D5Q;
  wire [0:0] CLBLM_R_X7Y153_SLICE_X9Y153_D6;
  wire [0:0] CLBLM_R_X7Y153_SLICE_X9Y153_DMUX;
  wire [0:0] CLBLM_R_X7Y153_SLICE_X9Y153_DO5;
  wire [0:0] CLBLM_R_X7Y153_SLICE_X9Y153_DO6;
  wire [0:0] CLBLM_R_X7Y153_SLICE_X9Y153_DQ;
  wire [0:0] CLBLM_R_X7Y153_SLICE_X9Y153_D_CY;
  wire [0:0] CLBLM_R_X7Y153_SLICE_X9Y153_D_XOR;
  wire [0:0] CLBLM_R_X7Y154_SLICE_X8Y154_A;
  wire [0:0] CLBLM_R_X7Y154_SLICE_X8Y154_A1;
  wire [0:0] CLBLM_R_X7Y154_SLICE_X8Y154_A2;
  wire [0:0] CLBLM_R_X7Y154_SLICE_X8Y154_A3;
  wire [0:0] CLBLM_R_X7Y154_SLICE_X8Y154_A4;
  wire [0:0] CLBLM_R_X7Y154_SLICE_X8Y154_A5;
  wire [0:0] CLBLM_R_X7Y154_SLICE_X8Y154_A6;
  wire [0:0] CLBLM_R_X7Y154_SLICE_X8Y154_AO5;
  wire [0:0] CLBLM_R_X7Y154_SLICE_X8Y154_AO6;
  wire [0:0] CLBLM_R_X7Y154_SLICE_X8Y154_AQ;
  wire [0:0] CLBLM_R_X7Y154_SLICE_X8Y154_A_CY;
  wire [0:0] CLBLM_R_X7Y154_SLICE_X8Y154_A_XOR;
  wire [0:0] CLBLM_R_X7Y154_SLICE_X8Y154_B;
  wire [0:0] CLBLM_R_X7Y154_SLICE_X8Y154_B1;
  wire [0:0] CLBLM_R_X7Y154_SLICE_X8Y154_B2;
  wire [0:0] CLBLM_R_X7Y154_SLICE_X8Y154_B3;
  wire [0:0] CLBLM_R_X7Y154_SLICE_X8Y154_B4;
  wire [0:0] CLBLM_R_X7Y154_SLICE_X8Y154_B5;
  wire [0:0] CLBLM_R_X7Y154_SLICE_X8Y154_B6;
  wire [0:0] CLBLM_R_X7Y154_SLICE_X8Y154_BO5;
  wire [0:0] CLBLM_R_X7Y154_SLICE_X8Y154_BO6;
  wire [0:0] CLBLM_R_X7Y154_SLICE_X8Y154_BQ;
  wire [0:0] CLBLM_R_X7Y154_SLICE_X8Y154_B_CY;
  wire [0:0] CLBLM_R_X7Y154_SLICE_X8Y154_B_XOR;
  wire [0:0] CLBLM_R_X7Y154_SLICE_X8Y154_C;
  wire [0:0] CLBLM_R_X7Y154_SLICE_X8Y154_C1;
  wire [0:0] CLBLM_R_X7Y154_SLICE_X8Y154_C2;
  wire [0:0] CLBLM_R_X7Y154_SLICE_X8Y154_C3;
  wire [0:0] CLBLM_R_X7Y154_SLICE_X8Y154_C4;
  wire [0:0] CLBLM_R_X7Y154_SLICE_X8Y154_C5;
  wire [0:0] CLBLM_R_X7Y154_SLICE_X8Y154_C6;
  wire [0:0] CLBLM_R_X7Y154_SLICE_X8Y154_CLK;
  wire [0:0] CLBLM_R_X7Y154_SLICE_X8Y154_CMUX;
  wire [0:0] CLBLM_R_X7Y154_SLICE_X8Y154_CO5;
  wire [0:0] CLBLM_R_X7Y154_SLICE_X8Y154_CO6;
  wire [0:0] CLBLM_R_X7Y154_SLICE_X8Y154_C_CY;
  wire [0:0] CLBLM_R_X7Y154_SLICE_X8Y154_C_XOR;
  wire [0:0] CLBLM_R_X7Y154_SLICE_X8Y154_D;
  wire [0:0] CLBLM_R_X7Y154_SLICE_X8Y154_D1;
  wire [0:0] CLBLM_R_X7Y154_SLICE_X8Y154_D2;
  wire [0:0] CLBLM_R_X7Y154_SLICE_X8Y154_D3;
  wire [0:0] CLBLM_R_X7Y154_SLICE_X8Y154_D4;
  wire [0:0] CLBLM_R_X7Y154_SLICE_X8Y154_D5;
  wire [0:0] CLBLM_R_X7Y154_SLICE_X8Y154_D6;
  wire [0:0] CLBLM_R_X7Y154_SLICE_X8Y154_DO5;
  wire [0:0] CLBLM_R_X7Y154_SLICE_X8Y154_DO6;
  wire [0:0] CLBLM_R_X7Y154_SLICE_X8Y154_D_CY;
  wire [0:0] CLBLM_R_X7Y154_SLICE_X8Y154_D_XOR;
  wire [0:0] CLBLM_R_X7Y154_SLICE_X9Y154_A;
  wire [0:0] CLBLM_R_X7Y154_SLICE_X9Y154_A1;
  wire [0:0] CLBLM_R_X7Y154_SLICE_X9Y154_A2;
  wire [0:0] CLBLM_R_X7Y154_SLICE_X9Y154_A3;
  wire [0:0] CLBLM_R_X7Y154_SLICE_X9Y154_A4;
  wire [0:0] CLBLM_R_X7Y154_SLICE_X9Y154_A5;
  wire [0:0] CLBLM_R_X7Y154_SLICE_X9Y154_A6;
  wire [0:0] CLBLM_R_X7Y154_SLICE_X9Y154_AO5;
  wire [0:0] CLBLM_R_X7Y154_SLICE_X9Y154_AO6;
  wire [0:0] CLBLM_R_X7Y154_SLICE_X9Y154_AQ;
  wire [0:0] CLBLM_R_X7Y154_SLICE_X9Y154_A_CY;
  wire [0:0] CLBLM_R_X7Y154_SLICE_X9Y154_A_XOR;
  wire [0:0] CLBLM_R_X7Y154_SLICE_X9Y154_B;
  wire [0:0] CLBLM_R_X7Y154_SLICE_X9Y154_B1;
  wire [0:0] CLBLM_R_X7Y154_SLICE_X9Y154_B2;
  wire [0:0] CLBLM_R_X7Y154_SLICE_X9Y154_B3;
  wire [0:0] CLBLM_R_X7Y154_SLICE_X9Y154_B4;
  wire [0:0] CLBLM_R_X7Y154_SLICE_X9Y154_B5;
  wire [0:0] CLBLM_R_X7Y154_SLICE_X9Y154_B6;
  wire [0:0] CLBLM_R_X7Y154_SLICE_X9Y154_BO5;
  wire [0:0] CLBLM_R_X7Y154_SLICE_X9Y154_BO6;
  wire [0:0] CLBLM_R_X7Y154_SLICE_X9Y154_BQ;
  wire [0:0] CLBLM_R_X7Y154_SLICE_X9Y154_B_CY;
  wire [0:0] CLBLM_R_X7Y154_SLICE_X9Y154_B_XOR;
  wire [0:0] CLBLM_R_X7Y154_SLICE_X9Y154_C;
  wire [0:0] CLBLM_R_X7Y154_SLICE_X9Y154_C1;
  wire [0:0] CLBLM_R_X7Y154_SLICE_X9Y154_C2;
  wire [0:0] CLBLM_R_X7Y154_SLICE_X9Y154_C3;
  wire [0:0] CLBLM_R_X7Y154_SLICE_X9Y154_C4;
  wire [0:0] CLBLM_R_X7Y154_SLICE_X9Y154_C5;
  wire [0:0] CLBLM_R_X7Y154_SLICE_X9Y154_C6;
  wire [0:0] CLBLM_R_X7Y154_SLICE_X9Y154_CLK;
  wire [0:0] CLBLM_R_X7Y154_SLICE_X9Y154_CMUX;
  wire [0:0] CLBLM_R_X7Y154_SLICE_X9Y154_CO5;
  wire [0:0] CLBLM_R_X7Y154_SLICE_X9Y154_CO6;
  wire [0:0] CLBLM_R_X7Y154_SLICE_X9Y154_C_CY;
  wire [0:0] CLBLM_R_X7Y154_SLICE_X9Y154_C_XOR;
  wire [0:0] CLBLM_R_X7Y154_SLICE_X9Y154_D;
  wire [0:0] CLBLM_R_X7Y154_SLICE_X9Y154_D1;
  wire [0:0] CLBLM_R_X7Y154_SLICE_X9Y154_D2;
  wire [0:0] CLBLM_R_X7Y154_SLICE_X9Y154_D3;
  wire [0:0] CLBLM_R_X7Y154_SLICE_X9Y154_D4;
  wire [0:0] CLBLM_R_X7Y154_SLICE_X9Y154_D5;
  wire [0:0] CLBLM_R_X7Y154_SLICE_X9Y154_D6;
  wire [0:0] CLBLM_R_X7Y154_SLICE_X9Y154_DO5;
  wire [0:0] CLBLM_R_X7Y154_SLICE_X9Y154_DO6;
  wire [0:0] CLBLM_R_X7Y154_SLICE_X9Y154_D_CY;
  wire [0:0] CLBLM_R_X7Y154_SLICE_X9Y154_D_XOR;
  wire [0:0] CLBLM_R_X7Y155_SLICE_X8Y155_A;
  wire [0:0] CLBLM_R_X7Y155_SLICE_X8Y155_A1;
  wire [0:0] CLBLM_R_X7Y155_SLICE_X8Y155_A2;
  wire [0:0] CLBLM_R_X7Y155_SLICE_X8Y155_A3;
  wire [0:0] CLBLM_R_X7Y155_SLICE_X8Y155_A4;
  wire [0:0] CLBLM_R_X7Y155_SLICE_X8Y155_A5;
  wire [0:0] CLBLM_R_X7Y155_SLICE_X8Y155_A5Q;
  wire [0:0] CLBLM_R_X7Y155_SLICE_X8Y155_A6;
  wire [0:0] CLBLM_R_X7Y155_SLICE_X8Y155_AMUX;
  wire [0:0] CLBLM_R_X7Y155_SLICE_X8Y155_AO5;
  wire [0:0] CLBLM_R_X7Y155_SLICE_X8Y155_AO6;
  wire [0:0] CLBLM_R_X7Y155_SLICE_X8Y155_AQ;
  wire [0:0] CLBLM_R_X7Y155_SLICE_X8Y155_AX;
  wire [0:0] CLBLM_R_X7Y155_SLICE_X8Y155_A_CY;
  wire [0:0] CLBLM_R_X7Y155_SLICE_X8Y155_A_XOR;
  wire [0:0] CLBLM_R_X7Y155_SLICE_X8Y155_B;
  wire [0:0] CLBLM_R_X7Y155_SLICE_X8Y155_B1;
  wire [0:0] CLBLM_R_X7Y155_SLICE_X8Y155_B2;
  wire [0:0] CLBLM_R_X7Y155_SLICE_X8Y155_B3;
  wire [0:0] CLBLM_R_X7Y155_SLICE_X8Y155_B4;
  wire [0:0] CLBLM_R_X7Y155_SLICE_X8Y155_B5;
  wire [0:0] CLBLM_R_X7Y155_SLICE_X8Y155_B6;
  wire [0:0] CLBLM_R_X7Y155_SLICE_X8Y155_BMUX;
  wire [0:0] CLBLM_R_X7Y155_SLICE_X8Y155_BO5;
  wire [0:0] CLBLM_R_X7Y155_SLICE_X8Y155_BO6;
  wire [0:0] CLBLM_R_X7Y155_SLICE_X8Y155_B_CY;
  wire [0:0] CLBLM_R_X7Y155_SLICE_X8Y155_B_XOR;
  wire [0:0] CLBLM_R_X7Y155_SLICE_X8Y155_C;
  wire [0:0] CLBLM_R_X7Y155_SLICE_X8Y155_C1;
  wire [0:0] CLBLM_R_X7Y155_SLICE_X8Y155_C2;
  wire [0:0] CLBLM_R_X7Y155_SLICE_X8Y155_C3;
  wire [0:0] CLBLM_R_X7Y155_SLICE_X8Y155_C4;
  wire [0:0] CLBLM_R_X7Y155_SLICE_X8Y155_C5;
  wire [0:0] CLBLM_R_X7Y155_SLICE_X8Y155_C6;
  wire [0:0] CLBLM_R_X7Y155_SLICE_X8Y155_CLK;
  wire [0:0] CLBLM_R_X7Y155_SLICE_X8Y155_CO5;
  wire [0:0] CLBLM_R_X7Y155_SLICE_X8Y155_CO6;
  wire [0:0] CLBLM_R_X7Y155_SLICE_X8Y155_C_CY;
  wire [0:0] CLBLM_R_X7Y155_SLICE_X8Y155_C_XOR;
  wire [0:0] CLBLM_R_X7Y155_SLICE_X8Y155_D;
  wire [0:0] CLBLM_R_X7Y155_SLICE_X8Y155_D1;
  wire [0:0] CLBLM_R_X7Y155_SLICE_X8Y155_D2;
  wire [0:0] CLBLM_R_X7Y155_SLICE_X8Y155_D3;
  wire [0:0] CLBLM_R_X7Y155_SLICE_X8Y155_D4;
  wire [0:0] CLBLM_R_X7Y155_SLICE_X8Y155_D5;
  wire [0:0] CLBLM_R_X7Y155_SLICE_X8Y155_D6;
  wire [0:0] CLBLM_R_X7Y155_SLICE_X8Y155_DO5;
  wire [0:0] CLBLM_R_X7Y155_SLICE_X8Y155_DO6;
  wire [0:0] CLBLM_R_X7Y155_SLICE_X8Y155_D_CY;
  wire [0:0] CLBLM_R_X7Y155_SLICE_X8Y155_D_XOR;
  wire [0:0] CLBLM_R_X7Y155_SLICE_X9Y155_A;
  wire [0:0] CLBLM_R_X7Y155_SLICE_X9Y155_A1;
  wire [0:0] CLBLM_R_X7Y155_SLICE_X9Y155_A2;
  wire [0:0] CLBLM_R_X7Y155_SLICE_X9Y155_A3;
  wire [0:0] CLBLM_R_X7Y155_SLICE_X9Y155_A4;
  wire [0:0] CLBLM_R_X7Y155_SLICE_X9Y155_A5;
  wire [0:0] CLBLM_R_X7Y155_SLICE_X9Y155_A6;
  wire [0:0] CLBLM_R_X7Y155_SLICE_X9Y155_AO5;
  wire [0:0] CLBLM_R_X7Y155_SLICE_X9Y155_AO6;
  wire [0:0] CLBLM_R_X7Y155_SLICE_X9Y155_A_CY;
  wire [0:0] CLBLM_R_X7Y155_SLICE_X9Y155_A_XOR;
  wire [0:0] CLBLM_R_X7Y155_SLICE_X9Y155_B;
  wire [0:0] CLBLM_R_X7Y155_SLICE_X9Y155_B1;
  wire [0:0] CLBLM_R_X7Y155_SLICE_X9Y155_B2;
  wire [0:0] CLBLM_R_X7Y155_SLICE_X9Y155_B3;
  wire [0:0] CLBLM_R_X7Y155_SLICE_X9Y155_B4;
  wire [0:0] CLBLM_R_X7Y155_SLICE_X9Y155_B5;
  wire [0:0] CLBLM_R_X7Y155_SLICE_X9Y155_B6;
  wire [0:0] CLBLM_R_X7Y155_SLICE_X9Y155_BO5;
  wire [0:0] CLBLM_R_X7Y155_SLICE_X9Y155_BO6;
  wire [0:0] CLBLM_R_X7Y155_SLICE_X9Y155_B_CY;
  wire [0:0] CLBLM_R_X7Y155_SLICE_X9Y155_B_XOR;
  wire [0:0] CLBLM_R_X7Y155_SLICE_X9Y155_C;
  wire [0:0] CLBLM_R_X7Y155_SLICE_X9Y155_C1;
  wire [0:0] CLBLM_R_X7Y155_SLICE_X9Y155_C2;
  wire [0:0] CLBLM_R_X7Y155_SLICE_X9Y155_C3;
  wire [0:0] CLBLM_R_X7Y155_SLICE_X9Y155_C4;
  wire [0:0] CLBLM_R_X7Y155_SLICE_X9Y155_C5;
  wire [0:0] CLBLM_R_X7Y155_SLICE_X9Y155_C6;
  wire [0:0] CLBLM_R_X7Y155_SLICE_X9Y155_CO5;
  wire [0:0] CLBLM_R_X7Y155_SLICE_X9Y155_CO6;
  wire [0:0] CLBLM_R_X7Y155_SLICE_X9Y155_C_CY;
  wire [0:0] CLBLM_R_X7Y155_SLICE_X9Y155_C_XOR;
  wire [0:0] CLBLM_R_X7Y155_SLICE_X9Y155_D;
  wire [0:0] CLBLM_R_X7Y155_SLICE_X9Y155_D1;
  wire [0:0] CLBLM_R_X7Y155_SLICE_X9Y155_D2;
  wire [0:0] CLBLM_R_X7Y155_SLICE_X9Y155_D3;
  wire [0:0] CLBLM_R_X7Y155_SLICE_X9Y155_D4;
  wire [0:0] CLBLM_R_X7Y155_SLICE_X9Y155_D5;
  wire [0:0] CLBLM_R_X7Y155_SLICE_X9Y155_D6;
  wire [0:0] CLBLM_R_X7Y155_SLICE_X9Y155_DO5;
  wire [0:0] CLBLM_R_X7Y155_SLICE_X9Y155_DO6;
  wire [0:0] CLBLM_R_X7Y155_SLICE_X9Y155_D_CY;
  wire [0:0] CLBLM_R_X7Y155_SLICE_X9Y155_D_XOR;
  wire [0:0] CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_CE0;
  wire [0:0] CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_CE1;
  wire [0:0] CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_I0;
  wire [0:0] CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_I1;
  wire [0:0] CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_IGNORE0;
  wire [0:0] CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_IGNORE1;
  wire [0:0] CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_O;
  wire [0:0] CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_S0;
  wire [0:0] CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_S1;
  wire [0:0] CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_CE;
  wire [0:0] CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_I;
  wire [0:0] CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  wire [0:0] CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_CE;
  wire [0:0] CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_I;
  wire [0:0] CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O;
  wire [0:0] LIOB33_SING_X0Y100_IOB_X0Y100_O;
  wire [0:0] LIOB33_SING_X0Y149_IOB_X0Y149_O;
  wire [0:0] LIOB33_SING_X0Y150_IOB_X0Y150_O;
  wire [0:0] LIOB33_SING_X0Y199_IOB_X0Y199_O;
  wire [0:0] LIOB33_SING_X0Y50_IOB_X0Y50_I;
  wire [0:0] LIOB33_X0Y101_IOB_X0Y101_O;
  wire [0:0] LIOB33_X0Y101_IOB_X0Y102_O;
  wire [0:0] LIOB33_X0Y103_IOB_X0Y103_O;
  wire [0:0] LIOB33_X0Y103_IOB_X0Y104_O;
  wire [0:0] LIOB33_X0Y105_IOB_X0Y105_O;
  wire [0:0] LIOB33_X0Y105_IOB_X0Y106_O;
  wire [0:0] LIOB33_X0Y107_IOB_X0Y107_O;
  wire [0:0] LIOB33_X0Y107_IOB_X0Y108_O;
  wire [0:0] LIOB33_X0Y109_IOB_X0Y109_O;
  wire [0:0] LIOB33_X0Y109_IOB_X0Y110_O;
  wire [0:0] LIOB33_X0Y111_IOB_X0Y111_O;
  wire [0:0] LIOB33_X0Y111_IOB_X0Y112_O;
  wire [0:0] LIOB33_X0Y113_IOB_X0Y113_O;
  wire [0:0] LIOB33_X0Y113_IOB_X0Y114_O;
  wire [0:0] LIOB33_X0Y115_IOB_X0Y115_O;
  wire [0:0] LIOB33_X0Y115_IOB_X0Y116_O;
  wire [0:0] LIOB33_X0Y117_IOB_X0Y117_O;
  wire [0:0] LIOB33_X0Y117_IOB_X0Y118_O;
  wire [0:0] LIOB33_X0Y119_IOB_X0Y119_O;
  wire [0:0] LIOB33_X0Y119_IOB_X0Y120_O;
  wire [0:0] LIOB33_X0Y121_IOB_X0Y121_O;
  wire [0:0] LIOB33_X0Y121_IOB_X0Y122_O;
  wire [0:0] LIOB33_X0Y123_IOB_X0Y123_O;
  wire [0:0] LIOB33_X0Y123_IOB_X0Y124_O;
  wire [0:0] LIOB33_X0Y125_IOB_X0Y125_O;
  wire [0:0] LIOB33_X0Y125_IOB_X0Y126_O;
  wire [0:0] LIOB33_X0Y127_IOB_X0Y127_O;
  wire [0:0] LIOB33_X0Y127_IOB_X0Y128_O;
  wire [0:0] LIOB33_X0Y129_IOB_X0Y129_O;
  wire [0:0] LIOB33_X0Y129_IOB_X0Y130_O;
  wire [0:0] LIOB33_X0Y131_IOB_X0Y131_O;
  wire [0:0] LIOB33_X0Y131_IOB_X0Y132_O;
  wire [0:0] LIOB33_X0Y133_IOB_X0Y133_O;
  wire [0:0] LIOB33_X0Y133_IOB_X0Y134_O;
  wire [0:0] LIOB33_X0Y135_IOB_X0Y135_O;
  wire [0:0] LIOB33_X0Y135_IOB_X0Y136_O;
  wire [0:0] LIOB33_X0Y137_IOB_X0Y137_O;
  wire [0:0] LIOB33_X0Y137_IOB_X0Y138_O;
  wire [0:0] LIOB33_X0Y139_IOB_X0Y139_O;
  wire [0:0] LIOB33_X0Y139_IOB_X0Y140_O;
  wire [0:0] LIOB33_X0Y141_IOB_X0Y141_O;
  wire [0:0] LIOB33_X0Y141_IOB_X0Y142_O;
  wire [0:0] LIOB33_X0Y143_IOB_X0Y143_O;
  wire [0:0] LIOB33_X0Y145_IOB_X0Y145_O;
  wire [0:0] LIOB33_X0Y145_IOB_X0Y146_O;
  wire [0:0] LIOB33_X0Y147_IOB_X0Y147_O;
  wire [0:0] LIOB33_X0Y147_IOB_X0Y148_O;
  wire [0:0] LIOB33_X0Y151_IOB_X0Y151_O;
  wire [0:0] LIOB33_X0Y151_IOB_X0Y152_O;
  wire [0:0] LIOB33_X0Y153_IOB_X0Y153_O;
  wire [0:0] LIOB33_X0Y153_IOB_X0Y154_O;
  wire [0:0] LIOB33_X0Y155_IOB_X0Y155_O;
  wire [0:0] LIOB33_X0Y155_IOB_X0Y156_O;
  wire [0:0] LIOB33_X0Y157_IOB_X0Y157_O;
  wire [0:0] LIOB33_X0Y157_IOB_X0Y158_O;
  wire [0:0] LIOB33_X0Y159_IOB_X0Y159_O;
  wire [0:0] LIOB33_X0Y159_IOB_X0Y160_O;
  wire [0:0] LIOB33_X0Y161_IOB_X0Y161_O;
  wire [0:0] LIOB33_X0Y161_IOB_X0Y162_O;
  wire [0:0] LIOB33_X0Y163_IOB_X0Y163_O;
  wire [0:0] LIOB33_X0Y163_IOB_X0Y164_O;
  wire [0:0] LIOB33_X0Y165_IOB_X0Y165_O;
  wire [0:0] LIOB33_X0Y165_IOB_X0Y166_O;
  wire [0:0] LIOB33_X0Y167_IOB_X0Y167_O;
  wire [0:0] LIOB33_X0Y167_IOB_X0Y168_O;
  wire [0:0] LIOB33_X0Y169_IOB_X0Y169_O;
  wire [0:0] LIOB33_X0Y169_IOB_X0Y170_O;
  wire [0:0] LIOB33_X0Y171_IOB_X0Y171_O;
  wire [0:0] LIOB33_X0Y171_IOB_X0Y172_O;
  wire [0:0] LIOB33_X0Y173_IOB_X0Y173_O;
  wire [0:0] LIOB33_X0Y173_IOB_X0Y174_O;
  wire [0:0] LIOB33_X0Y175_IOB_X0Y175_O;
  wire [0:0] LIOB33_X0Y175_IOB_X0Y176_O;
  wire [0:0] LIOB33_X0Y177_IOB_X0Y177_O;
  wire [0:0] LIOB33_X0Y177_IOB_X0Y178_O;
  wire [0:0] LIOB33_X0Y179_IOB_X0Y179_O;
  wire [0:0] LIOB33_X0Y179_IOB_X0Y180_O;
  wire [0:0] LIOB33_X0Y181_IOB_X0Y181_O;
  wire [0:0] LIOB33_X0Y181_IOB_X0Y182_O;
  wire [0:0] LIOB33_X0Y183_IOB_X0Y183_O;
  wire [0:0] LIOB33_X0Y183_IOB_X0Y184_O;
  wire [0:0] LIOB33_X0Y185_IOB_X0Y185_O;
  wire [0:0] LIOB33_X0Y185_IOB_X0Y186_O;
  wire [0:0] LIOB33_X0Y187_IOB_X0Y187_O;
  wire [0:0] LIOB33_X0Y187_IOB_X0Y188_O;
  wire [0:0] LIOB33_X0Y189_IOB_X0Y189_O;
  wire [0:0] LIOB33_X0Y189_IOB_X0Y190_O;
  wire [0:0] LIOB33_X0Y191_IOB_X0Y191_O;
  wire [0:0] LIOB33_X0Y191_IOB_X0Y192_O;
  wire [0:0] LIOB33_X0Y193_IOB_X0Y193_O;
  wire [0:0] LIOB33_X0Y193_IOB_X0Y194_O;
  wire [0:0] LIOB33_X0Y195_IOB_X0Y195_O;
  wire [0:0] LIOB33_X0Y195_IOB_X0Y196_O;
  wire [0:0] LIOB33_X0Y197_IOB_X0Y197_O;
  wire [0:0] LIOB33_X0Y197_IOB_X0Y198_O;
  wire [0:0] LIOB33_X0Y51_IOB_X0Y51_I;
  wire [0:0] LIOB33_X0Y51_IOB_X0Y52_I;
  wire [0:0] LIOB33_X0Y53_IOB_X0Y53_I;
  wire [0:0] LIOB33_X0Y53_IOB_X0Y54_I;
  wire [0:0] LIOB33_X0Y55_IOB_X0Y55_I;
  wire [0:0] LIOB33_X0Y55_IOB_X0Y56_I;
  wire [0:0] LIOB33_X0Y57_IOB_X0Y57_I;
  wire [0:0] LIOB33_X0Y57_IOB_X0Y58_I;
  wire [0:0] LIOB33_X0Y59_IOB_X0Y59_I;
  wire [0:0] LIOB33_X0Y59_IOB_X0Y60_I;
  wire [0:0] LIOB33_X0Y61_IOB_X0Y61_I;
  wire [0:0] LIOB33_X0Y61_IOB_X0Y62_I;
  wire [0:0] LIOB33_X0Y63_IOB_X0Y63_I;
  wire [0:0] LIOB33_X0Y63_IOB_X0Y64_O;
  wire [0:0] LIOB33_X0Y65_IOB_X0Y65_O;
  wire [0:0] LIOB33_X0Y65_IOB_X0Y66_O;
  wire [0:0] LIOB33_X0Y77_IOB_X0Y78_I;
  wire [0:0] LIOI3_SING_X0Y100_OLOGIC_X0Y100_D1;
  wire [0:0] LIOI3_SING_X0Y100_OLOGIC_X0Y100_OQ;
  wire [0:0] LIOI3_SING_X0Y100_OLOGIC_X0Y100_T1;
  wire [0:0] LIOI3_SING_X0Y100_OLOGIC_X0Y100_TQ;
  wire [0:0] LIOI3_SING_X0Y149_OLOGIC_X0Y149_D1;
  wire [0:0] LIOI3_SING_X0Y149_OLOGIC_X0Y149_OQ;
  wire [0:0] LIOI3_SING_X0Y149_OLOGIC_X0Y149_T1;
  wire [0:0] LIOI3_SING_X0Y149_OLOGIC_X0Y149_TQ;
  wire [0:0] LIOI3_SING_X0Y150_OLOGIC_X0Y150_D1;
  wire [0:0] LIOI3_SING_X0Y150_OLOGIC_X0Y150_OQ;
  wire [0:0] LIOI3_SING_X0Y150_OLOGIC_X0Y150_T1;
  wire [0:0] LIOI3_SING_X0Y150_OLOGIC_X0Y150_TQ;
  wire [0:0] LIOI3_SING_X0Y199_OLOGIC_X0Y199_D1;
  wire [0:0] LIOI3_SING_X0Y199_OLOGIC_X0Y199_OQ;
  wire [0:0] LIOI3_SING_X0Y199_OLOGIC_X0Y199_T1;
  wire [0:0] LIOI3_SING_X0Y199_OLOGIC_X0Y199_TQ;
  wire [0:0] LIOI3_SING_X0Y50_ILOGIC_X0Y50_D;
  wire [0:0] LIOI3_SING_X0Y50_ILOGIC_X0Y50_O;
  wire [0:0] LIOI3_TBYTESRC_X0Y107_OLOGIC_X0Y107_D1;
  wire [0:0] LIOI3_TBYTESRC_X0Y107_OLOGIC_X0Y107_OQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y107_OLOGIC_X0Y107_T1;
  wire [0:0] LIOI3_TBYTESRC_X0Y107_OLOGIC_X0Y107_TQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y107_OLOGIC_X0Y108_D1;
  wire [0:0] LIOI3_TBYTESRC_X0Y107_OLOGIC_X0Y108_OQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y107_OLOGIC_X0Y108_T1;
  wire [0:0] LIOI3_TBYTESRC_X0Y107_OLOGIC_X0Y108_TQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y119_OLOGIC_X0Y119_D1;
  wire [0:0] LIOI3_TBYTESRC_X0Y119_OLOGIC_X0Y119_OQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y119_OLOGIC_X0Y119_T1;
  wire [0:0] LIOI3_TBYTESRC_X0Y119_OLOGIC_X0Y119_TQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y119_OLOGIC_X0Y120_D1;
  wire [0:0] LIOI3_TBYTESRC_X0Y119_OLOGIC_X0Y120_OQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y119_OLOGIC_X0Y120_T1;
  wire [0:0] LIOI3_TBYTESRC_X0Y119_OLOGIC_X0Y120_TQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y131_OLOGIC_X0Y131_D1;
  wire [0:0] LIOI3_TBYTESRC_X0Y131_OLOGIC_X0Y131_OQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y131_OLOGIC_X0Y131_T1;
  wire [0:0] LIOI3_TBYTESRC_X0Y131_OLOGIC_X0Y131_TQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y131_OLOGIC_X0Y132_D1;
  wire [0:0] LIOI3_TBYTESRC_X0Y131_OLOGIC_X0Y132_OQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y131_OLOGIC_X0Y132_T1;
  wire [0:0] LIOI3_TBYTESRC_X0Y131_OLOGIC_X0Y132_TQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y143_OLOGIC_X0Y143_D1;
  wire [0:0] LIOI3_TBYTESRC_X0Y143_OLOGIC_X0Y143_OQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y143_OLOGIC_X0Y143_T1;
  wire [0:0] LIOI3_TBYTESRC_X0Y143_OLOGIC_X0Y143_TQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y143_OLOGIC_X0Y144_D1;
  wire [0:0] LIOI3_TBYTESRC_X0Y143_OLOGIC_X0Y144_OQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y143_OLOGIC_X0Y144_T1;
  wire [0:0] LIOI3_TBYTESRC_X0Y143_OLOGIC_X0Y144_TQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y157_OLOGIC_X0Y157_D1;
  wire [0:0] LIOI3_TBYTESRC_X0Y157_OLOGIC_X0Y157_OQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y157_OLOGIC_X0Y157_T1;
  wire [0:0] LIOI3_TBYTESRC_X0Y157_OLOGIC_X0Y157_TQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y157_OLOGIC_X0Y158_D1;
  wire [0:0] LIOI3_TBYTESRC_X0Y157_OLOGIC_X0Y158_OQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y157_OLOGIC_X0Y158_T1;
  wire [0:0] LIOI3_TBYTESRC_X0Y157_OLOGIC_X0Y158_TQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y169_OLOGIC_X0Y169_D1;
  wire [0:0] LIOI3_TBYTESRC_X0Y169_OLOGIC_X0Y169_OQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y169_OLOGIC_X0Y169_T1;
  wire [0:0] LIOI3_TBYTESRC_X0Y169_OLOGIC_X0Y169_TQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y169_OLOGIC_X0Y170_D1;
  wire [0:0] LIOI3_TBYTESRC_X0Y169_OLOGIC_X0Y170_OQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y169_OLOGIC_X0Y170_T1;
  wire [0:0] LIOI3_TBYTESRC_X0Y169_OLOGIC_X0Y170_TQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y181_OLOGIC_X0Y181_D1;
  wire [0:0] LIOI3_TBYTESRC_X0Y181_OLOGIC_X0Y181_OQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y181_OLOGIC_X0Y181_T1;
  wire [0:0] LIOI3_TBYTESRC_X0Y181_OLOGIC_X0Y181_TQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y181_OLOGIC_X0Y182_D1;
  wire [0:0] LIOI3_TBYTESRC_X0Y181_OLOGIC_X0Y182_OQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y181_OLOGIC_X0Y182_T1;
  wire [0:0] LIOI3_TBYTESRC_X0Y181_OLOGIC_X0Y182_TQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y193_OLOGIC_X0Y193_D1;
  wire [0:0] LIOI3_TBYTESRC_X0Y193_OLOGIC_X0Y193_OQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y193_OLOGIC_X0Y193_T1;
  wire [0:0] LIOI3_TBYTESRC_X0Y193_OLOGIC_X0Y193_TQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y193_OLOGIC_X0Y194_D1;
  wire [0:0] LIOI3_TBYTESRC_X0Y193_OLOGIC_X0Y194_OQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y193_OLOGIC_X0Y194_T1;
  wire [0:0] LIOI3_TBYTESRC_X0Y193_OLOGIC_X0Y194_TQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y57_ILOGIC_X0Y57_D;
  wire [0:0] LIOI3_TBYTESRC_X0Y57_ILOGIC_X0Y57_O;
  wire [0:0] LIOI3_TBYTESRC_X0Y57_ILOGIC_X0Y58_D;
  wire [0:0] LIOI3_TBYTESRC_X0Y57_ILOGIC_X0Y58_O;
  wire [0:0] LIOI3_TBYTETERM_X0Y113_OLOGIC_X0Y113_D1;
  wire [0:0] LIOI3_TBYTETERM_X0Y113_OLOGIC_X0Y113_OQ;
  wire [0:0] LIOI3_TBYTETERM_X0Y113_OLOGIC_X0Y113_T1;
  wire [0:0] LIOI3_TBYTETERM_X0Y113_OLOGIC_X0Y113_TQ;
  wire [0:0] LIOI3_TBYTETERM_X0Y113_OLOGIC_X0Y114_D1;
  wire [0:0] LIOI3_TBYTETERM_X0Y113_OLOGIC_X0Y114_OQ;
  wire [0:0] LIOI3_TBYTETERM_X0Y113_OLOGIC_X0Y114_T1;
  wire [0:0] LIOI3_TBYTETERM_X0Y113_OLOGIC_X0Y114_TQ;
  wire [0:0] LIOI3_TBYTETERM_X0Y137_OLOGIC_X0Y137_D1;
  wire [0:0] LIOI3_TBYTETERM_X0Y137_OLOGIC_X0Y137_OQ;
  wire [0:0] LIOI3_TBYTETERM_X0Y137_OLOGIC_X0Y137_T1;
  wire [0:0] LIOI3_TBYTETERM_X0Y137_OLOGIC_X0Y137_TQ;
  wire [0:0] LIOI3_TBYTETERM_X0Y137_OLOGIC_X0Y138_D1;
  wire [0:0] LIOI3_TBYTETERM_X0Y137_OLOGIC_X0Y138_OQ;
  wire [0:0] LIOI3_TBYTETERM_X0Y137_OLOGIC_X0Y138_T1;
  wire [0:0] LIOI3_TBYTETERM_X0Y137_OLOGIC_X0Y138_TQ;
  wire [0:0] LIOI3_TBYTETERM_X0Y163_OLOGIC_X0Y163_D1;
  wire [0:0] LIOI3_TBYTETERM_X0Y163_OLOGIC_X0Y163_OQ;
  wire [0:0] LIOI3_TBYTETERM_X0Y163_OLOGIC_X0Y163_T1;
  wire [0:0] LIOI3_TBYTETERM_X0Y163_OLOGIC_X0Y163_TQ;
  wire [0:0] LIOI3_TBYTETERM_X0Y163_OLOGIC_X0Y164_D1;
  wire [0:0] LIOI3_TBYTETERM_X0Y163_OLOGIC_X0Y164_OQ;
  wire [0:0] LIOI3_TBYTETERM_X0Y163_OLOGIC_X0Y164_T1;
  wire [0:0] LIOI3_TBYTETERM_X0Y163_OLOGIC_X0Y164_TQ;
  wire [0:0] LIOI3_TBYTETERM_X0Y187_OLOGIC_X0Y187_D1;
  wire [0:0] LIOI3_TBYTETERM_X0Y187_OLOGIC_X0Y187_OQ;
  wire [0:0] LIOI3_TBYTETERM_X0Y187_OLOGIC_X0Y187_T1;
  wire [0:0] LIOI3_TBYTETERM_X0Y187_OLOGIC_X0Y187_TQ;
  wire [0:0] LIOI3_TBYTETERM_X0Y187_OLOGIC_X0Y188_D1;
  wire [0:0] LIOI3_TBYTETERM_X0Y187_OLOGIC_X0Y188_OQ;
  wire [0:0] LIOI3_TBYTETERM_X0Y187_OLOGIC_X0Y188_T1;
  wire [0:0] LIOI3_TBYTETERM_X0Y187_OLOGIC_X0Y188_TQ;
  wire [0:0] LIOI3_TBYTETERM_X0Y63_ILOGIC_X0Y63_D;
  wire [0:0] LIOI3_TBYTETERM_X0Y63_ILOGIC_X0Y63_O;
  wire [0:0] LIOI3_TBYTETERM_X0Y63_OLOGIC_X0Y64_D1;
  wire [0:0] LIOI3_TBYTETERM_X0Y63_OLOGIC_X0Y64_OQ;
  wire [0:0] LIOI3_TBYTETERM_X0Y63_OLOGIC_X0Y64_T1;
  wire [0:0] LIOI3_TBYTETERM_X0Y63_OLOGIC_X0Y64_TQ;
  wire [0:0] LIOI3_X0Y101_OLOGIC_X0Y101_D1;
  wire [0:0] LIOI3_X0Y101_OLOGIC_X0Y101_OQ;
  wire [0:0] LIOI3_X0Y101_OLOGIC_X0Y101_T1;
  wire [0:0] LIOI3_X0Y101_OLOGIC_X0Y101_TQ;
  wire [0:0] LIOI3_X0Y101_OLOGIC_X0Y102_D1;
  wire [0:0] LIOI3_X0Y101_OLOGIC_X0Y102_OQ;
  wire [0:0] LIOI3_X0Y101_OLOGIC_X0Y102_T1;
  wire [0:0] LIOI3_X0Y101_OLOGIC_X0Y102_TQ;
  wire [0:0] LIOI3_X0Y103_OLOGIC_X0Y103_D1;
  wire [0:0] LIOI3_X0Y103_OLOGIC_X0Y103_OQ;
  wire [0:0] LIOI3_X0Y103_OLOGIC_X0Y103_T1;
  wire [0:0] LIOI3_X0Y103_OLOGIC_X0Y103_TQ;
  wire [0:0] LIOI3_X0Y103_OLOGIC_X0Y104_D1;
  wire [0:0] LIOI3_X0Y103_OLOGIC_X0Y104_OQ;
  wire [0:0] LIOI3_X0Y103_OLOGIC_X0Y104_T1;
  wire [0:0] LIOI3_X0Y103_OLOGIC_X0Y104_TQ;
  wire [0:0] LIOI3_X0Y105_OLOGIC_X0Y105_D1;
  wire [0:0] LIOI3_X0Y105_OLOGIC_X0Y105_OQ;
  wire [0:0] LIOI3_X0Y105_OLOGIC_X0Y105_T1;
  wire [0:0] LIOI3_X0Y105_OLOGIC_X0Y105_TQ;
  wire [0:0] LIOI3_X0Y105_OLOGIC_X0Y106_D1;
  wire [0:0] LIOI3_X0Y105_OLOGIC_X0Y106_OQ;
  wire [0:0] LIOI3_X0Y105_OLOGIC_X0Y106_T1;
  wire [0:0] LIOI3_X0Y105_OLOGIC_X0Y106_TQ;
  wire [0:0] LIOI3_X0Y109_OLOGIC_X0Y109_D1;
  wire [0:0] LIOI3_X0Y109_OLOGIC_X0Y109_OQ;
  wire [0:0] LIOI3_X0Y109_OLOGIC_X0Y109_T1;
  wire [0:0] LIOI3_X0Y109_OLOGIC_X0Y109_TQ;
  wire [0:0] LIOI3_X0Y109_OLOGIC_X0Y110_D1;
  wire [0:0] LIOI3_X0Y109_OLOGIC_X0Y110_OQ;
  wire [0:0] LIOI3_X0Y109_OLOGIC_X0Y110_T1;
  wire [0:0] LIOI3_X0Y109_OLOGIC_X0Y110_TQ;
  wire [0:0] LIOI3_X0Y111_OLOGIC_X0Y111_D1;
  wire [0:0] LIOI3_X0Y111_OLOGIC_X0Y111_OQ;
  wire [0:0] LIOI3_X0Y111_OLOGIC_X0Y111_T1;
  wire [0:0] LIOI3_X0Y111_OLOGIC_X0Y111_TQ;
  wire [0:0] LIOI3_X0Y111_OLOGIC_X0Y112_D1;
  wire [0:0] LIOI3_X0Y111_OLOGIC_X0Y112_OQ;
  wire [0:0] LIOI3_X0Y111_OLOGIC_X0Y112_T1;
  wire [0:0] LIOI3_X0Y111_OLOGIC_X0Y112_TQ;
  wire [0:0] LIOI3_X0Y115_OLOGIC_X0Y115_D1;
  wire [0:0] LIOI3_X0Y115_OLOGIC_X0Y115_OQ;
  wire [0:0] LIOI3_X0Y115_OLOGIC_X0Y115_T1;
  wire [0:0] LIOI3_X0Y115_OLOGIC_X0Y115_TQ;
  wire [0:0] LIOI3_X0Y115_OLOGIC_X0Y116_D1;
  wire [0:0] LIOI3_X0Y115_OLOGIC_X0Y116_OQ;
  wire [0:0] LIOI3_X0Y115_OLOGIC_X0Y116_T1;
  wire [0:0] LIOI3_X0Y115_OLOGIC_X0Y116_TQ;
  wire [0:0] LIOI3_X0Y117_OLOGIC_X0Y117_D1;
  wire [0:0] LIOI3_X0Y117_OLOGIC_X0Y117_OQ;
  wire [0:0] LIOI3_X0Y117_OLOGIC_X0Y117_T1;
  wire [0:0] LIOI3_X0Y117_OLOGIC_X0Y117_TQ;
  wire [0:0] LIOI3_X0Y117_OLOGIC_X0Y118_D1;
  wire [0:0] LIOI3_X0Y117_OLOGIC_X0Y118_OQ;
  wire [0:0] LIOI3_X0Y117_OLOGIC_X0Y118_T1;
  wire [0:0] LIOI3_X0Y117_OLOGIC_X0Y118_TQ;
  wire [0:0] LIOI3_X0Y121_OLOGIC_X0Y121_D1;
  wire [0:0] LIOI3_X0Y121_OLOGIC_X0Y121_OQ;
  wire [0:0] LIOI3_X0Y121_OLOGIC_X0Y121_T1;
  wire [0:0] LIOI3_X0Y121_OLOGIC_X0Y121_TQ;
  wire [0:0] LIOI3_X0Y121_OLOGIC_X0Y122_D1;
  wire [0:0] LIOI3_X0Y121_OLOGIC_X0Y122_OQ;
  wire [0:0] LIOI3_X0Y121_OLOGIC_X0Y122_T1;
  wire [0:0] LIOI3_X0Y121_OLOGIC_X0Y122_TQ;
  wire [0:0] LIOI3_X0Y123_OLOGIC_X0Y123_D1;
  wire [0:0] LIOI3_X0Y123_OLOGIC_X0Y123_OQ;
  wire [0:0] LIOI3_X0Y123_OLOGIC_X0Y123_T1;
  wire [0:0] LIOI3_X0Y123_OLOGIC_X0Y123_TQ;
  wire [0:0] LIOI3_X0Y123_OLOGIC_X0Y124_D1;
  wire [0:0] LIOI3_X0Y123_OLOGIC_X0Y124_OQ;
  wire [0:0] LIOI3_X0Y123_OLOGIC_X0Y124_T1;
  wire [0:0] LIOI3_X0Y123_OLOGIC_X0Y124_TQ;
  wire [0:0] LIOI3_X0Y125_OLOGIC_X0Y125_D1;
  wire [0:0] LIOI3_X0Y125_OLOGIC_X0Y125_OQ;
  wire [0:0] LIOI3_X0Y125_OLOGIC_X0Y125_T1;
  wire [0:0] LIOI3_X0Y125_OLOGIC_X0Y125_TQ;
  wire [0:0] LIOI3_X0Y125_OLOGIC_X0Y126_D1;
  wire [0:0] LIOI3_X0Y125_OLOGIC_X0Y126_OQ;
  wire [0:0] LIOI3_X0Y125_OLOGIC_X0Y126_T1;
  wire [0:0] LIOI3_X0Y125_OLOGIC_X0Y126_TQ;
  wire [0:0] LIOI3_X0Y127_OLOGIC_X0Y127_D1;
  wire [0:0] LIOI3_X0Y127_OLOGIC_X0Y127_OQ;
  wire [0:0] LIOI3_X0Y127_OLOGIC_X0Y127_T1;
  wire [0:0] LIOI3_X0Y127_OLOGIC_X0Y127_TQ;
  wire [0:0] LIOI3_X0Y127_OLOGIC_X0Y128_D1;
  wire [0:0] LIOI3_X0Y127_OLOGIC_X0Y128_OQ;
  wire [0:0] LIOI3_X0Y127_OLOGIC_X0Y128_T1;
  wire [0:0] LIOI3_X0Y127_OLOGIC_X0Y128_TQ;
  wire [0:0] LIOI3_X0Y129_OLOGIC_X0Y129_D1;
  wire [0:0] LIOI3_X0Y129_OLOGIC_X0Y129_OQ;
  wire [0:0] LIOI3_X0Y129_OLOGIC_X0Y129_T1;
  wire [0:0] LIOI3_X0Y129_OLOGIC_X0Y129_TQ;
  wire [0:0] LIOI3_X0Y129_OLOGIC_X0Y130_D1;
  wire [0:0] LIOI3_X0Y129_OLOGIC_X0Y130_OQ;
  wire [0:0] LIOI3_X0Y129_OLOGIC_X0Y130_T1;
  wire [0:0] LIOI3_X0Y129_OLOGIC_X0Y130_TQ;
  wire [0:0] LIOI3_X0Y133_OLOGIC_X0Y133_D1;
  wire [0:0] LIOI3_X0Y133_OLOGIC_X0Y133_OQ;
  wire [0:0] LIOI3_X0Y133_OLOGIC_X0Y133_T1;
  wire [0:0] LIOI3_X0Y133_OLOGIC_X0Y133_TQ;
  wire [0:0] LIOI3_X0Y133_OLOGIC_X0Y134_D1;
  wire [0:0] LIOI3_X0Y133_OLOGIC_X0Y134_OQ;
  wire [0:0] LIOI3_X0Y133_OLOGIC_X0Y134_T1;
  wire [0:0] LIOI3_X0Y133_OLOGIC_X0Y134_TQ;
  wire [0:0] LIOI3_X0Y135_OLOGIC_X0Y135_D1;
  wire [0:0] LIOI3_X0Y135_OLOGIC_X0Y135_OQ;
  wire [0:0] LIOI3_X0Y135_OLOGIC_X0Y135_T1;
  wire [0:0] LIOI3_X0Y135_OLOGIC_X0Y135_TQ;
  wire [0:0] LIOI3_X0Y135_OLOGIC_X0Y136_D1;
  wire [0:0] LIOI3_X0Y135_OLOGIC_X0Y136_OQ;
  wire [0:0] LIOI3_X0Y135_OLOGIC_X0Y136_T1;
  wire [0:0] LIOI3_X0Y135_OLOGIC_X0Y136_TQ;
  wire [0:0] LIOI3_X0Y139_OLOGIC_X0Y139_D1;
  wire [0:0] LIOI3_X0Y139_OLOGIC_X0Y139_OQ;
  wire [0:0] LIOI3_X0Y139_OLOGIC_X0Y139_T1;
  wire [0:0] LIOI3_X0Y139_OLOGIC_X0Y139_TQ;
  wire [0:0] LIOI3_X0Y139_OLOGIC_X0Y140_D1;
  wire [0:0] LIOI3_X0Y139_OLOGIC_X0Y140_OQ;
  wire [0:0] LIOI3_X0Y139_OLOGIC_X0Y140_T1;
  wire [0:0] LIOI3_X0Y139_OLOGIC_X0Y140_TQ;
  wire [0:0] LIOI3_X0Y141_OLOGIC_X0Y141_D1;
  wire [0:0] LIOI3_X0Y141_OLOGIC_X0Y141_OQ;
  wire [0:0] LIOI3_X0Y141_OLOGIC_X0Y141_T1;
  wire [0:0] LIOI3_X0Y141_OLOGIC_X0Y141_TQ;
  wire [0:0] LIOI3_X0Y141_OLOGIC_X0Y142_D1;
  wire [0:0] LIOI3_X0Y141_OLOGIC_X0Y142_OQ;
  wire [0:0] LIOI3_X0Y141_OLOGIC_X0Y142_T1;
  wire [0:0] LIOI3_X0Y141_OLOGIC_X0Y142_TQ;
  wire [0:0] LIOI3_X0Y145_OLOGIC_X0Y145_D1;
  wire [0:0] LIOI3_X0Y145_OLOGIC_X0Y145_OQ;
  wire [0:0] LIOI3_X0Y145_OLOGIC_X0Y145_T1;
  wire [0:0] LIOI3_X0Y145_OLOGIC_X0Y145_TQ;
  wire [0:0] LIOI3_X0Y145_OLOGIC_X0Y146_D1;
  wire [0:0] LIOI3_X0Y145_OLOGIC_X0Y146_OQ;
  wire [0:0] LIOI3_X0Y145_OLOGIC_X0Y146_T1;
  wire [0:0] LIOI3_X0Y145_OLOGIC_X0Y146_TQ;
  wire [0:0] LIOI3_X0Y147_OLOGIC_X0Y147_D1;
  wire [0:0] LIOI3_X0Y147_OLOGIC_X0Y147_OQ;
  wire [0:0] LIOI3_X0Y147_OLOGIC_X0Y147_T1;
  wire [0:0] LIOI3_X0Y147_OLOGIC_X0Y147_TQ;
  wire [0:0] LIOI3_X0Y147_OLOGIC_X0Y148_D1;
  wire [0:0] LIOI3_X0Y147_OLOGIC_X0Y148_OQ;
  wire [0:0] LIOI3_X0Y147_OLOGIC_X0Y148_T1;
  wire [0:0] LIOI3_X0Y147_OLOGIC_X0Y148_TQ;
  wire [0:0] LIOI3_X0Y151_OLOGIC_X0Y151_D1;
  wire [0:0] LIOI3_X0Y151_OLOGIC_X0Y151_OQ;
  wire [0:0] LIOI3_X0Y151_OLOGIC_X0Y151_T1;
  wire [0:0] LIOI3_X0Y151_OLOGIC_X0Y151_TQ;
  wire [0:0] LIOI3_X0Y151_OLOGIC_X0Y152_D1;
  wire [0:0] LIOI3_X0Y151_OLOGIC_X0Y152_OQ;
  wire [0:0] LIOI3_X0Y151_OLOGIC_X0Y152_T1;
  wire [0:0] LIOI3_X0Y151_OLOGIC_X0Y152_TQ;
  wire [0:0] LIOI3_X0Y153_OLOGIC_X0Y153_D1;
  wire [0:0] LIOI3_X0Y153_OLOGIC_X0Y153_OQ;
  wire [0:0] LIOI3_X0Y153_OLOGIC_X0Y153_T1;
  wire [0:0] LIOI3_X0Y153_OLOGIC_X0Y153_TQ;
  wire [0:0] LIOI3_X0Y153_OLOGIC_X0Y154_D1;
  wire [0:0] LIOI3_X0Y153_OLOGIC_X0Y154_OQ;
  wire [0:0] LIOI3_X0Y153_OLOGIC_X0Y154_T1;
  wire [0:0] LIOI3_X0Y153_OLOGIC_X0Y154_TQ;
  wire [0:0] LIOI3_X0Y155_OLOGIC_X0Y155_D1;
  wire [0:0] LIOI3_X0Y155_OLOGIC_X0Y155_OQ;
  wire [0:0] LIOI3_X0Y155_OLOGIC_X0Y155_T1;
  wire [0:0] LIOI3_X0Y155_OLOGIC_X0Y155_TQ;
  wire [0:0] LIOI3_X0Y155_OLOGIC_X0Y156_D1;
  wire [0:0] LIOI3_X0Y155_OLOGIC_X0Y156_OQ;
  wire [0:0] LIOI3_X0Y155_OLOGIC_X0Y156_T1;
  wire [0:0] LIOI3_X0Y155_OLOGIC_X0Y156_TQ;
  wire [0:0] LIOI3_X0Y159_OLOGIC_X0Y159_D1;
  wire [0:0] LIOI3_X0Y159_OLOGIC_X0Y159_OQ;
  wire [0:0] LIOI3_X0Y159_OLOGIC_X0Y159_T1;
  wire [0:0] LIOI3_X0Y159_OLOGIC_X0Y159_TQ;
  wire [0:0] LIOI3_X0Y159_OLOGIC_X0Y160_D1;
  wire [0:0] LIOI3_X0Y159_OLOGIC_X0Y160_OQ;
  wire [0:0] LIOI3_X0Y159_OLOGIC_X0Y160_T1;
  wire [0:0] LIOI3_X0Y159_OLOGIC_X0Y160_TQ;
  wire [0:0] LIOI3_X0Y161_OLOGIC_X0Y161_D1;
  wire [0:0] LIOI3_X0Y161_OLOGIC_X0Y161_OQ;
  wire [0:0] LIOI3_X0Y161_OLOGIC_X0Y161_T1;
  wire [0:0] LIOI3_X0Y161_OLOGIC_X0Y161_TQ;
  wire [0:0] LIOI3_X0Y161_OLOGIC_X0Y162_D1;
  wire [0:0] LIOI3_X0Y161_OLOGIC_X0Y162_OQ;
  wire [0:0] LIOI3_X0Y161_OLOGIC_X0Y162_T1;
  wire [0:0] LIOI3_X0Y161_OLOGIC_X0Y162_TQ;
  wire [0:0] LIOI3_X0Y165_OLOGIC_X0Y165_D1;
  wire [0:0] LIOI3_X0Y165_OLOGIC_X0Y165_OQ;
  wire [0:0] LIOI3_X0Y165_OLOGIC_X0Y165_T1;
  wire [0:0] LIOI3_X0Y165_OLOGIC_X0Y165_TQ;
  wire [0:0] LIOI3_X0Y165_OLOGIC_X0Y166_D1;
  wire [0:0] LIOI3_X0Y165_OLOGIC_X0Y166_OQ;
  wire [0:0] LIOI3_X0Y165_OLOGIC_X0Y166_T1;
  wire [0:0] LIOI3_X0Y165_OLOGIC_X0Y166_TQ;
  wire [0:0] LIOI3_X0Y167_OLOGIC_X0Y167_D1;
  wire [0:0] LIOI3_X0Y167_OLOGIC_X0Y167_OQ;
  wire [0:0] LIOI3_X0Y167_OLOGIC_X0Y167_T1;
  wire [0:0] LIOI3_X0Y167_OLOGIC_X0Y167_TQ;
  wire [0:0] LIOI3_X0Y167_OLOGIC_X0Y168_D1;
  wire [0:0] LIOI3_X0Y167_OLOGIC_X0Y168_OQ;
  wire [0:0] LIOI3_X0Y167_OLOGIC_X0Y168_T1;
  wire [0:0] LIOI3_X0Y167_OLOGIC_X0Y168_TQ;
  wire [0:0] LIOI3_X0Y171_OLOGIC_X0Y171_D1;
  wire [0:0] LIOI3_X0Y171_OLOGIC_X0Y171_OQ;
  wire [0:0] LIOI3_X0Y171_OLOGIC_X0Y171_T1;
  wire [0:0] LIOI3_X0Y171_OLOGIC_X0Y171_TQ;
  wire [0:0] LIOI3_X0Y171_OLOGIC_X0Y172_D1;
  wire [0:0] LIOI3_X0Y171_OLOGIC_X0Y172_OQ;
  wire [0:0] LIOI3_X0Y171_OLOGIC_X0Y172_T1;
  wire [0:0] LIOI3_X0Y171_OLOGIC_X0Y172_TQ;
  wire [0:0] LIOI3_X0Y173_OLOGIC_X0Y173_D1;
  wire [0:0] LIOI3_X0Y173_OLOGIC_X0Y173_OQ;
  wire [0:0] LIOI3_X0Y173_OLOGIC_X0Y173_T1;
  wire [0:0] LIOI3_X0Y173_OLOGIC_X0Y173_TQ;
  wire [0:0] LIOI3_X0Y173_OLOGIC_X0Y174_D1;
  wire [0:0] LIOI3_X0Y173_OLOGIC_X0Y174_OQ;
  wire [0:0] LIOI3_X0Y173_OLOGIC_X0Y174_T1;
  wire [0:0] LIOI3_X0Y173_OLOGIC_X0Y174_TQ;
  wire [0:0] LIOI3_X0Y175_OLOGIC_X0Y175_D1;
  wire [0:0] LIOI3_X0Y175_OLOGIC_X0Y175_OQ;
  wire [0:0] LIOI3_X0Y175_OLOGIC_X0Y175_T1;
  wire [0:0] LIOI3_X0Y175_OLOGIC_X0Y175_TQ;
  wire [0:0] LIOI3_X0Y175_OLOGIC_X0Y176_D1;
  wire [0:0] LIOI3_X0Y175_OLOGIC_X0Y176_OQ;
  wire [0:0] LIOI3_X0Y175_OLOGIC_X0Y176_T1;
  wire [0:0] LIOI3_X0Y175_OLOGIC_X0Y176_TQ;
  wire [0:0] LIOI3_X0Y177_OLOGIC_X0Y177_D1;
  wire [0:0] LIOI3_X0Y177_OLOGIC_X0Y177_OQ;
  wire [0:0] LIOI3_X0Y177_OLOGIC_X0Y177_T1;
  wire [0:0] LIOI3_X0Y177_OLOGIC_X0Y177_TQ;
  wire [0:0] LIOI3_X0Y177_OLOGIC_X0Y178_D1;
  wire [0:0] LIOI3_X0Y177_OLOGIC_X0Y178_OQ;
  wire [0:0] LIOI3_X0Y177_OLOGIC_X0Y178_T1;
  wire [0:0] LIOI3_X0Y177_OLOGIC_X0Y178_TQ;
  wire [0:0] LIOI3_X0Y179_OLOGIC_X0Y179_D1;
  wire [0:0] LIOI3_X0Y179_OLOGIC_X0Y179_OQ;
  wire [0:0] LIOI3_X0Y179_OLOGIC_X0Y179_T1;
  wire [0:0] LIOI3_X0Y179_OLOGIC_X0Y179_TQ;
  wire [0:0] LIOI3_X0Y179_OLOGIC_X0Y180_D1;
  wire [0:0] LIOI3_X0Y179_OLOGIC_X0Y180_OQ;
  wire [0:0] LIOI3_X0Y179_OLOGIC_X0Y180_T1;
  wire [0:0] LIOI3_X0Y179_OLOGIC_X0Y180_TQ;
  wire [0:0] LIOI3_X0Y183_OLOGIC_X0Y183_D1;
  wire [0:0] LIOI3_X0Y183_OLOGIC_X0Y183_OQ;
  wire [0:0] LIOI3_X0Y183_OLOGIC_X0Y183_T1;
  wire [0:0] LIOI3_X0Y183_OLOGIC_X0Y183_TQ;
  wire [0:0] LIOI3_X0Y183_OLOGIC_X0Y184_D1;
  wire [0:0] LIOI3_X0Y183_OLOGIC_X0Y184_OQ;
  wire [0:0] LIOI3_X0Y183_OLOGIC_X0Y184_T1;
  wire [0:0] LIOI3_X0Y183_OLOGIC_X0Y184_TQ;
  wire [0:0] LIOI3_X0Y185_OLOGIC_X0Y185_D1;
  wire [0:0] LIOI3_X0Y185_OLOGIC_X0Y185_OQ;
  wire [0:0] LIOI3_X0Y185_OLOGIC_X0Y185_T1;
  wire [0:0] LIOI3_X0Y185_OLOGIC_X0Y185_TQ;
  wire [0:0] LIOI3_X0Y185_OLOGIC_X0Y186_D1;
  wire [0:0] LIOI3_X0Y185_OLOGIC_X0Y186_OQ;
  wire [0:0] LIOI3_X0Y185_OLOGIC_X0Y186_T1;
  wire [0:0] LIOI3_X0Y185_OLOGIC_X0Y186_TQ;
  wire [0:0] LIOI3_X0Y189_OLOGIC_X0Y189_D1;
  wire [0:0] LIOI3_X0Y189_OLOGIC_X0Y189_OQ;
  wire [0:0] LIOI3_X0Y189_OLOGIC_X0Y189_T1;
  wire [0:0] LIOI3_X0Y189_OLOGIC_X0Y189_TQ;
  wire [0:0] LIOI3_X0Y189_OLOGIC_X0Y190_D1;
  wire [0:0] LIOI3_X0Y189_OLOGIC_X0Y190_OQ;
  wire [0:0] LIOI3_X0Y189_OLOGIC_X0Y190_T1;
  wire [0:0] LIOI3_X0Y189_OLOGIC_X0Y190_TQ;
  wire [0:0] LIOI3_X0Y191_OLOGIC_X0Y191_D1;
  wire [0:0] LIOI3_X0Y191_OLOGIC_X0Y191_OQ;
  wire [0:0] LIOI3_X0Y191_OLOGIC_X0Y191_T1;
  wire [0:0] LIOI3_X0Y191_OLOGIC_X0Y191_TQ;
  wire [0:0] LIOI3_X0Y191_OLOGIC_X0Y192_D1;
  wire [0:0] LIOI3_X0Y191_OLOGIC_X0Y192_OQ;
  wire [0:0] LIOI3_X0Y191_OLOGIC_X0Y192_T1;
  wire [0:0] LIOI3_X0Y191_OLOGIC_X0Y192_TQ;
  wire [0:0] LIOI3_X0Y195_OLOGIC_X0Y195_D1;
  wire [0:0] LIOI3_X0Y195_OLOGIC_X0Y195_OQ;
  wire [0:0] LIOI3_X0Y195_OLOGIC_X0Y195_T1;
  wire [0:0] LIOI3_X0Y195_OLOGIC_X0Y195_TQ;
  wire [0:0] LIOI3_X0Y195_OLOGIC_X0Y196_D1;
  wire [0:0] LIOI3_X0Y195_OLOGIC_X0Y196_OQ;
  wire [0:0] LIOI3_X0Y195_OLOGIC_X0Y196_T1;
  wire [0:0] LIOI3_X0Y195_OLOGIC_X0Y196_TQ;
  wire [0:0] LIOI3_X0Y197_OLOGIC_X0Y197_D1;
  wire [0:0] LIOI3_X0Y197_OLOGIC_X0Y197_OQ;
  wire [0:0] LIOI3_X0Y197_OLOGIC_X0Y197_T1;
  wire [0:0] LIOI3_X0Y197_OLOGIC_X0Y197_TQ;
  wire [0:0] LIOI3_X0Y197_OLOGIC_X0Y198_D1;
  wire [0:0] LIOI3_X0Y197_OLOGIC_X0Y198_OQ;
  wire [0:0] LIOI3_X0Y197_OLOGIC_X0Y198_T1;
  wire [0:0] LIOI3_X0Y197_OLOGIC_X0Y198_TQ;
  wire [0:0] LIOI3_X0Y51_ILOGIC_X0Y51_D;
  wire [0:0] LIOI3_X0Y51_ILOGIC_X0Y51_O;
  wire [0:0] LIOI3_X0Y51_ILOGIC_X0Y52_D;
  wire [0:0] LIOI3_X0Y51_ILOGIC_X0Y52_O;
  wire [0:0] LIOI3_X0Y53_ILOGIC_X0Y53_D;
  wire [0:0] LIOI3_X0Y53_ILOGIC_X0Y53_O;
  wire [0:0] LIOI3_X0Y53_ILOGIC_X0Y54_D;
  wire [0:0] LIOI3_X0Y53_ILOGIC_X0Y54_O;
  wire [0:0] LIOI3_X0Y55_ILOGIC_X0Y55_D;
  wire [0:0] LIOI3_X0Y55_ILOGIC_X0Y55_O;
  wire [0:0] LIOI3_X0Y55_ILOGIC_X0Y56_D;
  wire [0:0] LIOI3_X0Y55_ILOGIC_X0Y56_O;
  wire [0:0] LIOI3_X0Y59_ILOGIC_X0Y59_D;
  wire [0:0] LIOI3_X0Y59_ILOGIC_X0Y59_O;
  wire [0:0] LIOI3_X0Y59_ILOGIC_X0Y60_D;
  wire [0:0] LIOI3_X0Y59_ILOGIC_X0Y60_O;
  wire [0:0] LIOI3_X0Y61_ILOGIC_X0Y61_D;
  wire [0:0] LIOI3_X0Y61_ILOGIC_X0Y61_O;
  wire [0:0] LIOI3_X0Y61_ILOGIC_X0Y62_D;
  wire [0:0] LIOI3_X0Y61_ILOGIC_X0Y62_O;
  wire [0:0] LIOI3_X0Y65_OLOGIC_X0Y65_D1;
  wire [0:0] LIOI3_X0Y65_OLOGIC_X0Y65_OQ;
  wire [0:0] LIOI3_X0Y65_OLOGIC_X0Y65_T1;
  wire [0:0] LIOI3_X0Y65_OLOGIC_X0Y65_TQ;
  wire [0:0] LIOI3_X0Y65_OLOGIC_X0Y66_D1;
  wire [0:0] LIOI3_X0Y65_OLOGIC_X0Y66_OQ;
  wire [0:0] LIOI3_X0Y65_OLOGIC_X0Y66_T1;
  wire [0:0] LIOI3_X0Y65_OLOGIC_X0Y66_TQ;
  wire [0:0] LIOI3_X0Y77_ILOGIC_X0Y78_D;
  wire [0:0] LIOI3_X0Y77_ILOGIC_X0Y78_O;
  wire [0:0] RIOB33_SING_X105Y100_IOB_X1Y100_I;
  wire [0:0] RIOB33_SING_X105Y149_IOB_X1Y149_I;
  wire [0:0] RIOB33_SING_X105Y150_IOB_X1Y150_O;
  wire [0:0] RIOB33_SING_X105Y199_IOB_X1Y199_O;
  wire [0:0] RIOB33_X105Y101_IOB_X1Y101_I;
  wire [0:0] RIOB33_X105Y101_IOB_X1Y102_I;
  wire [0:0] RIOB33_X105Y103_IOB_X1Y103_I;
  wire [0:0] RIOB33_X105Y103_IOB_X1Y104_I;
  wire [0:0] RIOB33_X105Y105_IOB_X1Y105_I;
  wire [0:0] RIOB33_X105Y105_IOB_X1Y106_I;
  wire [0:0] RIOB33_X105Y107_IOB_X1Y107_I;
  wire [0:0] RIOB33_X105Y107_IOB_X1Y108_I;
  wire [0:0] RIOB33_X105Y109_IOB_X1Y109_I;
  wire [0:0] RIOB33_X105Y109_IOB_X1Y110_I;
  wire [0:0] RIOB33_X105Y111_IOB_X1Y111_I;
  wire [0:0] RIOB33_X105Y111_IOB_X1Y112_I;
  wire [0:0] RIOB33_X105Y113_IOB_X1Y113_I;
  wire [0:0] RIOB33_X105Y113_IOB_X1Y114_I;
  wire [0:0] RIOB33_X105Y115_IOB_X1Y115_I;
  wire [0:0] RIOB33_X105Y115_IOB_X1Y116_I;
  wire [0:0] RIOB33_X105Y117_IOB_X1Y117_I;
  wire [0:0] RIOB33_X105Y117_IOB_X1Y118_I;
  wire [0:0] RIOB33_X105Y119_IOB_X1Y119_I;
  wire [0:0] RIOB33_X105Y119_IOB_X1Y120_I;
  wire [0:0] RIOB33_X105Y121_IOB_X1Y121_I;
  wire [0:0] RIOB33_X105Y121_IOB_X1Y122_I;
  wire [0:0] RIOB33_X105Y123_IOB_X1Y123_I;
  wire [0:0] RIOB33_X105Y123_IOB_X1Y124_I;
  wire [0:0] RIOB33_X105Y125_IOB_X1Y125_I;
  wire [0:0] RIOB33_X105Y125_IOB_X1Y126_I;
  wire [0:0] RIOB33_X105Y127_IOB_X1Y127_I;
  wire [0:0] RIOB33_X105Y127_IOB_X1Y128_I;
  wire [0:0] RIOB33_X105Y129_IOB_X1Y129_I;
  wire [0:0] RIOB33_X105Y129_IOB_X1Y130_I;
  wire [0:0] RIOB33_X105Y131_IOB_X1Y131_I;
  wire [0:0] RIOB33_X105Y131_IOB_X1Y132_I;
  wire [0:0] RIOB33_X105Y133_IOB_X1Y133_I;
  wire [0:0] RIOB33_X105Y133_IOB_X1Y134_I;
  wire [0:0] RIOB33_X105Y135_IOB_X1Y135_I;
  wire [0:0] RIOB33_X105Y135_IOB_X1Y136_I;
  wire [0:0] RIOB33_X105Y137_IOB_X1Y137_I;
  wire [0:0] RIOB33_X105Y137_IOB_X1Y138_I;
  wire [0:0] RIOB33_X105Y139_IOB_X1Y139_I;
  wire [0:0] RIOB33_X105Y139_IOB_X1Y140_I;
  wire [0:0] RIOB33_X105Y141_IOB_X1Y141_I;
  wire [0:0] RIOB33_X105Y141_IOB_X1Y142_I;
  wire [0:0] RIOB33_X105Y143_IOB_X1Y143_I;
  wire [0:0] RIOB33_X105Y143_IOB_X1Y144_I;
  wire [0:0] RIOB33_X105Y145_IOB_X1Y145_I;
  wire [0:0] RIOB33_X105Y145_IOB_X1Y146_I;
  wire [0:0] RIOB33_X105Y147_IOB_X1Y147_I;
  wire [0:0] RIOB33_X105Y147_IOB_X1Y148_I;
  wire [0:0] RIOB33_X105Y151_IOB_X1Y151_O;
  wire [0:0] RIOB33_X105Y151_IOB_X1Y152_O;
  wire [0:0] RIOB33_X105Y153_IOB_X1Y153_O;
  wire [0:0] RIOB33_X105Y153_IOB_X1Y154_O;
  wire [0:0] RIOB33_X105Y155_IOB_X1Y155_O;
  wire [0:0] RIOB33_X105Y155_IOB_X1Y156_O;
  wire [0:0] RIOB33_X105Y157_IOB_X1Y157_O;
  wire [0:0] RIOB33_X105Y157_IOB_X1Y158_O;
  wire [0:0] RIOB33_X105Y159_IOB_X1Y159_O;
  wire [0:0] RIOB33_X105Y159_IOB_X1Y160_O;
  wire [0:0] RIOB33_X105Y161_IOB_X1Y161_O;
  wire [0:0] RIOB33_X105Y161_IOB_X1Y162_O;
  wire [0:0] RIOB33_X105Y163_IOB_X1Y163_O;
  wire [0:0] RIOB33_X105Y163_IOB_X1Y164_O;
  wire [0:0] RIOB33_X105Y165_IOB_X1Y165_O;
  wire [0:0] RIOB33_X105Y165_IOB_X1Y166_O;
  wire [0:0] RIOB33_X105Y167_IOB_X1Y167_O;
  wire [0:0] RIOB33_X105Y167_IOB_X1Y168_O;
  wire [0:0] RIOB33_X105Y169_IOB_X1Y169_O;
  wire [0:0] RIOB33_X105Y169_IOB_X1Y170_O;
  wire [0:0] RIOB33_X105Y171_IOB_X1Y171_O;
  wire [0:0] RIOB33_X105Y171_IOB_X1Y172_O;
  wire [0:0] RIOB33_X105Y173_IOB_X1Y173_O;
  wire [0:0] RIOB33_X105Y173_IOB_X1Y174_O;
  wire [0:0] RIOB33_X105Y175_IOB_X1Y175_O;
  wire [0:0] RIOB33_X105Y175_IOB_X1Y176_O;
  wire [0:0] RIOB33_X105Y177_IOB_X1Y177_O;
  wire [0:0] RIOB33_X105Y177_IOB_X1Y178_O;
  wire [0:0] RIOB33_X105Y179_IOB_X1Y179_O;
  wire [0:0] RIOB33_X105Y179_IOB_X1Y180_O;
  wire [0:0] RIOB33_X105Y181_IOB_X1Y181_O;
  wire [0:0] RIOB33_X105Y181_IOB_X1Y182_O;
  wire [0:0] RIOB33_X105Y183_IOB_X1Y183_O;
  wire [0:0] RIOB33_X105Y183_IOB_X1Y184_O;
  wire [0:0] RIOB33_X105Y185_IOB_X1Y185_O;
  wire [0:0] RIOB33_X105Y185_IOB_X1Y186_O;
  wire [0:0] RIOB33_X105Y187_IOB_X1Y187_O;
  wire [0:0] RIOB33_X105Y187_IOB_X1Y188_O;
  wire [0:0] RIOB33_X105Y189_IOB_X1Y189_O;
  wire [0:0] RIOB33_X105Y189_IOB_X1Y190_O;
  wire [0:0] RIOB33_X105Y191_IOB_X1Y191_O;
  wire [0:0] RIOB33_X105Y191_IOB_X1Y192_O;
  wire [0:0] RIOB33_X105Y193_IOB_X1Y193_O;
  wire [0:0] RIOB33_X105Y193_IOB_X1Y194_O;
  wire [0:0] RIOB33_X105Y195_IOB_X1Y195_O;
  wire [0:0] RIOB33_X105Y195_IOB_X1Y196_O;
  wire [0:0] RIOB33_X105Y197_IOB_X1Y197_O;
  wire [0:0] RIOB33_X105Y197_IOB_X1Y198_O;
  wire [0:0] RIOI3_SING_X105Y100_ILOGIC_X1Y100_D;
  wire [0:0] RIOI3_SING_X105Y100_ILOGIC_X1Y100_O;
  wire [0:0] RIOI3_SING_X105Y149_ILOGIC_X1Y149_D;
  wire [0:0] RIOI3_SING_X105Y149_ILOGIC_X1Y149_O;
  wire [0:0] RIOI3_SING_X105Y150_OLOGIC_X1Y150_D1;
  wire [0:0] RIOI3_SING_X105Y150_OLOGIC_X1Y150_OQ;
  wire [0:0] RIOI3_SING_X105Y150_OLOGIC_X1Y150_T1;
  wire [0:0] RIOI3_SING_X105Y150_OLOGIC_X1Y150_TQ;
  wire [0:0] RIOI3_SING_X105Y199_OLOGIC_X1Y199_D1;
  wire [0:0] RIOI3_SING_X105Y199_OLOGIC_X1Y199_OQ;
  wire [0:0] RIOI3_SING_X105Y199_OLOGIC_X1Y199_T1;
  wire [0:0] RIOI3_SING_X105Y199_OLOGIC_X1Y199_TQ;
  wire [0:0] RIOI3_TBYTESRC_X105Y107_ILOGIC_X1Y107_D;
  wire [0:0] RIOI3_TBYTESRC_X105Y107_ILOGIC_X1Y107_O;
  wire [0:0] RIOI3_TBYTESRC_X105Y107_ILOGIC_X1Y108_D;
  wire [0:0] RIOI3_TBYTESRC_X105Y107_ILOGIC_X1Y108_O;
  wire [0:0] RIOI3_TBYTESRC_X105Y119_ILOGIC_X1Y119_D;
  wire [0:0] RIOI3_TBYTESRC_X105Y119_ILOGIC_X1Y119_O;
  wire [0:0] RIOI3_TBYTESRC_X105Y119_ILOGIC_X1Y120_D;
  wire [0:0] RIOI3_TBYTESRC_X105Y119_ILOGIC_X1Y120_O;
  wire [0:0] RIOI3_TBYTESRC_X105Y131_ILOGIC_X1Y131_D;
  wire [0:0] RIOI3_TBYTESRC_X105Y131_ILOGIC_X1Y131_O;
  wire [0:0] RIOI3_TBYTESRC_X105Y131_ILOGIC_X1Y132_D;
  wire [0:0] RIOI3_TBYTESRC_X105Y131_ILOGIC_X1Y132_O;
  wire [0:0] RIOI3_TBYTESRC_X105Y143_ILOGIC_X1Y143_D;
  wire [0:0] RIOI3_TBYTESRC_X105Y143_ILOGIC_X1Y143_O;
  wire [0:0] RIOI3_TBYTESRC_X105Y143_ILOGIC_X1Y144_D;
  wire [0:0] RIOI3_TBYTESRC_X105Y143_ILOGIC_X1Y144_O;
  wire [0:0] RIOI3_TBYTESRC_X105Y157_OLOGIC_X1Y157_D1;
  wire [0:0] RIOI3_TBYTESRC_X105Y157_OLOGIC_X1Y157_OQ;
  wire [0:0] RIOI3_TBYTESRC_X105Y157_OLOGIC_X1Y157_T1;
  wire [0:0] RIOI3_TBYTESRC_X105Y157_OLOGIC_X1Y157_TQ;
  wire [0:0] RIOI3_TBYTESRC_X105Y157_OLOGIC_X1Y158_D1;
  wire [0:0] RIOI3_TBYTESRC_X105Y157_OLOGIC_X1Y158_OQ;
  wire [0:0] RIOI3_TBYTESRC_X105Y157_OLOGIC_X1Y158_T1;
  wire [0:0] RIOI3_TBYTESRC_X105Y157_OLOGIC_X1Y158_TQ;
  wire [0:0] RIOI3_TBYTESRC_X105Y169_OLOGIC_X1Y169_D1;
  wire [0:0] RIOI3_TBYTESRC_X105Y169_OLOGIC_X1Y169_OQ;
  wire [0:0] RIOI3_TBYTESRC_X105Y169_OLOGIC_X1Y169_T1;
  wire [0:0] RIOI3_TBYTESRC_X105Y169_OLOGIC_X1Y169_TQ;
  wire [0:0] RIOI3_TBYTESRC_X105Y169_OLOGIC_X1Y170_D1;
  wire [0:0] RIOI3_TBYTESRC_X105Y169_OLOGIC_X1Y170_OQ;
  wire [0:0] RIOI3_TBYTESRC_X105Y169_OLOGIC_X1Y170_T1;
  wire [0:0] RIOI3_TBYTESRC_X105Y169_OLOGIC_X1Y170_TQ;
  wire [0:0] RIOI3_TBYTESRC_X105Y181_OLOGIC_X1Y181_D1;
  wire [0:0] RIOI3_TBYTESRC_X105Y181_OLOGIC_X1Y181_OQ;
  wire [0:0] RIOI3_TBYTESRC_X105Y181_OLOGIC_X1Y181_T1;
  wire [0:0] RIOI3_TBYTESRC_X105Y181_OLOGIC_X1Y181_TQ;
  wire [0:0] RIOI3_TBYTESRC_X105Y181_OLOGIC_X1Y182_D1;
  wire [0:0] RIOI3_TBYTESRC_X105Y181_OLOGIC_X1Y182_OQ;
  wire [0:0] RIOI3_TBYTESRC_X105Y181_OLOGIC_X1Y182_T1;
  wire [0:0] RIOI3_TBYTESRC_X105Y181_OLOGIC_X1Y182_TQ;
  wire [0:0] RIOI3_TBYTESRC_X105Y193_OLOGIC_X1Y193_D1;
  wire [0:0] RIOI3_TBYTESRC_X105Y193_OLOGIC_X1Y193_OQ;
  wire [0:0] RIOI3_TBYTESRC_X105Y193_OLOGIC_X1Y193_T1;
  wire [0:0] RIOI3_TBYTESRC_X105Y193_OLOGIC_X1Y193_TQ;
  wire [0:0] RIOI3_TBYTESRC_X105Y193_OLOGIC_X1Y194_D1;
  wire [0:0] RIOI3_TBYTESRC_X105Y193_OLOGIC_X1Y194_OQ;
  wire [0:0] RIOI3_TBYTESRC_X105Y193_OLOGIC_X1Y194_T1;
  wire [0:0] RIOI3_TBYTESRC_X105Y193_OLOGIC_X1Y194_TQ;
  wire [0:0] RIOI3_TBYTETERM_X105Y113_ILOGIC_X1Y113_D;
  wire [0:0] RIOI3_TBYTETERM_X105Y113_ILOGIC_X1Y113_O;
  wire [0:0] RIOI3_TBYTETERM_X105Y137_ILOGIC_X1Y137_D;
  wire [0:0] RIOI3_TBYTETERM_X105Y137_ILOGIC_X1Y137_O;
  wire [0:0] RIOI3_TBYTETERM_X105Y137_ILOGIC_X1Y138_D;
  wire [0:0] RIOI3_TBYTETERM_X105Y137_ILOGIC_X1Y138_O;
  wire [0:0] RIOI3_TBYTETERM_X105Y163_OLOGIC_X1Y163_D1;
  wire [0:0] RIOI3_TBYTETERM_X105Y163_OLOGIC_X1Y163_OQ;
  wire [0:0] RIOI3_TBYTETERM_X105Y163_OLOGIC_X1Y163_T1;
  wire [0:0] RIOI3_TBYTETERM_X105Y163_OLOGIC_X1Y163_TQ;
  wire [0:0] RIOI3_TBYTETERM_X105Y163_OLOGIC_X1Y164_D1;
  wire [0:0] RIOI3_TBYTETERM_X105Y163_OLOGIC_X1Y164_OQ;
  wire [0:0] RIOI3_TBYTETERM_X105Y163_OLOGIC_X1Y164_T1;
  wire [0:0] RIOI3_TBYTETERM_X105Y163_OLOGIC_X1Y164_TQ;
  wire [0:0] RIOI3_TBYTETERM_X105Y187_OLOGIC_X1Y187_D1;
  wire [0:0] RIOI3_TBYTETERM_X105Y187_OLOGIC_X1Y187_OQ;
  wire [0:0] RIOI3_TBYTETERM_X105Y187_OLOGIC_X1Y187_T1;
  wire [0:0] RIOI3_TBYTETERM_X105Y187_OLOGIC_X1Y187_TQ;
  wire [0:0] RIOI3_TBYTETERM_X105Y187_OLOGIC_X1Y188_D1;
  wire [0:0] RIOI3_TBYTETERM_X105Y187_OLOGIC_X1Y188_OQ;
  wire [0:0] RIOI3_TBYTETERM_X105Y187_OLOGIC_X1Y188_T1;
  wire [0:0] RIOI3_TBYTETERM_X105Y187_OLOGIC_X1Y188_TQ;
  wire [0:0] RIOI3_X105Y101_ILOGIC_X1Y101_D;
  wire [0:0] RIOI3_X105Y101_ILOGIC_X1Y101_O;
  wire [0:0] RIOI3_X105Y101_ILOGIC_X1Y102_D;
  wire [0:0] RIOI3_X105Y101_ILOGIC_X1Y102_O;
  wire [0:0] RIOI3_X105Y103_ILOGIC_X1Y103_D;
  wire [0:0] RIOI3_X105Y103_ILOGIC_X1Y103_O;
  wire [0:0] RIOI3_X105Y103_ILOGIC_X1Y104_D;
  wire [0:0] RIOI3_X105Y103_ILOGIC_X1Y104_O;
  wire [0:0] RIOI3_X105Y105_ILOGIC_X1Y105_D;
  wire [0:0] RIOI3_X105Y105_ILOGIC_X1Y105_O;
  wire [0:0] RIOI3_X105Y105_ILOGIC_X1Y106_D;
  wire [0:0] RIOI3_X105Y105_ILOGIC_X1Y106_O;
  wire [0:0] RIOI3_X105Y109_ILOGIC_X1Y109_D;
  wire [0:0] RIOI3_X105Y109_ILOGIC_X1Y109_O;
  wire [0:0] RIOI3_X105Y109_ILOGIC_X1Y110_D;
  wire [0:0] RIOI3_X105Y109_ILOGIC_X1Y110_O;
  wire [0:0] RIOI3_X105Y111_ILOGIC_X1Y111_D;
  wire [0:0] RIOI3_X105Y111_ILOGIC_X1Y111_O;
  wire [0:0] RIOI3_X105Y111_ILOGIC_X1Y112_D;
  wire [0:0] RIOI3_X105Y111_ILOGIC_X1Y112_O;
  wire [0:0] RIOI3_X105Y115_ILOGIC_X1Y115_D;
  wire [0:0] RIOI3_X105Y115_ILOGIC_X1Y115_O;
  wire [0:0] RIOI3_X105Y115_ILOGIC_X1Y116_D;
  wire [0:0] RIOI3_X105Y115_ILOGIC_X1Y116_O;
  wire [0:0] RIOI3_X105Y117_ILOGIC_X1Y117_D;
  wire [0:0] RIOI3_X105Y117_ILOGIC_X1Y117_O;
  wire [0:0] RIOI3_X105Y117_ILOGIC_X1Y118_D;
  wire [0:0] RIOI3_X105Y117_ILOGIC_X1Y118_O;
  wire [0:0] RIOI3_X105Y121_ILOGIC_X1Y121_D;
  wire [0:0] RIOI3_X105Y121_ILOGIC_X1Y121_O;
  wire [0:0] RIOI3_X105Y121_ILOGIC_X1Y122_D;
  wire [0:0] RIOI3_X105Y121_ILOGIC_X1Y122_O;
  wire [0:0] RIOI3_X105Y123_ILOGIC_X1Y123_D;
  wire [0:0] RIOI3_X105Y123_ILOGIC_X1Y123_O;
  wire [0:0] RIOI3_X105Y123_ILOGIC_X1Y124_D;
  wire [0:0] RIOI3_X105Y123_ILOGIC_X1Y124_O;
  wire [0:0] RIOI3_X105Y125_ILOGIC_X1Y125_D;
  wire [0:0] RIOI3_X105Y125_ILOGIC_X1Y125_O;
  wire [0:0] RIOI3_X105Y125_ILOGIC_X1Y126_D;
  wire [0:0] RIOI3_X105Y125_ILOGIC_X1Y126_O;
  wire [0:0] RIOI3_X105Y127_ILOGIC_X1Y127_D;
  wire [0:0] RIOI3_X105Y127_ILOGIC_X1Y127_O;
  wire [0:0] RIOI3_X105Y127_ILOGIC_X1Y128_D;
  wire [0:0] RIOI3_X105Y127_ILOGIC_X1Y128_O;
  wire [0:0] RIOI3_X105Y129_ILOGIC_X1Y129_D;
  wire [0:0] RIOI3_X105Y129_ILOGIC_X1Y129_O;
  wire [0:0] RIOI3_X105Y129_ILOGIC_X1Y130_D;
  wire [0:0] RIOI3_X105Y129_ILOGIC_X1Y130_O;
  wire [0:0] RIOI3_X105Y133_ILOGIC_X1Y133_D;
  wire [0:0] RIOI3_X105Y133_ILOGIC_X1Y133_O;
  wire [0:0] RIOI3_X105Y133_ILOGIC_X1Y134_D;
  wire [0:0] RIOI3_X105Y133_ILOGIC_X1Y134_O;
  wire [0:0] RIOI3_X105Y135_ILOGIC_X1Y135_D;
  wire [0:0] RIOI3_X105Y135_ILOGIC_X1Y135_O;
  wire [0:0] RIOI3_X105Y135_ILOGIC_X1Y136_D;
  wire [0:0] RIOI3_X105Y135_ILOGIC_X1Y136_O;
  wire [0:0] RIOI3_X105Y139_ILOGIC_X1Y139_D;
  wire [0:0] RIOI3_X105Y139_ILOGIC_X1Y139_O;
  wire [0:0] RIOI3_X105Y139_ILOGIC_X1Y140_D;
  wire [0:0] RIOI3_X105Y139_ILOGIC_X1Y140_O;
  wire [0:0] RIOI3_X105Y141_ILOGIC_X1Y141_D;
  wire [0:0] RIOI3_X105Y141_ILOGIC_X1Y141_O;
  wire [0:0] RIOI3_X105Y141_ILOGIC_X1Y142_D;
  wire [0:0] RIOI3_X105Y141_ILOGIC_X1Y142_O;
  wire [0:0] RIOI3_X105Y145_ILOGIC_X1Y145_D;
  wire [0:0] RIOI3_X105Y145_ILOGIC_X1Y145_O;
  wire [0:0] RIOI3_X105Y145_ILOGIC_X1Y146_D;
  wire [0:0] RIOI3_X105Y145_ILOGIC_X1Y146_O;
  wire [0:0] RIOI3_X105Y147_ILOGIC_X1Y147_D;
  wire [0:0] RIOI3_X105Y147_ILOGIC_X1Y147_O;
  wire [0:0] RIOI3_X105Y147_ILOGIC_X1Y148_D;
  wire [0:0] RIOI3_X105Y147_ILOGIC_X1Y148_O;
  wire [0:0] RIOI3_X105Y151_OLOGIC_X1Y151_D1;
  wire [0:0] RIOI3_X105Y151_OLOGIC_X1Y151_OQ;
  wire [0:0] RIOI3_X105Y151_OLOGIC_X1Y151_T1;
  wire [0:0] RIOI3_X105Y151_OLOGIC_X1Y151_TQ;
  wire [0:0] RIOI3_X105Y151_OLOGIC_X1Y152_D1;
  wire [0:0] RIOI3_X105Y151_OLOGIC_X1Y152_OQ;
  wire [0:0] RIOI3_X105Y151_OLOGIC_X1Y152_T1;
  wire [0:0] RIOI3_X105Y151_OLOGIC_X1Y152_TQ;
  wire [0:0] RIOI3_X105Y153_OLOGIC_X1Y153_D1;
  wire [0:0] RIOI3_X105Y153_OLOGIC_X1Y153_OQ;
  wire [0:0] RIOI3_X105Y153_OLOGIC_X1Y153_T1;
  wire [0:0] RIOI3_X105Y153_OLOGIC_X1Y153_TQ;
  wire [0:0] RIOI3_X105Y153_OLOGIC_X1Y154_D1;
  wire [0:0] RIOI3_X105Y153_OLOGIC_X1Y154_OQ;
  wire [0:0] RIOI3_X105Y153_OLOGIC_X1Y154_T1;
  wire [0:0] RIOI3_X105Y153_OLOGIC_X1Y154_TQ;
  wire [0:0] RIOI3_X105Y155_OLOGIC_X1Y155_D1;
  wire [0:0] RIOI3_X105Y155_OLOGIC_X1Y155_OQ;
  wire [0:0] RIOI3_X105Y155_OLOGIC_X1Y155_T1;
  wire [0:0] RIOI3_X105Y155_OLOGIC_X1Y155_TQ;
  wire [0:0] RIOI3_X105Y155_OLOGIC_X1Y156_D1;
  wire [0:0] RIOI3_X105Y155_OLOGIC_X1Y156_OQ;
  wire [0:0] RIOI3_X105Y155_OLOGIC_X1Y156_T1;
  wire [0:0] RIOI3_X105Y155_OLOGIC_X1Y156_TQ;
  wire [0:0] RIOI3_X105Y159_OLOGIC_X1Y159_D1;
  wire [0:0] RIOI3_X105Y159_OLOGIC_X1Y159_OQ;
  wire [0:0] RIOI3_X105Y159_OLOGIC_X1Y159_T1;
  wire [0:0] RIOI3_X105Y159_OLOGIC_X1Y159_TQ;
  wire [0:0] RIOI3_X105Y159_OLOGIC_X1Y160_D1;
  wire [0:0] RIOI3_X105Y159_OLOGIC_X1Y160_OQ;
  wire [0:0] RIOI3_X105Y159_OLOGIC_X1Y160_T1;
  wire [0:0] RIOI3_X105Y159_OLOGIC_X1Y160_TQ;
  wire [0:0] RIOI3_X105Y161_OLOGIC_X1Y161_D1;
  wire [0:0] RIOI3_X105Y161_OLOGIC_X1Y161_OQ;
  wire [0:0] RIOI3_X105Y161_OLOGIC_X1Y161_T1;
  wire [0:0] RIOI3_X105Y161_OLOGIC_X1Y161_TQ;
  wire [0:0] RIOI3_X105Y161_OLOGIC_X1Y162_D1;
  wire [0:0] RIOI3_X105Y161_OLOGIC_X1Y162_OQ;
  wire [0:0] RIOI3_X105Y161_OLOGIC_X1Y162_T1;
  wire [0:0] RIOI3_X105Y161_OLOGIC_X1Y162_TQ;
  wire [0:0] RIOI3_X105Y165_OLOGIC_X1Y165_D1;
  wire [0:0] RIOI3_X105Y165_OLOGIC_X1Y165_OQ;
  wire [0:0] RIOI3_X105Y165_OLOGIC_X1Y165_T1;
  wire [0:0] RIOI3_X105Y165_OLOGIC_X1Y165_TQ;
  wire [0:0] RIOI3_X105Y165_OLOGIC_X1Y166_D1;
  wire [0:0] RIOI3_X105Y165_OLOGIC_X1Y166_OQ;
  wire [0:0] RIOI3_X105Y165_OLOGIC_X1Y166_T1;
  wire [0:0] RIOI3_X105Y165_OLOGIC_X1Y166_TQ;
  wire [0:0] RIOI3_X105Y167_OLOGIC_X1Y167_D1;
  wire [0:0] RIOI3_X105Y167_OLOGIC_X1Y167_OQ;
  wire [0:0] RIOI3_X105Y167_OLOGIC_X1Y167_T1;
  wire [0:0] RIOI3_X105Y167_OLOGIC_X1Y167_TQ;
  wire [0:0] RIOI3_X105Y167_OLOGIC_X1Y168_D1;
  wire [0:0] RIOI3_X105Y167_OLOGIC_X1Y168_OQ;
  wire [0:0] RIOI3_X105Y167_OLOGIC_X1Y168_T1;
  wire [0:0] RIOI3_X105Y167_OLOGIC_X1Y168_TQ;
  wire [0:0] RIOI3_X105Y171_OLOGIC_X1Y171_D1;
  wire [0:0] RIOI3_X105Y171_OLOGIC_X1Y171_OQ;
  wire [0:0] RIOI3_X105Y171_OLOGIC_X1Y171_T1;
  wire [0:0] RIOI3_X105Y171_OLOGIC_X1Y171_TQ;
  wire [0:0] RIOI3_X105Y171_OLOGIC_X1Y172_D1;
  wire [0:0] RIOI3_X105Y171_OLOGIC_X1Y172_OQ;
  wire [0:0] RIOI3_X105Y171_OLOGIC_X1Y172_T1;
  wire [0:0] RIOI3_X105Y171_OLOGIC_X1Y172_TQ;
  wire [0:0] RIOI3_X105Y173_OLOGIC_X1Y173_D1;
  wire [0:0] RIOI3_X105Y173_OLOGIC_X1Y173_OQ;
  wire [0:0] RIOI3_X105Y173_OLOGIC_X1Y173_T1;
  wire [0:0] RIOI3_X105Y173_OLOGIC_X1Y173_TQ;
  wire [0:0] RIOI3_X105Y173_OLOGIC_X1Y174_D1;
  wire [0:0] RIOI3_X105Y173_OLOGIC_X1Y174_OQ;
  wire [0:0] RIOI3_X105Y173_OLOGIC_X1Y174_T1;
  wire [0:0] RIOI3_X105Y173_OLOGIC_X1Y174_TQ;
  wire [0:0] RIOI3_X105Y175_OLOGIC_X1Y175_D1;
  wire [0:0] RIOI3_X105Y175_OLOGIC_X1Y175_OQ;
  wire [0:0] RIOI3_X105Y175_OLOGIC_X1Y175_T1;
  wire [0:0] RIOI3_X105Y175_OLOGIC_X1Y175_TQ;
  wire [0:0] RIOI3_X105Y175_OLOGIC_X1Y176_D1;
  wire [0:0] RIOI3_X105Y175_OLOGIC_X1Y176_OQ;
  wire [0:0] RIOI3_X105Y175_OLOGIC_X1Y176_T1;
  wire [0:0] RIOI3_X105Y175_OLOGIC_X1Y176_TQ;
  wire [0:0] RIOI3_X105Y177_OLOGIC_X1Y177_D1;
  wire [0:0] RIOI3_X105Y177_OLOGIC_X1Y177_OQ;
  wire [0:0] RIOI3_X105Y177_OLOGIC_X1Y177_T1;
  wire [0:0] RIOI3_X105Y177_OLOGIC_X1Y177_TQ;
  wire [0:0] RIOI3_X105Y177_OLOGIC_X1Y178_D1;
  wire [0:0] RIOI3_X105Y177_OLOGIC_X1Y178_OQ;
  wire [0:0] RIOI3_X105Y177_OLOGIC_X1Y178_T1;
  wire [0:0] RIOI3_X105Y177_OLOGIC_X1Y178_TQ;
  wire [0:0] RIOI3_X105Y179_OLOGIC_X1Y179_D1;
  wire [0:0] RIOI3_X105Y179_OLOGIC_X1Y179_OQ;
  wire [0:0] RIOI3_X105Y179_OLOGIC_X1Y179_T1;
  wire [0:0] RIOI3_X105Y179_OLOGIC_X1Y179_TQ;
  wire [0:0] RIOI3_X105Y179_OLOGIC_X1Y180_D1;
  wire [0:0] RIOI3_X105Y179_OLOGIC_X1Y180_OQ;
  wire [0:0] RIOI3_X105Y179_OLOGIC_X1Y180_T1;
  wire [0:0] RIOI3_X105Y179_OLOGIC_X1Y180_TQ;
  wire [0:0] RIOI3_X105Y183_OLOGIC_X1Y183_D1;
  wire [0:0] RIOI3_X105Y183_OLOGIC_X1Y183_OQ;
  wire [0:0] RIOI3_X105Y183_OLOGIC_X1Y183_T1;
  wire [0:0] RIOI3_X105Y183_OLOGIC_X1Y183_TQ;
  wire [0:0] RIOI3_X105Y183_OLOGIC_X1Y184_D1;
  wire [0:0] RIOI3_X105Y183_OLOGIC_X1Y184_OQ;
  wire [0:0] RIOI3_X105Y183_OLOGIC_X1Y184_T1;
  wire [0:0] RIOI3_X105Y183_OLOGIC_X1Y184_TQ;
  wire [0:0] RIOI3_X105Y185_OLOGIC_X1Y185_D1;
  wire [0:0] RIOI3_X105Y185_OLOGIC_X1Y185_OQ;
  wire [0:0] RIOI3_X105Y185_OLOGIC_X1Y185_T1;
  wire [0:0] RIOI3_X105Y185_OLOGIC_X1Y185_TQ;
  wire [0:0] RIOI3_X105Y185_OLOGIC_X1Y186_D1;
  wire [0:0] RIOI3_X105Y185_OLOGIC_X1Y186_OQ;
  wire [0:0] RIOI3_X105Y185_OLOGIC_X1Y186_T1;
  wire [0:0] RIOI3_X105Y185_OLOGIC_X1Y186_TQ;
  wire [0:0] RIOI3_X105Y189_OLOGIC_X1Y189_D1;
  wire [0:0] RIOI3_X105Y189_OLOGIC_X1Y189_OQ;
  wire [0:0] RIOI3_X105Y189_OLOGIC_X1Y189_T1;
  wire [0:0] RIOI3_X105Y189_OLOGIC_X1Y189_TQ;
  wire [0:0] RIOI3_X105Y189_OLOGIC_X1Y190_D1;
  wire [0:0] RIOI3_X105Y189_OLOGIC_X1Y190_OQ;
  wire [0:0] RIOI3_X105Y189_OLOGIC_X1Y190_T1;
  wire [0:0] RIOI3_X105Y189_OLOGIC_X1Y190_TQ;
  wire [0:0] RIOI3_X105Y191_OLOGIC_X1Y191_D1;
  wire [0:0] RIOI3_X105Y191_OLOGIC_X1Y191_OQ;
  wire [0:0] RIOI3_X105Y191_OLOGIC_X1Y191_T1;
  wire [0:0] RIOI3_X105Y191_OLOGIC_X1Y191_TQ;
  wire [0:0] RIOI3_X105Y191_OLOGIC_X1Y192_D1;
  wire [0:0] RIOI3_X105Y191_OLOGIC_X1Y192_OQ;
  wire [0:0] RIOI3_X105Y191_OLOGIC_X1Y192_T1;
  wire [0:0] RIOI3_X105Y191_OLOGIC_X1Y192_TQ;
  wire [0:0] RIOI3_X105Y195_OLOGIC_X1Y195_D1;
  wire [0:0] RIOI3_X105Y195_OLOGIC_X1Y195_OQ;
  wire [0:0] RIOI3_X105Y195_OLOGIC_X1Y195_T1;
  wire [0:0] RIOI3_X105Y195_OLOGIC_X1Y195_TQ;
  wire [0:0] RIOI3_X105Y195_OLOGIC_X1Y196_D1;
  wire [0:0] RIOI3_X105Y195_OLOGIC_X1Y196_OQ;
  wire [0:0] RIOI3_X105Y195_OLOGIC_X1Y196_T1;
  wire [0:0] RIOI3_X105Y195_OLOGIC_X1Y196_TQ;
  wire [0:0] RIOI3_X105Y197_OLOGIC_X1Y197_D1;
  wire [0:0] RIOI3_X105Y197_OLOGIC_X1Y197_OQ;
  wire [0:0] RIOI3_X105Y197_OLOGIC_X1Y197_T1;
  wire [0:0] RIOI3_X105Y197_OLOGIC_X1Y197_TQ;
  wire [0:0] RIOI3_X105Y197_OLOGIC_X1Y198_D1;
  wire [0:0] RIOI3_X105Y197_OLOGIC_X1Y198_OQ;
  wire [0:0] RIOI3_X105Y197_OLOGIC_X1Y198_T1;
  wire [0:0] RIOI3_X105Y197_OLOGIC_X1Y198_TQ;


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y75_SLICE_X0Y75_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y75_SLICE_X0Y75_DO5),
.O6(CLBLL_L_X2Y75_SLICE_X0Y75_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y75_SLICE_X0Y75_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y75_SLICE_X0Y75_CO5),
.O6(CLBLL_L_X2Y75_SLICE_X0Y75_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y75_SLICE_X0Y75_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y75_SLICE_X0Y75_BO5),
.O6(CLBLL_L_X2Y75_SLICE_X0Y75_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0f0f0f0f0f0f0f0f)
  ) CLBLL_L_X2Y75_SLICE_X0Y75_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(LIOB33_X0Y55_IOB_X0Y56_I),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y75_SLICE_X0Y75_AO5),
.O6(CLBLL_L_X2Y75_SLICE_X0Y75_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y75_SLICE_X1Y75_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y75_SLICE_X1Y75_DO5),
.O6(CLBLL_L_X2Y75_SLICE_X1Y75_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y75_SLICE_X1Y75_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y75_SLICE_X1Y75_CO5),
.O6(CLBLL_L_X2Y75_SLICE_X1Y75_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y75_SLICE_X1Y75_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y75_SLICE_X1Y75_BO5),
.O6(CLBLL_L_X2Y75_SLICE_X1Y75_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y75_SLICE_X1Y75_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y75_SLICE_X1Y75_AO5),
.O6(CLBLL_L_X2Y75_SLICE_X1Y75_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y144_SLICE_X0Y144_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y144_SLICE_X0Y144_DO5),
.O6(CLBLL_L_X2Y144_SLICE_X0Y144_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y144_SLICE_X0Y144_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y144_SLICE_X0Y144_CO5),
.O6(CLBLL_L_X2Y144_SLICE_X0Y144_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y144_SLICE_X0Y144_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y144_SLICE_X0Y144_BO5),
.O6(CLBLL_L_X2Y144_SLICE_X0Y144_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y144_SLICE_X0Y144_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y144_SLICE_X0Y144_AO5),
.O6(CLBLL_L_X2Y144_SLICE_X0Y144_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y144_SLICE_X1Y144_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y144_SLICE_X1Y144_DO5),
.O6(CLBLL_L_X2Y144_SLICE_X1Y144_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y144_SLICE_X1Y144_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y144_SLICE_X1Y144_CO5),
.O6(CLBLL_L_X2Y144_SLICE_X1Y144_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y144_SLICE_X1Y144_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y144_SLICE_X1Y144_BO5),
.O6(CLBLL_L_X2Y144_SLICE_X1Y144_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffffffffff77)
  ) CLBLL_L_X2Y144_SLICE_X1Y144_ALUT (
.I0(CLBLM_R_X3Y145_SLICE_X3Y145_CQ),
.I1(CLBLL_L_X2Y146_SLICE_X1Y146_B5Q),
.I2(1'b1),
.I3(CLBLM_R_X3Y144_SLICE_X3Y144_AQ),
.I4(CLBLL_L_X2Y146_SLICE_X0Y146_DQ),
.I5(CLBLM_R_X5Y143_SLICE_X6Y143_D5Q),
.O5(CLBLL_L_X2Y144_SLICE_X1Y144_AO5),
.O6(CLBLL_L_X2Y144_SLICE_X1Y144_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X2Y145_SLICE_X0Y145_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X2Y145_SLICE_X0Y145_AO6),
.Q(CLBLL_L_X2Y145_SLICE_X0Y145_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X2Y145_SLICE_X0Y145_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X2Y145_SLICE_X0Y145_BO6),
.Q(CLBLL_L_X2Y145_SLICE_X0Y145_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y145_SLICE_X0Y145_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y145_SLICE_X0Y145_DO5),
.O6(CLBLL_L_X2Y145_SLICE_X0Y145_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y145_SLICE_X0Y145_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y145_SLICE_X0Y145_CO5),
.O6(CLBLL_L_X2Y145_SLICE_X0Y145_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff300000003000)
  ) CLBLL_L_X2Y145_SLICE_X0Y145_BLUT (
.I0(1'b1),
.I1(CLBLL_L_X2Y146_SLICE_X0Y146_BQ),
.I2(CLBLL_L_X2Y145_SLICE_X0Y145_AQ),
.I3(CLBLL_L_X2Y146_SLICE_X0Y146_AQ),
.I4(LIOB33_X0Y61_IOB_X0Y62_I),
.I5(CLBLM_R_X5Y144_SLICE_X7Y144_B5Q),
.O5(CLBLL_L_X2Y145_SLICE_X0Y145_BO5),
.O6(CLBLL_L_X2Y145_SLICE_X0Y145_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaaffffaaaacf0f)
  ) CLBLL_L_X2Y145_SLICE_X0Y145_ALUT (
.I0(CLBLM_R_X5Y142_SLICE_X6Y142_D5Q),
.I1(CLBLL_L_X2Y146_SLICE_X0Y146_BQ),
.I2(CLBLL_L_X2Y145_SLICE_X0Y145_AQ),
.I3(CLBLL_L_X2Y146_SLICE_X0Y146_AQ),
.I4(LIOB33_X0Y61_IOB_X0Y62_I),
.I5(CLBLM_R_X3Y146_SLICE_X2Y146_CQ),
.O5(CLBLL_L_X2Y145_SLICE_X0Y145_AO5),
.O6(CLBLL_L_X2Y145_SLICE_X0Y145_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X2Y145_SLICE_X1Y145_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X2Y145_SLICE_X1Y145_AO6),
.Q(CLBLL_L_X2Y145_SLICE_X1Y145_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X2Y145_SLICE_X1Y145_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X2Y145_SLICE_X1Y145_BO6),
.Q(CLBLL_L_X2Y145_SLICE_X1Y145_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X2Y145_SLICE_X1Y145_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X2Y145_SLICE_X1Y145_CO6),
.Q(CLBLL_L_X2Y145_SLICE_X1Y145_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hf000000088000000)
  ) CLBLL_L_X2Y145_SLICE_X1Y145_DLUT (
.I0(CLBLL_L_X2Y145_SLICE_X1Y145_BQ),
.I1(CLBLL_L_X2Y145_SLICE_X1Y145_CQ),
.I2(CLBLL_L_X2Y146_SLICE_X1Y146_DO6),
.I3(CLBLL_L_X2Y145_SLICE_X1Y145_AQ),
.I4(CLBLM_R_X3Y146_SLICE_X2Y146_BQ),
.I5(1'b1),
.O5(CLBLL_L_X2Y145_SLICE_X1Y145_DO5),
.O6(CLBLL_L_X2Y145_SLICE_X1Y145_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f0fffff0f0eebb)
  ) CLBLL_L_X2Y145_SLICE_X1Y145_CLUT (
.I0(CLBLL_L_X4Y143_SLICE_X4Y143_D5Q),
.I1(CLBLL_L_X2Y145_SLICE_X1Y145_CQ),
.I2(CLBLL_L_X4Y145_SLICE_X4Y145_C5Q),
.I3(CLBLL_L_X2Y146_SLICE_X1Y146_CO6),
.I4(LIOB33_X0Y61_IOB_X0Y62_I),
.I5(CLBLL_L_X2Y145_SLICE_X1Y145_DO5),
.O5(CLBLL_L_X2Y145_SLICE_X1Y145_CO5),
.O6(CLBLL_L_X2Y145_SLICE_X1Y145_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hc0c5c0cac0c5c0ca)
  ) CLBLL_L_X2Y145_SLICE_X1Y145_BLUT (
.I0(CLBLL_L_X2Y145_SLICE_X1Y145_DO6),
.I1(CLBLL_L_X2Y146_SLICE_X0Y146_AQ),
.I2(LIOB33_X0Y61_IOB_X0Y62_I),
.I3(CLBLL_L_X4Y143_SLICE_X4Y143_D5Q),
.I4(CLBLL_L_X2Y145_SLICE_X1Y145_BQ),
.I5(1'b1),
.O5(CLBLL_L_X2Y145_SLICE_X1Y145_BO5),
.O6(CLBLL_L_X2Y145_SLICE_X1Y145_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff000000780078)
  ) CLBLL_L_X2Y145_SLICE_X1Y145_ALUT (
.I0(CLBLL_L_X2Y146_SLICE_X1Y146_DO6),
.I1(CLBLM_R_X3Y146_SLICE_X2Y146_BQ),
.I2(CLBLL_L_X2Y145_SLICE_X1Y145_AQ),
.I3(CLBLL_L_X4Y143_SLICE_X4Y143_D5Q),
.I4(CLBLM_R_X5Y143_SLICE_X6Y143_C5Q),
.I5(LIOB33_X0Y61_IOB_X0Y62_I),
.O5(CLBLL_L_X2Y145_SLICE_X1Y145_AO5),
.O6(CLBLL_L_X2Y145_SLICE_X1Y145_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X2Y146_SLICE_X0Y146_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X2Y146_SLICE_X0Y146_AO6),
.Q(CLBLL_L_X2Y146_SLICE_X0Y146_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X2Y146_SLICE_X0Y146_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X2Y146_SLICE_X0Y146_BO6),
.Q(CLBLL_L_X2Y146_SLICE_X0Y146_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X2Y146_SLICE_X0Y146_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X2Y146_SLICE_X0Y146_CO6),
.Q(CLBLL_L_X2Y146_SLICE_X0Y146_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X2Y146_SLICE_X0Y146_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X2Y146_SLICE_X0Y146_DO6),
.Q(CLBLL_L_X2Y146_SLICE_X0Y146_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hdccccccc10000000)
  ) CLBLL_L_X2Y146_SLICE_X0Y146_DLUT (
.I0(CLBLM_R_X3Y144_SLICE_X3Y144_AQ),
.I1(LIOB33_X0Y61_IOB_X0Y62_I),
.I2(CLBLL_L_X2Y146_SLICE_X1Y146_B5Q),
.I3(CLBLM_R_X3Y145_SLICE_X3Y145_CQ),
.I4(CLBLM_R_X5Y153_SLICE_X6Y153_B5Q),
.I5(CLBLM_R_X5Y145_SLICE_X6Y145_BQ),
.O5(CLBLL_L_X2Y146_SLICE_X0Y146_DO5),
.O6(CLBLL_L_X2Y146_SLICE_X0Y146_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hcdcccdcc01000100)
  ) CLBLL_L_X2Y146_SLICE_X0Y146_CLUT (
.I0(CLBLL_L_X2Y145_SLICE_X0Y145_AQ),
.I1(LIOB33_X0Y61_IOB_X0Y62_I),
.I2(CLBLL_L_X2Y146_SLICE_X0Y146_AQ),
.I3(CLBLL_L_X2Y146_SLICE_X0Y146_BQ),
.I4(1'b1),
.I5(CLBLL_L_X4Y149_SLICE_X4Y149_D5Q),
.O5(CLBLL_L_X2Y146_SLICE_X0Y146_CO5),
.O6(CLBLL_L_X2Y146_SLICE_X0Y146_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'haabbaaae00110004)
  ) CLBLL_L_X2Y146_SLICE_X0Y146_BLUT (
.I0(LIOB33_X0Y61_IOB_X0Y62_I),
.I1(CLBLL_L_X2Y146_SLICE_X0Y146_BQ),
.I2(CLBLL_L_X2Y146_SLICE_X0Y146_AQ),
.I3(CLBLM_R_X3Y146_SLICE_X2Y146_CQ),
.I4(CLBLL_L_X2Y145_SLICE_X0Y145_AQ),
.I5(CLBLM_R_X3Y147_SLICE_X2Y147_BQ),
.O5(CLBLL_L_X2Y146_SLICE_X0Y146_BO5),
.O6(CLBLL_L_X2Y146_SLICE_X0Y146_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaaaaaa003c0030)
  ) CLBLL_L_X2Y146_SLICE_X0Y146_ALUT (
.I0(CLBLL_L_X4Y146_SLICE_X4Y146_B5Q),
.I1(CLBLL_L_X2Y146_SLICE_X0Y146_BQ),
.I2(CLBLL_L_X2Y146_SLICE_X0Y146_AQ),
.I3(CLBLM_R_X3Y146_SLICE_X2Y146_CQ),
.I4(CLBLL_L_X2Y145_SLICE_X0Y145_AQ),
.I5(LIOB33_X0Y61_IOB_X0Y62_I),
.O5(CLBLL_L_X2Y146_SLICE_X0Y146_AO5),
.O6(CLBLL_L_X2Y146_SLICE_X0Y146_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X2Y146_SLICE_X1Y146_B5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X2Y146_SLICE_X1Y146_BO5),
.Q(CLBLL_L_X2Y146_SLICE_X1Y146_B5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X2Y146_SLICE_X1Y146_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X2Y146_SLICE_X1Y146_AO6),
.Q(CLBLL_L_X2Y146_SLICE_X1Y146_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X2Y146_SLICE_X1Y146_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X2Y146_SLICE_X1Y146_BO6),
.Q(CLBLL_L_X2Y146_SLICE_X1Y146_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h8000000000000000)
  ) CLBLL_L_X2Y146_SLICE_X1Y146_DLUT (
.I0(CLBLL_L_X2Y145_SLICE_X1Y145_CQ),
.I1(CLBLL_L_X4Y149_SLICE_X5Y149_CQ),
.I2(CLBLL_L_X4Y149_SLICE_X4Y149_AQ),
.I3(CLBLM_R_X3Y147_SLICE_X2Y147_CQ),
.I4(CLBLL_L_X2Y146_SLICE_X1Y146_AQ),
.I5(CLBLM_R_X3Y149_SLICE_X2Y149_BQ),
.O5(CLBLL_L_X2Y146_SLICE_X1Y146_DO5),
.O6(CLBLL_L_X2Y146_SLICE_X1Y146_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h7fffffff7f7fffff)
  ) CLBLL_L_X2Y146_SLICE_X1Y146_CLUT (
.I0(CLBLL_L_X2Y146_SLICE_X1Y146_AQ),
.I1(CLBLM_R_X3Y149_SLICE_X2Y149_BQ),
.I2(CLBLL_L_X4Y149_SLICE_X4Y149_AQ),
.I3(CLBLL_L_X4Y149_SLICE_X5Y149_CQ),
.I4(CLBLM_R_X3Y147_SLICE_X2Y147_CQ),
.I5(1'b1),
.O5(CLBLL_L_X2Y146_SLICE_X1Y146_CO5),
.O6(CLBLL_L_X2Y146_SLICE_X1Y146_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hdddd8888f5a0f5a0)
  ) CLBLL_L_X2Y146_SLICE_X1Y146_BLUT (
.I0(LIOB33_X0Y61_IOB_X0Y62_I),
.I1(CLBLM_R_X5Y150_SLICE_X6Y150_AQ),
.I2(CLBLL_L_X4Y147_SLICE_X4Y147_CQ),
.I3(CLBLM_R_X3Y144_SLICE_X2Y144_CO6),
.I4(CLBLL_L_X2Y148_SLICE_X1Y148_AO6),
.I5(1'b1),
.O5(CLBLL_L_X2Y146_SLICE_X1Y146_BO5),
.O6(CLBLL_L_X2Y146_SLICE_X1Y146_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hab01ab01ba10ba10)
  ) CLBLL_L_X2Y146_SLICE_X1Y146_ALUT (
.I0(LIOB33_X0Y61_IOB_X0Y62_I),
.I1(CLBLL_L_X4Y143_SLICE_X4Y143_D5Q),
.I2(CLBLL_L_X2Y146_SLICE_X1Y146_AQ),
.I3(CLBLM_L_X8Y144_SLICE_X11Y144_BQ),
.I4(1'b1),
.I5(CLBLL_L_X4Y149_SLICE_X5Y149_CQ),
.O5(CLBLL_L_X2Y146_SLICE_X1Y146_AO5),
.O6(CLBLL_L_X2Y146_SLICE_X1Y146_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y147_SLICE_X0Y147_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y147_SLICE_X0Y147_DO5),
.O6(CLBLL_L_X2Y147_SLICE_X0Y147_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y147_SLICE_X0Y147_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y147_SLICE_X0Y147_CO5),
.O6(CLBLL_L_X2Y147_SLICE_X0Y147_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y147_SLICE_X0Y147_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y147_SLICE_X0Y147_BO5),
.O6(CLBLL_L_X2Y147_SLICE_X0Y147_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y147_SLICE_X0Y147_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y147_SLICE_X0Y147_AO5),
.O6(CLBLL_L_X2Y147_SLICE_X0Y147_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y147_SLICE_X1Y147_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y147_SLICE_X1Y147_DO5),
.O6(CLBLL_L_X2Y147_SLICE_X1Y147_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y147_SLICE_X1Y147_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y147_SLICE_X1Y147_CO5),
.O6(CLBLL_L_X2Y147_SLICE_X1Y147_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y147_SLICE_X1Y147_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y147_SLICE_X1Y147_BO5),
.O6(CLBLL_L_X2Y147_SLICE_X1Y147_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h00000000cccccccc)
  ) CLBLL_L_X2Y147_SLICE_X1Y147_ALUT (
.I0(1'b1),
.I1(CLBLM_R_X5Y147_SLICE_X7Y147_BQ),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(CLBLL_L_X4Y147_SLICE_X4Y147_C5Q),
.O5(CLBLL_L_X2Y147_SLICE_X1Y147_AO5),
.O6(CLBLL_L_X2Y147_SLICE_X1Y147_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X2Y148_SLICE_X0Y148_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(LIOB33_X0Y61_IOB_X0Y62_I),
.D(CLBLM_R_X3Y145_SLICE_X3Y145_CQ),
.Q(CLBLL_L_X2Y148_SLICE_X0Y148_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y148_SLICE_X0Y148_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y148_SLICE_X0Y148_DO5),
.O6(CLBLL_L_X2Y148_SLICE_X0Y148_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y148_SLICE_X0Y148_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y148_SLICE_X0Y148_CO5),
.O6(CLBLL_L_X2Y148_SLICE_X0Y148_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y148_SLICE_X0Y148_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y148_SLICE_X0Y148_BO5),
.O6(CLBLL_L_X2Y148_SLICE_X0Y148_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y148_SLICE_X0Y148_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y148_SLICE_X0Y148_AO5),
.O6(CLBLL_L_X2Y148_SLICE_X0Y148_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y148_SLICE_X1Y148_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y148_SLICE_X1Y148_DO5),
.O6(CLBLL_L_X2Y148_SLICE_X1Y148_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000001100000000)
  ) CLBLL_L_X2Y148_SLICE_X1Y148_CLUT (
.I0(CLBLL_L_X2Y146_SLICE_X1Y146_B5Q),
.I1(CLBLL_L_X4Y148_SLICE_X5Y148_BQ),
.I2(1'b1),
.I3(CLBLM_R_X3Y145_SLICE_X3Y145_CQ),
.I4(CLBLM_R_X3Y144_SLICE_X3Y144_AQ),
.I5(CLBLM_R_X5Y145_SLICE_X7Y145_CO6),
.O5(CLBLL_L_X2Y148_SLICE_X1Y148_CO5),
.O6(CLBLL_L_X2Y148_SLICE_X1Y148_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h6aaaaaaaaaaaaaaa)
  ) CLBLL_L_X2Y148_SLICE_X1Y148_BLUT (
.I0(LIOB33_X0Y55_IOB_X0Y55_I),
.I1(CLBLM_R_X3Y148_SLICE_X2Y148_BQ),
.I2(CLBLL_L_X4Y149_SLICE_X4Y149_D5Q),
.I3(CLBLL_L_X2Y146_SLICE_X1Y146_BQ),
.I4(CLBLM_R_X3Y149_SLICE_X2Y149_DQ),
.I5(CLBLL_L_X4Y149_SLICE_X4Y149_DQ),
.O5(CLBLL_L_X2Y148_SLICE_X1Y148_BO5),
.O6(CLBLL_L_X2Y148_SLICE_X1Y148_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h8ff00ff0ff00ff00)
  ) CLBLL_L_X2Y148_SLICE_X1Y148_ALUT (
.I0(LIOB33_X0Y55_IOB_X0Y55_I),
.I1(CLBLM_R_X3Y148_SLICE_X2Y148_BQ),
.I2(CLBLL_L_X4Y149_SLICE_X4Y149_D5Q),
.I3(CLBLL_L_X2Y146_SLICE_X1Y146_BQ),
.I4(CLBLM_R_X3Y149_SLICE_X2Y149_DQ),
.I5(CLBLL_L_X4Y149_SLICE_X4Y149_DQ),
.O5(CLBLL_L_X2Y148_SLICE_X1Y148_AO5),
.O6(CLBLL_L_X2Y148_SLICE_X1Y148_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y150_SLICE_X0Y150_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y150_SLICE_X0Y150_DO5),
.O6(CLBLL_L_X2Y150_SLICE_X0Y150_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y150_SLICE_X0Y150_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y150_SLICE_X0Y150_CO5),
.O6(CLBLL_L_X2Y150_SLICE_X0Y150_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y150_SLICE_X0Y150_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y150_SLICE_X0Y150_BO5),
.O6(CLBLL_L_X2Y150_SLICE_X0Y150_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y150_SLICE_X0Y150_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y150_SLICE_X0Y150_AO5),
.O6(CLBLL_L_X2Y150_SLICE_X0Y150_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X2Y150_SLICE_X1Y150_A_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLL_L_X2Y150_SLICE_X1Y150_AO6),
.Q(CLBLL_L_X2Y150_SLICE_X1Y150_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y150_SLICE_X1Y150_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y150_SLICE_X1Y150_DO5),
.O6(CLBLL_L_X2Y150_SLICE_X1Y150_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y150_SLICE_X1Y150_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y150_SLICE_X1Y150_CO5),
.O6(CLBLL_L_X2Y150_SLICE_X1Y150_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y150_SLICE_X1Y150_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y150_SLICE_X1Y150_BO5),
.O6(CLBLL_L_X2Y150_SLICE_X1Y150_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffbbffbb55115511)
  ) CLBLL_L_X2Y150_SLICE_X1Y150_ALUT (
.I0(LIOB33_X0Y61_IOB_X0Y62_I),
.I1(CLBLL_L_X4Y146_SLICE_X5Y146_BQ),
.I2(1'b1),
.I3(CLBLL_L_X4Y150_SLICE_X4Y150_DO6),
.I4(1'b1),
.I5(CLBLM_R_X5Y153_SLICE_X6Y153_DQ),
.O5(CLBLL_L_X2Y150_SLICE_X1Y150_AO5),
.O6(CLBLL_L_X2Y150_SLICE_X1Y150_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y166_SLICE_X0Y166_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y166_SLICE_X0Y166_DO5),
.O6(CLBLL_L_X2Y166_SLICE_X0Y166_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y166_SLICE_X0Y166_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y166_SLICE_X0Y166_CO5),
.O6(CLBLL_L_X2Y166_SLICE_X0Y166_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y166_SLICE_X0Y166_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y166_SLICE_X0Y166_BO5),
.O6(CLBLL_L_X2Y166_SLICE_X0Y166_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0f0f0f0f0f0f0f0f)
  ) CLBLL_L_X2Y166_SLICE_X0Y166_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(CLBLM_L_X12Y146_SLICE_X17Y146_AQ),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y166_SLICE_X0Y166_AO5),
.O6(CLBLL_L_X2Y166_SLICE_X0Y166_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y166_SLICE_X1Y166_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y166_SLICE_X1Y166_DO5),
.O6(CLBLL_L_X2Y166_SLICE_X1Y166_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y166_SLICE_X1Y166_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y166_SLICE_X1Y166_CO5),
.O6(CLBLL_L_X2Y166_SLICE_X1Y166_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y166_SLICE_X1Y166_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y166_SLICE_X1Y166_BO5),
.O6(CLBLL_L_X2Y166_SLICE_X1Y166_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y166_SLICE_X1Y166_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y166_SLICE_X1Y166_AO5),
.O6(CLBLL_L_X2Y166_SLICE_X1Y166_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y140_SLICE_X4Y140_A5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y140_SLICE_X4Y140_BO6),
.Q(CLBLL_L_X4Y140_SLICE_X4Y140_A5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y140_SLICE_X4Y140_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y140_SLICE_X4Y140_AO6),
.Q(CLBLL_L_X4Y140_SLICE_X4Y140_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X4Y140_SLICE_X4Y140_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y140_SLICE_X4Y140_DO5),
.O6(CLBLL_L_X4Y140_SLICE_X4Y140_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0f0f00000f0f0000)
  ) CLBLL_L_X4Y140_SLICE_X4Y140_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(CLBLL_L_X4Y140_SLICE_X5Y140_DO6),
.I3(1'b1),
.I4(LIOB33_X0Y53_IOB_X0Y54_I),
.I5(1'b1),
.O5(CLBLL_L_X4Y140_SLICE_X4Y140_CO5),
.O6(CLBLL_L_X4Y140_SLICE_X4Y140_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf707f80855555555)
  ) CLBLL_L_X4Y140_SLICE_X4Y140_BLUT (
.I0(LIOB33_X0Y59_IOB_X0Y60_I),
.I1(CLBLL_L_X4Y142_SLICE_X4Y142_CQ),
.I2(LIOB33_X0Y61_IOB_X0Y62_I),
.I3(CLBLM_R_X3Y149_SLICE_X3Y149_D5Q),
.I4(CLBLL_L_X4Y140_SLICE_X4Y140_A5Q),
.I5(1'b1),
.O5(CLBLL_L_X4Y140_SLICE_X4Y140_BO5),
.O6(CLBLL_L_X4Y140_SLICE_X4Y140_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hcc0fcc0fcc00cc00)
  ) CLBLL_L_X4Y140_SLICE_X4Y140_ALUT (
.I0(1'b1),
.I1(CLBLL_L_X4Y148_SLICE_X4Y148_AQ),
.I2(CLBLL_L_X4Y140_SLICE_X4Y140_AQ),
.I3(LIOB33_X0Y61_IOB_X0Y62_I),
.I4(1'b1),
.I5(CLBLL_L_X4Y140_SLICE_X4Y140_CO6),
.O5(CLBLL_L_X4Y140_SLICE_X4Y140_AO5),
.O6(CLBLL_L_X4Y140_SLICE_X4Y140_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y140_SLICE_X5Y140_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y140_SLICE_X5Y140_AO6),
.Q(CLBLL_L_X4Y140_SLICE_X5Y140_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y140_SLICE_X5Y140_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y140_SLICE_X5Y140_BO6),
.Q(CLBLL_L_X4Y140_SLICE_X5Y140_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h8000000000000000)
  ) CLBLL_L_X4Y140_SLICE_X5Y140_DLUT (
.I0(CLBLL_L_X4Y140_SLICE_X4Y140_AQ),
.I1(CLBLM_R_X5Y140_SLICE_X6Y140_BQ),
.I2(CLBLL_L_X4Y140_SLICE_X5Y140_BQ),
.I3(CLBLM_R_X5Y140_SLICE_X6Y140_CQ),
.I4(CLBLL_L_X4Y140_SLICE_X5Y140_AQ),
.I5(CLBLM_R_X5Y140_SLICE_X6Y140_AQ),
.O5(CLBLL_L_X4Y140_SLICE_X5Y140_DO5),
.O6(CLBLL_L_X4Y140_SLICE_X5Y140_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h8080000080000000)
  ) CLBLL_L_X4Y140_SLICE_X5Y140_CLUT (
.I0(CLBLL_L_X4Y140_SLICE_X4Y140_AQ),
.I1(CLBLM_R_X5Y140_SLICE_X6Y140_BQ),
.I2(CLBLM_R_X5Y140_SLICE_X6Y140_CQ),
.I3(CLBLL_L_X4Y140_SLICE_X5Y140_BQ),
.I4(CLBLM_R_X5Y140_SLICE_X6Y140_AQ),
.I5(1'b1),
.O5(CLBLL_L_X4Y140_SLICE_X5Y140_CO5),
.O6(CLBLL_L_X4Y140_SLICE_X5Y140_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'haaee0044eeaa4400)
  ) CLBLL_L_X4Y140_SLICE_X5Y140_BLUT (
.I0(LIOB33_X0Y61_IOB_X0Y62_I),
.I1(LIOB33_X0Y53_IOB_X0Y54_I),
.I2(1'b1),
.I3(CLBLL_L_X4Y140_SLICE_X5Y140_BQ),
.I4(CLBLL_L_X4Y140_SLICE_X4Y140_AQ),
.I5(CLBLL_L_X4Y140_SLICE_X5Y140_CO6),
.O5(CLBLL_L_X4Y140_SLICE_X5Y140_BO5),
.O6(CLBLL_L_X4Y140_SLICE_X5Y140_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h8d8dd8d888888888)
  ) CLBLL_L_X4Y140_SLICE_X5Y140_ALUT (
.I0(LIOB33_X0Y61_IOB_X0Y62_I),
.I1(CLBLM_R_X5Y152_SLICE_X6Y152_AQ),
.I2(CLBLL_L_X4Y140_SLICE_X5Y140_AQ),
.I3(1'b1),
.I4(CLBLL_L_X4Y140_SLICE_X5Y140_CO5),
.I5(LIOB33_X0Y53_IOB_X0Y54_I),
.O5(CLBLL_L_X4Y140_SLICE_X5Y140_AO5),
.O6(CLBLL_L_X4Y140_SLICE_X5Y140_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y142_SLICE_X4Y142_A5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y143_SLICE_X5Y143_CO6),
.Q(CLBLL_L_X4Y142_SLICE_X4Y142_A5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y142_SLICE_X4Y142_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y142_SLICE_X4Y142_AO6),
.Q(CLBLL_L_X4Y142_SLICE_X4Y142_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y142_SLICE_X4Y142_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y142_SLICE_X4Y142_BO6),
.Q(CLBLL_L_X4Y142_SLICE_X4Y142_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y142_SLICE_X4Y142_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y142_SLICE_X4Y142_CO6),
.Q(CLBLL_L_X4Y142_SLICE_X4Y142_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X4Y142_SLICE_X4Y142_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y142_SLICE_X4Y142_DO5),
.O6(CLBLL_L_X4Y142_SLICE_X4Y142_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hff3c003cff3c003c)
  ) CLBLL_L_X4Y142_SLICE_X4Y142_CLUT (
.I0(1'b1),
.I1(CLBLL_L_X4Y142_SLICE_X4Y142_CQ),
.I2(LIOB33_X0Y59_IOB_X0Y60_I),
.I3(LIOB33_X0Y61_IOB_X0Y62_I),
.I4(CLBLM_R_X7Y142_SLICE_X8Y142_DQ),
.I5(1'b1),
.O5(CLBLL_L_X4Y142_SLICE_X4Y142_CO5),
.O6(CLBLL_L_X4Y142_SLICE_X4Y142_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hea40ba10ea40ea40)
  ) CLBLL_L_X4Y142_SLICE_X4Y142_BLUT (
.I0(LIOB33_X0Y61_IOB_X0Y62_I),
.I1(CLBLL_L_X4Y142_SLICE_X4Y142_BQ),
.I2(CLBLM_L_X10Y144_SLICE_X12Y144_AO6),
.I3(CLBLL_L_X4Y143_SLICE_X4Y143_C5Q),
.I4(CLBLM_R_X5Y147_SLICE_X6Y147_AQ),
.I5(CLBLM_R_X3Y142_SLICE_X3Y142_AQ),
.O5(CLBLL_L_X4Y142_SLICE_X4Y142_BO5),
.O6(CLBLL_L_X4Y142_SLICE_X4Y142_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hff00ff004c4ccccc)
  ) CLBLL_L_X4Y142_SLICE_X4Y142_ALUT (
.I0(LIOB33_X0Y59_IOB_X0Y60_I),
.I1(CLBLM_R_X3Y151_SLICE_X2Y151_BO5),
.I2(CLBLL_L_X4Y142_SLICE_X4Y142_CQ),
.I3(CLBLL_L_X4Y144_SLICE_X5Y144_BQ),
.I4(CLBLL_L_X4Y140_SLICE_X4Y140_A5Q),
.I5(LIOB33_X0Y61_IOB_X0Y62_I),
.O5(CLBLL_L_X4Y142_SLICE_X4Y142_AO5),
.O6(CLBLL_L_X4Y142_SLICE_X4Y142_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y142_SLICE_X5Y142_C5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y142_SLICE_X5Y142_CO5),
.Q(CLBLL_L_X4Y142_SLICE_X5Y142_C5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y142_SLICE_X5Y142_D5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y142_SLICE_X5Y142_DO5),
.Q(CLBLL_L_X4Y142_SLICE_X5Y142_D5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y142_SLICE_X5Y142_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y142_SLICE_X5Y142_AO6),
.Q(CLBLL_L_X4Y142_SLICE_X5Y142_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y142_SLICE_X5Y142_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y142_SLICE_X5Y142_BO6),
.Q(CLBLL_L_X4Y142_SLICE_X5Y142_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y142_SLICE_X5Y142_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y142_SLICE_X5Y142_CO6),
.Q(CLBLL_L_X4Y142_SLICE_X5Y142_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y142_SLICE_X5Y142_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y142_SLICE_X5Y142_DO6),
.Q(CLBLL_L_X4Y142_SLICE_X5Y142_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hf5a0f5a0eeee4444)
  ) CLBLL_L_X4Y142_SLICE_X5Y142_DLUT (
.I0(LIOB33_X0Y61_IOB_X0Y62_I),
.I1(CLBLM_R_X7Y142_SLICE_X9Y142_BQ),
.I2(CLBLL_L_X4Y142_SLICE_X5Y142_BQ),
.I3(CLBLL_L_X4Y147_SLICE_X5Y147_CQ),
.I4(CLBLL_L_X4Y148_SLICE_X4Y148_CQ),
.I5(1'b1),
.O5(CLBLL_L_X4Y142_SLICE_X5Y142_DO5),
.O6(CLBLL_L_X4Y142_SLICE_X5Y142_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hfff000f0ccf0ccf0)
  ) CLBLL_L_X4Y142_SLICE_X5Y142_CLUT (
.I0(1'b1),
.I1(CLBLM_R_X5Y140_SLICE_X6Y140_BQ),
.I2(CLBLL_L_X4Y143_SLICE_X4Y143_DQ),
.I3(LIOB33_X0Y61_IOB_X0Y62_I),
.I4(CLBLL_L_X4Y142_SLICE_X4Y142_BQ),
.I5(1'b1),
.O5(CLBLL_L_X4Y142_SLICE_X5Y142_CO5),
.O6(CLBLL_L_X4Y142_SLICE_X5Y142_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hffcaffcc00ca00cc)
  ) CLBLL_L_X4Y142_SLICE_X5Y142_BLUT (
.I0(CLBLL_L_X4Y147_SLICE_X4Y147_BQ),
.I1(CLBLL_L_X4Y142_SLICE_X5Y142_BQ),
.I2(CLBLM_L_X8Y147_SLICE_X10Y147_C5Q),
.I3(LIOB33_X0Y61_IOB_X0Y62_I),
.I4(CLBLM_L_X10Y144_SLICE_X13Y144_CQ),
.I5(CLBLM_L_X12Y145_SLICE_X16Y145_AQ),
.O5(CLBLL_L_X4Y142_SLICE_X5Y142_BO5),
.O6(CLBLL_L_X4Y142_SLICE_X5Y142_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hff00ff00acacaaaa)
  ) CLBLL_L_X4Y142_SLICE_X5Y142_ALUT (
.I0(CLBLL_L_X4Y142_SLICE_X5Y142_AQ),
.I1(CLBLL_L_X4Y143_SLICE_X4Y143_CQ),
.I2(CLBLM_L_X8Y147_SLICE_X10Y147_C5Q),
.I3(CLBLL_L_X4Y140_SLICE_X5Y140_BQ),
.I4(CLBLM_L_X10Y144_SLICE_X13Y144_CQ),
.I5(LIOB33_X0Y61_IOB_X0Y62_I),
.O5(CLBLL_L_X4Y142_SLICE_X5Y142_AO5),
.O6(CLBLL_L_X4Y142_SLICE_X5Y142_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y143_SLICE_X4Y143_A5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y143_SLICE_X2Y143_CO6),
.Q(CLBLL_L_X4Y143_SLICE_X4Y143_A5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "C5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y143_SLICE_X4Y143_C5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y143_SLICE_X4Y143_CO5),
.Q(CLBLL_L_X4Y143_SLICE_X4Y143_C5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y143_SLICE_X4Y143_D5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y143_SLICE_X4Y143_DO5),
.Q(CLBLL_L_X4Y143_SLICE_X4Y143_D5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y143_SLICE_X4Y143_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y143_SLICE_X4Y143_AO6),
.Q(CLBLL_L_X4Y143_SLICE_X4Y143_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y143_SLICE_X4Y143_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y143_SLICE_X4Y143_BO6),
.Q(CLBLL_L_X4Y143_SLICE_X4Y143_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y143_SLICE_X4Y143_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y143_SLICE_X4Y143_CO6),
.Q(CLBLL_L_X4Y143_SLICE_X4Y143_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y143_SLICE_X4Y143_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y143_SLICE_X4Y143_DO6),
.Q(CLBLL_L_X4Y143_SLICE_X4Y143_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hccffcc00f0aaf0aa)
  ) CLBLL_L_X4Y143_SLICE_X4Y143_DLUT (
.I0(CLBLM_R_X7Y149_SLICE_X9Y149_AQ),
.I1(CLBLM_R_X5Y146_SLICE_X7Y146_C5Q),
.I2(CLBLL_L_X4Y143_SLICE_X4Y143_DQ),
.I3(LIOB33_X0Y61_IOB_X0Y62_I),
.I4(CLBLM_R_X5Y141_SLICE_X6Y141_BQ),
.I5(1'b1),
.O5(CLBLL_L_X4Y143_SLICE_X4Y143_DO5),
.O6(CLBLL_L_X4Y143_SLICE_X4Y143_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hfff000f0ccaaccaa)
  ) CLBLL_L_X4Y143_SLICE_X4Y143_CLUT (
.I0(RIOB33_X105Y121_IOB_X1Y122_I),
.I1(CLBLL_L_X4Y143_SLICE_X4Y143_CQ),
.I2(CLBLL_L_X2Y145_SLICE_X1Y145_AQ),
.I3(LIOB33_X0Y61_IOB_X0Y62_I),
.I4(CLBLL_L_X4Y146_SLICE_X4Y146_CQ),
.I5(1'b1),
.O5(CLBLL_L_X4Y143_SLICE_X4Y143_CO5),
.O6(CLBLL_L_X4Y143_SLICE_X4Y143_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hafa3afaccccc0000)
  ) CLBLL_L_X4Y143_SLICE_X4Y143_BLUT (
.I0(CLBLM_R_X5Y143_SLICE_X6Y143_CQ),
.I1(CLBLL_L_X4Y143_SLICE_X4Y143_BQ),
.I2(LIOB33_X0Y61_IOB_X0Y62_I),
.I3(CLBLM_R_X3Y145_SLICE_X2Y145_CQ),
.I4(CLBLM_R_X5Y145_SLICE_X6Y145_D5Q),
.I5(1'b1),
.O5(CLBLL_L_X4Y143_SLICE_X4Y143_BO5),
.O6(CLBLL_L_X4Y143_SLICE_X4Y143_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hcccccccc005a0000)
  ) CLBLL_L_X4Y143_SLICE_X4Y143_ALUT (
.I0(CLBLL_L_X4Y143_SLICE_X4Y143_BO5),
.I1(CLBLM_R_X5Y148_SLICE_X6Y148_BQ),
.I2(CLBLL_L_X4Y143_SLICE_X4Y143_AQ),
.I3(CLBLM_R_X3Y145_SLICE_X2Y145_CQ),
.I4(CLBLL_L_X4Y147_SLICE_X4Y147_AQ),
.I5(LIOB33_X0Y61_IOB_X0Y62_I),
.O5(CLBLL_L_X4Y143_SLICE_X4Y143_AO5),
.O6(CLBLL_L_X4Y143_SLICE_X4Y143_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y143_SLICE_X5Y143_B5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y143_SLICE_X5Y143_BO5),
.Q(CLBLL_L_X4Y143_SLICE_X5Y143_B5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y143_SLICE_X5Y143_D5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y143_SLICE_X5Y143_DO5),
.Q(CLBLL_L_X4Y143_SLICE_X5Y143_D5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y143_SLICE_X5Y143_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y143_SLICE_X5Y143_AO6),
.Q(CLBLL_L_X4Y143_SLICE_X5Y143_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y143_SLICE_X5Y143_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y143_SLICE_X5Y143_BO6),
.Q(CLBLL_L_X4Y143_SLICE_X5Y143_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y143_SLICE_X5Y143_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y143_SLICE_X5Y143_DO6),
.Q(CLBLL_L_X4Y143_SLICE_X5Y143_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hf3c0f3c0ffcc3300)
  ) CLBLL_L_X4Y143_SLICE_X5Y143_DLUT (
.I0(1'b1),
.I1(LIOB33_X0Y61_IOB_X0Y62_I),
.I2(LIOB33_X0Y63_IOB_X0Y63_I),
.I3(CLBLL_L_X4Y151_SLICE_X4Y151_AQ),
.I4(CLBLL_L_X4Y144_SLICE_X5Y144_DQ),
.I5(1'b1),
.O5(CLBLL_L_X4Y143_SLICE_X5Y143_DO5),
.O6(CLBLL_L_X4Y143_SLICE_X5Y143_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0fff00088880000)
  ) CLBLL_L_X4Y143_SLICE_X5Y143_CLUT (
.I0(CLBLL_L_X4Y143_SLICE_X4Y143_AQ),
.I1(CLBLM_R_X5Y145_SLICE_X6Y145_D5Q),
.I2(CLBLL_L_X4Y148_SLICE_X5Y148_DQ),
.I3(LIOB33_X0Y61_IOB_X0Y62_I),
.I4(CLBLL_L_X4Y143_SLICE_X4Y143_BQ),
.I5(1'b1),
.O5(CLBLL_L_X4Y143_SLICE_X5Y143_CO5),
.O6(CLBLL_L_X4Y143_SLICE_X5Y143_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hccccf0f0ff00aaaa)
  ) CLBLL_L_X4Y143_SLICE_X5Y143_BLUT (
.I0(LIOB33_X0Y59_IOB_X0Y59_I),
.I1(CLBLM_R_X5Y144_SLICE_X7Y144_BQ),
.I2(CLBLM_R_X7Y151_SLICE_X8Y151_C5Q),
.I3(CLBLM_R_X5Y143_SLICE_X7Y143_BQ),
.I4(LIOB33_X0Y61_IOB_X0Y62_I),
.I5(1'b1),
.O5(CLBLL_L_X4Y143_SLICE_X5Y143_BO5),
.O6(CLBLL_L_X4Y143_SLICE_X5Y143_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff0000c8fac8fa)
  ) CLBLL_L_X4Y143_SLICE_X5Y143_ALUT (
.I0(CLBLL_L_X4Y144_SLICE_X5Y144_DQ),
.I1(CLBLL_L_X4Y151_SLICE_X4Y151_BQ),
.I2(CLBLL_L_X4Y143_SLICE_X5Y143_AQ),
.I3(CLBLM_R_X3Y145_SLICE_X3Y145_D5Q),
.I4(CLBLL_L_X4Y143_SLICE_X5Y143_B5Q),
.I5(LIOB33_X0Y61_IOB_X0Y62_I),
.O5(CLBLL_L_X4Y143_SLICE_X5Y143_AO5),
.O6(CLBLL_L_X4Y143_SLICE_X5Y143_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y144_SLICE_X4Y144_B5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y144_SLICE_X4Y144_BO5),
.Q(CLBLL_L_X4Y144_SLICE_X4Y144_B5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "C5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y144_SLICE_X4Y144_C5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y144_SLICE_X4Y144_CO5),
.Q(CLBLL_L_X4Y144_SLICE_X4Y144_C5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y144_SLICE_X4Y144_D5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y144_SLICE_X4Y144_DO5),
.Q(CLBLL_L_X4Y144_SLICE_X4Y144_D5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y144_SLICE_X4Y144_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y144_SLICE_X4Y144_AO6),
.Q(CLBLL_L_X4Y144_SLICE_X4Y144_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y144_SLICE_X4Y144_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y144_SLICE_X4Y144_BO6),
.Q(CLBLL_L_X4Y144_SLICE_X4Y144_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y144_SLICE_X4Y144_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y144_SLICE_X4Y144_CO6),
.Q(CLBLL_L_X4Y144_SLICE_X4Y144_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y144_SLICE_X4Y144_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y144_SLICE_X4Y144_DO6),
.Q(CLBLL_L_X4Y144_SLICE_X4Y144_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0fff000aaffaa00)
  ) CLBLL_L_X4Y144_SLICE_X4Y144_DLUT (
.I0(CLBLL_L_X4Y140_SLICE_X5Y140_AQ),
.I1(1'b1),
.I2(CLBLM_R_X3Y146_SLICE_X2Y146_CQ),
.I3(LIOB33_X0Y61_IOB_X0Y62_I),
.I4(CLBLM_L_X12Y151_SLICE_X16Y151_AQ),
.I5(1'b1),
.O5(CLBLL_L_X4Y144_SLICE_X4Y144_DO5),
.O6(CLBLL_L_X4Y144_SLICE_X4Y144_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'haaffaa00f0ccf0cc)
  ) CLBLL_L_X4Y144_SLICE_X4Y144_CLUT (
.I0(CLBLM_L_X8Y145_SLICE_X11Y145_C5Q),
.I1(CLBLL_L_X4Y144_SLICE_X5Y144_BQ),
.I2(CLBLL_L_X4Y147_SLICE_X4Y147_BQ),
.I3(LIOB33_X0Y61_IOB_X0Y62_I),
.I4(CLBLL_L_X4Y147_SLICE_X5Y147_B5Q),
.I5(1'b1),
.O5(CLBLL_L_X4Y144_SLICE_X4Y144_CO5),
.O6(CLBLL_L_X4Y144_SLICE_X4Y144_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0ccf0ccaa33aacc)
  ) CLBLL_L_X4Y144_SLICE_X4Y144_BLUT (
.I0(CLBLM_R_X5Y145_SLICE_X6Y145_B5Q),
.I1(CLBLL_L_X4Y150_SLICE_X4Y150_B5Q),
.I2(CLBLL_L_X4Y144_SLICE_X4Y144_CQ),
.I3(LIOB33_X0Y61_IOB_X0Y62_I),
.I4(CLBLM_R_X5Y144_SLICE_X7Y144_BQ),
.I5(1'b1),
.O5(CLBLL_L_X4Y144_SLICE_X4Y144_BO5),
.O6(CLBLL_L_X4Y144_SLICE_X4Y144_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaaaaaaccf0cccc)
  ) CLBLL_L_X4Y144_SLICE_X4Y144_ALUT (
.I0(CLBLL_L_X2Y145_SLICE_X0Y145_BQ),
.I1(CLBLL_L_X4Y144_SLICE_X4Y144_BQ),
.I2(CLBLL_L_X4Y144_SLICE_X4Y144_AQ),
.I3(CLBLM_R_X7Y152_SLICE_X8Y152_D5Q),
.I4(CLBLM_R_X7Y142_SLICE_X8Y142_C5Q),
.I5(LIOB33_X0Y61_IOB_X0Y62_I),
.O5(CLBLL_L_X4Y144_SLICE_X4Y144_AO5),
.O6(CLBLL_L_X4Y144_SLICE_X4Y144_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y144_SLICE_X5Y144_D5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y144_SLICE_X5Y144_DO5),
.Q(CLBLL_L_X4Y144_SLICE_X5Y144_D5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y144_SLICE_X5Y144_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y144_SLICE_X5Y144_AO6),
.Q(CLBLL_L_X4Y144_SLICE_X5Y144_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y144_SLICE_X5Y144_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y144_SLICE_X5Y144_BO6),
.Q(CLBLL_L_X4Y144_SLICE_X5Y144_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y144_SLICE_X5Y144_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y144_SLICE_X5Y144_CO6),
.Q(CLBLL_L_X4Y144_SLICE_X5Y144_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y144_SLICE_X5Y144_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y144_SLICE_X5Y144_DO6),
.Q(CLBLL_L_X4Y144_SLICE_X5Y144_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hbb88bb88ffcc3300)
  ) CLBLL_L_X4Y144_SLICE_X5Y144_DLUT (
.I0(CLBLM_L_X10Y145_SLICE_X12Y145_AQ),
.I1(LIOB33_X0Y61_IOB_X0Y62_I),
.I2(1'b1),
.I3(CLBLL_L_X4Y145_SLICE_X5Y145_BQ),
.I4(CLBLL_L_X4Y144_SLICE_X5Y144_AQ),
.I5(1'b1),
.O5(CLBLL_L_X4Y144_SLICE_X5Y144_DO5),
.O6(CLBLL_L_X4Y144_SLICE_X5Y144_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff443400004434)
  ) CLBLL_L_X4Y144_SLICE_X5Y144_CLUT (
.I0(CLBLL_L_X4Y147_SLICE_X5Y147_BQ),
.I1(CLBLL_L_X4Y144_SLICE_X5Y144_CQ),
.I2(CLBLM_R_X5Y145_SLICE_X6Y145_B5Q),
.I3(CLBLM_R_X11Y146_SLICE_X15Y146_AO6),
.I4(LIOB33_X0Y61_IOB_X0Y62_I),
.I5(CLBLM_R_X3Y145_SLICE_X3Y145_D5Q),
.O5(CLBLL_L_X4Y144_SLICE_X5Y144_CO5),
.O6(CLBLL_L_X4Y144_SLICE_X5Y144_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff0000f444f444)
  ) CLBLL_L_X4Y144_SLICE_X5Y144_BLUT (
.I0(CLBLM_R_X11Y146_SLICE_X15Y146_AO6),
.I1(CLBLL_L_X4Y152_SLICE_X4Y152_B5Q),
.I2(CLBLL_L_X4Y147_SLICE_X5Y147_BQ),
.I3(CLBLL_L_X4Y144_SLICE_X5Y144_CQ),
.I4(CLBLM_L_X8Y148_SLICE_X11Y148_AQ),
.I5(LIOB33_X0Y61_IOB_X0Y62_I),
.O5(CLBLL_L_X4Y144_SLICE_X5Y144_BO5),
.O6(CLBLL_L_X4Y144_SLICE_X5Y144_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hff00ff00fcfc5454)
  ) CLBLL_L_X4Y144_SLICE_X5Y144_ALUT (
.I0(CLBLL_L_X4Y142_SLICE_X5Y142_DQ),
.I1(CLBLL_L_X4Y148_SLICE_X5Y148_DQ),
.I2(CLBLL_L_X4Y144_SLICE_X5Y144_AQ),
.I3(CLBLL_L_X4Y142_SLICE_X5Y142_D5Q),
.I4(CLBLL_L_X4Y147_SLICE_X5Y147_CQ),
.I5(LIOB33_X0Y61_IOB_X0Y62_I),
.O5(CLBLL_L_X4Y144_SLICE_X5Y144_AO5),
.O6(CLBLL_L_X4Y144_SLICE_X5Y144_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y145_SLICE_X4Y145_B5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y145_SLICE_X4Y145_BO5),
.Q(CLBLL_L_X4Y145_SLICE_X4Y145_B5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "C5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y145_SLICE_X4Y145_C5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y145_SLICE_X4Y145_CO5),
.Q(CLBLL_L_X4Y145_SLICE_X4Y145_C5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y145_SLICE_X4Y145_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y145_SLICE_X4Y145_AO6),
.Q(CLBLL_L_X4Y145_SLICE_X4Y145_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y145_SLICE_X4Y145_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y145_SLICE_X4Y145_BO6),
.Q(CLBLL_L_X4Y145_SLICE_X4Y145_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y145_SLICE_X4Y145_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y145_SLICE_X4Y145_CO6),
.Q(CLBLL_L_X4Y145_SLICE_X4Y145_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h7fffffff7f7f7f7f)
  ) CLBLL_L_X4Y145_SLICE_X4Y145_DLUT (
.I0(CLBLL_L_X4Y143_SLICE_X4Y143_AQ),
.I1(CLBLL_L_X4Y151_SLICE_X4Y151_AQ),
.I2(CLBLL_L_X4Y151_SLICE_X5Y151_CQ),
.I3(CLBLM_R_X5Y145_SLICE_X6Y145_D5Q),
.I4(CLBLL_L_X4Y143_SLICE_X4Y143_BQ),
.I5(1'b1),
.O5(CLBLL_L_X4Y145_SLICE_X4Y145_DO5),
.O6(CLBLL_L_X4Y145_SLICE_X4Y145_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0fff000ccaaccaa)
  ) CLBLL_L_X4Y145_SLICE_X4Y145_CLUT (
.I0(CLBLM_R_X3Y148_SLICE_X2Y148_A5Q),
.I1(CLBLL_L_X4Y145_SLICE_X4Y145_CQ),
.I2(CLBLM_R_X5Y148_SLICE_X6Y148_CQ),
.I3(LIOB33_X0Y61_IOB_X0Y62_I),
.I4(CLBLM_L_X10Y153_SLICE_X13Y153_A5Q),
.I5(1'b1),
.O5(CLBLL_L_X4Y145_SLICE_X4Y145_CO5),
.O6(CLBLL_L_X4Y145_SLICE_X4Y145_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'he2e2e2e2ee22ee22)
  ) CLBLL_L_X4Y145_SLICE_X4Y145_BLUT (
.I0(CLBLL_L_X4Y151_SLICE_X5Y151_CQ),
.I1(LIOB33_X0Y61_IOB_X0Y62_I),
.I2(CLBLL_L_X4Y146_SLICE_X4Y146_AQ),
.I3(CLBLM_R_X5Y141_SLICE_X6Y141_B5Q),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y145_SLICE_X4Y145_BO5),
.O6(CLBLL_L_X4Y145_SLICE_X4Y145_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfefe5454aafe0054)
  ) CLBLL_L_X4Y145_SLICE_X4Y145_ALUT (
.I0(LIOB33_X0Y61_IOB_X0Y62_I),
.I1(CLBLL_L_X4Y145_SLICE_X4Y145_BQ),
.I2(CLBLL_L_X4Y145_SLICE_X4Y145_AQ),
.I3(CLBLM_R_X7Y142_SLICE_X8Y142_C5Q),
.I4(CLBLM_L_X8Y149_SLICE_X11Y149_AQ),
.I5(CLBLM_R_X7Y152_SLICE_X8Y152_D5Q),
.O5(CLBLL_L_X4Y145_SLICE_X4Y145_AO5),
.O6(CLBLL_L_X4Y145_SLICE_X4Y145_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y145_SLICE_X5Y145_C5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y145_SLICE_X5Y145_CO5),
.Q(CLBLL_L_X4Y145_SLICE_X5Y145_C5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y145_SLICE_X5Y145_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y145_SLICE_X5Y145_AO6),
.Q(CLBLL_L_X4Y145_SLICE_X5Y145_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y145_SLICE_X5Y145_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y145_SLICE_X5Y145_BO6),
.Q(CLBLL_L_X4Y145_SLICE_X5Y145_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y145_SLICE_X5Y145_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y145_SLICE_X5Y145_CO6),
.Q(CLBLL_L_X4Y145_SLICE_X5Y145_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h8000000000000000)
  ) CLBLL_L_X4Y145_SLICE_X5Y145_DLUT (
.I0(CLBLM_R_X3Y145_SLICE_X3Y145_BQ),
.I1(CLBLM_R_X5Y152_SLICE_X6Y152_DQ),
.I2(CLBLL_L_X4Y151_SLICE_X5Y151_CQ),
.I3(CLBLL_L_X4Y143_SLICE_X5Y143_CO5),
.I4(CLBLM_R_X5Y152_SLICE_X6Y152_CQ),
.I5(CLBLL_L_X4Y151_SLICE_X4Y151_AQ),
.O5(CLBLL_L_X4Y145_SLICE_X5Y145_DO5),
.O6(CLBLL_L_X4Y145_SLICE_X5Y145_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'haaccaaccfff000f0)
  ) CLBLL_L_X4Y145_SLICE_X5Y145_CLUT (
.I0(CLBLM_R_X5Y147_SLICE_X6Y147_C5Q),
.I1(CLBLL_L_X4Y145_SLICE_X4Y145_C5Q),
.I2(CLBLM_R_X5Y146_SLICE_X7Y146_DQ),
.I3(LIOB33_X0Y61_IOB_X0Y62_I),
.I4(CLBLM_R_X7Y153_SLICE_X9Y153_CQ),
.I5(1'b1),
.O5(CLBLL_L_X4Y145_SLICE_X5Y145_CO5),
.O6(CLBLL_L_X4Y145_SLICE_X5Y145_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hff00ff00ffffe0e0)
  ) CLBLL_L_X4Y145_SLICE_X5Y145_BLUT (
.I0(CLBLL_L_X4Y145_SLICE_X5Y145_DO6),
.I1(CLBLL_L_X4Y145_SLICE_X5Y145_BQ),
.I2(CLBLL_L_X4Y147_SLICE_X5Y147_DO6),
.I3(CLBLM_R_X5Y145_SLICE_X7Y145_AQ),
.I4(CLBLM_R_X3Y145_SLICE_X2Y145_CQ),
.I5(LIOB33_X0Y61_IOB_X0Y62_I),
.O5(CLBLL_L_X4Y145_SLICE_X5Y145_BO5),
.O6(CLBLL_L_X4Y145_SLICE_X5Y145_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hff00ff00f0f0b8b8)
  ) CLBLL_L_X4Y145_SLICE_X5Y145_ALUT (
.I0(CLBLM_R_X3Y146_SLICE_X2Y146_DQ),
.I1(CLBLM_L_X10Y144_SLICE_X13Y144_CQ),
.I2(CLBLL_L_X4Y145_SLICE_X5Y145_AQ),
.I3(CLBLM_R_X7Y145_SLICE_X8Y145_C5Q),
.I4(CLBLM_L_X8Y147_SLICE_X10Y147_C5Q),
.I5(LIOB33_X0Y61_IOB_X0Y62_I),
.O5(CLBLL_L_X4Y145_SLICE_X5Y145_AO5),
.O6(CLBLL_L_X4Y145_SLICE_X5Y145_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y146_SLICE_X4Y146_B5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y146_SLICE_X4Y146_BO5),
.Q(CLBLL_L_X4Y146_SLICE_X4Y146_B5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "C5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y146_SLICE_X4Y146_C5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y146_SLICE_X4Y146_CO5),
.Q(CLBLL_L_X4Y146_SLICE_X4Y146_C5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y146_SLICE_X4Y146_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y146_SLICE_X4Y146_AO6),
.Q(CLBLL_L_X4Y146_SLICE_X4Y146_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y146_SLICE_X4Y146_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y146_SLICE_X4Y146_BO6),
.Q(CLBLL_L_X4Y146_SLICE_X4Y146_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y146_SLICE_X4Y146_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y146_SLICE_X4Y146_CO6),
.Q(CLBLL_L_X4Y146_SLICE_X4Y146_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h880088005ff5affa)
  ) CLBLL_L_X4Y146_SLICE_X4Y146_DLUT (
.I0(CLBLL_L_X2Y146_SLICE_X1Y146_AQ),
.I1(CLBLL_L_X4Y149_SLICE_X5Y149_CQ),
.I2(CLBLM_R_X7Y144_SLICE_X8Y144_DQ),
.I3(CLBLM_R_X3Y147_SLICE_X2Y147_CQ),
.I4(CLBLM_R_X5Y146_SLICE_X7Y146_C5Q),
.I5(1'b1),
.O5(CLBLL_L_X4Y146_SLICE_X4Y146_DO5),
.O6(CLBLL_L_X4Y146_SLICE_X4Y146_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'ha0f5a0f5fafa5050)
  ) CLBLL_L_X4Y146_SLICE_X4Y146_CLUT (
.I0(LIOB33_X0Y61_IOB_X0Y62_I),
.I1(1'b1),
.I2(CLBLM_R_X3Y147_SLICE_X3Y147_C5Q),
.I3(CLBLM_L_X12Y151_SLICE_X16Y151_AQ),
.I4(CLBLM_R_X3Y149_SLICE_X3Y149_CQ),
.I5(1'b1),
.O5(CLBLL_L_X4Y146_SLICE_X4Y146_CO5),
.O6(CLBLL_L_X4Y146_SLICE_X4Y146_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f0aaaaff006666)
  ) CLBLL_L_X4Y146_SLICE_X4Y146_BLUT (
.I0(CLBLM_R_X3Y151_SLICE_X3Y151_AQ),
.I1(CLBLL_L_X4Y145_SLICE_X4Y145_CQ),
.I2(CLBLM_R_X3Y147_SLICE_X2Y147_AQ),
.I3(CLBLL_L_X4Y144_SLICE_X4Y144_D5Q),
.I4(LIOB33_X0Y61_IOB_X0Y62_I),
.I5(1'b1),
.O5(CLBLL_L_X4Y146_SLICE_X4Y146_BO5),
.O6(CLBLL_L_X4Y146_SLICE_X4Y146_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaaccffaaaac0f0)
  ) CLBLL_L_X4Y146_SLICE_X4Y146_ALUT (
.I0(CLBLL_L_X4Y144_SLICE_X4Y144_DQ),
.I1(CLBLM_L_X10Y145_SLICE_X12Y145_AQ),
.I2(CLBLL_L_X4Y146_SLICE_X4Y146_AQ),
.I3(CLBLM_R_X5Y142_SLICE_X7Y142_BQ),
.I4(LIOB33_X0Y61_IOB_X0Y62_I),
.I5(CLBLL_L_X4Y149_SLICE_X4Y149_BQ),
.O5(CLBLL_L_X4Y146_SLICE_X4Y146_AO5),
.O6(CLBLL_L_X4Y146_SLICE_X4Y146_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y146_SLICE_X5Y146_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y146_SLICE_X5Y146_AO6),
.Q(CLBLL_L_X4Y146_SLICE_X5Y146_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y146_SLICE_X5Y146_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y146_SLICE_X5Y146_BO6),
.Q(CLBLL_L_X4Y146_SLICE_X5Y146_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y146_SLICE_X5Y146_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y146_SLICE_X5Y146_CO6),
.Q(CLBLL_L_X4Y146_SLICE_X5Y146_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y146_SLICE_X5Y146_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y146_SLICE_X5Y146_DO6),
.Q(CLBLL_L_X4Y146_SLICE_X5Y146_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hefabffaa45015500)
  ) CLBLL_L_X4Y146_SLICE_X5Y146_DLUT (
.I0(LIOB33_X0Y61_IOB_X0Y62_I),
.I1(CLBLL_L_X4Y142_SLICE_X4Y142_AQ),
.I2(CLBLM_L_X10Y151_SLICE_X13Y151_AQ),
.I3(CLBLL_L_X4Y148_SLICE_X4Y148_AQ),
.I4(CLBLM_R_X3Y143_SLICE_X3Y143_BQ),
.I5(CLBLL_L_X4Y146_SLICE_X5Y146_CQ),
.O5(CLBLL_L_X4Y146_SLICE_X5Y146_DO5),
.O6(CLBLL_L_X4Y146_SLICE_X5Y146_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h888888888d8d8888)
  ) CLBLL_L_X4Y146_SLICE_X5Y146_CLUT (
.I0(LIOB33_X0Y61_IOB_X0Y62_I),
.I1(CLBLM_L_X8Y142_SLICE_X10Y142_CQ),
.I2(CLBLL_L_X4Y153_SLICE_X4Y153_AQ),
.I3(1'b1),
.I4(CLBLL_L_X4Y146_SLICE_X5Y146_AQ),
.I5(CLBLL_L_X4Y146_SLICE_X5Y146_CQ),
.O5(CLBLL_L_X4Y146_SLICE_X5Y146_CO5),
.O6(CLBLL_L_X4Y146_SLICE_X5Y146_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f3f0f000030000)
  ) CLBLL_L_X4Y146_SLICE_X5Y146_BLUT (
.I0(1'b1),
.I1(CLBLL_L_X4Y145_SLICE_X4Y145_DO5),
.I2(LIOB33_X0Y61_IOB_X0Y62_I),
.I3(CLBLM_R_X5Y145_SLICE_X6Y145_D5Q),
.I4(CLBLL_L_X4Y143_SLICE_X4Y143_BQ),
.I5(CLBLL_L_X4Y146_SLICE_X5Y146_DQ),
.O5(CLBLL_L_X4Y146_SLICE_X5Y146_BO5),
.O6(CLBLL_L_X4Y146_SLICE_X5Y146_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'heeef222300500050)
  ) CLBLL_L_X4Y146_SLICE_X5Y146_ALUT (
.I0(CLBLL_L_X4Y153_SLICE_X4Y153_AQ),
.I1(LIOB33_X0Y61_IOB_X0Y62_I),
.I2(CLBLL_L_X4Y146_SLICE_X5Y146_AQ),
.I3(CLBLL_L_X4Y146_SLICE_X5Y146_CQ),
.I4(CLBLM_L_X8Y146_SLICE_X11Y146_C5Q),
.I5(1'b1),
.O5(CLBLL_L_X4Y146_SLICE_X5Y146_AO5),
.O6(CLBLL_L_X4Y146_SLICE_X5Y146_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y147_SLICE_X4Y147_B5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y147_SLICE_X4Y147_BO5),
.Q(CLBLL_L_X4Y147_SLICE_X4Y147_B5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "C5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y147_SLICE_X4Y147_C5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y147_SLICE_X4Y147_CO5),
.Q(CLBLL_L_X4Y147_SLICE_X4Y147_C5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y147_SLICE_X4Y147_D5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y147_SLICE_X4Y147_DO5),
.Q(CLBLL_L_X4Y147_SLICE_X4Y147_D5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y147_SLICE_X4Y147_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y147_SLICE_X4Y147_AO6),
.Q(CLBLL_L_X4Y147_SLICE_X4Y147_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y147_SLICE_X4Y147_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y147_SLICE_X4Y147_BO6),
.Q(CLBLL_L_X4Y147_SLICE_X4Y147_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y147_SLICE_X4Y147_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y147_SLICE_X4Y147_CO6),
.Q(CLBLL_L_X4Y147_SLICE_X4Y147_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y147_SLICE_X4Y147_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y147_SLICE_X4Y147_DO6),
.Q(CLBLL_L_X4Y147_SLICE_X4Y147_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hff00eeeef0f0ff00)
  ) CLBLL_L_X4Y147_SLICE_X4Y147_DLUT (
.I0(CLBLM_R_X3Y146_SLICE_X3Y146_AQ),
.I1(CLBLM_R_X7Y153_SLICE_X9Y153_DQ),
.I2(CLBLL_L_X4Y144_SLICE_X4Y144_AQ),
.I3(CLBLM_R_X3Y147_SLICE_X3Y147_B5Q),
.I4(LIOB33_X0Y61_IOB_X0Y62_I),
.I5(1'b1),
.O5(CLBLL_L_X4Y147_SLICE_X4Y147_DO5),
.O6(CLBLL_L_X4Y147_SLICE_X4Y147_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f0aaaaff00f0f0)
  ) CLBLL_L_X4Y147_SLICE_X4Y147_CLUT (
.I0(CLBLM_L_X10Y149_SLICE_X13Y149_AQ),
.I1(1'b1),
.I2(CLBLL_L_X4Y147_SLICE_X4Y147_DQ),
.I3(CLBLM_R_X7Y149_SLICE_X9Y149_A5Q),
.I4(LIOB33_X0Y61_IOB_X0Y62_I),
.I5(1'b1),
.O5(CLBLL_L_X4Y147_SLICE_X4Y147_CO5),
.O6(CLBLL_L_X4Y147_SLICE_X4Y147_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hb8b8b8b8f3c0f3c0)
  ) CLBLL_L_X4Y147_SLICE_X4Y147_BLUT (
.I0(CLBLM_R_X5Y150_SLICE_X6Y150_B5Q),
.I1(LIOB33_X0Y61_IOB_X0Y62_I),
.I2(CLBLL_L_X2Y146_SLICE_X1Y146_AQ),
.I3(CLBLM_R_X7Y143_SLICE_X9Y143_B5Q),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y147_SLICE_X4Y147_BO5),
.O6(CLBLL_L_X4Y147_SLICE_X4Y147_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hef23ef23ef23ef23)
  ) CLBLL_L_X4Y147_SLICE_X4Y147_ALUT (
.I0(CLBLL_L_X4Y150_SLICE_X4Y150_DO6),
.I1(LIOB33_X0Y61_IOB_X0Y62_I),
.I2(CLBLM_R_X5Y146_SLICE_X7Y146_BQ),
.I3(CLBLL_L_X4Y143_SLICE_X5Y143_BQ),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y147_SLICE_X4Y147_AO5),
.O6(CLBLL_L_X4Y147_SLICE_X4Y147_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y147_SLICE_X5Y147_B5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y147_SLICE_X5Y147_BO5),
.Q(CLBLL_L_X4Y147_SLICE_X5Y147_B5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "C5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y147_SLICE_X5Y147_C5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y147_SLICE_X5Y147_CO5),
.Q(CLBLL_L_X4Y147_SLICE_X5Y147_C5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y147_SLICE_X5Y147_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y147_SLICE_X5Y147_AO6),
.Q(CLBLL_L_X4Y147_SLICE_X5Y147_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y147_SLICE_X5Y147_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y147_SLICE_X5Y147_BO6),
.Q(CLBLL_L_X4Y147_SLICE_X5Y147_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y147_SLICE_X5Y147_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y147_SLICE_X5Y147_CO6),
.Q(CLBLL_L_X4Y147_SLICE_X5Y147_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffffdfffdfff)
  ) CLBLL_L_X4Y147_SLICE_X5Y147_DLUT (
.I0(CLBLM_R_X5Y145_SLICE_X6Y145_D5Q),
.I1(CLBLL_L_X4Y150_SLICE_X5Y150_CO5),
.I2(CLBLL_L_X4Y143_SLICE_X4Y143_BQ),
.I3(CLBLL_L_X4Y145_SLICE_X5Y145_BQ),
.I4(1'b1),
.I5(CLBLL_L_X4Y145_SLICE_X4Y145_DO5),
.O5(CLBLL_L_X4Y147_SLICE_X5Y147_DO5),
.O6(CLBLL_L_X4Y147_SLICE_X5Y147_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hff55aa00e4e4e4e4)
  ) CLBLL_L_X4Y147_SLICE_X5Y147_CLUT (
.I0(LIOB33_X0Y61_IOB_X0Y62_I),
.I1(CLBLM_R_X7Y143_SLICE_X9Y143_B5Q),
.I2(CLBLL_L_X4Y148_SLICE_X5Y148_CQ),
.I3(CLBLM_R_X5Y147_SLICE_X6Y147_B5Q),
.I4(RIOB33_X105Y109_IOB_X1Y109_I),
.I5(1'b1),
.O5(CLBLL_L_X4Y147_SLICE_X5Y147_CO5),
.O6(CLBLL_L_X4Y147_SLICE_X5Y147_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hcfcfc0c0afa0afa0)
  ) CLBLL_L_X4Y147_SLICE_X5Y147_BLUT (
.I0(CLBLM_R_X3Y148_SLICE_X2Y148_B5Q),
.I1(CLBLL_L_X4Y148_SLICE_X5Y148_D5Q),
.I2(LIOB33_X0Y61_IOB_X0Y62_I),
.I3(CLBLM_R_X7Y153_SLICE_X9Y153_DQ),
.I4(CLBLM_L_X8Y153_SLICE_X11Y153_CO6),
.I5(1'b1),
.O5(CLBLL_L_X4Y147_SLICE_X5Y147_BO5),
.O6(CLBLL_L_X4Y147_SLICE_X5Y147_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfedcefcd32102301)
  ) CLBLL_L_X4Y147_SLICE_X5Y147_ALUT (
.I0(CLBLM_L_X8Y149_SLICE_X11Y149_AQ),
.I1(LIOB33_X0Y61_IOB_X0Y62_I),
.I2(CLBLL_L_X4Y147_SLICE_X5Y147_AQ),
.I3(CLBLL_L_X4Y143_SLICE_X5Y143_BQ),
.I4(CLBLM_R_X5Y148_SLICE_X6Y148_AO6),
.I5(CLBLM_R_X5Y147_SLICE_X7Y147_BQ),
.O5(CLBLL_L_X4Y147_SLICE_X5Y147_AO5),
.O6(CLBLL_L_X4Y147_SLICE_X5Y147_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y148_SLICE_X4Y148_C5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y148_SLICE_X4Y148_CO5),
.Q(CLBLL_L_X4Y148_SLICE_X4Y148_C5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y148_SLICE_X4Y148_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y148_SLICE_X4Y148_AO6),
.Q(CLBLL_L_X4Y148_SLICE_X4Y148_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y148_SLICE_X4Y148_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y148_SLICE_X4Y148_BO6),
.Q(CLBLL_L_X4Y148_SLICE_X4Y148_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y148_SLICE_X4Y148_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y148_SLICE_X4Y148_CO6),
.Q(CLBLL_L_X4Y148_SLICE_X4Y148_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h8000000000000000)
  ) CLBLL_L_X4Y148_SLICE_X4Y148_DLUT (
.I0(CLBLL_L_X4Y151_SLICE_X4Y151_AQ),
.I1(CLBLM_R_X5Y145_SLICE_X6Y145_D5Q),
.I2(CLBLL_L_X4Y143_SLICE_X4Y143_AQ),
.I3(CLBLL_L_X4Y143_SLICE_X4Y143_BQ),
.I4(CLBLL_L_X4Y151_SLICE_X5Y151_CQ),
.I5(CLBLM_R_X3Y145_SLICE_X3Y145_BQ),
.O5(CLBLL_L_X4Y148_SLICE_X4Y148_DO5),
.O6(CLBLL_L_X4Y148_SLICE_X4Y148_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'ha0a0f5f5d8d8d8d8)
  ) CLBLL_L_X4Y148_SLICE_X4Y148_CLUT (
.I0(LIOB33_X0Y61_IOB_X0Y62_I),
.I1(CLBLL_L_X4Y148_SLICE_X5Y148_A5Q),
.I2(CLBLL_L_X4Y143_SLICE_X4Y143_A5Q),
.I3(1'b1),
.I4(CLBLM_L_X10Y153_SLICE_X13Y153_A5Q),
.I5(1'b1),
.O5(CLBLL_L_X4Y148_SLICE_X4Y148_CO5),
.O6(CLBLL_L_X4Y148_SLICE_X4Y148_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f0f0f0aaaaee22)
  ) CLBLL_L_X4Y148_SLICE_X4Y148_BLUT (
.I0(CLBLL_L_X4Y149_SLICE_X5Y149_BQ),
.I1(CLBLM_R_X3Y143_SLICE_X3Y143_BQ),
.I2(CLBLL_L_X4Y147_SLICE_X4Y147_C5Q),
.I3(CLBLM_L_X10Y149_SLICE_X13Y149_AQ),
.I4(CLBLL_L_X4Y142_SLICE_X4Y142_AQ),
.I5(LIOB33_X0Y61_IOB_X0Y62_I),
.O5(CLBLL_L_X4Y148_SLICE_X4Y148_BO5),
.O6(CLBLL_L_X4Y148_SLICE_X4Y148_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfcfcf5fc0c0c050c)
  ) CLBLL_L_X4Y148_SLICE_X4Y148_ALUT (
.I0(CLBLM_R_X3Y146_SLICE_X2Y146_D5Q),
.I1(CLBLL_L_X4Y148_SLICE_X4Y148_BQ),
.I2(LIOB33_X0Y61_IOB_X0Y62_I),
.I3(CLBLM_R_X3Y143_SLICE_X3Y143_BQ),
.I4(CLBLL_L_X4Y142_SLICE_X4Y142_AQ),
.I5(CLBLM_R_X3Y152_SLICE_X3Y152_CQ),
.O5(CLBLL_L_X4Y148_SLICE_X4Y148_AO5),
.O6(CLBLL_L_X4Y148_SLICE_X4Y148_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y148_SLICE_X5Y148_A5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y148_SLICE_X5Y148_AO5),
.Q(CLBLL_L_X4Y148_SLICE_X5Y148_A5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y148_SLICE_X5Y148_B5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y148_SLICE_X5Y148_BO5),
.Q(CLBLL_L_X4Y148_SLICE_X5Y148_B5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y148_SLICE_X5Y148_D5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y148_SLICE_X5Y148_DO5),
.Q(CLBLL_L_X4Y148_SLICE_X5Y148_D5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y148_SLICE_X5Y148_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y148_SLICE_X5Y148_AO6),
.Q(CLBLL_L_X4Y148_SLICE_X5Y148_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y148_SLICE_X5Y148_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y148_SLICE_X5Y148_BO6),
.Q(CLBLL_L_X4Y148_SLICE_X5Y148_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y148_SLICE_X5Y148_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y148_SLICE_X5Y148_CO6),
.Q(CLBLL_L_X4Y148_SLICE_X5Y148_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y148_SLICE_X5Y148_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y148_SLICE_X5Y148_DO6),
.Q(CLBLL_L_X4Y148_SLICE_X5Y148_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hee44ee44e4e4e4e4)
  ) CLBLL_L_X4Y148_SLICE_X5Y148_DLUT (
.I0(LIOB33_X0Y61_IOB_X0Y62_I),
.I1(CLBLM_R_X5Y152_SLICE_X6Y152_DQ),
.I2(CLBLM_R_X3Y148_SLICE_X3Y148_C5Q),
.I3(CLBLM_R_X5Y149_SLICE_X6Y149_CQ),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y148_SLICE_X5Y148_DO5),
.O6(CLBLL_L_X4Y148_SLICE_X5Y148_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hffee00eeffee00ee)
  ) CLBLL_L_X4Y148_SLICE_X5Y148_CLUT (
.I0(CLBLM_R_X7Y153_SLICE_X9Y153_AQ),
.I1(CLBLM_R_X5Y148_SLICE_X6Y148_BO6),
.I2(1'b1),
.I3(LIOB33_X0Y61_IOB_X0Y62_I),
.I4(CLBLL_L_X4Y148_SLICE_X5Y148_B5Q),
.I5(1'b1),
.O5(CLBLL_L_X4Y148_SLICE_X5Y148_CO5),
.O6(CLBLL_L_X4Y148_SLICE_X5Y148_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf606f606fff00f00)
  ) CLBLL_L_X4Y148_SLICE_X5Y148_BLUT (
.I0(CLBLL_L_X4Y140_SLICE_X5Y140_DO6),
.I1(CLBLL_L_X4Y148_SLICE_X5Y148_BQ),
.I2(LIOB33_X0Y61_IOB_X0Y62_I),
.I3(CLBLL_L_X4Y153_SLICE_X5Y153_A5Q),
.I4(CLBLM_R_X5Y152_SLICE_X7Y152_BQ),
.I5(1'b1),
.O5(CLBLL_L_X4Y148_SLICE_X5Y148_BO5),
.O6(CLBLL_L_X4Y148_SLICE_X5Y148_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfafa0a0acfc0cfc0)
  ) CLBLL_L_X4Y148_SLICE_X5Y148_ALUT (
.I0(CLBLL_L_X4Y148_SLICE_X5Y148_CQ),
.I1(CLBLL_L_X4Y153_SLICE_X5Y153_AQ),
.I2(LIOB33_X0Y61_IOB_X0Y62_I),
.I3(RIOB33_X105Y117_IOB_X1Y117_I),
.I4(CLBLM_R_X5Y145_SLICE_X7Y145_B5Q),
.I5(1'b1),
.O5(CLBLL_L_X4Y148_SLICE_X5Y148_AO5),
.O6(CLBLL_L_X4Y148_SLICE_X5Y148_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y149_SLICE_X4Y149_B5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y149_SLICE_X4Y149_BO5),
.Q(CLBLL_L_X4Y149_SLICE_X4Y149_B5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y149_SLICE_X4Y149_D5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y149_SLICE_X4Y149_DO5),
.Q(CLBLL_L_X4Y149_SLICE_X4Y149_D5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y149_SLICE_X4Y149_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y149_SLICE_X4Y149_AO6),
.Q(CLBLL_L_X4Y149_SLICE_X4Y149_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y149_SLICE_X4Y149_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y149_SLICE_X4Y149_BO6),
.Q(CLBLL_L_X4Y149_SLICE_X4Y149_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y149_SLICE_X4Y149_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y149_SLICE_X4Y149_CO6),
.Q(CLBLL_L_X4Y149_SLICE_X4Y149_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y149_SLICE_X4Y149_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y149_SLICE_X4Y149_DO6),
.Q(CLBLL_L_X4Y149_SLICE_X4Y149_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h8d8dd8d8aa00ff55)
  ) CLBLL_L_X4Y149_SLICE_X4Y149_DLUT (
.I0(LIOB33_X0Y61_IOB_X0Y62_I),
.I1(CLBLM_L_X10Y151_SLICE_X12Y151_DQ),
.I2(CLBLL_L_X4Y149_SLICE_X4Y149_DQ),
.I3(CLBLM_L_X10Y148_SLICE_X13Y148_AQ),
.I4(CLBLL_L_X4Y149_SLICE_X4Y149_D5Q),
.I5(1'b1),
.O5(CLBLL_L_X4Y149_SLICE_X4Y149_DO5),
.O6(CLBLL_L_X4Y149_SLICE_X4Y149_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'he2f3e2f3e2e2e2e2)
  ) CLBLL_L_X4Y149_SLICE_X4Y149_CLUT (
.I0(CLBLL_L_X4Y147_SLICE_X5Y147_C5Q),
.I1(LIOB33_X0Y61_IOB_X0Y62_I),
.I2(CLBLL_L_X4Y149_SLICE_X4Y149_DQ),
.I3(CLBLM_L_X8Y145_SLICE_X11Y145_DQ),
.I4(1'b1),
.I5(CLBLM_L_X8Y151_SLICE_X10Y151_AQ),
.O5(CLBLL_L_X4Y149_SLICE_X4Y149_CO5),
.O6(CLBLL_L_X4Y149_SLICE_X4Y149_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaaf0f0ccccff00)
  ) CLBLL_L_X4Y149_SLICE_X4Y149_BLUT (
.I0(CLBLM_R_X3Y149_SLICE_X2Y149_AQ),
.I1(CLBLL_L_X4Y149_SLICE_X4Y149_BQ),
.I2(CLBLM_R_X5Y152_SLICE_X6Y152_DQ),
.I3(CLBLM_L_X8Y147_SLICE_X10Y147_BQ),
.I4(LIOB33_X0Y61_IOB_X0Y62_I),
.I5(1'b1),
.O5(CLBLL_L_X4Y149_SLICE_X4Y149_BO5),
.O6(CLBLL_L_X4Y149_SLICE_X4Y149_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hff00ff5a0000005a)
  ) CLBLL_L_X4Y149_SLICE_X4Y149_ALUT (
.I0(CLBLL_L_X4Y146_SLICE_X4Y146_DO6),
.I1(1'b1),
.I2(CLBLL_L_X4Y149_SLICE_X4Y149_AQ),
.I3(LIOB33_X0Y61_IOB_X0Y62_I),
.I4(CLBLL_L_X4Y143_SLICE_X4Y143_D5Q),
.I5(CLBLM_R_X5Y149_SLICE_X6Y149_AQ),
.O5(CLBLL_L_X4Y149_SLICE_X4Y149_AO5),
.O6(CLBLL_L_X4Y149_SLICE_X4Y149_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y149_SLICE_X5Y149_C5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y149_SLICE_X5Y149_CO5),
.Q(CLBLL_L_X4Y149_SLICE_X5Y149_C5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y149_SLICE_X5Y149_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y149_SLICE_X5Y149_AO6),
.Q(CLBLL_L_X4Y149_SLICE_X5Y149_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y149_SLICE_X5Y149_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y149_SLICE_X5Y149_BO6),
.Q(CLBLL_L_X4Y149_SLICE_X5Y149_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y149_SLICE_X5Y149_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y149_SLICE_X5Y149_CO6),
.Q(CLBLL_L_X4Y149_SLICE_X5Y149_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y149_SLICE_X5Y149_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y149_SLICE_X5Y149_DO6),
.Q(CLBLL_L_X4Y149_SLICE_X5Y149_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff0000ffbfffbf)
  ) CLBLL_L_X4Y149_SLICE_X5Y149_DLUT (
.I0(CLBLL_L_X4Y151_SLICE_X4Y151_AQ),
.I1(CLBLL_L_X4Y143_SLICE_X4Y143_AQ),
.I2(CLBLL_L_X4Y143_SLICE_X4Y143_BQ),
.I3(CLBLL_L_X4Y151_SLICE_X5Y151_CQ),
.I4(CLBLL_L_X2Y145_SLICE_X0Y145_AQ),
.I5(LIOB33_X0Y61_IOB_X0Y62_I),
.O5(CLBLL_L_X4Y149_SLICE_X5Y149_DO5),
.O6(CLBLL_L_X4Y149_SLICE_X5Y149_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hcf03cf03c0c0f3f3)
  ) CLBLL_L_X4Y149_SLICE_X5Y149_CLUT (
.I0(1'b1),
.I1(LIOB33_X0Y61_IOB_X0Y62_I),
.I2(CLBLM_R_X5Y150_SLICE_X6Y150_C5Q),
.I3(CLBLM_R_X5Y149_SLICE_X6Y149_C5Q),
.I4(CLBLM_L_X8Y149_SLICE_X11Y149_BO6),
.I5(1'b1),
.O5(CLBLL_L_X4Y149_SLICE_X5Y149_CO5),
.O6(CLBLL_L_X4Y149_SLICE_X5Y149_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hd8d8d8d8ddd888d8)
  ) CLBLL_L_X4Y149_SLICE_X5Y149_BLUT (
.I0(LIOB33_X0Y61_IOB_X0Y62_I),
.I1(CLBLM_R_X7Y148_SLICE_X9Y148_BQ),
.I2(CLBLL_L_X4Y149_SLICE_X5Y149_AQ),
.I3(CLBLM_R_X3Y143_SLICE_X3Y143_BQ),
.I4(CLBLL_L_X4Y149_SLICE_X5Y149_C5Q),
.I5(CLBLL_L_X4Y142_SLICE_X4Y142_AQ),
.O5(CLBLL_L_X4Y149_SLICE_X5Y149_BO5),
.O6(CLBLL_L_X4Y149_SLICE_X5Y149_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffff300ff00f3)
  ) CLBLL_L_X4Y149_SLICE_X5Y149_ALUT (
.I0(1'b1),
.I1(CLBLM_R_X3Y143_SLICE_X3Y143_BQ),
.I2(CLBLL_L_X4Y142_SLICE_X4Y142_AQ),
.I3(LIOB33_X0Y61_IOB_X0Y62_I),
.I4(CLBLM_L_X10Y151_SLICE_X13Y151_A5Q),
.I5(CLBLM_R_X7Y142_SLICE_X8Y142_C5Q),
.O5(CLBLL_L_X4Y149_SLICE_X5Y149_AO5),
.O6(CLBLL_L_X4Y149_SLICE_X5Y149_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y150_SLICE_X4Y150_A5_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLL_L_X4Y150_SLICE_X4Y150_AO5),
.Q(CLBLL_L_X4Y150_SLICE_X4Y150_A5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y150_SLICE_X4Y150_B5_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLL_L_X4Y150_SLICE_X4Y150_BO5),
.Q(CLBLL_L_X4Y150_SLICE_X4Y150_B5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "C5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y150_SLICE_X4Y150_C5_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLL_L_X4Y150_SLICE_X4Y150_CO5),
.Q(CLBLL_L_X4Y150_SLICE_X4Y150_C5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y150_SLICE_X4Y150_A_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLL_L_X4Y150_SLICE_X4Y150_AO6),
.Q(CLBLL_L_X4Y150_SLICE_X4Y150_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y150_SLICE_X4Y150_B_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLL_L_X4Y150_SLICE_X4Y150_BO6),
.Q(CLBLL_L_X4Y150_SLICE_X4Y150_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y150_SLICE_X4Y150_C_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLL_L_X4Y150_SLICE_X4Y150_CO6),
.Q(CLBLL_L_X4Y150_SLICE_X4Y150_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffffff7ffffff)
  ) CLBLL_L_X4Y150_SLICE_X4Y150_DLUT (
.I0(CLBLM_R_X3Y151_SLICE_X3Y151_AQ),
.I1(CLBLL_L_X4Y145_SLICE_X5Y145_BQ),
.I2(CLBLL_L_X4Y150_SLICE_X5Y150_CO5),
.I3(CLBLM_R_X3Y151_SLICE_X3Y151_CQ),
.I4(CLBLL_L_X4Y150_SLICE_X4Y150_B5Q),
.I5(CLBLM_R_X3Y151_SLICE_X3Y151_BQ),
.O5(CLBLL_L_X4Y150_SLICE_X4Y150_DO5),
.O6(CLBLL_L_X4Y150_SLICE_X4Y150_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f05555ccccf0f0)
  ) CLBLL_L_X4Y150_SLICE_X4Y150_CLUT (
.I0(CLBLM_L_X10Y149_SLICE_X12Y149_BQ),
.I1(CLBLL_L_X4Y150_SLICE_X5Y150_BQ),
.I2(CLBLL_L_X4Y150_SLICE_X4Y150_BQ),
.I3(1'b1),
.I4(LIOB33_X0Y61_IOB_X0Y62_I),
.I5(1'b1),
.O5(CLBLL_L_X4Y150_SLICE_X4Y150_CO5),
.O6(CLBLL_L_X4Y150_SLICE_X4Y150_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f0ccccff00eeee)
  ) CLBLL_L_X4Y150_SLICE_X4Y150_BLUT (
.I0(CLBLM_R_X3Y151_SLICE_X2Y151_CO6),
.I1(CLBLM_R_X3Y145_SLICE_X2Y145_CQ),
.I2(CLBLL_L_X4Y149_SLICE_X5Y149_BQ),
.I3(CLBLM_R_X5Y143_SLICE_X7Y143_AQ),
.I4(LIOB33_X0Y61_IOB_X0Y62_I),
.I5(1'b1),
.O5(CLBLL_L_X4Y150_SLICE_X4Y150_BO5),
.O6(CLBLL_L_X4Y150_SLICE_X4Y150_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hcf03cf038b8b8b8b)
  ) CLBLL_L_X4Y150_SLICE_X4Y150_ALUT (
.I0(CLBLL_L_X4Y153_SLICE_X4Y153_B5Q),
.I1(LIOB33_X0Y61_IOB_X0Y62_I),
.I2(CLBLM_L_X10Y149_SLICE_X12Y149_BQ),
.I3(CLBLL_L_X4Y145_SLICE_X4Y145_BQ),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y150_SLICE_X4Y150_AO5),
.O6(CLBLL_L_X4Y150_SLICE_X4Y150_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y150_SLICE_X5Y150_A5_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLL_L_X4Y153_SLICE_X4Y153_CO6),
.Q(CLBLL_L_X4Y150_SLICE_X5Y150_A5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y150_SLICE_X5Y150_A_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLL_L_X4Y150_SLICE_X5Y150_AO6),
.Q(CLBLL_L_X4Y150_SLICE_X5Y150_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y150_SLICE_X5Y150_B_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLL_L_X4Y150_SLICE_X5Y150_BO6),
.Q(CLBLL_L_X4Y150_SLICE_X5Y150_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffffffeeffee)
  ) CLBLL_L_X4Y150_SLICE_X5Y150_DLUT (
.I0(CLBLL_L_X4Y145_SLICE_X5Y145_BQ),
.I1(CLBLM_R_X3Y151_SLICE_X3Y151_CQ),
.I2(1'b1),
.I3(CLBLM_R_X5Y152_SLICE_X6Y152_CQ),
.I4(1'b1),
.I5(CLBLM_R_X3Y151_SLICE_X3Y151_BQ),
.O5(CLBLL_L_X4Y150_SLICE_X5Y150_DO5),
.O6(CLBLL_L_X4Y150_SLICE_X5Y150_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffefe33ffffff)
  ) CLBLL_L_X4Y150_SLICE_X5Y150_CLUT (
.I0(CLBLM_R_X3Y151_SLICE_X3Y151_AQ),
.I1(CLBLM_R_X3Y145_SLICE_X3Y145_BQ),
.I2(CLBLL_L_X4Y150_SLICE_X4Y150_B5Q),
.I3(CLBLM_R_X5Y152_SLICE_X6Y152_CQ),
.I4(CLBLM_R_X5Y152_SLICE_X6Y152_DQ),
.I5(1'b1),
.O5(CLBLL_L_X4Y150_SLICE_X5Y150_CO5),
.O6(CLBLL_L_X4Y150_SLICE_X5Y150_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffaf8c0000af8c)
  ) CLBLL_L_X4Y150_SLICE_X5Y150_BLUT (
.I0(CLBLM_R_X7Y152_SLICE_X8Y152_D5Q),
.I1(CLBLL_L_X4Y150_SLICE_X5Y150_BQ),
.I2(CLBLM_R_X7Y142_SLICE_X8Y142_C5Q),
.I3(CLBLL_L_X4Y148_SLICE_X5Y148_D5Q),
.I4(LIOB33_X0Y61_IOB_X0Y62_I),
.I5(CLBLM_R_X5Y151_SLICE_X6Y151_BQ),
.O5(CLBLL_L_X4Y150_SLICE_X5Y150_BO5),
.O6(CLBLL_L_X4Y150_SLICE_X5Y150_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hccffccffccaaccaa)
  ) CLBLL_L_X4Y150_SLICE_X5Y150_ALUT (
.I0(CLBLL_L_X4Y150_SLICE_X5Y150_DO6),
.I1(CLBLM_R_X5Y145_SLICE_X6Y145_CQ),
.I2(1'b1),
.I3(LIOB33_X0Y61_IOB_X0Y62_I),
.I4(1'b1),
.I5(CLBLL_L_X4Y150_SLICE_X5Y150_CO6),
.O5(CLBLL_L_X4Y150_SLICE_X5Y150_AO5),
.O6(CLBLL_L_X4Y150_SLICE_X5Y150_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y151_SLICE_X4Y151_A5_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_R_X3Y151_SLICE_X3Y151_DO6),
.Q(CLBLL_L_X4Y151_SLICE_X4Y151_A5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y151_SLICE_X4Y151_B5_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLL_L_X4Y151_SLICE_X4Y151_BO5),
.Q(CLBLL_L_X4Y151_SLICE_X4Y151_B5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "C5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y151_SLICE_X4Y151_C5_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLL_L_X4Y151_SLICE_X4Y151_CO5),
.Q(CLBLL_L_X4Y151_SLICE_X4Y151_C5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y151_SLICE_X4Y151_A_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLL_L_X4Y151_SLICE_X4Y151_AO6),
.Q(CLBLL_L_X4Y151_SLICE_X4Y151_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y151_SLICE_X4Y151_B_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLL_L_X4Y151_SLICE_X4Y151_BO6),
.Q(CLBLL_L_X4Y151_SLICE_X4Y151_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y151_SLICE_X4Y151_C_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLL_L_X4Y151_SLICE_X4Y151_CO6),
.Q(CLBLL_L_X4Y151_SLICE_X4Y151_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y151_SLICE_X4Y151_D_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLL_L_X4Y151_SLICE_X4Y151_DO6),
.Q(CLBLL_L_X4Y151_SLICE_X4Y151_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffbf100000bf10)
  ) CLBLL_L_X4Y151_SLICE_X4Y151_DLUT (
.I0(CLBLL_L_X4Y142_SLICE_X4Y142_AQ),
.I1(CLBLM_L_X12Y151_SLICE_X16Y151_AQ),
.I2(CLBLM_R_X3Y143_SLICE_X3Y143_BQ),
.I3(CLBLL_L_X4Y152_SLICE_X4Y152_AQ),
.I4(LIOB33_X0Y61_IOB_X0Y62_I),
.I5(CLBLM_R_X7Y153_SLICE_X8Y153_CQ),
.O5(CLBLL_L_X4Y151_SLICE_X4Y151_DO5),
.O6(CLBLL_L_X4Y151_SLICE_X4Y151_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hffaa5500e4e4e4e4)
  ) CLBLL_L_X4Y151_SLICE_X4Y151_CLUT (
.I0(LIOB33_X0Y61_IOB_X0Y62_I),
.I1(CLBLL_L_X4Y143_SLICE_X4Y143_AQ),
.I2(CLBLM_R_X3Y147_SLICE_X3Y147_CQ),
.I3(CLBLM_L_X10Y150_SLICE_X12Y150_AQ),
.I4(CLBLM_R_X5Y152_SLICE_X7Y152_DQ),
.I5(1'b1),
.O5(CLBLL_L_X4Y151_SLICE_X4Y151_CO5),
.O6(CLBLL_L_X4Y151_SLICE_X4Y151_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf3f3c0c0bbbb8888)
  ) CLBLL_L_X4Y151_SLICE_X4Y151_BLUT (
.I0(CLBLM_R_X3Y151_SLICE_X3Y151_A5Q),
.I1(LIOB33_X0Y61_IOB_X0Y62_I),
.I2(CLBLM_L_X10Y153_SLICE_X13Y153_A5Q),
.I3(1'b1),
.I4(RIOB33_X105Y107_IOB_X1Y107_I),
.I5(1'b1),
.O5(CLBLL_L_X4Y151_SLICE_X4Y151_BO5),
.O6(CLBLL_L_X4Y151_SLICE_X4Y151_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffcffffc00cf00fc)
  ) CLBLL_L_X4Y151_SLICE_X4Y151_ALUT (
.I0(1'b1),
.I1(CLBLM_R_X3Y145_SLICE_X2Y145_CQ),
.I2(CLBLL_L_X4Y151_SLICE_X4Y151_AQ),
.I3(LIOB33_X0Y61_IOB_X0Y62_I),
.I4(CLBLL_L_X4Y143_SLICE_X5Y143_CO5),
.I5(CLBLL_L_X4Y150_SLICE_X4Y150_A5Q),
.O5(CLBLL_L_X4Y151_SLICE_X4Y151_AO5),
.O6(CLBLL_L_X4Y151_SLICE_X4Y151_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y151_SLICE_X5Y151_B5_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLL_L_X4Y151_SLICE_X5Y151_BO5),
.Q(CLBLL_L_X4Y151_SLICE_X5Y151_B5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y151_SLICE_X5Y151_D5_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLL_L_X4Y151_SLICE_X5Y151_DO5),
.Q(CLBLL_L_X4Y151_SLICE_X5Y151_D5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y151_SLICE_X5Y151_A_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLL_L_X4Y151_SLICE_X5Y151_AO6),
.Q(CLBLL_L_X4Y151_SLICE_X5Y151_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y151_SLICE_X5Y151_B_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLL_L_X4Y151_SLICE_X5Y151_BO6),
.Q(CLBLL_L_X4Y151_SLICE_X5Y151_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y151_SLICE_X5Y151_C_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLL_L_X4Y151_SLICE_X5Y151_CO6),
.Q(CLBLL_L_X4Y151_SLICE_X5Y151_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y151_SLICE_X5Y151_D_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLL_L_X4Y151_SLICE_X5Y151_DO6),
.Q(CLBLL_L_X4Y151_SLICE_X5Y151_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hdd88dd88f5f5a0a0)
  ) CLBLL_L_X4Y151_SLICE_X5Y151_DLUT (
.I0(LIOB33_X0Y61_IOB_X0Y62_I),
.I1(CLBLM_R_X5Y144_SLICE_X7Y144_CQ),
.I2(CLBLL_L_X4Y151_SLICE_X5Y151_DQ),
.I3(CLBLM_R_X3Y151_SLICE_X3Y151_BQ),
.I4(CLBLM_R_X3Y149_SLICE_X2Y149_C5Q),
.I5(1'b1),
.O5(CLBLL_L_X4Y151_SLICE_X5Y151_DO5),
.O6(CLBLL_L_X4Y151_SLICE_X5Y151_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hfff60f06fffc0f0c)
  ) CLBLL_L_X4Y151_SLICE_X5Y151_CLUT (
.I0(CLBLL_L_X4Y151_SLICE_X4Y151_AQ),
.I1(CLBLL_L_X4Y151_SLICE_X5Y151_CQ),
.I2(LIOB33_X0Y61_IOB_X0Y62_I),
.I3(CLBLM_R_X3Y145_SLICE_X2Y145_CQ),
.I4(CLBLL_L_X4Y151_SLICE_X5Y151_B5Q),
.I5(CLBLL_L_X4Y143_SLICE_X5Y143_CO5),
.O5(CLBLL_L_X4Y151_SLICE_X5Y151_CO5),
.O6(CLBLL_L_X4Y151_SLICE_X5Y151_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hc0c0cfcfa3aca3ac)
  ) CLBLL_L_X4Y151_SLICE_X5Y151_BLUT (
.I0(CLBLL_L_X4Y145_SLICE_X5Y145_AQ),
.I1(CLBLL_L_X4Y145_SLICE_X5Y145_BQ),
.I2(LIOB33_X0Y61_IOB_X0Y62_I),
.I3(CLBLL_L_X4Y146_SLICE_X4Y146_CQ),
.I4(CLBLM_L_X10Y153_SLICE_X13Y153_A5Q),
.I5(1'b1),
.O5(CLBLL_L_X4Y151_SLICE_X5Y151_BO5),
.O6(CLBLL_L_X4Y151_SLICE_X5Y151_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hee44fa50ee44ee44)
  ) CLBLL_L_X4Y151_SLICE_X5Y151_ALUT (
.I0(LIOB33_X0Y61_IOB_X0Y62_I),
.I1(CLBLL_L_X4Y151_SLICE_X5Y151_DQ),
.I2(CLBLL_L_X4Y151_SLICE_X5Y151_AQ),
.I3(CLBLM_R_X7Y150_SLICE_X8Y150_AQ),
.I4(CLBLM_R_X7Y152_SLICE_X8Y152_D5Q),
.I5(CLBLM_R_X7Y142_SLICE_X8Y142_C5Q),
.O5(CLBLL_L_X4Y151_SLICE_X5Y151_AO5),
.O6(CLBLL_L_X4Y151_SLICE_X5Y151_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y152_SLICE_X4Y152_B5_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLL_L_X4Y152_SLICE_X4Y152_BO5),
.Q(CLBLL_L_X4Y152_SLICE_X4Y152_B5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y152_SLICE_X4Y152_A_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLL_L_X4Y152_SLICE_X4Y152_AO6),
.Q(CLBLL_L_X4Y152_SLICE_X4Y152_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y152_SLICE_X4Y152_B_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLL_L_X4Y152_SLICE_X4Y152_BO6),
.Q(CLBLL_L_X4Y152_SLICE_X4Y152_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y152_SLICE_X4Y152_C_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLL_L_X4Y152_SLICE_X4Y152_CO6),
.Q(CLBLL_L_X4Y152_SLICE_X4Y152_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y152_SLICE_X4Y152_D_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLL_L_X4Y152_SLICE_X4Y152_DO6),
.Q(CLBLL_L_X4Y152_SLICE_X4Y152_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaaaabf00000015)
  ) CLBLL_L_X4Y152_SLICE_X4Y152_DLUT (
.I0(LIOB33_X0Y61_IOB_X0Y62_I),
.I1(CLBLL_L_X4Y152_SLICE_X4Y152_CQ),
.I2(CLBLL_L_X4Y152_SLICE_X4Y152_DQ),
.I3(CLBLL_L_X4Y152_SLICE_X4Y152_BQ),
.I4(CLBLM_R_X5Y153_SLICE_X6Y153_DQ),
.I5(CLBLM_R_X5Y152_SLICE_X7Y152_A5Q),
.O5(CLBLL_L_X4Y152_SLICE_X4Y152_DO5),
.O6(CLBLL_L_X4Y152_SLICE_X4Y152_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hddddddd8ddddddd8)
  ) CLBLL_L_X4Y152_SLICE_X4Y152_CLUT (
.I0(LIOB33_X0Y61_IOB_X0Y62_I),
.I1(CLBLM_R_X7Y152_SLICE_X8Y152_DQ),
.I2(CLBLL_L_X4Y152_SLICE_X4Y152_DQ),
.I3(CLBLL_L_X4Y152_SLICE_X4Y152_BQ),
.I4(CLBLM_R_X5Y153_SLICE_X6Y153_DQ),
.I5(1'b1),
.O5(CLBLL_L_X4Y152_SLICE_X4Y152_CO5),
.O6(CLBLL_L_X4Y152_SLICE_X4Y152_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f0aaaaff00cccc)
  ) CLBLL_L_X4Y152_SLICE_X4Y152_BLUT (
.I0(CLBLL_L_X4Y147_SLICE_X4Y147_B5Q),
.I1(CLBLM_R_X3Y145_SLICE_X2Y145_DO6),
.I2(CLBLL_L_X4Y151_SLICE_X4Y151_B5Q),
.I3(CLBLL_L_X4Y152_SLICE_X5Y152_BQ),
.I4(LIOB33_X0Y61_IOB_X0Y62_I),
.I5(1'b1),
.O5(CLBLL_L_X4Y152_SLICE_X4Y152_BO5),
.O6(CLBLL_L_X4Y152_SLICE_X4Y152_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffccdfce33001302)
  ) CLBLL_L_X4Y152_SLICE_X4Y152_ALUT (
.I0(CLBLM_R_X3Y143_SLICE_X3Y143_BQ),
.I1(LIOB33_X0Y61_IOB_X0Y62_I),
.I2(CLBLM_L_X10Y149_SLICE_X12Y149_BQ),
.I3(CLBLL_L_X4Y152_SLICE_X5Y152_BQ),
.I4(CLBLL_L_X4Y142_SLICE_X4Y142_AQ),
.I5(CLBLM_L_X8Y152_SLICE_X11Y152_BQ),
.O5(CLBLL_L_X4Y152_SLICE_X4Y152_AO5),
.O6(CLBLL_L_X4Y152_SLICE_X4Y152_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y152_SLICE_X5Y152_A5_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLL_L_X4Y152_SLICE_X5Y152_CO5),
.Q(CLBLL_L_X4Y152_SLICE_X5Y152_A5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y152_SLICE_X5Y152_A_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLL_L_X4Y152_SLICE_X5Y152_AO6),
.Q(CLBLL_L_X4Y152_SLICE_X5Y152_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y152_SLICE_X5Y152_B_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLL_L_X4Y152_SLICE_X5Y152_BO6),
.Q(CLBLL_L_X4Y152_SLICE_X5Y152_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h8000000000000000)
  ) CLBLL_L_X4Y152_SLICE_X5Y152_DLUT (
.I0(CLBLM_R_X5Y154_SLICE_X6Y154_AQ),
.I1(CLBLL_L_X4Y153_SLICE_X5Y153_AQ),
.I2(CLBLM_R_X7Y153_SLICE_X9Y153_AQ),
.I3(CLBLM_R_X3Y149_SLICE_X3Y149_AQ),
.I4(CLBLM_R_X3Y149_SLICE_X2Y149_AQ),
.I5(CLBLM_R_X5Y154_SLICE_X6Y154_BQ),
.O5(CLBLL_L_X4Y152_SLICE_X5Y152_DO5),
.O6(CLBLL_L_X4Y152_SLICE_X5Y152_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hff00000088d8d888)
  ) CLBLL_L_X4Y152_SLICE_X5Y152_CLUT (
.I0(LIOB33_X0Y61_IOB_X0Y62_I),
.I1(CLBLM_R_X5Y152_SLICE_X6Y152_BQ),
.I2(CLBLL_L_X2Y150_SLICE_X1Y150_AQ),
.I3(CLBLL_L_X4Y152_SLICE_X5Y152_A5Q),
.I4(CLBLL_L_X4Y152_SLICE_X5Y152_DO6),
.I5(1'b1),
.O5(CLBLL_L_X4Y152_SLICE_X5Y152_CO5),
.O6(CLBLL_L_X4Y152_SLICE_X5Y152_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hff00ff00f0f07474)
  ) CLBLL_L_X4Y152_SLICE_X5Y152_BLUT (
.I0(CLBLM_L_X10Y153_SLICE_X13Y153_A5Q),
.I1(CLBLM_R_X3Y143_SLICE_X3Y143_BQ),
.I2(CLBLL_L_X4Y146_SLICE_X5Y146_DQ),
.I3(CLBLM_R_X5Y153_SLICE_X7Y153_BQ),
.I4(CLBLL_L_X4Y142_SLICE_X4Y142_AQ),
.I5(LIOB33_X0Y61_IOB_X0Y62_I),
.O5(CLBLL_L_X4Y152_SLICE_X5Y152_BO5),
.O6(CLBLL_L_X4Y152_SLICE_X5Y152_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hff280028ffa000a0)
  ) CLBLL_L_X4Y152_SLICE_X5Y152_ALUT (
.I0(CLBLL_L_X2Y150_SLICE_X1Y150_AQ),
.I1(CLBLM_R_X3Y152_SLICE_X3Y152_AQ),
.I2(CLBLL_L_X4Y152_SLICE_X5Y152_AQ),
.I3(LIOB33_X0Y61_IOB_X0Y62_I),
.I4(CLBLL_L_X4Y144_SLICE_X4Y144_C5Q),
.I5(CLBLL_L_X4Y152_SLICE_X5Y152_CO6),
.O5(CLBLL_L_X4Y152_SLICE_X5Y152_AO5),
.O6(CLBLL_L_X4Y152_SLICE_X5Y152_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y153_SLICE_X4Y153_A5_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLL_L_X4Y153_SLICE_X4Y153_AO5),
.Q(CLBLL_L_X4Y153_SLICE_X4Y153_A5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y153_SLICE_X4Y153_B5_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLL_L_X4Y153_SLICE_X4Y153_BO5),
.Q(CLBLL_L_X4Y153_SLICE_X4Y153_B5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y153_SLICE_X4Y153_A_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLL_L_X4Y153_SLICE_X4Y153_AO6),
.Q(CLBLL_L_X4Y153_SLICE_X4Y153_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y153_SLICE_X4Y153_B_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLL_L_X4Y153_SLICE_X4Y153_BO6),
.Q(CLBLL_L_X4Y153_SLICE_X4Y153_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaa300000ff00ff)
  ) CLBLL_L_X4Y153_SLICE_X4Y153_DLUT (
.I0(CLBLM_R_X5Y147_SLICE_X7Y147_AQ),
.I1(CLBLL_L_X4Y153_SLICE_X5Y153_A5Q),
.I2(CLBLM_R_X7Y145_SLICE_X8Y145_A5Q),
.I3(RIOB33_X105Y131_IOB_X1Y131_I),
.I4(LIOB33_X0Y61_IOB_X0Y62_I),
.I5(1'b1),
.O5(CLBLL_L_X4Y153_SLICE_X4Y153_DO5),
.O6(CLBLL_L_X4Y153_SLICE_X4Y153_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h88b88888000000ff)
  ) CLBLL_L_X4Y153_SLICE_X4Y153_CLUT (
.I0(CLBLL_L_X4Y142_SLICE_X4Y142_AQ),
.I1(LIOB33_X0Y61_IOB_X0Y62_I),
.I2(RIOB33_X105Y131_IOB_X1Y131_I),
.I3(CLBLM_R_X5Y142_SLICE_X7Y142_CO6),
.I4(RIOB33_SING_X105Y100_IOB_X1Y100_I),
.I5(1'b1),
.O5(CLBLL_L_X4Y153_SLICE_X4Y153_CO5),
.O6(CLBLL_L_X4Y153_SLICE_X4Y153_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hbb88bb88cf03cf03)
  ) CLBLL_L_X4Y153_SLICE_X4Y153_BLUT (
.I0(CLBLM_L_X10Y152_SLICE_X13Y152_AQ),
.I1(LIOB33_X0Y61_IOB_X0Y62_I),
.I2(CLBLM_L_X10Y153_SLICE_X13Y153_A5Q),
.I3(CLBLL_L_X4Y149_SLICE_X4Y149_CQ),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y153_SLICE_X4Y153_BO5),
.O6(CLBLL_L_X4Y153_SLICE_X4Y153_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'haa00aaffccffcc00)
  ) CLBLL_L_X4Y153_SLICE_X4Y153_ALUT (
.I0(CLBLM_R_X5Y154_SLICE_X7Y154_AQ),
.I1(CLBLL_L_X4Y152_SLICE_X4Y152_BQ),
.I2(1'b1),
.I3(LIOB33_X0Y61_IOB_X0Y62_I),
.I4(CLBLM_R_X5Y150_SLICE_X6Y150_C5Q),
.I5(1'b1),
.O5(CLBLL_L_X4Y153_SLICE_X4Y153_AO5),
.O6(CLBLL_L_X4Y153_SLICE_X4Y153_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y153_SLICE_X5Y153_A5_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLL_L_X4Y153_SLICE_X4Y153_DO6),
.Q(CLBLL_L_X4Y153_SLICE_X5Y153_A5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y153_SLICE_X5Y153_A_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLL_L_X4Y153_SLICE_X5Y153_AO6),
.Q(CLBLL_L_X4Y153_SLICE_X5Y153_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X4Y153_SLICE_X5Y153_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y153_SLICE_X5Y153_DO5),
.O6(CLBLL_L_X4Y153_SLICE_X5Y153_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X4Y153_SLICE_X5Y153_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y153_SLICE_X5Y153_CO5),
.O6(CLBLL_L_X4Y153_SLICE_X5Y153_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h8000000080808080)
  ) CLBLL_L_X4Y153_SLICE_X5Y153_BLUT (
.I0(CLBLM_R_X3Y149_SLICE_X2Y149_AQ),
.I1(CLBLM_R_X3Y149_SLICE_X3Y149_AQ),
.I2(CLBLM_R_X7Y153_SLICE_X9Y153_AQ),
.I3(CLBLM_R_X5Y154_SLICE_X6Y154_BQ),
.I4(CLBLM_R_X5Y154_SLICE_X6Y154_AQ),
.I5(1'b1),
.O5(CLBLL_L_X4Y153_SLICE_X5Y153_BO5),
.O6(CLBLL_L_X4Y153_SLICE_X5Y153_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hceec0220ceec0220)
  ) CLBLL_L_X4Y153_SLICE_X5Y153_ALUT (
.I0(CLBLL_L_X2Y150_SLICE_X1Y150_AQ),
.I1(LIOB33_X0Y61_IOB_X0Y62_I),
.I2(CLBLL_L_X4Y153_SLICE_X5Y153_AQ),
.I3(CLBLL_L_X4Y153_SLICE_X5Y153_BO6),
.I4(CLBLL_L_X4Y148_SLICE_X5Y148_AQ),
.I5(1'b1),
.O5(CLBLL_L_X4Y153_SLICE_X5Y153_AO5),
.O6(CLBLL_L_X4Y153_SLICE_X5Y153_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y142_SLICE_X10Y142_A5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y142_SLICE_X11Y142_CO6),
.Q(CLBLM_L_X8Y142_SLICE_X10Y142_A5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y142_SLICE_X10Y142_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y142_SLICE_X10Y142_AO6),
.Q(CLBLM_L_X8Y142_SLICE_X10Y142_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y142_SLICE_X10Y142_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y142_SLICE_X10Y142_BO6),
.Q(CLBLM_L_X8Y142_SLICE_X10Y142_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y142_SLICE_X10Y142_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y142_SLICE_X10Y142_CO6),
.Q(CLBLM_L_X8Y142_SLICE_X10Y142_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hffeef0e0f0e0f0e0)
  ) CLBLM_L_X8Y142_SLICE_X10Y142_DLUT (
.I0(CLBLM_R_X7Y141_SLICE_X9Y141_AQ),
.I1(CLBLM_L_X8Y142_SLICE_X10Y142_CQ),
.I2(CLBLM_L_X10Y142_SLICE_X12Y142_CO6),
.I3(CLBLM_R_X7Y143_SLICE_X9Y143_CQ),
.I4(CLBLM_L_X8Y145_SLICE_X11Y145_DQ),
.I5(RIOB33_X105Y131_IOB_X1Y131_I),
.O5(CLBLM_L_X8Y142_SLICE_X10Y142_DO5),
.O6(CLBLM_L_X8Y142_SLICE_X10Y142_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hf000f000f909f000)
  ) CLBLM_L_X8Y142_SLICE_X10Y142_CLUT (
.I0(CLBLM_R_X7Y141_SLICE_X9Y141_AQ),
.I1(CLBLM_L_X8Y142_SLICE_X10Y142_CQ),
.I2(LIOB33_X0Y61_IOB_X0Y62_I),
.I3(CLBLM_R_X5Y142_SLICE_X7Y142_BQ),
.I4(CLBLM_L_X8Y142_SLICE_X10Y142_DO6),
.I5(CLBLL_L_X4Y151_SLICE_X4Y151_CQ),
.O5(CLBLM_L_X8Y142_SLICE_X10Y142_CO5),
.O6(CLBLM_L_X8Y142_SLICE_X10Y142_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hbb11ee44aa00aa00)
  ) CLBLM_L_X8Y142_SLICE_X10Y142_BLUT (
.I0(LIOB33_X0Y61_IOB_X0Y62_I),
.I1(CLBLM_L_X8Y142_SLICE_X10Y142_BQ),
.I2(1'b1),
.I3(CLBLM_R_X5Y143_SLICE_X6Y143_BQ),
.I4(CLBLM_L_X8Y144_SLICE_X10Y144_AO6),
.I5(CLBLM_L_X10Y144_SLICE_X12Y144_AO6),
.O5(CLBLM_L_X8Y142_SLICE_X10Y142_BO5),
.O6(CLBLM_L_X8Y142_SLICE_X10Y142_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'heeea4440fffa5550)
  ) CLBLM_L_X8Y142_SLICE_X10Y142_ALUT (
.I0(LIOB33_X0Y61_IOB_X0Y62_I),
.I1(CLBLM_L_X10Y145_SLICE_X12Y145_AQ),
.I2(CLBLM_L_X8Y142_SLICE_X10Y142_AQ),
.I3(CLBLM_R_X7Y142_SLICE_X8Y142_CQ),
.I4(CLBLM_L_X8Y143_SLICE_X11Y143_CQ),
.I5(CLBLM_R_X5Y142_SLICE_X7Y142_BQ),
.O5(CLBLM_L_X8Y142_SLICE_X10Y142_AO5),
.O6(CLBLM_L_X8Y142_SLICE_X10Y142_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y142_SLICE_X11Y142_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y142_SLICE_X11Y142_AO6),
.Q(CLBLM_L_X8Y142_SLICE_X11Y142_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y142_SLICE_X11Y142_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y142_SLICE_X11Y142_BO6),
.Q(CLBLM_L_X8Y142_SLICE_X11Y142_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h2020202020ff2020)
  ) CLBLM_L_X8Y142_SLICE_X11Y142_DLUT (
.I0(CLBLM_L_X8Y142_SLICE_X11Y142_BQ),
.I1(CLBLL_L_X4Y151_SLICE_X4Y151_CQ),
.I2(RIOB33_X105Y131_IOB_X1Y131_I),
.I3(CLBLM_L_X8Y142_SLICE_X10Y142_CQ),
.I4(CLBLM_R_X7Y141_SLICE_X9Y141_AQ),
.I5(CLBLM_R_X7Y143_SLICE_X9Y143_CQ),
.O5(CLBLM_L_X8Y142_SLICE_X11Y142_DO5),
.O6(CLBLM_L_X8Y142_SLICE_X11Y142_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'haca0a0a0cc000000)
  ) CLBLM_L_X8Y142_SLICE_X11Y142_CLUT (
.I0(CLBLM_L_X10Y142_SLICE_X13Y142_AQ),
.I1(RIOB33_X105Y131_IOB_X1Y131_I),
.I2(LIOB33_X0Y61_IOB_X0Y62_I),
.I3(CLBLL_L_X4Y150_SLICE_X5Y150_A5Q),
.I4(CLBLM_R_X5Y142_SLICE_X7Y142_CO6),
.I5(1'b1),
.O5(CLBLM_L_X8Y142_SLICE_X11Y142_CO5),
.O6(CLBLM_L_X8Y142_SLICE_X11Y142_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaaffee00005544)
  ) CLBLM_L_X8Y142_SLICE_X11Y142_BLUT (
.I0(LIOB33_X0Y61_IOB_X0Y62_I),
.I1(CLBLM_L_X10Y144_SLICE_X12Y144_CO6),
.I2(1'b1),
.I3(CLBLM_L_X8Y142_SLICE_X11Y142_DO6),
.I4(CLBLM_L_X8Y142_SLICE_X11Y142_CO5),
.I5(CLBLL_L_X4Y150_SLICE_X4Y150_B5Q),
.O5(CLBLM_L_X8Y142_SLICE_X11Y142_BO5),
.O6(CLBLM_L_X8Y142_SLICE_X11Y142_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffbbfaba55115010)
  ) CLBLM_L_X8Y142_SLICE_X11Y142_ALUT (
.I0(LIOB33_X0Y61_IOB_X0Y62_I),
.I1(CLBLM_R_X3Y145_SLICE_X3Y145_D5Q),
.I2(CLBLM_L_X8Y142_SLICE_X11Y142_AQ),
.I3(CLBLL_L_X4Y151_SLICE_X4Y151_BQ),
.I4(CLBLL_L_X4Y142_SLICE_X4Y142_A5Q),
.I5(CLBLM_L_X8Y144_SLICE_X11Y144_CQ),
.O5(CLBLM_L_X8Y142_SLICE_X11Y142_AO5),
.O6(CLBLM_L_X8Y142_SLICE_X11Y142_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y143_SLICE_X10Y143_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y143_SLICE_X10Y143_AO6),
.Q(CLBLM_L_X8Y143_SLICE_X10Y143_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y143_SLICE_X10Y143_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y143_SLICE_X10Y143_BO6),
.Q(CLBLM_L_X8Y143_SLICE_X10Y143_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y143_SLICE_X10Y143_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y143_SLICE_X10Y143_CO6),
.Q(CLBLM_L_X8Y143_SLICE_X10Y143_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y143_SLICE_X10Y143_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y143_SLICE_X10Y143_DO6),
.Q(CLBLM_L_X8Y143_SLICE_X10Y143_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hff00ff00bbbbb0b0)
  ) CLBLM_L_X8Y143_SLICE_X10Y143_DLUT (
.I0(CLBLL_L_X4Y151_SLICE_X4Y151_BQ),
.I1(CLBLM_R_X3Y145_SLICE_X3Y145_D5Q),
.I2(CLBLM_L_X8Y143_SLICE_X10Y143_DQ),
.I3(CLBLM_R_X5Y146_SLICE_X7Y146_DQ),
.I4(CLBLM_R_X7Y148_SLICE_X9Y148_C5Q),
.I5(LIOB33_X0Y61_IOB_X0Y62_I),
.O5(CLBLM_L_X8Y143_SLICE_X10Y143_DO5),
.O6(CLBLM_L_X8Y143_SLICE_X10Y143_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'haaffaa00aacfaac0)
  ) CLBLM_L_X8Y143_SLICE_X10Y143_CLUT (
.I0(CLBLM_L_X8Y142_SLICE_X10Y142_AQ),
.I1(CLBLM_L_X8Y143_SLICE_X10Y143_CQ),
.I2(CLBLL_L_X4Y142_SLICE_X5Y142_DQ),
.I3(LIOB33_X0Y61_IOB_X0Y62_I),
.I4(CLBLM_R_X5Y143_SLICE_X7Y143_CQ),
.I5(CLBLL_L_X4Y147_SLICE_X5Y147_CQ),
.O5(CLBLM_L_X8Y143_SLICE_X10Y143_CO5),
.O6(CLBLM_L_X8Y143_SLICE_X10Y143_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf5f5e4b1a0a0e4b1)
  ) CLBLM_L_X8Y143_SLICE_X10Y143_BLUT (
.I0(LIOB33_X0Y61_IOB_X0Y62_I),
.I1(CLBLM_L_X8Y143_SLICE_X10Y143_BQ),
.I2(CLBLM_L_X10Y144_SLICE_X13Y144_CQ),
.I3(CLBLM_L_X10Y143_SLICE_X12Y143_CO6),
.I4(CLBLM_L_X8Y149_SLICE_X11Y149_AQ),
.I5(CLBLM_L_X8Y151_SLICE_X10Y151_CQ),
.O5(CLBLM_L_X8Y143_SLICE_X10Y143_BO5),
.O6(CLBLM_L_X8Y143_SLICE_X10Y143_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hccccf000cccc5a00)
  ) CLBLM_L_X8Y143_SLICE_X10Y143_ALUT (
.I0(CLBLM_L_X10Y144_SLICE_X13Y144_A5Q),
.I1(CLBLM_L_X8Y151_SLICE_X10Y151_BQ),
.I2(CLBLM_L_X8Y143_SLICE_X10Y143_AQ),
.I3(CLBLM_L_X10Y144_SLICE_X12Y144_AO6),
.I4(LIOB33_X0Y61_IOB_X0Y62_I),
.I5(CLBLM_R_X3Y142_SLICE_X2Y142_BO5),
.O5(CLBLM_L_X8Y143_SLICE_X10Y143_AO5),
.O6(CLBLM_L_X8Y143_SLICE_X10Y143_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y143_SLICE_X11Y143_D5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y143_SLICE_X11Y143_DO5),
.Q(CLBLM_L_X8Y143_SLICE_X11Y143_D5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y143_SLICE_X11Y143_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y143_SLICE_X11Y143_AO6),
.Q(CLBLM_L_X8Y143_SLICE_X11Y143_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y143_SLICE_X11Y143_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y143_SLICE_X11Y143_BO6),
.Q(CLBLM_L_X8Y143_SLICE_X11Y143_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y143_SLICE_X11Y143_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y143_SLICE_X11Y143_CO6),
.Q(CLBLM_L_X8Y143_SLICE_X11Y143_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y143_SLICE_X11Y143_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y143_SLICE_X11Y143_DO6),
.Q(CLBLM_L_X8Y143_SLICE_X11Y143_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hfafa0a0acacacaca)
  ) CLBLM_L_X8Y143_SLICE_X11Y143_DLUT (
.I0(CLBLL_L_X4Y143_SLICE_X4Y143_AQ),
.I1(CLBLM_L_X10Y143_SLICE_X13Y143_BQ),
.I2(LIOB33_X0Y61_IOB_X0Y62_I),
.I3(1'b1),
.I4(CLBLM_L_X8Y143_SLICE_X10Y143_DQ),
.I5(1'b1),
.O5(CLBLM_L_X8Y143_SLICE_X11Y143_DO5),
.O6(CLBLM_L_X8Y143_SLICE_X11Y143_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hafaca0acafaca0ac)
  ) CLBLM_L_X8Y143_SLICE_X11Y143_CLUT (
.I0(CLBLL_L_X4Y149_SLICE_X5Y149_C5Q),
.I1(CLBLM_L_X8Y143_SLICE_X11Y143_CQ),
.I2(LIOB33_X0Y61_IOB_X0Y62_I),
.I3(CLBLM_L_X12Y149_SLICE_X17Y149_CO6),
.I4(CLBLM_L_X8Y143_SLICE_X10Y143_DQ),
.I5(1'b1),
.O5(CLBLM_L_X8Y143_SLICE_X11Y143_CO5),
.O6(CLBLM_L_X8Y143_SLICE_X11Y143_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hffdd3311eecc2200)
  ) CLBLM_L_X8Y143_SLICE_X11Y143_BLUT (
.I0(CLBLM_R_X13Y149_SLICE_X18Y149_AO6),
.I1(LIOB33_X0Y61_IOB_X0Y62_I),
.I2(1'b1),
.I3(CLBLM_L_X8Y145_SLICE_X11Y145_BQ),
.I4(CLBLM_R_X7Y141_SLICE_X9Y141_AQ),
.I5(CLBLM_L_X8Y143_SLICE_X11Y143_BQ),
.O5(CLBLM_L_X8Y143_SLICE_X11Y143_BO5),
.O6(CLBLM_L_X8Y143_SLICE_X11Y143_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hee22ff33ec20fc30)
  ) CLBLM_L_X8Y143_SLICE_X11Y143_ALUT (
.I0(CLBLM_R_X7Y152_SLICE_X8Y152_D5Q),
.I1(LIOB33_X0Y61_IOB_X0Y62_I),
.I2(CLBLM_L_X8Y143_SLICE_X11Y143_AQ),
.I3(CLBLM_L_X10Y143_SLICE_X12Y143_AQ),
.I4(CLBLM_R_X7Y142_SLICE_X8Y142_C5Q),
.I5(CLBLM_R_X7Y145_SLICE_X8Y145_D5Q),
.O5(CLBLM_L_X8Y143_SLICE_X11Y143_AO5),
.O6(CLBLM_L_X8Y143_SLICE_X11Y143_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y144_SLICE_X10Y144_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(LIOB33_X0Y61_IOB_X0Y62_I),
.D(CLBLM_R_X7Y144_SLICE_X8Y144_DQ),
.Q(CLBLM_L_X8Y144_SLICE_X10Y144_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y144_SLICE_X10Y144_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(LIOB33_X0Y61_IOB_X0Y62_I),
.D(CLBLM_R_X7Y142_SLICE_X9Y142_AQ),
.Q(CLBLM_L_X8Y144_SLICE_X10Y144_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h003088b800000000)
  ) CLBLM_L_X8Y144_SLICE_X10Y144_DLUT (
.I0(CLBLM_L_X8Y143_SLICE_X11Y143_BQ),
.I1(CLBLM_R_X7Y153_SLICE_X8Y153_A5Q),
.I2(CLBLM_L_X8Y144_SLICE_X11Y144_B5Q),
.I3(CLBLM_R_X11Y144_SLICE_X14Y144_AO6),
.I4(CLBLM_R_X11Y144_SLICE_X14Y144_CO6),
.I5(CLBLM_R_X7Y144_SLICE_X9Y144_B5Q),
.O5(CLBLM_L_X8Y144_SLICE_X10Y144_DO5),
.O6(CLBLM_L_X8Y144_SLICE_X10Y144_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h222222222f222222)
  ) CLBLM_L_X8Y144_SLICE_X10Y144_CLUT (
.I0(CLBLM_R_X7Y144_SLICE_X8Y144_CQ),
.I1(CLBLM_R_X7Y146_SLICE_X9Y146_DO6),
.I2(CLBLM_R_X11Y144_SLICE_X14Y144_BO6),
.I3(CLBLM_R_X7Y153_SLICE_X8Y153_A5Q),
.I4(CLBLL_L_X4Y144_SLICE_X4Y144_DQ),
.I5(CLBLM_R_X7Y144_SLICE_X9Y144_B5Q),
.O5(CLBLM_L_X8Y144_SLICE_X10Y144_CO5),
.O6(CLBLM_L_X8Y144_SLICE_X10Y144_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h3cc3c33cbb11bb11)
  ) CLBLM_L_X8Y144_SLICE_X10Y144_BLUT (
.I0(LIOB33_X0Y61_IOB_X0Y62_I),
.I1(CLBLM_L_X12Y151_SLICE_X16Y151_AQ),
.I2(CLBLM_L_X10Y149_SLICE_X12Y149_BQ),
.I3(CLBLM_L_X10Y151_SLICE_X13Y151_AQ),
.I4(CLBLM_R_X3Y146_SLICE_X2Y146_D5Q),
.I5(1'b1),
.O5(CLBLM_L_X8Y144_SLICE_X10Y144_BO5),
.O6(CLBLM_L_X8Y144_SLICE_X10Y144_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0a0000005a555555)
  ) CLBLM_L_X8Y144_SLICE_X10Y144_ALUT (
.I0(CLBLM_R_X5Y145_SLICE_X7Y145_B5Q),
.I1(1'b1),
.I2(CLBLM_R_X3Y142_SLICE_X2Y142_BO5),
.I3(CLBLM_L_X8Y143_SLICE_X10Y143_AQ),
.I4(CLBLM_L_X10Y144_SLICE_X13Y144_A5Q),
.I5(1'b1),
.O5(CLBLM_L_X8Y144_SLICE_X10Y144_AO5),
.O6(CLBLM_L_X8Y144_SLICE_X10Y144_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y144_SLICE_X11Y144_B5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y144_SLICE_X11Y144_BO5),
.Q(CLBLM_L_X8Y144_SLICE_X11Y144_B5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y144_SLICE_X11Y144_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y144_SLICE_X11Y144_AO6),
.Q(CLBLM_L_X8Y144_SLICE_X11Y144_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y144_SLICE_X11Y144_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y144_SLICE_X11Y144_BO6),
.Q(CLBLM_L_X8Y144_SLICE_X11Y144_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y144_SLICE_X11Y144_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y144_SLICE_X11Y144_CO6),
.Q(CLBLM_L_X8Y144_SLICE_X11Y144_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y144_SLICE_X11Y144_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y144_SLICE_X11Y144_DO6),
.Q(CLBLM_L_X8Y144_SLICE_X11Y144_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hbbb8bbb888888888)
  ) CLBLM_L_X8Y144_SLICE_X11Y144_DLUT (
.I0(CLBLM_L_X8Y142_SLICE_X11Y142_BQ),
.I1(LIOB33_X0Y61_IOB_X0Y62_I),
.I2(CLBLM_L_X8Y144_SLICE_X11Y144_DQ),
.I3(CLBLM_R_X7Y142_SLICE_X9Y142_AQ),
.I4(1'b1),
.I5(CLBLM_L_X12Y149_SLICE_X17Y149_CO6),
.O5(CLBLM_L_X8Y144_SLICE_X11Y144_DO5),
.O6(CLBLM_L_X8Y144_SLICE_X11Y144_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hffac00acffac00ac)
  ) CLBLM_L_X8Y144_SLICE_X11Y144_CLUT (
.I0(CLBLL_L_X4Y142_SLICE_X5Y142_AQ),
.I1(CLBLM_L_X8Y144_SLICE_X11Y144_CQ),
.I2(CLBLM_R_X13Y149_SLICE_X18Y149_AO6),
.I3(LIOB33_X0Y61_IOB_X0Y62_I),
.I4(CLBLM_L_X10Y146_SLICE_X12Y146_DQ),
.I5(1'b1),
.O5(CLBLM_L_X8Y144_SLICE_X11Y144_CO5),
.O6(CLBLM_L_X8Y144_SLICE_X11Y144_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hbbbb8888f3f3c0c0)
  ) CLBLM_L_X8Y144_SLICE_X11Y144_BLUT (
.I0(CLBLM_L_X10Y142_SLICE_X12Y142_AQ),
.I1(LIOB33_X0Y61_IOB_X0Y62_I),
.I2(CLBLM_R_X7Y143_SLICE_X9Y143_AQ),
.I3(1'b1),
.I4(CLBLM_L_X10Y149_SLICE_X13Y149_AQ),
.I5(1'b1),
.O5(CLBLM_L_X8Y144_SLICE_X11Y144_BO5),
.O6(CLBLM_L_X8Y144_SLICE_X11Y144_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h8dd888888dd88888)
  ) CLBLM_L_X8Y144_SLICE_X11Y144_ALUT (
.I0(LIOB33_X0Y61_IOB_X0Y62_I),
.I1(CLBLM_R_X7Y146_SLICE_X9Y146_AQ),
.I2(CLBLM_L_X8Y144_SLICE_X11Y144_AQ),
.I3(CLBLM_L_X10Y143_SLICE_X13Y143_DO6),
.I4(CLBLM_L_X10Y144_SLICE_X12Y144_AO6),
.I5(1'b1),
.O5(CLBLM_L_X8Y144_SLICE_X11Y144_AO5),
.O6(CLBLM_L_X8Y144_SLICE_X11Y144_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y145_SLICE_X10Y145_A5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y145_SLICE_X10Y145_AO5),
.Q(CLBLM_L_X8Y145_SLICE_X10Y145_A5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y145_SLICE_X10Y145_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y145_SLICE_X10Y145_AO6),
.Q(CLBLM_L_X8Y145_SLICE_X10Y145_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hf3f0f7f5f3f0f3f0)
  ) CLBLM_L_X8Y145_SLICE_X10Y145_DLUT (
.I0(CLBLL_L_X4Y148_SLICE_X4Y148_CQ),
.I1(CLBLM_L_X10Y148_SLICE_X12Y148_AO5),
.I2(CLBLM_R_X7Y145_SLICE_X9Y145_CO6),
.I3(CLBLM_R_X7Y142_SLICE_X8Y142_DQ),
.I4(CLBLM_L_X12Y146_SLICE_X16Y146_CO6),
.I5(CLBLL_L_X4Y149_SLICE_X5Y149_C5Q),
.O5(CLBLM_L_X8Y145_SLICE_X10Y145_DO5),
.O6(CLBLM_L_X8Y145_SLICE_X10Y145_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hcecececececeffce)
  ) CLBLM_L_X8Y145_SLICE_X10Y145_CLUT (
.I0(CLBLM_L_X8Y144_SLICE_X11Y144_BQ),
.I1(CLBLM_R_X7Y145_SLICE_X9Y145_BO6),
.I2(CLBLM_L_X10Y148_SLICE_X12Y148_AO5),
.I3(CLBLM_L_X10Y149_SLICE_X13Y149_AQ),
.I4(CLBLM_L_X12Y146_SLICE_X16Y146_CO6),
.I5(CLBLL_L_X4Y148_SLICE_X4Y148_CQ),
.O5(CLBLM_L_X8Y145_SLICE_X10Y145_CO5),
.O6(CLBLM_L_X8Y145_SLICE_X10Y145_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffffaaeeafef)
  ) CLBLM_L_X8Y145_SLICE_X10Y145_BLUT (
.I0(CLBLM_R_X7Y144_SLICE_X9Y144_DO6),
.I1(CLBLM_R_X7Y144_SLICE_X9Y144_BQ),
.I2(CLBLM_L_X8Y146_SLICE_X10Y146_AO6),
.I3(CLBLM_L_X10Y148_SLICE_X12Y148_AO5),
.I4(CLBLM_L_X12Y151_SLICE_X16Y151_AQ),
.I5(CLBLM_L_X8Y144_SLICE_X10Y144_CO6),
.O5(CLBLM_L_X8Y145_SLICE_X10Y145_BO5),
.O6(CLBLM_L_X8Y145_SLICE_X10Y145_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hff00f0f0aaaa3c3c)
  ) CLBLM_L_X8Y145_SLICE_X10Y145_ALUT (
.I0(CLBLM_L_X10Y143_SLICE_X12Y143_BQ),
.I1(CLBLM_L_X8Y144_SLICE_X11Y144_B5Q),
.I2(CLBLM_R_X3Y145_SLICE_X3Y145_BQ),
.I3(CLBLL_L_X4Y146_SLICE_X5Y146_AQ),
.I4(LIOB33_X0Y61_IOB_X0Y62_I),
.I5(1'b1),
.O5(CLBLM_L_X8Y145_SLICE_X10Y145_AO5),
.O6(CLBLM_L_X8Y145_SLICE_X10Y145_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y145_SLICE_X11Y145_C5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y145_SLICE_X11Y145_CO5),
.Q(CLBLM_L_X8Y145_SLICE_X11Y145_C5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y145_SLICE_X11Y145_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y145_SLICE_X11Y145_AO6),
.Q(CLBLM_L_X8Y145_SLICE_X11Y145_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y145_SLICE_X11Y145_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y145_SLICE_X11Y145_BO6),
.Q(CLBLM_L_X8Y145_SLICE_X11Y145_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y145_SLICE_X11Y145_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y145_SLICE_X11Y145_CO6),
.Q(CLBLM_L_X8Y145_SLICE_X11Y145_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y145_SLICE_X11Y145_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y145_SLICE_X11Y145_DO6),
.Q(CLBLM_L_X8Y145_SLICE_X11Y145_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hfefecccc32320000)
  ) CLBLM_L_X8Y145_SLICE_X11Y145_DLUT (
.I0(CLBLM_L_X10Y144_SLICE_X12Y144_CO6),
.I1(LIOB33_X0Y61_IOB_X0Y62_I),
.I2(CLBLM_L_X8Y145_SLICE_X11Y145_DQ),
.I3(1'b1),
.I4(CLBLM_R_X7Y152_SLICE_X9Y152_DO6),
.I5(CLBLM_L_X8Y145_SLICE_X11Y145_AQ),
.O5(CLBLM_L_X8Y145_SLICE_X11Y145_DO5),
.O6(CLBLM_L_X8Y145_SLICE_X11Y145_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hffcc00ccf0aaf0aa)
  ) CLBLM_L_X8Y145_SLICE_X11Y145_CLUT (
.I0(RIOB33_X105Y117_IOB_X1Y118_I),
.I1(CLBLM_L_X10Y149_SLICE_X13Y149_AQ),
.I2(CLBLM_L_X8Y144_SLICE_X11Y144_DQ),
.I3(LIOB33_X0Y61_IOB_X0Y62_I),
.I4(CLBLM_L_X8Y153_SLICE_X10Y153_D5Q),
.I5(1'b1),
.O5(CLBLM_L_X8Y145_SLICE_X11Y145_CO5),
.O6(CLBLM_L_X8Y145_SLICE_X11Y145_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfc0cfe0efc0cf404)
  ) CLBLM_L_X8Y145_SLICE_X11Y145_BLUT (
.I0(CLBLM_L_X10Y144_SLICE_X13Y144_CQ),
.I1(CLBLM_L_X8Y145_SLICE_X11Y145_BQ),
.I2(LIOB33_X0Y61_IOB_X0Y62_I),
.I3(CLBLL_L_X4Y146_SLICE_X5Y146_BQ),
.I4(CLBLM_L_X8Y147_SLICE_X10Y147_C5Q),
.I5(CLBLM_R_X3Y145_SLICE_X3Y145_DQ),
.O5(CLBLM_L_X8Y145_SLICE_X11Y145_BO5),
.O6(CLBLM_L_X8Y145_SLICE_X11Y145_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hacacafafaca0afa0)
  ) CLBLM_L_X8Y145_SLICE_X11Y145_ALUT (
.I0(CLBLM_R_X7Y145_SLICE_X8Y145_D5Q),
.I1(CLBLM_R_X7Y152_SLICE_X8Y152_D5Q),
.I2(LIOB33_X0Y61_IOB_X0Y62_I),
.I3(CLBLM_L_X8Y145_SLICE_X11Y145_AQ),
.I4(CLBLM_R_X7Y142_SLICE_X8Y142_C5Q),
.I5(CLBLM_L_X8Y145_SLICE_X10Y145_AQ),
.O5(CLBLM_L_X8Y145_SLICE_X11Y145_AO5),
.O6(CLBLM_L_X8Y145_SLICE_X11Y145_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y146_SLICE_X10Y146_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(LIOB33_X0Y61_IOB_X0Y62_I),
.D(CLBLM_R_X5Y142_SLICE_X7Y142_A5Q),
.Q(CLBLM_L_X8Y146_SLICE_X10Y146_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y146_SLICE_X10Y146_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(LIOB33_X0Y61_IOB_X0Y62_I),
.D(CLBLM_L_X8Y145_SLICE_X10Y145_A5Q),
.Q(CLBLM_L_X8Y146_SLICE_X10Y146_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0fcf00ccafefaaee)
  ) CLBLM_L_X8Y146_SLICE_X10Y146_DLUT (
.I0(CLBLM_R_X5Y140_SLICE_X6Y140_A5Q),
.I1(CLBLM_R_X5Y150_SLICE_X7Y150_A5Q),
.I2(CLBLM_R_X11Y146_SLICE_X14Y146_CO6),
.I3(CLBLM_L_X8Y146_SLICE_X10Y146_AO5),
.I4(CLBLM_R_X5Y143_SLICE_X6Y143_CQ),
.I5(CLBLM_R_X7Y146_SLICE_X9Y146_DO6),
.O5(CLBLM_L_X8Y146_SLICE_X10Y146_DO5),
.O6(CLBLM_L_X8Y146_SLICE_X10Y146_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h3bff3b3b0aff0a0a)
  ) CLBLM_L_X8Y146_SLICE_X10Y146_CLUT (
.I0(CLBLM_L_X8Y144_SLICE_X10Y144_AQ),
.I1(CLBLM_L_X8Y146_SLICE_X10Y146_AO6),
.I2(CLBLM_R_X11Y146_SLICE_X14Y146_CO6),
.I3(CLBLM_L_X10Y148_SLICE_X12Y148_AO5),
.I4(CLBLM_R_X7Y148_SLICE_X9Y148_A5Q),
.I5(CLBLM_L_X10Y149_SLICE_X12Y149_BQ),
.O5(CLBLM_L_X8Y146_SLICE_X10Y146_CO5),
.O6(CLBLM_L_X8Y146_SLICE_X10Y146_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff0ace0ace0ace)
  ) CLBLM_L_X8Y146_SLICE_X10Y146_BLUT (
.I0(CLBLM_R_X7Y144_SLICE_X8Y144_DQ),
.I1(CLBLL_L_X4Y142_SLICE_X5Y142_C5Q),
.I2(CLBLM_L_X8Y146_SLICE_X10Y146_AO5),
.I3(CLBLM_R_X7Y146_SLICE_X9Y146_DO6),
.I4(CLBLM_L_X8Y146_SLICE_X10Y146_CO6),
.I5(1'b1),
.O5(CLBLM_L_X8Y146_SLICE_X10Y146_BO5),
.O6(CLBLM_L_X8Y146_SLICE_X10Y146_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffbfffffeffffff)
  ) CLBLM_L_X8Y146_SLICE_X10Y146_ALUT (
.I0(CLBLM_R_X7Y153_SLICE_X8Y153_A5Q),
.I1(CLBLM_R_X7Y149_SLICE_X8Y149_AQ),
.I2(CLBLM_R_X7Y146_SLICE_X9Y146_CO6),
.I3(CLBLL_L_X4Y148_SLICE_X4Y148_CQ),
.I4(CLBLM_R_X7Y144_SLICE_X9Y144_B5Q),
.I5(1'b1),
.O5(CLBLM_L_X8Y146_SLICE_X10Y146_AO5),
.O6(CLBLM_L_X8Y146_SLICE_X10Y146_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y146_SLICE_X11Y146_B5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y146_SLICE_X11Y146_BO5),
.Q(CLBLM_L_X8Y146_SLICE_X11Y146_B5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "C5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y146_SLICE_X11Y146_C5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y146_SLICE_X11Y146_CO5),
.Q(CLBLM_L_X8Y146_SLICE_X11Y146_C5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y146_SLICE_X11Y146_D5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y146_SLICE_X11Y146_DO5),
.Q(CLBLM_L_X8Y146_SLICE_X11Y146_D5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y146_SLICE_X11Y146_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y146_SLICE_X11Y146_AO6),
.Q(CLBLM_L_X8Y146_SLICE_X11Y146_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y146_SLICE_X11Y146_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y146_SLICE_X11Y146_BO6),
.Q(CLBLM_L_X8Y146_SLICE_X11Y146_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y146_SLICE_X11Y146_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y146_SLICE_X11Y146_CO6),
.Q(CLBLM_L_X8Y146_SLICE_X11Y146_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y146_SLICE_X11Y146_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y146_SLICE_X11Y146_DO6),
.Q(CLBLM_L_X8Y146_SLICE_X11Y146_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hff006666f0f0cccc)
  ) CLBLM_L_X8Y146_SLICE_X11Y146_DLUT (
.I0(CLBLM_L_X8Y148_SLICE_X11Y148_BQ),
.I1(CLBLM_R_X5Y152_SLICE_X6Y152_CQ),
.I2(CLBLL_L_X4Y142_SLICE_X5Y142_AQ),
.I3(CLBLM_L_X10Y146_SLICE_X13Y146_CQ),
.I4(LIOB33_X0Y61_IOB_X0Y62_I),
.I5(1'b1),
.O5(CLBLM_L_X8Y146_SLICE_X11Y146_DO5),
.O6(CLBLM_L_X8Y146_SLICE_X11Y146_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0ccf0ccccf0ccaa)
  ) CLBLM_L_X8Y146_SLICE_X11Y146_CLUT (
.I0(CLBLM_L_X8Y146_SLICE_X11Y146_C5Q),
.I1(CLBLM_R_X3Y145_SLICE_X3Y145_BQ),
.I2(CLBLM_L_X8Y143_SLICE_X11Y143_AQ),
.I3(LIOB33_X0Y61_IOB_X0Y62_I),
.I4(CLBLM_R_X13Y149_SLICE_X18Y149_AO6),
.I5(1'b1),
.O5(CLBLM_L_X8Y146_SLICE_X11Y146_CO5),
.O6(CLBLM_L_X8Y146_SLICE_X11Y146_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hdddd8888e4e4e4e4)
  ) CLBLM_L_X8Y146_SLICE_X11Y146_BLUT (
.I0(LIOB33_X0Y61_IOB_X0Y62_I),
.I1(CLBLM_L_X8Y147_SLICE_X11Y147_C5Q),
.I2(CLBLM_R_X7Y146_SLICE_X8Y146_D5Q),
.I3(1'b1),
.I4(CLBLM_R_X7Y153_SLICE_X9Y153_C5Q),
.I5(1'b1),
.O5(CLBLM_L_X8Y146_SLICE_X11Y146_BO5),
.O6(CLBLM_L_X8Y146_SLICE_X11Y146_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hdddd8888d8d8d8d8)
  ) CLBLM_L_X8Y146_SLICE_X11Y146_ALUT (
.I0(LIOB33_X0Y61_IOB_X0Y62_I),
.I1(CLBLM_L_X8Y146_SLICE_X11Y146_BQ),
.I2(CLBLM_L_X8Y146_SLICE_X11Y146_AQ),
.I3(1'b1),
.I4(CLBLM_R_X7Y146_SLICE_X9Y146_AQ),
.I5(CLBLM_R_X11Y146_SLICE_X14Y146_DO6),
.O5(CLBLM_L_X8Y146_SLICE_X11Y146_AO5),
.O6(CLBLM_L_X8Y146_SLICE_X11Y146_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y147_SLICE_X10Y147_C5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y147_SLICE_X10Y147_CO5),
.Q(CLBLM_L_X8Y147_SLICE_X10Y147_C5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y147_SLICE_X10Y147_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y147_SLICE_X10Y147_AO6),
.Q(CLBLM_L_X8Y147_SLICE_X10Y147_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y147_SLICE_X10Y147_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y147_SLICE_X10Y147_BO6),
.Q(CLBLM_L_X8Y147_SLICE_X10Y147_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y147_SLICE_X10Y147_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y147_SLICE_X10Y147_CO6),
.Q(CLBLM_L_X8Y147_SLICE_X10Y147_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffff00aaccee)
  ) CLBLM_L_X8Y147_SLICE_X10Y147_DLUT (
.I0(CLBLM_R_X7Y146_SLICE_X8Y146_B5Q),
.I1(CLBLM_L_X8Y147_SLICE_X10Y147_AQ),
.I2(1'b1),
.I3(CLBLM_R_X7Y148_SLICE_X8Y148_AO5),
.I4(CLBLM_L_X8Y150_SLICE_X11Y150_BO5),
.I5(CLBLM_L_X8Y144_SLICE_X10Y144_DO6),
.O5(CLBLM_L_X8Y147_SLICE_X10Y147_DO5),
.O6(CLBLM_L_X8Y147_SLICE_X10Y147_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'heeee2222ee22ee22)
  ) CLBLM_L_X8Y147_SLICE_X10Y147_CLUT (
.I0(RIOB33_X105Y111_IOB_X1Y112_I),
.I1(LIOB33_X0Y61_IOB_X0Y62_I),
.I2(1'b1),
.I3(CLBLM_L_X10Y146_SLICE_X12Y146_CQ),
.I4(CLBLM_L_X8Y151_SLICE_X10Y151_B5Q),
.I5(1'b1),
.O5(CLBLM_L_X8Y147_SLICE_X10Y147_CO5),
.O6(CLBLM_L_X8Y147_SLICE_X10Y147_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'haaffaaffaa00aaff)
  ) CLBLM_L_X8Y147_SLICE_X10Y147_BLUT (
.I0(CLBLM_L_X8Y147_SLICE_X11Y147_DQ),
.I1(1'b1),
.I2(1'b1),
.I3(LIOB33_X0Y61_IOB_X0Y62_I),
.I4(CLBLM_R_X5Y143_SLICE_X6Y143_BQ),
.I5(CLBLM_R_X3Y147_SLICE_X3Y147_DO6),
.O5(CLBLM_L_X8Y147_SLICE_X10Y147_BO5),
.O6(CLBLM_L_X8Y147_SLICE_X10Y147_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hccffcc00ccf0ccf0)
  ) CLBLM_L_X8Y147_SLICE_X10Y147_ALUT (
.I0(1'b1),
.I1(CLBLM_R_X7Y149_SLICE_X9Y149_BQ),
.I2(CLBLM_L_X8Y147_SLICE_X10Y147_AQ),
.I3(LIOB33_X0Y61_IOB_X0Y62_I),
.I4(CLBLM_L_X8Y145_SLICE_X11Y145_AQ),
.I5(CLBLM_R_X13Y149_SLICE_X18Y149_AO6),
.O5(CLBLM_L_X8Y147_SLICE_X10Y147_AO5),
.O6(CLBLM_L_X8Y147_SLICE_X10Y147_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y147_SLICE_X11Y147_C5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y147_SLICE_X11Y147_CO5),
.Q(CLBLM_L_X8Y147_SLICE_X11Y147_C5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y147_SLICE_X11Y147_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y147_SLICE_X11Y147_AO6),
.Q(CLBLM_L_X8Y147_SLICE_X11Y147_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y147_SLICE_X11Y147_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y147_SLICE_X11Y147_BO6),
.Q(CLBLM_L_X8Y147_SLICE_X11Y147_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y147_SLICE_X11Y147_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y147_SLICE_X11Y147_CO6),
.Q(CLBLM_L_X8Y147_SLICE_X11Y147_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y147_SLICE_X11Y147_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y147_SLICE_X11Y147_DO6),
.Q(CLBLM_L_X8Y147_SLICE_X11Y147_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hffaafff000aa00f0)
  ) CLBLM_L_X8Y147_SLICE_X11Y147_DLUT (
.I0(CLBLM_L_X10Y146_SLICE_X12Y146_BQ),
.I1(1'b1),
.I2(CLBLM_L_X8Y147_SLICE_X11Y147_DQ),
.I3(LIOB33_X0Y61_IOB_X0Y62_I),
.I4(CLBLM_R_X11Y148_SLICE_X15Y148_AO6),
.I5(CLBLL_L_X4Y144_SLICE_X5Y144_D5Q),
.O5(CLBLM_L_X8Y147_SLICE_X11Y147_DO5),
.O6(CLBLM_L_X8Y147_SLICE_X11Y147_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hdd11dd11dddd1111)
  ) CLBLM_L_X8Y147_SLICE_X11Y147_CLUT (
.I0(CLBLM_L_X10Y153_SLICE_X13Y153_A5Q),
.I1(LIOB33_X0Y61_IOB_X0Y62_I),
.I2(1'b1),
.I3(CLBLM_L_X8Y145_SLICE_X10Y145_AQ),
.I4(CLBLM_R_X7Y153_SLICE_X9Y153_A5Q),
.I5(1'b1),
.O5(CLBLM_L_X8Y147_SLICE_X11Y147_CO5),
.O6(CLBLM_L_X8Y147_SLICE_X11Y147_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hff00ff00eeee0e0e)
  ) CLBLM_L_X8Y147_SLICE_X11Y147_BLUT (
.I0(CLBLM_L_X8Y148_SLICE_X10Y148_B5Q),
.I1(CLBLM_L_X8Y147_SLICE_X11Y147_BQ),
.I2(CLBLM_R_X7Y142_SLICE_X8Y142_C5Q),
.I3(CLBLM_R_X5Y146_SLICE_X7Y146_BQ),
.I4(CLBLM_R_X7Y152_SLICE_X8Y152_D5Q),
.I5(LIOB33_X0Y61_IOB_X0Y62_I),
.O5(CLBLM_L_X8Y147_SLICE_X11Y147_BO5),
.O6(CLBLM_L_X8Y147_SLICE_X11Y147_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffb800b8ffb800b8)
  ) CLBLM_L_X8Y147_SLICE_X11Y147_ALUT (
.I0(CLBLM_R_X3Y148_SLICE_X3Y148_AQ),
.I1(CLBLM_R_X11Y146_SLICE_X14Y146_DO6),
.I2(CLBLM_L_X8Y147_SLICE_X11Y147_AQ),
.I3(LIOB33_X0Y61_IOB_X0Y62_I),
.I4(CLBLM_R_X5Y151_SLICE_X6Y151_AQ),
.I5(1'b1),
.O5(CLBLM_L_X8Y147_SLICE_X11Y147_AO5),
.O6(CLBLM_L_X8Y147_SLICE_X11Y147_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y148_SLICE_X10Y148_B5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y148_SLICE_X10Y148_BO5),
.Q(CLBLM_L_X8Y148_SLICE_X10Y148_B5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y148_SLICE_X10Y148_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y148_SLICE_X10Y148_AO6),
.Q(CLBLM_L_X8Y148_SLICE_X10Y148_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y148_SLICE_X10Y148_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y148_SLICE_X10Y148_BO6),
.Q(CLBLM_L_X8Y148_SLICE_X10Y148_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h30ff3030baffbaba)
  ) CLBLM_L_X8Y148_SLICE_X10Y148_DLUT (
.I0(CLBLM_R_X5Y151_SLICE_X6Y151_AQ),
.I1(CLBLM_R_X7Y148_SLICE_X8Y148_AO5),
.I2(CLBLM_L_X8Y153_SLICE_X10Y153_DQ),
.I3(CLBLM_R_X7Y148_SLICE_X8Y148_AO6),
.I4(CLBLM_L_X8Y153_SLICE_X10Y153_D5Q),
.I5(CLBLM_L_X8Y150_SLICE_X11Y150_BO6),
.O5(CLBLM_L_X8Y148_SLICE_X10Y148_DO5),
.O6(CLBLM_L_X8Y148_SLICE_X10Y148_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'habaaabaaffffabaa)
  ) CLBLM_L_X8Y148_SLICE_X10Y148_CLUT (
.I0(CLBLM_R_X7Y148_SLICE_X9Y148_DO6),
.I1(CLBLM_L_X12Y146_SLICE_X16Y146_CO6),
.I2(CLBLL_L_X4Y148_SLICE_X4Y148_CQ),
.I3(CLBLM_R_X3Y146_SLICE_X2Y146_D5Q),
.I4(CLBLM_R_X3Y149_SLICE_X3Y149_DQ),
.I5(CLBLM_L_X8Y146_SLICE_X10Y146_AO5),
.O5(CLBLM_L_X8Y148_SLICE_X10Y148_CO5),
.O6(CLBLM_L_X8Y148_SLICE_X10Y148_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h88bbbb88f3c0f3c0)
  ) CLBLM_L_X8Y148_SLICE_X10Y148_BLUT (
.I0(CLBLM_R_X7Y148_SLICE_X9Y148_CQ),
.I1(LIOB33_X0Y61_IOB_X0Y62_I),
.I2(CLBLM_L_X8Y147_SLICE_X10Y147_CQ),
.I3(CLBLM_R_X5Y152_SLICE_X6Y152_CQ),
.I4(CLBLM_R_X5Y146_SLICE_X6Y146_B5Q),
.I5(1'b1),
.O5(CLBLM_L_X8Y148_SLICE_X10Y148_BO5),
.O6(CLBLM_L_X8Y148_SLICE_X10Y148_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff0000c8c8c8c8)
  ) CLBLM_L_X8Y148_SLICE_X10Y148_ALUT (
.I0(CLBLM_L_X10Y146_SLICE_X12Y146_CQ),
.I1(CLBLM_R_X13Y149_SLICE_X18Y149_AO6),
.I2(CLBLM_L_X8Y148_SLICE_X10Y148_AQ),
.I3(1'b1),
.I4(CLBLL_L_X2Y148_SLICE_X0Y148_AQ),
.I5(LIOB33_X0Y61_IOB_X0Y62_I),
.O5(CLBLM_L_X8Y148_SLICE_X10Y148_AO5),
.O6(CLBLM_L_X8Y148_SLICE_X10Y148_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y148_SLICE_X11Y148_B5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y148_SLICE_X11Y148_BO5),
.Q(CLBLM_L_X8Y148_SLICE_X11Y148_B5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y148_SLICE_X11Y148_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y148_SLICE_X11Y148_AO6),
.Q(CLBLM_L_X8Y148_SLICE_X11Y148_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y148_SLICE_X11Y148_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y148_SLICE_X11Y148_BO6),
.Q(CLBLM_L_X8Y148_SLICE_X11Y148_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hccfcccfcffffccfc)
  ) CLBLM_L_X8Y148_SLICE_X11Y148_DLUT (
.I0(1'b1),
.I1(CLBLM_L_X10Y148_SLICE_X12Y148_BO6),
.I2(CLBLM_L_X8Y148_SLICE_X11Y148_BQ),
.I3(CLBLM_R_X7Y148_SLICE_X8Y148_AO5),
.I4(CLBLM_L_X8Y144_SLICE_X11Y144_CQ),
.I5(CLBLM_L_X8Y150_SLICE_X11Y150_BO6),
.O5(CLBLM_L_X8Y148_SLICE_X11Y148_DO5),
.O6(CLBLM_L_X8Y148_SLICE_X11Y148_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0fcf00ccafefaaee)
  ) CLBLM_L_X8Y148_SLICE_X11Y148_CLUT (
.I0(CLBLM_R_X5Y149_SLICE_X6Y149_BQ),
.I1(CLBLM_L_X8Y147_SLICE_X11Y147_DQ),
.I2(CLBLM_L_X12Y149_SLICE_X17Y149_BO5),
.I3(CLBLM_L_X10Y151_SLICE_X13Y151_BO6),
.I4(CLBLM_R_X7Y143_SLICE_X8Y143_BQ),
.I5(CLBLM_L_X10Y148_SLICE_X12Y148_AO6),
.O5(CLBLM_L_X8Y148_SLICE_X11Y148_CO5),
.O6(CLBLM_L_X8Y148_SLICE_X11Y148_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hffcc00ccf0aaf0aa)
  ) CLBLM_L_X8Y148_SLICE_X11Y148_BLUT (
.I0(CLBLM_R_X5Y153_SLICE_X6Y153_A5Q),
.I1(CLBLL_L_X4Y149_SLICE_X5Y149_C5Q),
.I2(CLBLM_L_X8Y147_SLICE_X11Y147_BQ),
.I3(LIOB33_X0Y61_IOB_X0Y62_I),
.I4(CLBLM_L_X8Y145_SLICE_X11Y145_BQ),
.I5(1'b1),
.O5(CLBLM_L_X8Y148_SLICE_X11Y148_BO5),
.O6(CLBLM_L_X8Y148_SLICE_X11Y148_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hcccccccca0aaaaa0)
  ) CLBLM_L_X8Y148_SLICE_X11Y148_ALUT (
.I0(CLBLM_R_X7Y151_SLICE_X9Y151_A5Q),
.I1(CLBLM_R_X7Y147_SLICE_X9Y147_D5Q),
.I2(CLBLM_L_X8Y148_SLICE_X11Y148_AQ),
.I3(RIOB33_X105Y111_IOB_X1Y112_I),
.I4(CLBLM_L_X8Y147_SLICE_X10Y147_CQ),
.I5(LIOB33_X0Y61_IOB_X0Y62_I),
.O5(CLBLM_L_X8Y148_SLICE_X11Y148_AO5),
.O6(CLBLM_L_X8Y148_SLICE_X11Y148_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y149_SLICE_X10Y149_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(LIOB33_X0Y61_IOB_X0Y62_I),
.D(CLBLM_R_X5Y149_SLICE_X6Y149_BQ),
.Q(CLBLM_L_X8Y149_SLICE_X10Y149_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffff00f0aafa)
  ) CLBLM_L_X8Y149_SLICE_X10Y149_DLUT (
.I0(CLBLM_L_X8Y148_SLICE_X10Y148_AQ),
.I1(1'b1),
.I2(CLBLL_L_X4Y150_SLICE_X4Y150_AQ),
.I3(CLBLM_L_X8Y150_SLICE_X10Y150_BO5),
.I4(CLBLM_L_X8Y150_SLICE_X11Y150_BO6),
.I5(CLBLM_R_X7Y149_SLICE_X9Y149_DO6),
.O5(CLBLM_L_X8Y149_SLICE_X10Y149_DO5),
.O6(CLBLM_L_X8Y149_SLICE_X10Y149_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0100313001000100)
  ) CLBLM_L_X8Y149_SLICE_X10Y149_CLUT (
.I0(CLBLM_R_X11Y144_SLICE_X14Y144_BO6),
.I1(CLBLM_R_X7Y144_SLICE_X9Y144_B5Q),
.I2(CLBLM_R_X7Y153_SLICE_X8Y153_A5Q),
.I3(CLBLM_R_X5Y145_SLICE_X7Y145_A5Q),
.I4(CLBLM_R_X11Y147_SLICE_X15Y147_BO6),
.I5(CLBLM_R_X7Y151_SLICE_X8Y151_C5Q),
.O5(CLBLM_L_X8Y149_SLICE_X10Y149_CO5),
.O6(CLBLM_L_X8Y149_SLICE_X10Y149_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000100000000)
  ) CLBLM_L_X8Y149_SLICE_X10Y149_BLUT (
.I0(CLBLM_R_X7Y144_SLICE_X9Y144_B5Q),
.I1(CLBLM_R_X7Y153_SLICE_X8Y153_A5Q),
.I2(CLBLM_L_X12Y147_SLICE_X16Y147_DO6),
.I3(CLBLM_R_X7Y149_SLICE_X8Y149_AQ),
.I4(CLBLM_L_X10Y146_SLICE_X13Y146_DO6),
.I5(CLBLL_L_X4Y148_SLICE_X4Y148_CQ),
.O5(CLBLM_L_X8Y149_SLICE_X10Y149_BO5),
.O6(CLBLM_L_X8Y149_SLICE_X10Y149_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0aff0a0aceffcece)
  ) CLBLM_L_X8Y149_SLICE_X10Y149_ALUT (
.I0(CLBLL_L_X4Y146_SLICE_X4Y146_CQ),
.I1(CLBLM_R_X5Y149_SLICE_X6Y149_C5Q),
.I2(CLBLM_L_X8Y150_SLICE_X10Y150_BO5),
.I3(CLBLM_L_X8Y149_SLICE_X10Y149_BO6),
.I4(CLBLL_L_X4Y143_SLICE_X5Y143_AQ),
.I5(CLBLM_L_X10Y150_SLICE_X12Y150_BO6),
.O5(CLBLM_L_X8Y149_SLICE_X10Y149_AO5),
.O6(CLBLM_L_X8Y149_SLICE_X10Y149_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y149_SLICE_X11Y149_A5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y149_SLICE_X11Y149_AO5),
.Q(CLBLM_L_X8Y149_SLICE_X11Y149_A5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y149_SLICE_X11Y149_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y149_SLICE_X11Y149_AO6),
.Q(CLBLM_L_X8Y149_SLICE_X11Y149_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f0fff0fafafffa)
  ) CLBLM_L_X8Y149_SLICE_X11Y149_DLUT (
.I0(CLBLM_L_X8Y143_SLICE_X10Y143_CQ),
.I1(1'b1),
.I2(CLBLM_L_X8Y151_SLICE_X10Y151_DO6),
.I3(CLBLM_L_X8Y144_SLICE_X11Y144_DQ),
.I4(CLBLM_L_X12Y149_SLICE_X17Y149_BO5),
.I5(CLBLM_R_X11Y148_SLICE_X15Y148_AO6),
.O5(CLBLM_L_X8Y149_SLICE_X11Y149_DO5),
.O6(CLBLM_L_X8Y149_SLICE_X11Y149_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hcceecceefcfefcfe)
  ) CLBLM_L_X8Y149_SLICE_X11Y149_CLUT (
.I0(CLBLM_R_X5Y148_SLICE_X6Y148_AQ),
.I1(CLBLM_L_X8Y149_SLICE_X10Y149_CO6),
.I2(CLBLM_L_X10Y151_SLICE_X12Y151_CQ),
.I3(CLBLM_L_X10Y151_SLICE_X13Y151_BO5),
.I4(1'b1),
.I5(CLBLM_L_X10Y151_SLICE_X13Y151_BO6),
.O5(CLBLM_L_X8Y149_SLICE_X11Y149_CO5),
.O6(CLBLM_L_X8Y149_SLICE_X11Y149_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000001000000033)
  ) CLBLM_L_X8Y149_SLICE_X11Y149_BLUT (
.I0(CLBLM_L_X8Y145_SLICE_X10Y145_DO6),
.I1(CLBLM_L_X8Y148_SLICE_X11Y148_DO6),
.I2(CLBLM_R_X11Y147_SLICE_X15Y147_DO6),
.I3(CLBLM_L_X8Y150_SLICE_X11Y150_CO6),
.I4(CLBLM_L_X8Y151_SLICE_X11Y151_DO6),
.I5(CLBLM_L_X12Y147_SLICE_X16Y147_DO6),
.O5(CLBLM_L_X8Y149_SLICE_X11Y149_BO5),
.O6(CLBLM_L_X8Y149_SLICE_X11Y149_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfafa0a0afc0cfc0c)
  ) CLBLM_L_X8Y149_SLICE_X11Y149_ALUT (
.I0(CLBLM_R_X7Y149_SLICE_X9Y149_B5Q),
.I1(RIOB33_SING_X105Y100_IOB_X1Y100_I),
.I2(LIOB33_X0Y61_IOB_X0Y62_I),
.I3(CLBLM_L_X8Y146_SLICE_X11Y146_CQ),
.I4(CLBLL_L_X4Y148_SLICE_X4Y148_BQ),
.I5(1'b1),
.O5(CLBLM_L_X8Y149_SLICE_X11Y149_AO5),
.O6(CLBLM_L_X8Y149_SLICE_X11Y149_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y150_SLICE_X10Y150_A_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_L_X8Y150_SLICE_X10Y150_AO6),
.Q(CLBLM_L_X8Y150_SLICE_X10Y150_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hafefafefaaeeaaee)
  ) CLBLM_L_X8Y150_SLICE_X10Y150_DLUT (
.I0(CLBLM_L_X8Y150_SLICE_X10Y150_CO6),
.I1(CLBLM_L_X8Y153_SLICE_X10Y153_BQ),
.I2(CLBLM_L_X8Y150_SLICE_X11Y150_BO5),
.I3(CLBLM_R_X7Y148_SLICE_X8Y148_AO5),
.I4(1'b1),
.I5(CLBLM_L_X8Y150_SLICE_X10Y150_AQ),
.O5(CLBLM_L_X8Y150_SLICE_X10Y150_DO5),
.O6(CLBLM_L_X8Y150_SLICE_X10Y150_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h000000000000f5a0)
  ) CLBLM_L_X8Y150_SLICE_X10Y150_CLUT (
.I0(CLBLM_R_X7Y144_SLICE_X9Y144_B5Q),
.I1(1'b1),
.I2(CLBLM_L_X8Y153_SLICE_X10Y153_B5Q),
.I3(CLBLL_L_X4Y145_SLICE_X4Y145_CQ),
.I4(CLBLM_R_X7Y153_SLICE_X8Y153_A5Q),
.I5(CLBLM_R_X11Y144_SLICE_X14Y144_AO6),
.O5(CLBLM_L_X8Y150_SLICE_X10Y150_CO5),
.O6(CLBLM_L_X8Y150_SLICE_X10Y150_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffffdffffff7f)
  ) CLBLM_L_X8Y150_SLICE_X10Y150_BLUT (
.I0(CLBLM_R_X7Y153_SLICE_X8Y153_A5Q),
.I1(CLBLL_L_X4Y148_SLICE_X4Y148_CQ),
.I2(CLBLM_R_X7Y149_SLICE_X8Y149_AQ),
.I3(CLBLM_R_X7Y144_SLICE_X9Y144_B5Q),
.I4(CLBLM_L_X12Y147_SLICE_X16Y147_DO6),
.I5(1'b1),
.O5(CLBLM_L_X8Y150_SLICE_X10Y150_BO5),
.O6(CLBLM_L_X8Y150_SLICE_X10Y150_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'haaccaaccaac0aac0)
  ) CLBLM_L_X8Y150_SLICE_X10Y150_ALUT (
.I0(CLBLM_L_X10Y146_SLICE_X12Y146_BQ),
.I1(CLBLM_R_X13Y149_SLICE_X18Y149_AO6),
.I2(CLBLM_L_X8Y150_SLICE_X10Y150_AQ),
.I3(LIOB33_X0Y61_IOB_X0Y62_I),
.I4(1'b1),
.I5(CLBLM_R_X7Y151_SLICE_X9Y151_AQ),
.O5(CLBLM_L_X8Y150_SLICE_X10Y150_AO5),
.O6(CLBLM_L_X8Y150_SLICE_X10Y150_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y150_SLICE_X11Y150_A_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_L_X8Y150_SLICE_X11Y150_AO6),
.Q(CLBLM_L_X8Y150_SLICE_X11Y150_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hbfbfbbbbafafaaaa)
  ) CLBLM_L_X8Y150_SLICE_X11Y150_DLUT (
.I0(CLBLM_R_X7Y150_SLICE_X9Y150_CO6),
.I1(CLBLM_R_X11Y148_SLICE_X15Y148_AO6),
.I2(CLBLM_L_X10Y151_SLICE_X13Y151_BO5),
.I3(1'b1),
.I4(CLBLM_L_X8Y146_SLICE_X10Y146_AQ),
.I5(CLBLM_L_X8Y152_SLICE_X11Y152_BQ),
.O5(CLBLM_L_X8Y150_SLICE_X11Y150_DO5),
.O6(CLBLM_L_X8Y150_SLICE_X11Y150_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0ace0aceffff0ace)
  ) CLBLM_L_X8Y150_SLICE_X11Y150_CLUT (
.I0(CLBLL_L_X2Y148_SLICE_X0Y148_AQ),
.I1(CLBLM_R_X7Y142_SLICE_X8Y142_D5Q),
.I2(CLBLM_L_X10Y151_SLICE_X13Y151_BO5),
.I3(CLBLM_L_X10Y150_SLICE_X12Y150_BO5),
.I4(CLBLM_L_X8Y143_SLICE_X11Y143_CQ),
.I5(CLBLM_L_X12Y149_SLICE_X17Y149_BO5),
.O5(CLBLM_L_X8Y150_SLICE_X11Y150_CO5),
.O6(CLBLM_L_X8Y150_SLICE_X11Y150_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffff7fffffffbf)
  ) CLBLM_L_X8Y150_SLICE_X11Y150_BLUT (
.I0(CLBLM_R_X7Y153_SLICE_X8Y153_A5Q),
.I1(CLBLM_R_X7Y144_SLICE_X9Y144_B5Q),
.I2(CLBLM_R_X7Y149_SLICE_X8Y149_AQ),
.I3(CLBLM_L_X12Y147_SLICE_X16Y147_DO6),
.I4(CLBLL_L_X4Y148_SLICE_X4Y148_CQ),
.I5(1'b1),
.O5(CLBLM_L_X8Y150_SLICE_X11Y150_BO5),
.O6(CLBLM_L_X8Y150_SLICE_X11Y150_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'heeee2222fcee3022)
  ) CLBLM_L_X8Y150_SLICE_X11Y150_ALUT (
.I0(CLBLM_R_X7Y148_SLICE_X9Y148_CQ),
.I1(LIOB33_X0Y61_IOB_X0Y62_I),
.I2(CLBLM_L_X8Y150_SLICE_X11Y150_AQ),
.I3(CLBLM_R_X3Y145_SLICE_X3Y145_D5Q),
.I4(CLBLM_R_X11Y151_SLICE_X15Y151_AQ),
.I5(CLBLL_L_X4Y151_SLICE_X4Y151_BQ),
.O5(CLBLM_L_X8Y150_SLICE_X11Y150_AO5),
.O6(CLBLM_L_X8Y150_SLICE_X11Y150_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y151_SLICE_X10Y151_A5_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_L_X8Y151_SLICE_X10Y151_AO5),
.Q(CLBLM_L_X8Y151_SLICE_X10Y151_A5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y151_SLICE_X10Y151_B5_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_L_X8Y151_SLICE_X10Y151_BO5),
.Q(CLBLM_L_X8Y151_SLICE_X10Y151_B5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "C5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y151_SLICE_X10Y151_C5_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_L_X8Y151_SLICE_X10Y151_CO5),
.Q(CLBLM_L_X8Y151_SLICE_X10Y151_C5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y151_SLICE_X10Y151_A_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_L_X8Y151_SLICE_X10Y151_AO6),
.Q(CLBLM_L_X8Y151_SLICE_X10Y151_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y151_SLICE_X10Y151_B_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_L_X8Y151_SLICE_X10Y151_BO6),
.Q(CLBLM_L_X8Y151_SLICE_X10Y151_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y151_SLICE_X10Y151_C_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_L_X8Y151_SLICE_X10Y151_CO6),
.Q(CLBLM_L_X8Y151_SLICE_X10Y151_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000040400000500)
  ) CLBLM_L_X8Y151_SLICE_X10Y151_DLUT (
.I0(CLBLM_R_X11Y146_SLICE_X15Y146_BO6),
.I1(CLBLM_R_X7Y153_SLICE_X8Y153_DQ),
.I2(CLBLM_L_X12Y147_SLICE_X16Y147_DO6),
.I3(CLBLM_L_X8Y152_SLICE_X11Y152_DQ),
.I4(CLBLM_R_X7Y149_SLICE_X8Y149_AQ),
.I5(CLBLL_L_X4Y148_SLICE_X4Y148_CQ),
.O5(CLBLM_L_X8Y151_SLICE_X10Y151_DO5),
.O6(CLBLM_L_X8Y151_SLICE_X10Y151_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hfa50fa50dddd8888)
  ) CLBLM_L_X8Y151_SLICE_X10Y151_CLUT (
.I0(LIOB33_X0Y61_IOB_X0Y62_I),
.I1(CLBLM_L_X8Y151_SLICE_X10Y151_CQ),
.I2(CLBLM_L_X8Y152_SLICE_X11Y152_DQ),
.I3(CLBLM_R_X7Y152_SLICE_X9Y152_C5Q),
.I4(CLBLM_R_X5Y145_SLICE_X6Y145_AQ),
.I5(1'b1),
.O5(CLBLM_L_X8Y151_SLICE_X10Y151_CO5),
.O6(CLBLM_L_X8Y151_SLICE_X10Y151_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hffaa00aaf0fff000)
  ) CLBLM_L_X8Y151_SLICE_X10Y151_BLUT (
.I0(CLBLM_R_X7Y152_SLICE_X9Y152_B5Q),
.I1(1'b1),
.I2(CLBLM_L_X10Y152_SLICE_X13Y152_BQ),
.I3(LIOB33_X0Y61_IOB_X0Y62_I),
.I4(CLBLL_L_X4Y149_SLICE_X4Y149_B5Q),
.I5(1'b1),
.O5(CLBLM_L_X8Y151_SLICE_X10Y151_BO5),
.O6(CLBLM_L_X8Y151_SLICE_X10Y151_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hcc50cc50f0fff000)
  ) CLBLM_L_X8Y151_SLICE_X10Y151_ALUT (
.I0(CLBLM_R_X7Y152_SLICE_X9Y152_BQ),
.I1(CLBLM_L_X8Y153_SLICE_X10Y153_C5Q),
.I2(CLBLM_L_X8Y151_SLICE_X10Y151_AQ),
.I3(LIOB33_X0Y61_IOB_X0Y62_I),
.I4(CLBLL_L_X4Y143_SLICE_X4Y143_BQ),
.I5(1'b1),
.O5(CLBLM_L_X8Y151_SLICE_X10Y151_AO5),
.O6(CLBLM_L_X8Y151_SLICE_X10Y151_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y151_SLICE_X11Y151_A_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_L_X8Y151_SLICE_X11Y151_AO6),
.Q(CLBLM_L_X8Y151_SLICE_X11Y151_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffff30ffffffba)
  ) CLBLM_L_X8Y151_SLICE_X11Y151_DLUT (
.I0(CLBLM_R_X5Y146_SLICE_X6Y146_BQ),
.I1(CLBLM_L_X10Y151_SLICE_X13Y151_BO6),
.I2(CLBLM_L_X10Y152_SLICE_X13Y152_CQ),
.I3(CLBLM_L_X8Y151_SLICE_X11Y151_CO6),
.I4(CLBLM_L_X10Y146_SLICE_X13Y146_DO6),
.I5(CLBLM_L_X10Y148_SLICE_X12Y148_AO6),
.O5(CLBLM_L_X8Y151_SLICE_X11Y151_DO5),
.O6(CLBLM_L_X8Y151_SLICE_X11Y151_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000400000000)
  ) CLBLM_L_X8Y151_SLICE_X11Y151_CLUT (
.I0(CLBLM_R_X7Y153_SLICE_X8Y153_A5Q),
.I1(CLBLM_R_X3Y148_SLICE_X3Y148_CQ),
.I2(CLBLM_R_X7Y149_SLICE_X8Y149_AQ),
.I3(CLBLL_L_X4Y148_SLICE_X4Y148_CQ),
.I4(CLBLM_L_X12Y147_SLICE_X16Y147_DO6),
.I5(CLBLM_R_X7Y144_SLICE_X9Y144_B5Q),
.O5(CLBLM_L_X8Y151_SLICE_X11Y151_CO5),
.O6(CLBLM_L_X8Y151_SLICE_X11Y151_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h3fbf33bb0faf00aa)
  ) CLBLM_L_X8Y151_SLICE_X11Y151_BLUT (
.I0(CLBLM_R_X7Y152_SLICE_X9Y152_B5Q),
.I1(CLBLM_L_X8Y150_SLICE_X11Y150_BO5),
.I2(CLBLM_L_X10Y151_SLICE_X13Y151_BO6),
.I3(CLBLM_L_X10Y150_SLICE_X12Y150_BO5),
.I4(CLBLM_R_X5Y153_SLICE_X7Y153_CQ),
.I5(CLBLM_L_X10Y152_SLICE_X12Y152_CQ),
.O5(CLBLM_L_X8Y151_SLICE_X11Y151_BO5),
.O6(CLBLM_L_X8Y151_SLICE_X11Y151_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffddffd000dd00d0)
  ) CLBLM_L_X8Y151_SLICE_X11Y151_ALUT (
.I0(CLBLM_R_X3Y145_SLICE_X3Y145_D5Q),
.I1(CLBLL_L_X4Y151_SLICE_X4Y151_BQ),
.I2(CLBLM_L_X8Y151_SLICE_X11Y151_AQ),
.I3(LIOB33_X0Y61_IOB_X0Y62_I),
.I4(CLBLL_L_X4Y151_SLICE_X4Y151_A5Q),
.I5(CLBLM_L_X8Y152_SLICE_X11Y152_DQ),
.O5(CLBLM_L_X8Y151_SLICE_X11Y151_AO5),
.O6(CLBLM_L_X8Y151_SLICE_X11Y151_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y152_SLICE_X10Y152_A5_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_L_X8Y154_SLICE_X10Y154_BO6),
.Q(CLBLM_L_X8Y152_SLICE_X10Y152_A5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "C5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y152_SLICE_X10Y152_C5_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_L_X8Y152_SLICE_X10Y152_CO5),
.Q(CLBLM_L_X8Y152_SLICE_X10Y152_C5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y152_SLICE_X10Y152_A_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_L_X8Y152_SLICE_X10Y152_AO6),
.Q(CLBLM_L_X8Y152_SLICE_X10Y152_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y152_SLICE_X10Y152_B_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_L_X8Y152_SLICE_X10Y152_BO6),
.Q(CLBLM_L_X8Y152_SLICE_X10Y152_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y152_SLICE_X10Y152_C_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_L_X8Y152_SLICE_X10Y152_CO6),
.Q(CLBLM_L_X8Y152_SLICE_X10Y152_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y152_SLICE_X10Y152_D_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_L_X8Y152_SLICE_X10Y152_DO6),
.Q(CLBLM_L_X8Y152_SLICE_X10Y152_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hccccfa00ccccfafa)
  ) CLBLM_L_X8Y152_SLICE_X10Y152_DLUT (
.I0(CLBLM_R_X7Y152_SLICE_X8Y152_B5Q),
.I1(CLBLM_R_X7Y152_SLICE_X9Y152_BQ),
.I2(CLBLM_L_X8Y152_SLICE_X10Y152_DQ),
.I3(CLBLM_R_X7Y152_SLICE_X8Y152_D5Q),
.I4(LIOB33_X0Y61_IOB_X0Y62_I),
.I5(CLBLM_R_X7Y142_SLICE_X8Y142_C5Q),
.O5(CLBLM_L_X8Y152_SLICE_X10Y152_DO5),
.O6(CLBLM_L_X8Y152_SLICE_X10Y152_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hf3f3c0c0ee22ee22)
  ) CLBLM_L_X8Y152_SLICE_X10Y152_CLUT (
.I0(CLBLM_L_X8Y142_SLICE_X10Y142_A5Q),
.I1(LIOB33_X0Y61_IOB_X0Y62_I),
.I2(CLBLM_R_X5Y153_SLICE_X7Y153_AQ),
.I3(CLBLM_L_X8Y151_SLICE_X10Y151_A5Q),
.I4(CLBLM_L_X10Y152_SLICE_X12Y152_DO6),
.I5(1'b1),
.O5(CLBLM_L_X8Y152_SLICE_X10Y152_CO5),
.O6(CLBLM_L_X8Y152_SLICE_X10Y152_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaa0033aaaa00cc)
  ) CLBLM_L_X8Y152_SLICE_X10Y152_BLUT (
.I0(CLBLM_R_X7Y148_SLICE_X9Y148_C5Q),
.I1(CLBLM_L_X8Y152_SLICE_X10Y152_BQ),
.I2(1'b1),
.I3(RIOB33_X105Y131_IOB_X1Y131_I),
.I4(LIOB33_X0Y61_IOB_X0Y62_I),
.I5(CLBLM_R_X7Y152_SLICE_X9Y152_AQ),
.O5(CLBLM_L_X8Y152_SLICE_X10Y152_BO5),
.O6(CLBLM_L_X8Y152_SLICE_X10Y152_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaa003caaaa00f0)
  ) CLBLM_L_X8Y152_SLICE_X10Y152_ALUT (
.I0(CLBLM_R_X11Y153_SLICE_X14Y153_AQ),
.I1(CLBLM_L_X8Y152_SLICE_X10Y152_BQ),
.I2(CLBLM_L_X8Y152_SLICE_X10Y152_AQ),
.I3(RIOB33_X105Y131_IOB_X1Y131_I),
.I4(LIOB33_X0Y61_IOB_X0Y62_I),
.I5(CLBLM_R_X7Y152_SLICE_X9Y152_AQ),
.O5(CLBLM_L_X8Y152_SLICE_X10Y152_AO5),
.O6(CLBLM_L_X8Y152_SLICE_X10Y152_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y152_SLICE_X11Y152_D5_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_L_X8Y152_SLICE_X11Y152_DO5),
.Q(CLBLM_L_X8Y152_SLICE_X11Y152_D5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y152_SLICE_X11Y152_A_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_L_X8Y152_SLICE_X11Y152_AO6),
.Q(CLBLM_L_X8Y152_SLICE_X11Y152_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y152_SLICE_X11Y152_B_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_L_X8Y152_SLICE_X11Y152_BO6),
.Q(CLBLM_L_X8Y152_SLICE_X11Y152_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y152_SLICE_X11Y152_C_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_L_X8Y152_SLICE_X11Y152_CO6),
.Q(CLBLM_L_X8Y152_SLICE_X11Y152_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y152_SLICE_X11Y152_D_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_L_X8Y152_SLICE_X11Y152_DO6),
.Q(CLBLM_L_X8Y152_SLICE_X11Y152_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hf000f0ffcc00ccff)
  ) CLBLM_L_X8Y152_SLICE_X11Y152_DLUT (
.I0(1'b1),
.I1(CLBLM_L_X8Y152_SLICE_X11Y152_CQ),
.I2(CLBLM_R_X7Y146_SLICE_X8Y146_C5Q),
.I3(LIOB33_X0Y61_IOB_X0Y62_I),
.I4(CLBLM_L_X10Y151_SLICE_X13Y151_AQ),
.I5(1'b1),
.O5(CLBLM_L_X8Y152_SLICE_X11Y152_DO5),
.O6(CLBLM_L_X8Y152_SLICE_X11Y152_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f0f0f0ee44ee44)
  ) CLBLM_L_X8Y152_SLICE_X11Y152_CLUT (
.I0(CLBLM_L_X12Y149_SLICE_X17Y149_CO6),
.I1(CLBLM_L_X8Y152_SLICE_X11Y152_CQ),
.I2(CLBLM_R_X5Y153_SLICE_X6Y153_B5Q),
.I3(CLBLM_L_X8Y153_SLICE_X11Y153_BQ),
.I4(1'b1),
.I5(LIOB33_X0Y61_IOB_X0Y62_I),
.O5(CLBLM_L_X8Y152_SLICE_X11Y152_CO5),
.O6(CLBLM_L_X8Y152_SLICE_X11Y152_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfaee5044fafa5050)
  ) CLBLM_L_X8Y152_SLICE_X11Y152_BLUT (
.I0(LIOB33_X0Y61_IOB_X0Y62_I),
.I1(CLBLM_L_X8Y152_SLICE_X11Y152_BQ),
.I2(CLBLM_R_X5Y150_SLICE_X7Y150_AQ),
.I3(CLBLL_L_X4Y147_SLICE_X5Y147_CQ),
.I4(CLBLM_R_X11Y153_SLICE_X15Y153_AQ),
.I5(CLBLL_L_X4Y142_SLICE_X5Y142_DQ),
.O5(CLBLM_L_X8Y152_SLICE_X11Y152_BO5),
.O6(CLBLM_L_X8Y152_SLICE_X11Y152_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hdddd88ddd8d888d8)
  ) CLBLM_L_X8Y152_SLICE_X11Y152_ALUT (
.I0(LIOB33_X0Y61_IOB_X0Y62_I),
.I1(CLBLM_R_X11Y150_SLICE_X14Y150_AQ),
.I2(CLBLM_L_X8Y152_SLICE_X11Y152_AQ),
.I3(CLBLM_R_X7Y142_SLICE_X8Y142_C5Q),
.I4(CLBLM_R_X7Y152_SLICE_X8Y152_D5Q),
.I5(CLBLM_L_X8Y151_SLICE_X10Y151_A5Q),
.O5(CLBLM_L_X8Y152_SLICE_X11Y152_AO5),
.O6(CLBLM_L_X8Y152_SLICE_X11Y152_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y153_SLICE_X10Y153_A5_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_L_X8Y153_SLICE_X10Y153_AO5),
.Q(CLBLM_L_X8Y153_SLICE_X10Y153_A5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y153_SLICE_X10Y153_B5_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_L_X8Y153_SLICE_X10Y153_BO5),
.Q(CLBLM_L_X8Y153_SLICE_X10Y153_B5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "C5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y153_SLICE_X10Y153_C5_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_L_X8Y153_SLICE_X10Y153_CO5),
.Q(CLBLM_L_X8Y153_SLICE_X10Y153_C5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y153_SLICE_X10Y153_D5_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_L_X8Y153_SLICE_X10Y153_DO5),
.Q(CLBLM_L_X8Y153_SLICE_X10Y153_D5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y153_SLICE_X10Y153_A_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_L_X8Y153_SLICE_X10Y153_AO6),
.Q(CLBLM_L_X8Y153_SLICE_X10Y153_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y153_SLICE_X10Y153_B_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_L_X8Y153_SLICE_X10Y153_BO6),
.Q(CLBLM_L_X8Y153_SLICE_X10Y153_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y153_SLICE_X10Y153_C_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_L_X8Y153_SLICE_X10Y153_CO6),
.Q(CLBLM_L_X8Y153_SLICE_X10Y153_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y153_SLICE_X10Y153_D_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_L_X8Y153_SLICE_X10Y153_DO6),
.Q(CLBLM_L_X8Y153_SLICE_X10Y153_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hfc0cfc0cfcfc0c0c)
  ) CLBLM_L_X8Y153_SLICE_X10Y153_DLUT (
.I0(1'b1),
.I1(CLBLM_L_X10Y151_SLICE_X13Y151_A5Q),
.I2(LIOB33_X0Y61_IOB_X0Y62_I),
.I3(CLBLM_L_X10Y145_SLICE_X12Y145_BQ),
.I4(CLBLM_R_X3Y149_SLICE_X3Y149_AQ),
.I5(1'b1),
.O5(CLBLM_L_X8Y153_SLICE_X10Y153_DO5),
.O6(CLBLM_L_X8Y153_SLICE_X10Y153_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hfc0cfc0ca3a3acac)
  ) CLBLM_L_X8Y153_SLICE_X10Y153_CLUT (
.I0(CLBLM_R_X3Y150_SLICE_X2Y150_D5Q),
.I1(CLBLL_L_X4Y143_SLICE_X4Y143_AQ),
.I2(LIOB33_X0Y61_IOB_X0Y62_I),
.I3(CLBLM_R_X7Y153_SLICE_X9Y153_BQ),
.I4(CLBLM_L_X8Y153_SLICE_X10Y153_B5Q),
.I5(1'b1),
.O5(CLBLM_L_X8Y153_SLICE_X10Y153_CO5),
.O6(CLBLM_L_X8Y153_SLICE_X10Y153_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'haa00ff558888dddd)
  ) CLBLM_L_X8Y153_SLICE_X10Y153_BLUT (
.I0(LIOB33_X0Y61_IOB_X0Y62_I),
.I1(CLBLM_L_X8Y153_SLICE_X10Y153_A5Q),
.I2(1'b1),
.I3(CLBLM_R_X7Y152_SLICE_X9Y152_CQ),
.I4(CLBLM_L_X10Y153_SLICE_X13Y153_A5Q),
.I5(1'b1),
.O5(CLBLM_L_X8Y153_SLICE_X10Y153_BO5),
.O6(CLBLM_L_X8Y153_SLICE_X10Y153_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hee22ee22fcfc3030)
  ) CLBLM_L_X8Y153_SLICE_X10Y153_ALUT (
.I0(CLBLM_R_X7Y155_SLICE_X8Y155_A5Q),
.I1(LIOB33_X0Y61_IOB_X0Y62_I),
.I2(CLBLM_R_X5Y153_SLICE_X7Y153_DO6),
.I3(CLBLM_L_X10Y152_SLICE_X12Y152_BQ),
.I4(CLBLM_L_X10Y147_SLICE_X13Y147_AQ),
.I5(1'b1),
.O5(CLBLM_L_X8Y153_SLICE_X10Y153_AO5),
.O6(CLBLM_L_X8Y153_SLICE_X10Y153_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y153_SLICE_X11Y153_A_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_L_X8Y153_SLICE_X11Y153_AO6),
.Q(CLBLM_L_X8Y153_SLICE_X11Y153_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y153_SLICE_X11Y153_B_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_L_X8Y153_SLICE_X11Y153_BO6),
.Q(CLBLM_L_X8Y153_SLICE_X11Y153_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hdddd0000ffff0000)
  ) CLBLM_L_X8Y153_SLICE_X11Y153_DLUT (
.I0(CLBLM_R_X7Y145_SLICE_X8Y145_A5Q),
.I1(CLBLL_L_X4Y153_SLICE_X5Y153_A5Q),
.I2(1'b1),
.I3(1'b1),
.I4(CLBLM_L_X8Y145_SLICE_X11Y145_DQ),
.I5(RIOB33_X105Y131_IOB_X1Y131_I),
.O5(CLBLM_L_X8Y153_SLICE_X11Y153_DO5),
.O6(CLBLM_L_X8Y153_SLICE_X11Y153_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffffffffffae)
  ) CLBLM_L_X8Y153_SLICE_X11Y153_CLUT (
.I0(CLBLM_R_X7Y153_SLICE_X9Y153_C5Q),
.I1(CLBLM_L_X10Y153_SLICE_X12Y153_BQ),
.I2(CLBLM_R_X7Y154_SLICE_X8Y154_DO6),
.I3(CLBLM_L_X10Y153_SLICE_X12Y153_AQ),
.I4(CLBLM_L_X8Y146_SLICE_X11Y146_BQ),
.I5(CLBLM_R_X7Y151_SLICE_X9Y151_D5Q),
.O5(CLBLM_L_X8Y153_SLICE_X11Y153_CO5),
.O6(CLBLM_L_X8Y153_SLICE_X11Y153_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hff55af05ee44ae04)
  ) CLBLM_L_X8Y153_SLICE_X11Y153_BLUT (
.I0(LIOB33_X0Y61_IOB_X0Y62_I),
.I1(CLBLM_L_X8Y153_SLICE_X11Y153_BQ),
.I2(CLBLM_R_X3Y145_SLICE_X3Y145_D5Q),
.I3(CLBLM_L_X10Y154_SLICE_X12Y154_A5Q),
.I4(CLBLL_L_X4Y151_SLICE_X4Y151_BQ),
.I5(CLBLM_L_X8Y153_SLICE_X10Y153_CQ),
.O5(CLBLM_L_X8Y153_SLICE_X11Y153_BO5),
.O6(CLBLM_L_X8Y153_SLICE_X11Y153_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h888888888dd8d8d8)
  ) CLBLM_L_X8Y153_SLICE_X11Y153_ALUT (
.I0(LIOB33_X0Y61_IOB_X0Y62_I),
.I1(CLBLM_R_X11Y153_SLICE_X14Y153_A5Q),
.I2(CLBLM_L_X8Y153_SLICE_X11Y153_AQ),
.I3(CLBLM_L_X10Y153_SLICE_X12Y153_CO5),
.I4(CLBLM_L_X8Y154_SLICE_X11Y154_AQ),
.I5(CLBLM_R_X5Y150_SLICE_X6Y150_B5Q),
.O5(CLBLM_L_X8Y153_SLICE_X11Y153_AO5),
.O6(CLBLM_L_X8Y153_SLICE_X11Y153_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y154_SLICE_X10Y154_A_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_L_X8Y154_SLICE_X10Y154_AO6),
.Q(CLBLM_L_X8Y154_SLICE_X10Y154_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X8Y154_SLICE_X10Y154_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X8Y154_SLICE_X10Y154_DO5),
.O6(CLBLM_L_X8Y154_SLICE_X10Y154_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X8Y154_SLICE_X10Y154_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X8Y154_SLICE_X10Y154_CO5),
.O6(CLBLM_L_X8Y154_SLICE_X10Y154_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hff33cc00a0a00000)
  ) CLBLM_L_X8Y154_SLICE_X10Y154_BLUT (
.I0(CLBLM_L_X10Y154_SLICE_X12Y154_B5Q),
.I1(LIOB33_X0Y61_IOB_X0Y62_I),
.I2(CLBLM_R_X5Y142_SLICE_X7Y142_CO6),
.I3(CLBLM_L_X8Y153_SLICE_X10Y153_B5Q),
.I4(RIOB33_X105Y131_IOB_X1Y131_I),
.I5(1'b1),
.O5(CLBLM_L_X8Y154_SLICE_X10Y154_BO5),
.O6(CLBLM_L_X8Y154_SLICE_X10Y154_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hccccffffcccc5af0)
  ) CLBLM_L_X8Y154_SLICE_X10Y154_ALUT (
.I0(CLBLM_R_X7Y155_SLICE_X8Y155_BO5),
.I1(CLBLM_L_X10Y154_SLICE_X13Y154_AQ),
.I2(CLBLM_L_X8Y154_SLICE_X10Y154_AQ),
.I3(CLBLM_R_X7Y154_SLICE_X8Y154_AQ),
.I4(LIOB33_X0Y61_IOB_X0Y62_I),
.I5(CLBLM_R_X5Y150_SLICE_X6Y150_B5Q),
.O5(CLBLM_L_X8Y154_SLICE_X10Y154_AO5),
.O6(CLBLM_L_X8Y154_SLICE_X10Y154_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y154_SLICE_X11Y154_A_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_L_X8Y154_SLICE_X11Y154_AO6),
.Q(CLBLM_L_X8Y154_SLICE_X11Y154_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X8Y154_SLICE_X11Y154_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X8Y154_SLICE_X11Y154_DO5),
.O6(CLBLM_L_X8Y154_SLICE_X11Y154_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X8Y154_SLICE_X11Y154_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X8Y154_SLICE_X11Y154_CO5),
.O6(CLBLM_L_X8Y154_SLICE_X11Y154_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X8Y154_SLICE_X11Y154_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X8Y154_SLICE_X11Y154_BO5),
.O6(CLBLM_L_X8Y154_SLICE_X11Y154_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hcc00cc00cc5accf0)
  ) CLBLM_L_X8Y154_SLICE_X11Y154_ALUT (
.I0(CLBLM_L_X10Y153_SLICE_X12Y153_A5Q),
.I1(CLBLM_L_X10Y155_SLICE_X12Y155_AQ),
.I2(CLBLM_L_X8Y154_SLICE_X11Y154_AQ),
.I3(LIOB33_X0Y61_IOB_X0Y62_I),
.I4(CLBLM_R_X5Y152_SLICE_X6Y152_BQ),
.I5(CLBLM_R_X5Y150_SLICE_X6Y150_B5Q),
.O5(CLBLM_L_X8Y154_SLICE_X11Y154_AO5),
.O6(CLBLM_L_X8Y154_SLICE_X11Y154_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y142_SLICE_X12Y142_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y142_SLICE_X12Y142_AO6),
.Q(CLBLM_L_X10Y142_SLICE_X12Y142_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X10Y142_SLICE_X12Y142_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X10Y142_SLICE_X12Y142_DO5),
.O6(CLBLM_L_X10Y142_SLICE_X12Y142_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h5500550000000000)
  ) CLBLM_L_X10Y142_SLICE_X12Y142_CLUT (
.I0(CLBLL_L_X4Y151_SLICE_X4Y151_CQ),
.I1(1'b1),
.I2(1'b1),
.I3(RIOB33_X105Y131_IOB_X1Y131_I),
.I4(1'b1),
.I5(CLBLM_L_X8Y142_SLICE_X11Y142_BQ),
.O5(CLBLM_L_X10Y142_SLICE_X12Y142_CO5),
.O6(CLBLM_L_X10Y142_SLICE_X12Y142_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000008000000000)
  ) CLBLM_L_X10Y142_SLICE_X12Y142_BLUT (
.I0(CLBLM_R_X7Y142_SLICE_X9Y142_CQ),
.I1(RIOB33_X105Y101_IOB_X1Y101_I),
.I2(RIOB33_SING_X105Y100_IOB_X1Y100_I),
.I3(RIOB33_X105Y103_IOB_X1Y104_I),
.I4(RIOB33_X105Y103_IOB_X1Y103_I),
.I5(RIOB33_X105Y131_IOB_X1Y131_I),
.O5(CLBLM_L_X10Y142_SLICE_X12Y142_BO5),
.O6(CLBLM_L_X10Y142_SLICE_X12Y142_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hcc00cc0acc00cc00)
  ) CLBLM_L_X10Y142_SLICE_X12Y142_ALUT (
.I0(CLBLM_L_X8Y148_SLICE_X11Y148_B5Q),
.I1(CLBLM_L_X8Y147_SLICE_X10Y147_C5Q),
.I2(RIOB33_X105Y101_IOB_X1Y102_I),
.I3(LIOB33_X0Y61_IOB_X0Y62_I),
.I4(RIOB33_SING_X105Y100_IOB_X1Y100_I),
.I5(CLBLM_L_X10Y147_SLICE_X12Y147_CO6),
.O5(CLBLM_L_X10Y142_SLICE_X12Y142_AO5),
.O6(CLBLM_L_X10Y142_SLICE_X12Y142_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y142_SLICE_X13Y142_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y142_SLICE_X13Y142_AO6),
.Q(CLBLM_L_X10Y142_SLICE_X13Y142_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X10Y142_SLICE_X13Y142_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X10Y142_SLICE_X13Y142_DO5),
.O6(CLBLM_L_X10Y142_SLICE_X13Y142_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h4444444444444444)
  ) CLBLM_L_X10Y142_SLICE_X13Y142_CLUT (
.I0(CLBLM_L_X10Y145_SLICE_X12Y145_AQ),
.I1(CLBLM_R_X5Y142_SLICE_X7Y142_BQ),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X10Y142_SLICE_X13Y142_CO5),
.O6(CLBLM_L_X10Y142_SLICE_X13Y142_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffffffffffff7)
  ) CLBLM_L_X10Y142_SLICE_X13Y142_BLUT (
.I0(CLBLM_L_X10Y144_SLICE_X13Y144_CQ),
.I1(RIOB33_X105Y105_IOB_X1Y105_I),
.I2(CLBLM_R_X7Y142_SLICE_X9Y142_BQ),
.I3(CLBLM_L_X10Y147_SLICE_X12Y147_AO5),
.I4(CLBLM_L_X8Y147_SLICE_X10Y147_C5Q),
.I5(CLBLM_L_X10Y142_SLICE_X13Y142_CO6),
.O5(CLBLM_L_X10Y142_SLICE_X13Y142_BO5),
.O6(CLBLM_L_X10Y142_SLICE_X13Y142_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'haa3caaf0aa00aa00)
  ) CLBLM_L_X10Y142_SLICE_X13Y142_ALUT (
.I0(CLBLM_R_X11Y146_SLICE_X14Y146_AQ),
.I1(CLBLM_L_X8Y142_SLICE_X10Y142_BQ),
.I2(CLBLM_L_X10Y142_SLICE_X13Y142_AQ),
.I3(LIOB33_X0Y61_IOB_X0Y62_I),
.I4(CLBLM_L_X8Y144_SLICE_X10Y144_AO6),
.I5(CLBLM_L_X10Y144_SLICE_X12Y144_AO6),
.O5(CLBLM_L_X10Y142_SLICE_X13Y142_AO5),
.O6(CLBLM_L_X10Y142_SLICE_X13Y142_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y143_SLICE_X12Y143_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y143_SLICE_X12Y143_AO6),
.Q(CLBLM_L_X10Y143_SLICE_X12Y143_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y143_SLICE_X12Y143_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y143_SLICE_X12Y143_BO6),
.Q(CLBLM_L_X10Y143_SLICE_X12Y143_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h2000000000000000)
  ) CLBLM_L_X10Y143_SLICE_X12Y143_DLUT (
.I0(CLBLM_L_X8Y143_SLICE_X10Y143_AQ),
.I1(CLBLM_R_X3Y142_SLICE_X2Y142_BO5),
.I2(CLBLM_R_X5Y145_SLICE_X7Y145_B5Q),
.I3(CLBLM_L_X10Y142_SLICE_X13Y142_AQ),
.I4(CLBLM_L_X10Y144_SLICE_X13Y144_A5Q),
.I5(CLBLM_L_X8Y142_SLICE_X10Y142_BQ),
.O5(CLBLM_L_X10Y143_SLICE_X12Y143_DO5),
.O6(CLBLM_L_X10Y143_SLICE_X12Y143_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h5fff5fff0fff0fff)
  ) CLBLM_L_X10Y143_SLICE_X12Y143_CLUT (
.I0(CLBLM_L_X10Y143_SLICE_X12Y143_BQ),
.I1(1'b1),
.I2(CLBLM_L_X10Y144_SLICE_X13Y144_DQ),
.I3(CLBLM_R_X7Y143_SLICE_X9Y143_AQ),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X10Y143_SLICE_X12Y143_CO5),
.O6(CLBLM_L_X10Y143_SLICE_X12Y143_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f0f0f0aaccaa33)
  ) CLBLM_L_X10Y143_SLICE_X12Y143_BLUT (
.I0(CLBLM_L_X8Y146_SLICE_X11Y146_B5Q),
.I1(CLBLM_L_X10Y143_SLICE_X12Y143_BQ),
.I2(CLBLM_R_X7Y153_SLICE_X9Y153_C5Q),
.I3(CLBLM_L_X8Y149_SLICE_X11Y149_AQ),
.I4(CLBLM_L_X10Y143_SLICE_X12Y143_CO5),
.I5(LIOB33_X0Y61_IOB_X0Y62_I),
.O5(CLBLM_L_X10Y143_SLICE_X12Y143_BO5),
.O6(CLBLM_L_X10Y143_SLICE_X12Y143_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff0000c4c8c4c8)
  ) CLBLM_L_X10Y143_SLICE_X12Y143_ALUT (
.I0(RIOB33_X105Y109_IOB_X1Y110_I),
.I1(CLBLM_R_X7Y151_SLICE_X9Y151_A5Q),
.I2(CLBLM_L_X10Y143_SLICE_X12Y143_AQ),
.I3(CLBLM_L_X10Y145_SLICE_X12Y145_A5Q),
.I4(CLBLM_L_X10Y144_SLICE_X12Y144_AQ),
.I5(LIOB33_X0Y61_IOB_X0Y62_I),
.O5(CLBLM_L_X10Y143_SLICE_X12Y143_AO5),
.O6(CLBLM_L_X10Y143_SLICE_X12Y143_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y143_SLICE_X13Y143_C5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y143_SLICE_X13Y143_CO5),
.Q(CLBLM_L_X10Y143_SLICE_X13Y143_C5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y143_SLICE_X13Y143_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y143_SLICE_X13Y143_AO6),
.Q(CLBLM_L_X10Y143_SLICE_X13Y143_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y143_SLICE_X13Y143_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y143_SLICE_X13Y143_BO6),
.Q(CLBLM_L_X10Y143_SLICE_X13Y143_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y143_SLICE_X13Y143_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y143_SLICE_X13Y143_CO6),
.Q(CLBLM_L_X10Y143_SLICE_X13Y143_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h880000003fffffff)
  ) CLBLM_L_X10Y143_SLICE_X13Y143_DLUT (
.I0(CLBLM_L_X8Y144_SLICE_X10Y144_AO6),
.I1(CLBLM_L_X10Y142_SLICE_X13Y142_AQ),
.I2(CLBLM_L_X8Y144_SLICE_X11Y144_AQ),
.I3(CLBLM_L_X10Y143_SLICE_X13Y143_BQ),
.I4(CLBLM_L_X8Y142_SLICE_X10Y142_BQ),
.I5(1'b1),
.O5(CLBLM_L_X10Y143_SLICE_X13Y143_DO5),
.O6(CLBLM_L_X10Y143_SLICE_X13Y143_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hff00aaaaccccf0f0)
  ) CLBLM_L_X10Y143_SLICE_X13Y143_CLUT (
.I0(CLBLM_L_X10Y143_SLICE_X12Y143_AQ),
.I1(CLBLM_L_X10Y143_SLICE_X13Y143_CQ),
.I2(RIOB33_X105Y127_IOB_X1Y128_I),
.I3(CLBLM_L_X10Y146_SLICE_X12Y146_D5Q),
.I4(LIOB33_X0Y61_IOB_X0Y62_I),
.I5(1'b1),
.O5(CLBLM_L_X10Y143_SLICE_X13Y143_CO5),
.O6(CLBLM_L_X10Y143_SLICE_X13Y143_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hff00ff0022228888)
  ) CLBLM_L_X10Y143_SLICE_X13Y143_BLUT (
.I0(CLBLM_L_X10Y144_SLICE_X12Y144_AO6),
.I1(CLBLM_L_X10Y143_SLICE_X13Y143_BQ),
.I2(1'b1),
.I3(CLBLM_L_X8Y143_SLICE_X11Y143_BQ),
.I4(CLBLM_L_X10Y143_SLICE_X12Y143_DO6),
.I5(LIOB33_X0Y61_IOB_X0Y62_I),
.O5(CLBLM_L_X10Y143_SLICE_X13Y143_BO5),
.O6(CLBLM_L_X10Y143_SLICE_X13Y143_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaaaaaafff000f0)
  ) CLBLM_L_X10Y143_SLICE_X13Y143_ALUT (
.I0(CLBLM_L_X8Y146_SLICE_X11Y146_B5Q),
.I1(1'b1),
.I2(CLBLM_L_X10Y143_SLICE_X13Y143_AQ),
.I3(CLBLM_R_X11Y146_SLICE_X14Y146_DO6),
.I4(CLBLM_L_X8Y142_SLICE_X10Y142_AQ),
.I5(LIOB33_X0Y61_IOB_X0Y62_I),
.O5(CLBLM_L_X10Y143_SLICE_X13Y143_AO5),
.O6(CLBLM_L_X10Y143_SLICE_X13Y143_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y144_SLICE_X12Y144_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(LIOB33_X0Y61_IOB_X0Y62_I),
.D(CLBLM_R_X3Y145_SLICE_X3Y145_C5Q),
.Q(CLBLM_L_X10Y144_SLICE_X12Y144_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X10Y144_SLICE_X12Y144_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X10Y144_SLICE_X12Y144_DO5),
.O6(CLBLM_L_X10Y144_SLICE_X12Y144_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffffffff0200)
  ) CLBLM_L_X10Y144_SLICE_X12Y144_CLUT (
.I0(CLBLM_L_X10Y142_SLICE_X12Y142_AQ),
.I1(RIOB33_X105Y101_IOB_X1Y102_I),
.I2(RIOB33_SING_X105Y100_IOB_X1Y100_I),
.I3(CLBLM_L_X8Y148_SLICE_X11Y148_B5Q),
.I4(CLBLM_L_X10Y142_SLICE_X12Y142_BO6),
.I5(CLBLM_L_X8Y154_SLICE_X10Y154_BO5),
.O5(CLBLM_L_X10Y144_SLICE_X12Y144_CO5),
.O6(CLBLM_L_X10Y144_SLICE_X12Y144_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h00ff00ffeb41aa00)
  ) CLBLM_L_X10Y144_SLICE_X12Y144_BLUT (
.I0(LIOB33_X0Y61_IOB_X0Y62_I),
.I1(CLBLM_R_X3Y142_SLICE_X2Y142_BO5),
.I2(CLBLM_L_X10Y144_SLICE_X13Y144_A5Q),
.I3(CLBLM_L_X10Y144_SLICE_X13Y144_BQ),
.I4(CLBLM_L_X10Y144_SLICE_X12Y144_AO6),
.I5(1'b1),
.O5(CLBLM_L_X10Y144_SLICE_X12Y144_BO5),
.O6(CLBLM_L_X10Y144_SLICE_X12Y144_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h00fb00bf44444444)
  ) CLBLM_L_X10Y144_SLICE_X12Y144_ALUT (
.I0(CLBLM_L_X8Y145_SLICE_X11Y145_DQ),
.I1(CLBLM_L_X10Y147_SLICE_X12Y147_BQ),
.I2(CLBLM_L_X10Y144_SLICE_X13Y144_C5Q),
.I3(CLBLM_L_X10Y145_SLICE_X12Y145_CO6),
.I4(CLBLM_L_X10Y143_SLICE_X13Y143_C5Q),
.I5(1'b1),
.O5(CLBLM_L_X10Y144_SLICE_X12Y144_AO5),
.O6(CLBLM_L_X10Y144_SLICE_X12Y144_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y144_SLICE_X13Y144_A5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y144_SLICE_X12Y144_BO5),
.Q(CLBLM_L_X10Y144_SLICE_X13Y144_A5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "C5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y144_SLICE_X13Y144_C5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y144_SLICE_X13Y144_CO5),
.Q(CLBLM_L_X10Y144_SLICE_X13Y144_C5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y144_SLICE_X13Y144_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y144_SLICE_X13Y144_AO6),
.Q(CLBLM_L_X10Y144_SLICE_X13Y144_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y144_SLICE_X13Y144_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y144_SLICE_X13Y144_BO6),
.Q(CLBLM_L_X10Y144_SLICE_X13Y144_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y144_SLICE_X13Y144_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y144_SLICE_X13Y144_CO6),
.Q(CLBLM_L_X10Y144_SLICE_X13Y144_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y144_SLICE_X13Y144_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y144_SLICE_X13Y144_DO6),
.Q(CLBLM_L_X10Y144_SLICE_X13Y144_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hffcc3300dede1212)
  ) CLBLM_L_X10Y144_SLICE_X13Y144_DLUT (
.I0(CLBLM_R_X7Y143_SLICE_X9Y143_AQ),
.I1(LIOB33_X0Y61_IOB_X0Y62_I),
.I2(CLBLM_L_X10Y144_SLICE_X13Y144_DQ),
.I3(CLBLM_L_X8Y151_SLICE_X10Y151_BQ),
.I4(CLBLM_L_X10Y144_SLICE_X13Y144_AQ),
.I5(CLBLM_L_X8Y149_SLICE_X11Y149_AQ),
.O5(CLBLM_L_X10Y144_SLICE_X13Y144_DO5),
.O6(CLBLM_L_X10Y144_SLICE_X13Y144_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hccf0ccf0aaccaacc)
  ) CLBLM_L_X10Y144_SLICE_X13Y144_CLUT (
.I0(CLBLM_L_X10Y143_SLICE_X13Y143_AQ),
.I1(CLBLM_L_X10Y143_SLICE_X13Y143_C5Q),
.I2(CLBLM_L_X8Y147_SLICE_X10Y147_C5Q),
.I3(LIOB33_X0Y61_IOB_X0Y62_I),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X10Y144_SLICE_X13Y144_CO5),
.O6(CLBLM_L_X10Y144_SLICE_X13Y144_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf1f4fbfe01040b0e)
  ) CLBLM_L_X10Y144_SLICE_X13Y144_BLUT (
.I0(CLBLM_L_X10Y144_SLICE_X12Y144_AO5),
.I1(CLBLM_L_X10Y144_SLICE_X13Y144_BQ),
.I2(LIOB33_X0Y61_IOB_X0Y62_I),
.I3(CLBLM_L_X10Y145_SLICE_X12Y145_CO6),
.I4(CLBLM_L_X10Y143_SLICE_X13Y143_C5Q),
.I5(CLBLM_R_X5Y148_SLICE_X7Y148_BQ),
.O5(CLBLM_L_X10Y144_SLICE_X13Y144_BO5),
.O6(CLBLM_L_X10Y144_SLICE_X13Y144_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaacc0caaaa33f3)
  ) CLBLM_L_X10Y144_SLICE_X13Y144_ALUT (
.I0(CLBLM_L_X10Y149_SLICE_X13Y149_AQ),
.I1(CLBLM_R_X7Y144_SLICE_X8Y144_C5Q),
.I2(RIOB33_X105Y131_IOB_X1Y132_I),
.I3(RIOB33_X105Y133_IOB_X1Y133_I),
.I4(LIOB33_X0Y61_IOB_X0Y62_I),
.I5(CLBLM_L_X10Y145_SLICE_X13Y145_CO6),
.O5(CLBLM_L_X10Y144_SLICE_X13Y144_AO5),
.O6(CLBLM_L_X10Y144_SLICE_X13Y144_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y145_SLICE_X12Y145_A5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y145_SLICE_X12Y145_AO5),
.Q(CLBLM_L_X10Y145_SLICE_X12Y145_A5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y145_SLICE_X12Y145_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y145_SLICE_X12Y145_AO6),
.Q(CLBLM_L_X10Y145_SLICE_X12Y145_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y145_SLICE_X12Y145_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y145_SLICE_X12Y145_BO6),
.Q(CLBLM_L_X10Y145_SLICE_X12Y145_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hf3f3f3fbf0f0f0fa)
  ) CLBLM_L_X10Y145_SLICE_X12Y145_DLUT (
.I0(CLBLM_L_X10Y151_SLICE_X13Y151_A5Q),
.I1(CLBLM_L_X10Y148_SLICE_X12Y148_AO5),
.I2(CLBLM_R_X7Y145_SLICE_X9Y145_DO6),
.I3(CLBLL_L_X4Y148_SLICE_X4Y148_CQ),
.I4(CLBLM_L_X12Y146_SLICE_X16Y146_CO6),
.I5(CLBLM_R_X3Y145_SLICE_X3Y145_C5Q),
.O5(CLBLM_L_X10Y145_SLICE_X12Y145_DO5),
.O6(CLBLM_L_X10Y145_SLICE_X12Y145_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0404040005050500)
  ) CLBLM_L_X10Y145_SLICE_X12Y145_CLUT (
.I0(CLBLM_R_X3Y142_SLICE_X2Y142_BO5),
.I1(CLBLM_L_X8Y145_SLICE_X11Y145_DQ),
.I2(CLBLM_L_X10Y145_SLICE_X13Y145_DO6),
.I3(CLBLM_R_X5Y145_SLICE_X7Y145_B5Q),
.I4(CLBLM_L_X8Y146_SLICE_X10Y146_AQ),
.I5(CLBLM_L_X10Y147_SLICE_X12Y147_BQ),
.O5(CLBLM_L_X10Y145_SLICE_X12Y145_CO5),
.O6(CLBLM_L_X10Y145_SLICE_X12Y145_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hcecccecc02000200)
  ) CLBLM_L_X10Y145_SLICE_X12Y145_BLUT (
.I0(CLBLM_L_X10Y142_SLICE_X12Y142_CO6),
.I1(LIOB33_X0Y61_IOB_X0Y62_I),
.I2(CLBLM_L_X10Y144_SLICE_X12Y144_AQ),
.I3(CLBLM_L_X8Y145_SLICE_X11Y145_DQ),
.I4(1'b1),
.I5(CLBLM_R_X3Y145_SLICE_X3Y145_DQ),
.O5(CLBLM_L_X10Y145_SLICE_X12Y145_BO5),
.O6(CLBLM_L_X10Y145_SLICE_X12Y145_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hd8d8d8d8fa50fa50)
  ) CLBLM_L_X10Y145_SLICE_X12Y145_ALUT (
.I0(LIOB33_X0Y61_IOB_X0Y62_I),
.I1(CLBLM_L_X8Y147_SLICE_X11Y147_AQ),
.I2(RIOB33_X105Y109_IOB_X1Y110_I),
.I3(CLBLM_L_X8Y153_SLICE_X10Y153_CQ),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X10Y145_SLICE_X12Y145_AO5),
.O6(CLBLM_L_X10Y145_SLICE_X12Y145_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y145_SLICE_X13Y145_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y145_SLICE_X13Y145_AO6),
.Q(CLBLM_L_X10Y145_SLICE_X13Y145_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffff3030f0f0)
  ) CLBLM_L_X10Y145_SLICE_X13Y145_DLUT (
.I0(1'b1),
.I1(CLBLM_L_X10Y144_SLICE_X13Y144_A5Q),
.I2(CLBLM_L_X8Y146_SLICE_X10Y146_AQ),
.I3(1'b1),
.I4(CLBLM_L_X10Y145_SLICE_X13Y145_AQ),
.I5(CLBLM_L_X10Y143_SLICE_X13Y143_DO5),
.O5(CLBLM_L_X10Y145_SLICE_X13Y145_DO5),
.O6(CLBLM_L_X10Y145_SLICE_X13Y145_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h9669966969966996)
  ) CLBLM_L_X10Y145_SLICE_X13Y145_CLUT (
.I0(CLBLM_L_X10Y153_SLICE_X13Y153_A5Q),
.I1(CLBLM_L_X10Y149_SLICE_X13Y149_AQ),
.I2(CLBLM_L_X8Y144_SLICE_X10Y144_BO6),
.I3(CLBLL_L_X4Y149_SLICE_X5Y149_C5Q),
.I4(1'b1),
.I5(CLBLM_L_X10Y151_SLICE_X13Y151_A5Q),
.O5(CLBLM_L_X10Y145_SLICE_X13Y145_CO5),
.O6(CLBLM_L_X10Y145_SLICE_X13Y145_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h9669699669969669)
  ) CLBLM_L_X10Y145_SLICE_X13Y145_BLUT (
.I0(CLBLM_L_X8Y144_SLICE_X10Y144_BO6),
.I1(CLBLM_L_X10Y149_SLICE_X13Y149_AQ),
.I2(CLBLM_L_X10Y151_SLICE_X13Y151_A5Q),
.I3(CLBLM_R_X7Y144_SLICE_X8Y144_C5Q),
.I4(CLBLM_L_X10Y153_SLICE_X13Y153_A5Q),
.I5(CLBLL_L_X4Y149_SLICE_X5Y149_C5Q),
.O5(CLBLM_L_X10Y145_SLICE_X13Y145_BO5),
.O6(CLBLM_L_X10Y145_SLICE_X13Y145_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hff00ff0078780000)
  ) CLBLM_L_X10Y145_SLICE_X13Y145_ALUT (
.I0(CLBLM_L_X10Y143_SLICE_X13Y143_DO6),
.I1(CLBLM_L_X8Y144_SLICE_X11Y144_AQ),
.I2(CLBLM_L_X10Y145_SLICE_X13Y145_AQ),
.I3(CLBLM_R_X5Y145_SLICE_X6Y145_DQ),
.I4(CLBLM_L_X10Y144_SLICE_X12Y144_AO6),
.I5(LIOB33_X0Y61_IOB_X0Y62_I),
.O5(CLBLM_L_X10Y145_SLICE_X13Y145_AO5),
.O6(CLBLM_L_X10Y145_SLICE_X13Y145_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y146_SLICE_X12Y146_D5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y146_SLICE_X12Y146_DO5),
.Q(CLBLM_L_X10Y146_SLICE_X12Y146_D5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y146_SLICE_X12Y146_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y146_SLICE_X12Y146_AO6),
.Q(CLBLM_L_X10Y146_SLICE_X12Y146_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y146_SLICE_X12Y146_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y146_SLICE_X12Y146_BO6),
.Q(CLBLM_L_X10Y146_SLICE_X12Y146_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y146_SLICE_X12Y146_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y146_SLICE_X12Y146_CO6),
.Q(CLBLM_L_X10Y146_SLICE_X12Y146_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y146_SLICE_X12Y146_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y146_SLICE_X12Y146_DO6),
.Q(CLBLM_L_X10Y146_SLICE_X12Y146_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hfff00f00cacacaca)
  ) CLBLM_L_X10Y146_SLICE_X12Y146_DLUT (
.I0(CLBLM_L_X8Y145_SLICE_X11Y145_CQ),
.I1(CLBLM_L_X10Y146_SLICE_X12Y146_AQ),
.I2(LIOB33_X0Y61_IOB_X0Y62_I),
.I3(CLBLL_L_X4Y149_SLICE_X5Y149_C5Q),
.I4(CLBLM_L_X8Y148_SLICE_X10Y148_B5Q),
.I5(1'b1),
.O5(CLBLM_L_X10Y146_SLICE_X12Y146_DO5),
.O6(CLBLM_L_X10Y146_SLICE_X12Y146_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hfd0dfc0cf808fc0c)
  ) CLBLM_L_X10Y146_SLICE_X12Y146_CLUT (
.I0(CLBLM_L_X8Y147_SLICE_X10Y147_C5Q),
.I1(CLBLM_L_X10Y146_SLICE_X12Y146_CQ),
.I2(LIOB33_X0Y61_IOB_X0Y62_I),
.I3(CLBLM_L_X10Y145_SLICE_X12Y145_A5Q),
.I4(CLBLM_L_X10Y144_SLICE_X13Y144_CQ),
.I5(CLBLM_R_X7Y146_SLICE_X8Y146_AQ),
.O5(CLBLM_L_X10Y146_SLICE_X12Y146_CO5),
.O6(CLBLM_L_X10Y146_SLICE_X12Y146_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hff0ffc0cf505f404)
  ) CLBLM_L_X10Y146_SLICE_X12Y146_BLUT (
.I0(CLBLL_L_X4Y142_SLICE_X5Y142_DQ),
.I1(CLBLM_L_X10Y146_SLICE_X12Y146_BQ),
.I2(LIOB33_X0Y61_IOB_X0Y62_I),
.I3(CLBLM_R_X7Y146_SLICE_X8Y146_AQ),
.I4(CLBLM_L_X10Y149_SLICE_X12Y149_AQ),
.I5(CLBLL_L_X4Y147_SLICE_X5Y147_CQ),
.O5(CLBLM_L_X10Y146_SLICE_X12Y146_BO5),
.O6(CLBLM_L_X10Y146_SLICE_X12Y146_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hff00aaaaff00e2e2)
  ) CLBLM_L_X10Y146_SLICE_X12Y146_ALUT (
.I0(CLBLM_R_X5Y145_SLICE_X6Y145_DQ),
.I1(CLBLL_L_X4Y142_SLICE_X5Y142_DQ),
.I2(CLBLM_L_X10Y146_SLICE_X12Y146_AQ),
.I3(CLBLM_L_X8Y142_SLICE_X11Y142_AQ),
.I4(LIOB33_X0Y61_IOB_X0Y62_I),
.I5(CLBLL_L_X4Y147_SLICE_X5Y147_CQ),
.O5(CLBLM_L_X10Y146_SLICE_X12Y146_AO5),
.O6(CLBLM_L_X10Y146_SLICE_X12Y146_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y146_SLICE_X13Y146_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y146_SLICE_X13Y146_AO6),
.Q(CLBLM_L_X10Y146_SLICE_X13Y146_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y146_SLICE_X13Y146_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y146_SLICE_X13Y146_BO6),
.Q(CLBLM_L_X10Y146_SLICE_X13Y146_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y146_SLICE_X13Y146_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y146_SLICE_X13Y146_CO6),
.Q(CLBLM_L_X10Y146_SLICE_X13Y146_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffefffefefefe)
  ) CLBLM_L_X10Y146_SLICE_X13Y146_DLUT (
.I0(RIOB33_X105Y133_IOB_X1Y133_I),
.I1(RIOB33_X105Y129_IOB_X1Y130_I),
.I2(RIOB33_X105Y129_IOB_X1Y129_I),
.I3(RIOB33_X105Y131_IOB_X1Y132_I),
.I4(CLBLM_L_X10Y144_SLICE_X13Y144_AQ),
.I5(1'b1),
.O5(CLBLM_L_X10Y146_SLICE_X13Y146_DO5),
.O6(CLBLM_L_X10Y146_SLICE_X13Y146_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hff00afafff008c8c)
  ) CLBLM_L_X10Y146_SLICE_X13Y146_CLUT (
.I0(CLBLM_L_X10Y145_SLICE_X12Y145_AQ),
.I1(CLBLM_L_X10Y146_SLICE_X13Y146_CQ),
.I2(CLBLM_R_X5Y142_SLICE_X7Y142_BQ),
.I3(CLBLM_L_X10Y146_SLICE_X13Y146_BQ),
.I4(LIOB33_X0Y61_IOB_X0Y62_I),
.I5(CLBLL_L_X4Y144_SLICE_X5Y144_D5Q),
.O5(CLBLM_L_X10Y146_SLICE_X13Y146_CO5),
.O6(CLBLM_L_X10Y146_SLICE_X13Y146_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaafc00aaaafcfc)
  ) CLBLM_L_X10Y146_SLICE_X13Y146_BLUT (
.I0(CLBLM_L_X10Y148_SLICE_X13Y148_CQ),
.I1(CLBLM_L_X10Y146_SLICE_X13Y146_BQ),
.I2(CLBLM_L_X8Y146_SLICE_X11Y146_CQ),
.I3(CLBLM_L_X10Y145_SLICE_X12Y145_AQ),
.I4(LIOB33_X0Y61_IOB_X0Y62_I),
.I5(CLBLM_R_X5Y142_SLICE_X7Y142_BQ),
.O5(CLBLM_L_X10Y146_SLICE_X13Y146_BO5),
.O6(CLBLM_L_X10Y146_SLICE_X13Y146_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffaff5000fa0050)
  ) CLBLM_L_X10Y146_SLICE_X13Y146_ALUT (
.I0(CLBLM_R_X11Y146_SLICE_X14Y146_DO6),
.I1(1'b1),
.I2(CLBLM_L_X10Y146_SLICE_X13Y146_AQ),
.I3(LIOB33_X0Y61_IOB_X0Y62_I),
.I4(CLBLL_L_X4Y146_SLICE_X4Y146_AQ),
.I5(CLBLL_L_X4Y150_SLICE_X5Y150_A5Q),
.O5(CLBLM_L_X10Y146_SLICE_X13Y146_AO5),
.O6(CLBLM_L_X10Y146_SLICE_X13Y146_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y147_SLICE_X12Y147_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(LIOB33_X0Y61_IOB_X0Y62_I),
.D(CLBLM_L_X8Y146_SLICE_X10Y146_AQ),
.Q(CLBLM_L_X10Y147_SLICE_X12Y147_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y147_SLICE_X12Y147_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(LIOB33_X0Y61_IOB_X0Y62_I),
.D(CLBLM_R_X7Y143_SLICE_X9Y143_BQ),
.Q(CLBLM_L_X10Y147_SLICE_X12Y147_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y147_SLICE_X12Y147_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(LIOB33_X0Y61_IOB_X0Y62_I),
.D(CLBLL_L_X4Y143_SLICE_X5Y143_AQ),
.Q(CLBLM_L_X10Y147_SLICE_X12Y147_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff01ffffff0101)
  ) CLBLM_L_X10Y147_SLICE_X12Y147_DLUT (
.I0(CLBLL_L_X4Y148_SLICE_X4Y148_CQ),
.I1(CLBLM_L_X10Y151_SLICE_X13Y151_AQ),
.I2(CLBLM_L_X12Y146_SLICE_X16Y146_CO6),
.I3(CLBLM_L_X10Y148_SLICE_X12Y148_AO5),
.I4(CLBLM_R_X7Y145_SLICE_X9Y145_AO6),
.I5(CLBLM_L_X8Y152_SLICE_X11Y152_D5Q),
.O5(CLBLM_L_X10Y147_SLICE_X12Y147_DO5),
.O6(CLBLM_L_X10Y147_SLICE_X12Y147_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000001300)
  ) CLBLM_L_X10Y147_SLICE_X12Y147_CLUT (
.I0(RIOB33_X105Y131_IOB_X1Y131_I),
.I1(CLBLL_L_X4Y153_SLICE_X5Y153_A5Q),
.I2(CLBLL_L_X4Y150_SLICE_X5Y150_A5Q),
.I3(CLBLM_R_X5Y142_SLICE_X7Y142_CO6),
.I4(CLBLM_L_X8Y145_SLICE_X11Y145_DQ),
.I5(CLBLM_L_X10Y149_SLICE_X12Y149_BO6),
.O5(CLBLM_L_X10Y147_SLICE_X12Y147_CO5),
.O6(CLBLM_L_X10Y147_SLICE_X12Y147_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'haaffaaff08050800)
  ) CLBLM_L_X10Y147_SLICE_X12Y147_BLUT (
.I0(CLBLM_R_X7Y153_SLICE_X8Y153_A5Q),
.I1(CLBLM_R_X7Y153_SLICE_X9Y153_A5Q),
.I2(CLBLM_R_X11Y147_SLICE_X15Y147_BO6),
.I3(CLBLM_R_X7Y144_SLICE_X9Y144_B5Q),
.I4(CLBLM_L_X10Y144_SLICE_X12Y144_AQ),
.I5(1'b1),
.O5(CLBLM_L_X10Y147_SLICE_X12Y147_BO5),
.O6(CLBLM_L_X10Y147_SLICE_X12Y147_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaa00ff22222222)
  ) CLBLM_L_X10Y147_SLICE_X12Y147_ALUT (
.I0(CLBLL_L_X4Y142_SLICE_X5Y142_DQ),
.I1(CLBLL_L_X4Y147_SLICE_X5Y147_CQ),
.I2(1'b1),
.I3(CLBLM_L_X10Y146_SLICE_X13Y146_DO6),
.I4(LIOB33_X0Y61_IOB_X0Y62_I),
.I5(1'b1),
.O5(CLBLM_L_X10Y147_SLICE_X12Y147_AO5),
.O6(CLBLM_L_X10Y147_SLICE_X12Y147_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y147_SLICE_X13Y147_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y147_SLICE_X13Y147_AO6),
.Q(CLBLM_L_X10Y147_SLICE_X13Y147_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h00000000a0a0c0c0)
  ) CLBLM_L_X10Y147_SLICE_X13Y147_DLUT (
.I0(CLBLM_L_X8Y147_SLICE_X11Y147_C5Q),
.I1(CLBLM_L_X10Y143_SLICE_X13Y143_CQ),
.I2(CLBLM_R_X7Y144_SLICE_X9Y144_B5Q),
.I3(1'b1),
.I4(CLBLM_R_X7Y153_SLICE_X8Y153_A5Q),
.I5(CLBLM_R_X11Y147_SLICE_X15Y147_BO6),
.O5(CLBLM_L_X10Y147_SLICE_X13Y147_DO5),
.O6(CLBLM_L_X10Y147_SLICE_X13Y147_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000001000000055)
  ) CLBLM_L_X10Y147_SLICE_X13Y147_CLUT (
.I0(CLBLM_L_X8Y148_SLICE_X11Y148_CO6),
.I1(CLBLM_L_X8Y145_SLICE_X10Y145_CO6),
.I2(CLBLM_R_X11Y145_SLICE_X14Y145_DO6),
.I3(CLBLM_L_X10Y150_SLICE_X13Y150_DO6),
.I4(CLBLM_L_X8Y147_SLICE_X10Y147_DO6),
.I5(CLBLM_L_X12Y147_SLICE_X16Y147_DO6),
.O5(CLBLM_L_X10Y147_SLICE_X13Y147_CO5),
.O6(CLBLM_L_X10Y147_SLICE_X13Y147_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffffffffeffff)
  ) CLBLM_L_X10Y147_SLICE_X13Y147_BLUT (
.I0(CLBLM_L_X10Y146_SLICE_X12Y146_DQ),
.I1(CLBLM_R_X5Y142_SLICE_X6Y142_D5Q),
.I2(CLBLM_R_X7Y151_SLICE_X8Y151_D5Q),
.I3(CLBLL_L_X4Y147_SLICE_X4Y147_CQ),
.I4(CLBLL_L_X4Y148_SLICE_X4Y148_CQ),
.I5(CLBLM_R_X7Y149_SLICE_X8Y149_AQ),
.O5(CLBLM_L_X10Y147_SLICE_X13Y147_BO5),
.O6(CLBLM_L_X10Y147_SLICE_X13Y147_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hff00ff00f0f0f4f4)
  ) CLBLM_L_X10Y147_SLICE_X13Y147_ALUT (
.I0(CLBLM_L_X10Y146_SLICE_X13Y146_DO5),
.I1(CLBLM_L_X10Y145_SLICE_X13Y145_BO6),
.I2(CLBLM_L_X10Y147_SLICE_X13Y147_AQ),
.I3(CLBLM_R_X7Y147_SLICE_X9Y147_A5Q),
.I4(RIOB33_X105Y131_IOB_X1Y132_I),
.I5(LIOB33_X0Y61_IOB_X0Y62_I),
.O5(CLBLM_L_X10Y147_SLICE_X13Y147_AO5),
.O6(CLBLM_L_X10Y147_SLICE_X13Y147_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y148_SLICE_X12Y148_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y147_SLICE_X12Y147_AO6),
.Q(CLBLM_L_X10Y148_SLICE_X12Y148_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h00aa00aa30ba30ba)
  ) CLBLM_L_X10Y148_SLICE_X12Y148_DLUT (
.I0(CLBLM_L_X8Y147_SLICE_X11Y147_CQ),
.I1(CLBLL_L_X4Y148_SLICE_X4Y148_CQ),
.I2(CLBLM_L_X10Y153_SLICE_X13Y153_A5Q),
.I3(CLBLM_L_X10Y148_SLICE_X12Y148_AO5),
.I4(1'b1),
.I5(CLBLM_L_X12Y146_SLICE_X16Y146_CO6),
.O5(CLBLM_L_X10Y148_SLICE_X12Y148_DO5),
.O6(CLBLM_L_X10Y148_SLICE_X12Y148_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hffcfffefffccffee)
  ) CLBLM_L_X10Y148_SLICE_X12Y148_CLUT (
.I0(CLBLM_R_X7Y148_SLICE_X9Y148_BQ),
.I1(CLBLM_L_X10Y149_SLICE_X13Y149_CO6),
.I2(CLBLM_L_X10Y151_SLICE_X13Y151_BO6),
.I3(CLBLM_L_X10Y147_SLICE_X12Y147_BO5),
.I4(CLBLM_L_X12Y149_SLICE_X17Y149_BO5),
.I5(CLBLM_R_X5Y146_SLICE_X6Y146_AQ),
.O5(CLBLM_L_X10Y148_SLICE_X12Y148_CO5),
.O6(CLBLM_L_X10Y148_SLICE_X12Y148_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000202000002200)
  ) CLBLM_L_X10Y148_SLICE_X12Y148_BLUT (
.I0(CLBLM_R_X7Y149_SLICE_X8Y149_AQ),
.I1(CLBLM_L_X12Y147_SLICE_X16Y147_DO6),
.I2(CLBLM_R_X5Y146_SLICE_X6Y146_B5Q),
.I3(CLBLM_L_X10Y148_SLICE_X13Y148_BQ),
.I4(CLBLM_L_X10Y147_SLICE_X12Y147_BO6),
.I5(CLBLL_L_X4Y148_SLICE_X4Y148_CQ),
.O5(CLBLM_L_X10Y148_SLICE_X12Y148_BO5),
.O6(CLBLM_L_X10Y148_SLICE_X12Y148_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffefffffffdffff)
  ) CLBLM_L_X10Y148_SLICE_X12Y148_ALUT (
.I0(CLBLM_R_X7Y153_SLICE_X8Y153_A5Q),
.I1(CLBLM_R_X7Y149_SLICE_X8Y149_AQ),
.I2(CLBLL_L_X4Y148_SLICE_X4Y148_CQ),
.I3(CLBLM_R_X7Y146_SLICE_X9Y146_CO6),
.I4(CLBLM_R_X7Y144_SLICE_X9Y144_B5Q),
.I5(1'b1),
.O5(CLBLM_L_X10Y148_SLICE_X12Y148_AO5),
.O6(CLBLM_L_X10Y148_SLICE_X12Y148_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y148_SLICE_X13Y148_C5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y148_SLICE_X13Y148_CO5),
.Q(CLBLM_L_X10Y148_SLICE_X13Y148_C5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y148_SLICE_X13Y148_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y148_SLICE_X13Y148_AO6),
.Q(CLBLM_L_X10Y148_SLICE_X13Y148_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y148_SLICE_X13Y148_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y148_SLICE_X13Y148_BO6),
.Q(CLBLM_L_X10Y148_SLICE_X13Y148_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y148_SLICE_X13Y148_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y148_SLICE_X13Y148_CO6),
.Q(CLBLM_L_X10Y148_SLICE_X13Y148_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffeffffffffffff)
  ) CLBLM_L_X10Y148_SLICE_X13Y148_DLUT (
.I0(CLBLM_L_X10Y142_SLICE_X13Y142_BO6),
.I1(CLBLM_L_X12Y145_SLICE_X17Y145_BO6),
.I2(CLBLM_R_X5Y148_SLICE_X6Y148_DO6),
.I3(CLBLM_R_X3Y142_SLICE_X2Y142_BO5),
.I4(CLBLM_L_X10Y144_SLICE_X13Y144_A5Q),
.I5(CLBLM_R_X11Y152_SLICE_X14Y152_AO6),
.O5(CLBLM_L_X10Y148_SLICE_X13Y148_DO5),
.O6(CLBLM_L_X10Y148_SLICE_X13Y148_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hee44ee44eeee4444)
  ) CLBLM_L_X10Y148_SLICE_X13Y148_CLUT (
.I0(LIOB33_X0Y61_IOB_X0Y62_I),
.I1(CLBLM_R_X3Y151_SLICE_X3Y151_CQ),
.I2(1'b1),
.I3(CLBLM_L_X8Y143_SLICE_X11Y143_D5Q),
.I4(CLBLM_L_X12Y146_SLICE_X16Y146_DQ),
.I5(1'b1),
.O5(CLBLM_L_X10Y148_SLICE_X13Y148_CO5),
.O6(CLBLM_L_X10Y148_SLICE_X13Y148_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfff0ffcc00f000cc)
  ) CLBLM_L_X10Y148_SLICE_X13Y148_BLUT (
.I0(1'b1),
.I1(CLBLM_L_X10Y148_SLICE_X13Y148_BQ),
.I2(CLBLM_L_X8Y147_SLICE_X11Y147_BQ),
.I3(LIOB33_X0Y61_IOB_X0Y62_I),
.I4(CLBLM_R_X13Y149_SLICE_X18Y149_AO6),
.I5(CLBLM_R_X7Y151_SLICE_X8Y151_BQ),
.O5(CLBLM_L_X10Y148_SLICE_X13Y148_BO5),
.O6(CLBLM_L_X10Y148_SLICE_X13Y148_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffc800c8fffa00fa)
  ) CLBLM_L_X10Y148_SLICE_X13Y148_ALUT (
.I0(CLBLM_L_X10Y148_SLICE_X13Y148_CQ),
.I1(CLBLM_L_X10Y145_SLICE_X12Y145_AQ),
.I2(CLBLM_L_X10Y148_SLICE_X13Y148_AQ),
.I3(LIOB33_X0Y61_IOB_X0Y62_I),
.I4(CLBLM_L_X10Y148_SLICE_X12Y148_AQ),
.I5(CLBLM_R_X5Y142_SLICE_X7Y142_BQ),
.O5(CLBLM_L_X10Y148_SLICE_X13Y148_AO5),
.O6(CLBLM_L_X10Y148_SLICE_X13Y148_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y149_SLICE_X12Y149_A5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y149_SLICE_X12Y149_AO5),
.Q(CLBLM_L_X10Y149_SLICE_X12Y149_A5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y149_SLICE_X12Y149_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y149_SLICE_X12Y149_AO6),
.Q(CLBLM_L_X10Y149_SLICE_X12Y149_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y149_SLICE_X12Y149_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X12Y149_SLICE_X17Y149_AO6),
.Q(CLBLM_L_X10Y149_SLICE_X12Y149_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffffffffffcc)
  ) CLBLM_L_X10Y149_SLICE_X12Y149_DLUT (
.I0(1'b1),
.I1(CLBLM_L_X10Y150_SLICE_X12Y150_AO5),
.I2(1'b1),
.I3(CLBLM_R_X7Y149_SLICE_X8Y149_DO6),
.I4(CLBLM_L_X8Y149_SLICE_X11Y149_DO6),
.I5(CLBLM_R_X7Y150_SLICE_X9Y150_BO6),
.O5(CLBLM_L_X10Y149_SLICE_X12Y149_DO5),
.O6(CLBLM_L_X10Y149_SLICE_X12Y149_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffffffffffa2)
  ) CLBLM_L_X10Y149_SLICE_X12Y149_CLUT (
.I0(CLBLM_L_X12Y147_SLICE_X16Y147_DO6),
.I1(CLBLM_R_X11Y148_SLICE_X15Y148_BO6),
.I2(CLBLM_L_X10Y147_SLICE_X12Y147_DO6),
.I3(CLBLM_R_X7Y149_SLICE_X8Y149_DO6),
.I4(CLBLM_L_X10Y150_SLICE_X12Y150_CO6),
.I5(CLBLM_R_X7Y150_SLICE_X9Y150_BO6),
.O5(CLBLM_L_X10Y149_SLICE_X12Y149_CO5),
.O6(CLBLM_L_X10Y149_SLICE_X12Y149_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hcfcccccc10111111)
  ) CLBLM_L_X10Y149_SLICE_X12Y149_BLUT (
.I0(CLBLM_L_X10Y145_SLICE_X12Y145_BQ),
.I1(CLBLM_L_X8Y154_SLICE_X10Y154_BO5),
.I2(CLBLL_L_X4Y153_SLICE_X5Y153_A5Q),
.I3(CLBLM_R_X7Y145_SLICE_X8Y145_A5Q),
.I4(RIOB33_X105Y131_IOB_X1Y131_I),
.I5(1'b1),
.O5(CLBLM_L_X10Y149_SLICE_X12Y149_BO5),
.O6(CLBLM_L_X10Y149_SLICE_X12Y149_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfafa5050ee44ee44)
  ) CLBLM_L_X10Y149_SLICE_X12Y149_ALUT (
.I0(LIOB33_X0Y61_IOB_X0Y62_I),
.I1(CLBLL_L_X4Y150_SLICE_X4Y150_B5Q),
.I2(CLBLM_R_X3Y145_SLICE_X3Y145_BQ),
.I3(CLBLM_L_X10Y152_SLICE_X12Y152_AQ),
.I4(CLBLM_L_X10Y146_SLICE_X13Y146_AQ),
.I5(1'b1),
.O5(CLBLM_L_X10Y149_SLICE_X12Y149_AO5),
.O6(CLBLM_L_X10Y149_SLICE_X12Y149_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y149_SLICE_X13Y149_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y149_SLICE_X13Y149_AO6),
.Q(CLBLM_L_X10Y149_SLICE_X13Y149_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hff0aff0affceffce)
  ) CLBLM_L_X10Y149_SLICE_X13Y149_DLUT (
.I0(CLBLM_R_X5Y149_SLICE_X7Y149_CQ),
.I1(CLBLM_R_X7Y151_SLICE_X8Y151_BQ),
.I2(CLBLM_L_X10Y148_SLICE_X12Y148_AO6),
.I3(CLBLM_L_X10Y147_SLICE_X13Y147_DO6),
.I4(1'b1),
.I5(CLBLM_L_X12Y149_SLICE_X17Y149_CO6),
.O5(CLBLM_L_X10Y149_SLICE_X13Y149_DO5),
.O6(CLBLM_L_X10Y149_SLICE_X13Y149_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff0000ffff44f4)
  ) CLBLM_L_X10Y149_SLICE_X13Y149_CLUT (
.I0(CLBLM_R_X11Y144_SLICE_X14Y144_CO6),
.I1(CLBLM_L_X10Y150_SLICE_X13Y150_AQ),
.I2(CLBLM_R_X7Y151_SLICE_X8Y151_DQ),
.I3(CLBLM_R_X11Y144_SLICE_X14Y144_BO6),
.I4(CLBLM_L_X10Y146_SLICE_X13Y146_DO6),
.I5(CLBLM_L_X10Y147_SLICE_X12Y147_BO6),
.O5(CLBLM_L_X10Y149_SLICE_X13Y149_CO5),
.O6(CLBLM_L_X10Y149_SLICE_X13Y149_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hdc00ffffcc00ffff)
  ) CLBLM_L_X10Y149_SLICE_X13Y149_BLUT (
.I0(CLBLL_L_X4Y151_SLICE_X4Y151_CQ),
.I1(RIOB33_X105Y101_IOB_X1Y101_I),
.I2(CLBLM_L_X8Y142_SLICE_X11Y142_BQ),
.I3(CLBLM_L_X10Y149_SLICE_X12Y149_BO5),
.I4(RIOB33_SING_X105Y100_IOB_X1Y100_I),
.I5(RIOB33_X105Y131_IOB_X1Y131_I),
.O5(CLBLM_L_X10Y149_SLICE_X13Y149_BO5),
.O6(CLBLM_L_X10Y149_SLICE_X13Y149_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hbb11bb113f3f3f3f)
  ) CLBLM_L_X10Y149_SLICE_X13Y149_ALUT (
.I0(LIOB33_X0Y61_IOB_X0Y62_I),
.I1(CLBLM_L_X10Y147_SLICE_X13Y147_CO6),
.I2(CLBLM_L_X10Y148_SLICE_X12Y148_AQ),
.I3(CLBLM_R_X7Y145_SLICE_X8Y145_AQ),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X10Y149_SLICE_X13Y149_AO5),
.O6(CLBLM_L_X10Y149_SLICE_X13Y149_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y150_SLICE_X12Y150_A_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(LIOB33_X0Y61_IOB_X0Y62_I),
.D(CLBLM_L_X10Y151_SLICE_X12Y151_BQ),
.Q(CLBLM_L_X10Y150_SLICE_X12Y150_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h00004c0c00004400)
  ) CLBLM_L_X10Y150_SLICE_X12Y150_DLUT (
.I0(CLBLM_R_X11Y144_SLICE_X14Y144_BO6),
.I1(CLBLM_R_X7Y144_SLICE_X9Y144_B5Q),
.I2(CLBLM_R_X11Y147_SLICE_X15Y147_BO6),
.I3(CLBLM_R_X7Y147_SLICE_X9Y147_D5Q),
.I4(CLBLM_R_X7Y153_SLICE_X8Y153_A5Q),
.I5(CLBLM_L_X8Y151_SLICE_X10Y151_C5Q),
.O5(CLBLM_L_X10Y150_SLICE_X12Y150_DO5),
.O6(CLBLM_L_X10Y150_SLICE_X12Y150_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hffafffaaffefffee)
  ) CLBLM_L_X10Y150_SLICE_X12Y150_CLUT (
.I0(CLBLM_L_X10Y150_SLICE_X12Y150_AO6),
.I1(CLBLM_L_X8Y151_SLICE_X10Y151_C5Q),
.I2(CLBLM_L_X10Y148_SLICE_X12Y148_AO6),
.I3(CLBLM_L_X8Y149_SLICE_X11Y149_DO6),
.I4(CLBLM_R_X7Y147_SLICE_X9Y147_D5Q),
.I5(CLBLM_L_X10Y150_SLICE_X12Y150_BO6),
.O5(CLBLM_L_X10Y150_SLICE_X12Y150_CO5),
.O6(CLBLM_L_X10Y150_SLICE_X12Y150_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffefffffffdffff)
  ) CLBLM_L_X10Y150_SLICE_X12Y150_BLUT (
.I0(CLBLM_R_X7Y153_SLICE_X8Y153_A5Q),
.I1(CLBLM_L_X12Y147_SLICE_X16Y147_DO6),
.I2(CLBLM_R_X7Y149_SLICE_X8Y149_AQ),
.I3(CLBLL_L_X4Y148_SLICE_X4Y148_CQ),
.I4(CLBLM_R_X7Y144_SLICE_X9Y144_B5Q),
.I5(1'b1),
.O5(CLBLM_L_X10Y150_SLICE_X12Y150_BO5),
.O6(CLBLM_L_X10Y150_SLICE_X12Y150_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h3f0f3300bfafbbaa)
  ) CLBLM_L_X10Y150_SLICE_X12Y150_ALUT (
.I0(CLBLM_L_X10Y150_SLICE_X12Y150_DO6),
.I1(CLBLM_L_X10Y151_SLICE_X13Y151_BO5),
.I2(CLBLM_L_X12Y149_SLICE_X17Y149_CO6),
.I3(CLBLM_L_X8Y151_SLICE_X10Y151_AQ),
.I4(CLBLM_L_X8Y150_SLICE_X11Y150_AQ),
.I5(1'b1),
.O5(CLBLM_L_X10Y150_SLICE_X12Y150_AO5),
.O6(CLBLM_L_X10Y150_SLICE_X12Y150_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y150_SLICE_X13Y150_A_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_L_X10Y150_SLICE_X13Y150_AO6),
.Q(CLBLM_L_X10Y150_SLICE_X13Y150_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hffceffceffffffce)
  ) CLBLM_L_X10Y150_SLICE_X13Y150_DLUT (
.I0(CLBLM_L_X8Y145_SLICE_X11Y145_CQ),
.I1(CLBLM_L_X10Y146_SLICE_X13Y146_DO6),
.I2(CLBLM_L_X10Y150_SLICE_X12Y150_BO5),
.I3(CLBLM_L_X10Y150_SLICE_X13Y150_CO6),
.I4(CLBLM_L_X10Y147_SLICE_X12Y147_BQ),
.I5(CLBLM_L_X10Y151_SLICE_X13Y151_BO5),
.O5(CLBLM_L_X10Y150_SLICE_X13Y150_DO5),
.O6(CLBLM_L_X10Y150_SLICE_X13Y150_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0001000000000000)
  ) CLBLM_L_X10Y150_SLICE_X13Y150_CLUT (
.I0(CLBLM_R_X7Y149_SLICE_X8Y149_AQ),
.I1(CLBLM_L_X12Y147_SLICE_X16Y147_DO6),
.I2(CLBLM_R_X7Y153_SLICE_X8Y153_A5Q),
.I3(CLBLL_L_X4Y148_SLICE_X4Y148_CQ),
.I4(CLBLM_R_X7Y144_SLICE_X9Y144_B5Q),
.I5(CLBLM_L_X8Y149_SLICE_X11Y149_A5Q),
.O5(CLBLM_L_X10Y150_SLICE_X13Y150_CO5),
.O6(CLBLM_L_X10Y150_SLICE_X13Y150_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h30ff3030baffbaba)
  ) CLBLM_L_X10Y150_SLICE_X13Y150_BLUT (
.I0(CLBLM_R_X11Y150_SLICE_X14Y150_DO6),
.I1(CLBLM_L_X10Y151_SLICE_X13Y151_BO6),
.I2(CLBLM_R_X5Y148_SLICE_X7Y148_BQ),
.I3(CLBLM_L_X10Y151_SLICE_X13Y151_BO5),
.I4(CLBLM_L_X10Y150_SLICE_X12Y150_AQ),
.I5(1'b1),
.O5(CLBLM_L_X10Y150_SLICE_X13Y150_BO5),
.O6(CLBLM_L_X10Y150_SLICE_X13Y150_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaaaaaaff00f0f0)
  ) CLBLM_L_X10Y150_SLICE_X13Y150_ALUT (
.I0(CLBLM_R_X7Y151_SLICE_X8Y151_DQ),
.I1(1'b1),
.I2(CLBLM_L_X10Y150_SLICE_X13Y150_AQ),
.I3(CLBLL_L_X4Y150_SLICE_X5Y150_BQ),
.I4(CLBLM_R_X13Y149_SLICE_X18Y149_AO6),
.I5(LIOB33_X0Y61_IOB_X0Y62_I),
.O5(CLBLM_L_X10Y150_SLICE_X13Y150_AO5),
.O6(CLBLM_L_X10Y150_SLICE_X13Y150_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y151_SLICE_X12Y151_A_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_L_X10Y151_SLICE_X12Y151_AO6),
.Q(CLBLM_L_X10Y151_SLICE_X12Y151_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y151_SLICE_X12Y151_B_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_L_X10Y151_SLICE_X12Y151_BO6),
.Q(CLBLM_L_X10Y151_SLICE_X12Y151_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y151_SLICE_X12Y151_C_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_L_X10Y151_SLICE_X12Y151_CO6),
.Q(CLBLM_L_X10Y151_SLICE_X12Y151_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y151_SLICE_X12Y151_D_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_L_X10Y151_SLICE_X12Y151_DO6),
.Q(CLBLM_L_X10Y151_SLICE_X12Y151_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaafff0aaaa00f0)
  ) CLBLM_L_X10Y151_SLICE_X12Y151_DLUT (
.I0(CLBLM_L_X8Y151_SLICE_X11Y151_AQ),
.I1(1'b1),
.I2(CLBLM_L_X10Y151_SLICE_X12Y151_DQ),
.I3(CLBLM_L_X12Y149_SLICE_X17Y149_CO6),
.I4(LIOB33_X0Y61_IOB_X0Y62_I),
.I5(CLBLM_L_X8Y142_SLICE_X11Y142_AQ),
.O5(CLBLM_L_X10Y151_SLICE_X12Y151_DO5),
.O6(CLBLM_L_X10Y151_SLICE_X12Y151_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaaf0ccaaaaf0cc)
  ) CLBLM_L_X10Y151_SLICE_X12Y151_CLUT (
.I0(CLBLM_L_X8Y152_SLICE_X11Y152_AQ),
.I1(CLBLM_L_X10Y151_SLICE_X12Y151_CQ),
.I2(CLBLM_L_X10Y151_SLICE_X12Y151_BQ),
.I3(CLBLM_R_X11Y148_SLICE_X15Y148_AO6),
.I4(LIOB33_X0Y61_IOB_X0Y62_I),
.I5(1'b1),
.O5(CLBLM_L_X10Y151_SLICE_X12Y151_CO5),
.O6(CLBLM_L_X10Y151_SLICE_X12Y151_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfaff5055eaee4044)
  ) CLBLM_L_X10Y151_SLICE_X12Y151_BLUT (
.I0(LIOB33_X0Y61_IOB_X0Y62_I),
.I1(CLBLM_L_X8Y143_SLICE_X11Y143_D5Q),
.I2(CLBLL_L_X4Y147_SLICE_X5Y147_CQ),
.I3(CLBLL_L_X4Y142_SLICE_X5Y142_DQ),
.I4(CLBLM_L_X8Y146_SLICE_X11Y146_D5Q),
.I5(CLBLM_L_X10Y151_SLICE_X12Y151_BQ),
.O5(CLBLM_L_X10Y151_SLICE_X12Y151_BO5),
.O6(CLBLM_L_X10Y151_SLICE_X12Y151_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hbbb88888bbb8bbb8)
  ) CLBLM_L_X10Y151_SLICE_X12Y151_ALUT (
.I0(CLBLM_L_X10Y152_SLICE_X13Y152_CQ),
.I1(LIOB33_X0Y61_IOB_X0Y62_I),
.I2(CLBLM_L_X10Y151_SLICE_X12Y151_AQ),
.I3(CLBLM_L_X10Y149_SLICE_X12Y149_A5Q),
.I4(CLBLM_L_X10Y145_SLICE_X12Y145_AQ),
.I5(CLBLM_R_X5Y142_SLICE_X7Y142_BQ),
.O5(CLBLM_L_X10Y151_SLICE_X12Y151_AO5),
.O6(CLBLM_L_X10Y151_SLICE_X12Y151_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y151_SLICE_X13Y151_A5_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_L_X10Y151_SLICE_X13Y151_AO5),
.Q(CLBLM_L_X10Y151_SLICE_X13Y151_A5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y151_SLICE_X13Y151_A_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_L_X10Y151_SLICE_X13Y151_AO6),
.Q(CLBLM_L_X10Y151_SLICE_X13Y151_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hababaaaaaaa8aaa8)
  ) CLBLM_L_X10Y151_SLICE_X13Y151_DLUT (
.I0(CLBLM_L_X8Y151_SLICE_X11Y151_AQ),
.I1(CLBLM_R_X7Y153_SLICE_X8Y153_A5Q),
.I2(CLBLM_L_X10Y147_SLICE_X13Y147_BO6),
.I3(CLBLM_L_X10Y146_SLICE_X13Y146_DO6),
.I4(CLBLM_L_X10Y151_SLICE_X12Y151_DQ),
.I5(CLBLM_R_X7Y144_SLICE_X9Y144_B5Q),
.O5(CLBLM_L_X10Y151_SLICE_X13Y151_DO5),
.O6(CLBLM_L_X10Y151_SLICE_X13Y151_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h00000000008000a0)
  ) CLBLM_L_X10Y151_SLICE_X13Y151_CLUT (
.I0(CLBLM_R_X3Y150_SLICE_X2Y150_AQ),
.I1(CLBLM_L_X12Y149_SLICE_X17Y149_CO6),
.I2(CLBLM_R_X5Y153_SLICE_X7Y153_DO6),
.I3(CLBLM_L_X10Y148_SLICE_X13Y148_DO6),
.I4(CLBLM_L_X10Y151_SLICE_X12Y151_DQ),
.I5(CLBLM_R_X13Y146_SLICE_X18Y146_BO6),
.O5(CLBLM_L_X10Y151_SLICE_X13Y151_CO5),
.O6(CLBLM_L_X10Y151_SLICE_X13Y151_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'heffffffffffffffe)
  ) CLBLM_L_X10Y151_SLICE_X13Y151_BLUT (
.I0(CLBLM_R_X7Y149_SLICE_X8Y149_AQ),
.I1(CLBLM_L_X12Y147_SLICE_X16Y147_DO6),
.I2(CLBLM_R_X7Y153_SLICE_X8Y153_A5Q),
.I3(CLBLL_L_X4Y148_SLICE_X4Y148_CQ),
.I4(CLBLM_R_X7Y144_SLICE_X9Y144_B5Q),
.I5(1'b1),
.O5(CLBLM_L_X10Y151_SLICE_X13Y151_BO5),
.O6(CLBLM_L_X10Y151_SLICE_X13Y151_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfafa5050bb11bb11)
  ) CLBLM_L_X10Y151_SLICE_X13Y151_ALUT (
.I0(LIOB33_X0Y61_IOB_X0Y62_I),
.I1(CLBLM_R_X11Y148_SLICE_X14Y148_BO6),
.I2(CLBLM_L_X10Y149_SLICE_X12Y149_CO6),
.I3(CLBLM_R_X7Y151_SLICE_X8Y151_CQ),
.I4(CLBLM_L_X10Y145_SLICE_X13Y145_AQ),
.I5(1'b1),
.O5(CLBLM_L_X10Y151_SLICE_X13Y151_AO5),
.O6(CLBLM_L_X10Y151_SLICE_X13Y151_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y152_SLICE_X12Y152_A_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_L_X10Y152_SLICE_X12Y152_AO6),
.Q(CLBLM_L_X10Y152_SLICE_X12Y152_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y152_SLICE_X12Y152_B_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_L_X10Y152_SLICE_X12Y152_BO6),
.Q(CLBLM_L_X10Y152_SLICE_X12Y152_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y152_SLICE_X12Y152_C_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_L_X10Y152_SLICE_X12Y152_CO6),
.Q(CLBLM_L_X10Y152_SLICE_X12Y152_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h5500f7085500f708)
  ) CLBLM_L_X10Y152_SLICE_X12Y152_DLUT (
.I0(CLBLM_R_X7Y146_SLICE_X8Y146_A5Q),
.I1(CLBLM_L_X10Y152_SLICE_X12Y152_AQ),
.I2(CLBLM_R_X5Y147_SLICE_X6Y147_AQ),
.I3(CLBLM_L_X8Y152_SLICE_X10Y152_CQ),
.I4(CLBLM_L_X10Y153_SLICE_X13Y153_CQ),
.I5(1'b1),
.O5(CLBLM_L_X10Y152_SLICE_X12Y152_DO5),
.O6(CLBLM_L_X10Y152_SLICE_X12Y152_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f0aaccf0f0aacc)
  ) CLBLM_L_X10Y152_SLICE_X12Y152_CLUT (
.I0(CLBLM_L_X8Y152_SLICE_X11Y152_AQ),
.I1(CLBLM_L_X10Y152_SLICE_X12Y152_CQ),
.I2(CLBLM_L_X10Y153_SLICE_X13Y153_AQ),
.I3(CLBLM_R_X13Y149_SLICE_X18Y149_AO6),
.I4(LIOB33_X0Y61_IOB_X0Y62_I),
.I5(1'b1),
.O5(CLBLM_L_X10Y152_SLICE_X12Y152_CO5),
.O6(CLBLM_L_X10Y152_SLICE_X12Y152_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffc00fcff540054)
  ) CLBLM_L_X10Y152_SLICE_X12Y152_BLUT (
.I0(CLBLL_L_X4Y142_SLICE_X5Y142_DQ),
.I1(CLBLM_L_X10Y152_SLICE_X12Y152_BQ),
.I2(CLBLM_L_X8Y146_SLICE_X11Y146_D5Q),
.I3(LIOB33_X0Y61_IOB_X0Y62_I),
.I4(CLBLM_R_X7Y146_SLICE_X8Y146_A5Q),
.I5(CLBLL_L_X4Y147_SLICE_X5Y147_CQ),
.O5(CLBLM_L_X10Y152_SLICE_X12Y152_BO5),
.O6(CLBLM_L_X10Y152_SLICE_X12Y152_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hcccc00f0cccca5f0)
  ) CLBLM_L_X10Y152_SLICE_X12Y152_ALUT (
.I0(CLBLM_R_X5Y147_SLICE_X6Y147_AQ),
.I1(CLBLM_L_X10Y149_SLICE_X12Y149_AQ),
.I2(CLBLM_L_X10Y152_SLICE_X12Y152_AQ),
.I3(CLBLM_R_X7Y146_SLICE_X8Y146_A5Q),
.I4(LIOB33_X0Y61_IOB_X0Y62_I),
.I5(CLBLM_L_X10Y153_SLICE_X13Y153_CQ),
.O5(CLBLM_L_X10Y152_SLICE_X12Y152_AO5),
.O6(CLBLM_L_X10Y152_SLICE_X12Y152_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y152_SLICE_X13Y152_A_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_L_X10Y152_SLICE_X13Y152_AO6),
.Q(CLBLM_L_X10Y152_SLICE_X13Y152_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y152_SLICE_X13Y152_B_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_L_X10Y152_SLICE_X13Y152_BO6),
.Q(CLBLM_L_X10Y152_SLICE_X13Y152_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y152_SLICE_X13Y152_C_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_L_X10Y152_SLICE_X13Y152_CO6),
.Q(CLBLM_L_X10Y152_SLICE_X13Y152_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000200000000000)
  ) CLBLM_L_X10Y152_SLICE_X13Y152_DLUT (
.I0(CLBLM_L_X10Y152_SLICE_X12Y152_AQ),
.I1(CLBLM_L_X10Y153_SLICE_X13Y153_CQ),
.I2(CLBLM_R_X11Y153_SLICE_X14Y153_AQ),
.I3(CLBLM_L_X8Y152_SLICE_X10Y152_CQ),
.I4(CLBLM_R_X5Y147_SLICE_X6Y147_AQ),
.I5(CLBLM_R_X7Y146_SLICE_X8Y146_A5Q),
.O5(CLBLM_L_X10Y152_SLICE_X13Y152_DO5),
.O6(CLBLM_L_X10Y152_SLICE_X13Y152_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f0ffccf0f000cc)
  ) CLBLM_L_X10Y152_SLICE_X13Y152_CLUT (
.I0(1'b1),
.I1(CLBLM_L_X10Y152_SLICE_X13Y152_CQ),
.I2(CLBLM_R_X5Y146_SLICE_X7Y146_AQ),
.I3(CLBLM_R_X11Y148_SLICE_X15Y148_AO6),
.I4(LIOB33_X0Y61_IOB_X0Y62_I),
.I5(CLBLM_L_X10Y152_SLICE_X12Y152_BQ),
.O5(CLBLM_L_X10Y152_SLICE_X13Y152_CO5),
.O6(CLBLM_L_X10Y152_SLICE_X13Y152_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfeee5444baaa1000)
  ) CLBLM_L_X10Y152_SLICE_X13Y152_BLUT (
.I0(LIOB33_X0Y61_IOB_X0Y62_I),
.I1(CLBLM_L_X10Y152_SLICE_X13Y152_BQ),
.I2(CLBLM_L_X10Y152_SLICE_X13Y152_AQ),
.I3(CLBLM_L_X10Y152_SLICE_X13Y152_DO6),
.I4(CLBLM_L_X8Y149_SLICE_X11Y149_A5Q),
.I5(CLBLM_L_X10Y153_SLICE_X13Y153_DO6),
.O5(CLBLM_L_X10Y152_SLICE_X13Y152_BO5),
.O6(CLBLM_L_X10Y152_SLICE_X13Y152_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hddd8ddd88d888d88)
  ) CLBLM_L_X10Y152_SLICE_X13Y152_ALUT (
.I0(LIOB33_X0Y61_IOB_X0Y62_I),
.I1(CLBLM_L_X8Y151_SLICE_X10Y151_C5Q),
.I2(CLBLM_L_X10Y152_SLICE_X13Y152_AQ),
.I3(CLBLM_L_X10Y152_SLICE_X13Y152_DO6),
.I4(1'b1),
.I5(CLBLM_L_X10Y153_SLICE_X13Y153_DO6),
.O5(CLBLM_L_X10Y152_SLICE_X13Y152_AO5),
.O6(CLBLM_L_X10Y152_SLICE_X13Y152_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y153_SLICE_X12Y153_A5_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_L_X10Y153_SLICE_X12Y153_CO6),
.Q(CLBLM_L_X10Y153_SLICE_X12Y153_A5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y153_SLICE_X12Y153_A_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_L_X10Y153_SLICE_X12Y153_AO6),
.Q(CLBLM_L_X10Y153_SLICE_X12Y153_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y153_SLICE_X12Y153_B_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_L_X10Y153_SLICE_X12Y153_BO6),
.Q(CLBLM_L_X10Y153_SLICE_X12Y153_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h1101ffff1111ffff)
  ) CLBLM_L_X10Y153_SLICE_X12Y153_DLUT (
.I0(CLBLM_L_X10Y145_SLICE_X12Y145_BQ),
.I1(CLBLM_L_X8Y154_SLICE_X10Y154_BO5),
.I2(RIOB33_X105Y131_IOB_X1Y131_I),
.I3(CLBLL_L_X4Y153_SLICE_X5Y153_A5Q),
.I4(RIOB33_SING_X105Y100_IOB_X1Y100_I),
.I5(CLBLM_R_X7Y145_SLICE_X8Y145_A5Q),
.O5(CLBLM_L_X10Y153_SLICE_X12Y153_DO5),
.O6(CLBLM_L_X10Y153_SLICE_X12Y153_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h888b88b8f0f00000)
  ) CLBLM_L_X10Y153_SLICE_X12Y153_CLUT (
.I0(CLBLM_L_X10Y147_SLICE_X12Y147_AQ),
.I1(LIOB33_X0Y61_IOB_X0Y62_I),
.I2(CLBLM_L_X10Y153_SLICE_X12Y153_A5Q),
.I3(CLBLM_R_X5Y150_SLICE_X6Y150_B5Q),
.I4(CLBLM_R_X5Y152_SLICE_X6Y152_BQ),
.I5(1'b1),
.O5(CLBLM_L_X10Y153_SLICE_X12Y153_CO5),
.O6(CLBLM_L_X10Y153_SLICE_X12Y153_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f00000f9fc090c)
  ) CLBLM_L_X10Y153_SLICE_X12Y153_BLUT (
.I0(CLBLM_R_X7Y154_SLICE_X8Y154_DO6),
.I1(CLBLM_L_X10Y153_SLICE_X12Y153_BQ),
.I2(LIOB33_X0Y61_IOB_X0Y62_I),
.I3(CLBLM_R_X5Y152_SLICE_X6Y152_BQ),
.I4(CLBLM_L_X12Y146_SLICE_X16Y146_BQ),
.I5(CLBLM_R_X5Y150_SLICE_X6Y150_B5Q),
.O5(CLBLM_L_X10Y153_SLICE_X12Y153_BO5),
.O6(CLBLM_L_X10Y153_SLICE_X12Y153_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hff00ff0044444444)
  ) CLBLM_L_X10Y153_SLICE_X12Y153_ALUT (
.I0(CLBLM_R_X7Y154_SLICE_X8Y154_DO6),
.I1(CLBLM_L_X10Y153_SLICE_X12Y153_BQ),
.I2(1'b1),
.I3(CLBLM_L_X10Y153_SLICE_X13Y153_BQ),
.I4(1'b1),
.I5(LIOB33_X0Y61_IOB_X0Y62_I),
.O5(CLBLM_L_X10Y153_SLICE_X12Y153_AO5),
.O6(CLBLM_L_X10Y153_SLICE_X12Y153_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y153_SLICE_X13Y153_A5_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_L_X12Y153_SLICE_X16Y153_AO5),
.Q(CLBLM_L_X10Y153_SLICE_X13Y153_A5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y153_SLICE_X13Y153_A_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_L_X10Y153_SLICE_X13Y153_AO6),
.Q(CLBLM_L_X10Y153_SLICE_X13Y153_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y153_SLICE_X13Y153_B_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_L_X10Y153_SLICE_X13Y153_BO6),
.Q(CLBLM_L_X10Y153_SLICE_X13Y153_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y153_SLICE_X13Y153_C_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_L_X10Y153_SLICE_X13Y153_CO6),
.Q(CLBLM_L_X10Y153_SLICE_X13Y153_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h1555555555555555)
  ) CLBLM_L_X10Y153_SLICE_X13Y153_DLUT (
.I0(CLBLM_L_X10Y155_SLICE_X12Y155_BO5),
.I1(CLBLM_L_X10Y155_SLICE_X13Y155_AO5),
.I2(CLBLM_L_X10Y152_SLICE_X13Y152_AQ),
.I3(CLBLM_L_X8Y152_SLICE_X10Y152_CQ),
.I4(CLBLM_L_X10Y152_SLICE_X12Y152_AQ),
.I5(CLBLM_R_X11Y153_SLICE_X14Y153_AQ),
.O5(CLBLM_L_X10Y153_SLICE_X13Y153_DO5),
.O6(CLBLM_L_X10Y153_SLICE_X13Y153_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaaaaaaff303030)
  ) CLBLM_L_X10Y153_SLICE_X13Y153_CLUT (
.I0(CLBLM_R_X5Y152_SLICE_X6Y152_DQ),
.I1(CLBLM_R_X7Y146_SLICE_X8Y146_A5Q),
.I2(CLBLM_L_X10Y153_SLICE_X13Y153_CQ),
.I3(CLBLM_L_X10Y154_SLICE_X13Y154_CO6),
.I4(CLBLM_L_X10Y153_SLICE_X13Y153_AQ),
.I5(LIOB33_X0Y61_IOB_X0Y62_I),
.O5(CLBLM_L_X10Y153_SLICE_X13Y153_CO5),
.O6(CLBLM_L_X10Y153_SLICE_X13Y153_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hff8b008bff880088)
  ) CLBLM_L_X10Y153_SLICE_X13Y153_BLUT (
.I0(CLBLM_R_X11Y153_SLICE_X15Y153_CO6),
.I1(CLBLM_L_X10Y153_SLICE_X13Y153_BQ),
.I2(CLBLM_R_X11Y153_SLICE_X15Y153_DO6),
.I3(LIOB33_X0Y61_IOB_X0Y62_I),
.I4(CLBLL_L_X4Y151_SLICE_X5Y151_BQ),
.I5(CLBLM_R_X11Y153_SLICE_X15Y153_BO5),
.O5(CLBLM_L_X10Y153_SLICE_X13Y153_BO5),
.O6(CLBLM_L_X10Y153_SLICE_X13Y153_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hcfef0323ccec0020)
  ) CLBLM_L_X10Y153_SLICE_X13Y153_ALUT (
.I0(CLBLM_L_X10Y154_SLICE_X13Y154_BO5),
.I1(LIOB33_X0Y61_IOB_X0Y62_I),
.I2(CLBLM_L_X10Y153_SLICE_X13Y153_AQ),
.I3(CLBLM_L_X10Y155_SLICE_X12Y155_BO5),
.I4(CLBLM_R_X7Y151_SLICE_X9Y151_BQ),
.I5(CLBLM_L_X10Y154_SLICE_X13Y154_CO6),
.O5(CLBLM_L_X10Y153_SLICE_X13Y153_AO5),
.O6(CLBLM_L_X10Y153_SLICE_X13Y153_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y154_SLICE_X12Y154_A5_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_L_X10Y154_SLICE_X12Y154_CO6),
.Q(CLBLM_L_X10Y154_SLICE_X12Y154_A5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y154_SLICE_X12Y154_B5_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_L_X10Y154_SLICE_X12Y154_DO6),
.Q(CLBLM_L_X10Y154_SLICE_X12Y154_B5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y154_SLICE_X12Y154_A_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_L_X10Y154_SLICE_X12Y154_AO6),
.Q(CLBLM_L_X10Y154_SLICE_X12Y154_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y154_SLICE_X12Y154_B_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_L_X10Y154_SLICE_X12Y154_BO6),
.Q(CLBLM_L_X10Y154_SLICE_X12Y154_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hff02000230303030)
  ) CLBLM_L_X10Y154_SLICE_X12Y154_DLUT (
.I0(RIOB33_X105Y131_IOB_X1Y131_I),
.I1(CLBLM_R_X5Y142_SLICE_X7Y142_CO6),
.I2(RIOB33_SING_X105Y100_IOB_X1Y100_I),
.I3(LIOB33_X0Y61_IOB_X0Y62_I),
.I4(CLBLM_L_X10Y154_SLICE_X12Y154_BQ),
.I5(1'b1),
.O5(CLBLM_L_X10Y154_SLICE_X12Y154_DO5),
.O6(CLBLM_L_X10Y154_SLICE_X12Y154_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f0aacc0f0f0f0f)
  ) CLBLM_L_X10Y154_SLICE_X12Y154_CLUT (
.I0(CLBLM_L_X10Y155_SLICE_X13Y155_BO6),
.I1(CLBLM_L_X10Y155_SLICE_X13Y155_CO6),
.I2(CLBLM_R_X3Y150_SLICE_X2Y150_BQ),
.I3(CLBLM_L_X10Y154_SLICE_X12Y154_A5Q),
.I4(LIOB33_X0Y61_IOB_X0Y62_I),
.I5(1'b1),
.O5(CLBLM_L_X10Y154_SLICE_X12Y154_CO5),
.O6(CLBLM_L_X10Y154_SLICE_X12Y154_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf5b1e4a0e4a0e4a0)
  ) CLBLM_L_X10Y154_SLICE_X12Y154_BLUT (
.I0(LIOB33_X0Y61_IOB_X0Y62_I),
.I1(CLBLM_L_X10Y154_SLICE_X12Y154_BQ),
.I2(CLBLM_R_X7Y152_SLICE_X8Y152_B5Q),
.I3(CLBLM_L_X10Y155_SLICE_X13Y155_BO6),
.I4(CLBLM_L_X10Y154_SLICE_X12Y154_A5Q),
.I5(CLBLM_L_X10Y155_SLICE_X13Y155_CO6),
.O5(CLBLM_L_X10Y154_SLICE_X12Y154_BO5),
.O6(CLBLM_L_X10Y154_SLICE_X12Y154_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfbfa5150abaa0100)
  ) CLBLM_L_X10Y154_SLICE_X12Y154_ALUT (
.I0(LIOB33_X0Y61_IOB_X0Y62_I),
.I1(CLBLM_L_X10Y154_SLICE_X13Y154_BO6),
.I2(CLBLM_L_X10Y154_SLICE_X12Y154_AQ),
.I3(CLBLM_L_X10Y155_SLICE_X13Y155_CO6),
.I4(CLBLM_R_X7Y154_SLICE_X9Y154_BQ),
.I5(CLBLM_L_X10Y154_SLICE_X13Y154_DO6),
.O5(CLBLM_L_X10Y154_SLICE_X12Y154_AO5),
.O6(CLBLM_L_X10Y154_SLICE_X12Y154_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y154_SLICE_X13Y154_A_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_L_X10Y154_SLICE_X13Y154_AO6),
.Q(CLBLM_L_X10Y154_SLICE_X13Y154_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h007f7f7f00ffffff)
  ) CLBLM_L_X10Y154_SLICE_X13Y154_DLUT (
.I0(CLBLM_L_X10Y154_SLICE_X12Y154_AQ),
.I1(CLBLM_L_X10Y154_SLICE_X12Y154_A5Q),
.I2(CLBLM_L_X10Y155_SLICE_X13Y155_AO6),
.I3(CLBLM_R_X7Y146_SLICE_X8Y146_A5Q),
.I4(CLBLM_L_X10Y153_SLICE_X13Y153_CQ),
.I5(CLBLM_L_X10Y154_SLICE_X12Y154_BQ),
.O5(CLBLM_L_X10Y154_SLICE_X13Y154_DO5),
.O6(CLBLM_L_X10Y154_SLICE_X13Y154_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h8000000080008000)
  ) CLBLM_L_X10Y154_SLICE_X13Y154_CLUT (
.I0(CLBLM_L_X10Y154_SLICE_X12Y154_AQ),
.I1(CLBLM_L_X10Y154_SLICE_X12Y154_A5Q),
.I2(CLBLM_L_X10Y154_SLICE_X12Y154_BQ),
.I3(CLBLM_L_X10Y155_SLICE_X13Y155_CO6),
.I4(CLBLM_L_X10Y154_SLICE_X13Y154_AQ),
.I5(1'b1),
.O5(CLBLM_L_X10Y154_SLICE_X13Y154_CO5),
.O6(CLBLM_L_X10Y154_SLICE_X13Y154_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0fff0fff7fffffff)
  ) CLBLM_L_X10Y154_SLICE_X13Y154_BLUT (
.I0(CLBLM_L_X10Y154_SLICE_X13Y154_AQ),
.I1(CLBLM_L_X10Y155_SLICE_X13Y155_AO6),
.I2(CLBLM_L_X10Y154_SLICE_X12Y154_A5Q),
.I3(CLBLM_L_X10Y154_SLICE_X12Y154_BQ),
.I4(CLBLM_L_X10Y154_SLICE_X12Y154_AQ),
.I5(1'b1),
.O5(CLBLM_L_X10Y154_SLICE_X13Y154_BO5),
.O6(CLBLM_L_X10Y154_SLICE_X13Y154_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffafffa000af00a0)
  ) CLBLM_L_X10Y154_SLICE_X13Y154_ALUT (
.I0(CLBLM_L_X10Y154_SLICE_X13Y154_DO6),
.I1(1'b1),
.I2(CLBLM_L_X10Y154_SLICE_X13Y154_AQ),
.I3(LIOB33_X0Y61_IOB_X0Y62_I),
.I4(CLBLM_L_X10Y154_SLICE_X13Y154_CO5),
.I5(CLBLM_L_X8Y145_SLICE_X11Y145_CQ),
.O5(CLBLM_L_X10Y154_SLICE_X13Y154_AO5),
.O6(CLBLM_L_X10Y154_SLICE_X13Y154_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y155_SLICE_X12Y155_A_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_L_X10Y155_SLICE_X12Y155_AO6),
.Q(CLBLM_L_X10Y155_SLICE_X12Y155_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X10Y155_SLICE_X12Y155_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X10Y155_SLICE_X12Y155_DO5),
.O6(CLBLM_L_X10Y155_SLICE_X12Y155_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X10Y155_SLICE_X12Y155_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X10Y155_SLICE_X12Y155_CO5),
.O6(CLBLM_L_X10Y155_SLICE_X12Y155_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffbffffff000000)
  ) CLBLM_L_X10Y155_SLICE_X12Y155_BLUT (
.I0(CLBLM_R_X5Y147_SLICE_X6Y147_AQ),
.I1(CLBLM_L_X10Y153_SLICE_X13Y153_BQ),
.I2(CLBLM_R_X11Y153_SLICE_X15Y153_DO6),
.I3(CLBLM_L_X10Y153_SLICE_X13Y153_CQ),
.I4(CLBLM_R_X7Y146_SLICE_X8Y146_A5Q),
.I5(1'b1),
.O5(CLBLM_L_X10Y155_SLICE_X12Y155_BO5),
.O6(CLBLM_L_X10Y155_SLICE_X12Y155_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'haaafbabf00051015)
  ) CLBLM_L_X10Y155_SLICE_X12Y155_ALUT (
.I0(LIOB33_X0Y61_IOB_X0Y62_I),
.I1(CLBLM_L_X10Y155_SLICE_X12Y155_BO5),
.I2(CLBLM_L_X10Y155_SLICE_X12Y155_AQ),
.I3(CLBLM_L_X10Y155_SLICE_X12Y155_BO6),
.I4(CLBLM_L_X10Y155_SLICE_X13Y155_AO6),
.I5(CLBLM_R_X5Y146_SLICE_X7Y146_CQ),
.O5(CLBLM_L_X10Y155_SLICE_X12Y155_AO5),
.O6(CLBLM_L_X10Y155_SLICE_X12Y155_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X10Y155_SLICE_X13Y155_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X10Y155_SLICE_X13Y155_DO5),
.O6(CLBLM_L_X10Y155_SLICE_X13Y155_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000020000000000)
  ) CLBLM_L_X10Y155_SLICE_X13Y155_CLUT (
.I0(CLBLM_L_X10Y155_SLICE_X12Y155_AQ),
.I1(CLBLM_L_X10Y153_SLICE_X13Y153_CQ),
.I2(CLBLM_R_X5Y147_SLICE_X6Y147_AQ),
.I3(CLBLM_L_X10Y153_SLICE_X13Y153_BQ),
.I4(CLBLM_R_X11Y153_SLICE_X15Y153_DO6),
.I5(CLBLM_R_X7Y146_SLICE_X8Y146_A5Q),
.O5(CLBLM_L_X10Y155_SLICE_X13Y155_CO5),
.O6(CLBLM_L_X10Y155_SLICE_X13Y155_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h00f700ff00ff00ff)
  ) CLBLM_L_X10Y155_SLICE_X13Y155_BLUT (
.I0(CLBLM_L_X10Y154_SLICE_X12Y154_A5Q),
.I1(CLBLM_L_X10Y153_SLICE_X13Y153_BQ),
.I2(CLBLM_R_X11Y153_SLICE_X15Y153_DO6),
.I3(CLBLM_L_X10Y155_SLICE_X12Y155_BO5),
.I4(CLBLM_L_X10Y155_SLICE_X12Y155_AQ),
.I5(CLBLM_L_X10Y155_SLICE_X13Y155_AO5),
.O5(CLBLM_L_X10Y155_SLICE_X13Y155_BO5),
.O6(CLBLM_L_X10Y155_SLICE_X13Y155_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0400000044444444)
  ) CLBLM_L_X10Y155_SLICE_X13Y155_ALUT (
.I0(CLBLM_R_X5Y147_SLICE_X6Y147_AQ),
.I1(CLBLM_R_X7Y146_SLICE_X8Y146_A5Q),
.I2(CLBLM_R_X11Y153_SLICE_X15Y153_DO6),
.I3(CLBLM_L_X10Y153_SLICE_X13Y153_BQ),
.I4(CLBLM_L_X10Y155_SLICE_X12Y155_AQ),
.I5(1'b1),
.O5(CLBLM_L_X10Y155_SLICE_X13Y155_AO5),
.O6(CLBLM_L_X10Y155_SLICE_X13Y155_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y145_SLICE_X16Y145_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(LIOB33_X0Y61_IOB_X0Y62_I),
.D(CLBLM_R_X11Y145_SLICE_X15Y145_AQ),
.Q(CLBLM_L_X12Y145_SLICE_X16Y145_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'heaeaeaeac0c0c0c0)
  ) CLBLM_L_X12Y145_SLICE_X16Y145_DLUT (
.I0(CLBLM_R_X7Y147_SLICE_X8Y147_AQ),
.I1(CLBLM_L_X12Y145_SLICE_X16Y145_AQ),
.I2(RIOB33_X105Y135_IOB_X1Y136_I),
.I3(1'b1),
.I4(1'b1),
.I5(RIOB33_X105Y137_IOB_X1Y137_I),
.O5(CLBLM_L_X12Y145_SLICE_X16Y145_DO5),
.O6(CLBLM_L_X12Y145_SLICE_X16Y145_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hbbaafbfabbaafbfa)
  ) CLBLM_L_X12Y145_SLICE_X16Y145_CLUT (
.I0(CLBLM_L_X12Y145_SLICE_X16Y145_AO6),
.I1(CLBLM_L_X12Y145_SLICE_X17Y145_AO5),
.I2(CLBLM_L_X10Y143_SLICE_X13Y143_AQ),
.I3(RIOB33_X105Y133_IOB_X1Y134_I),
.I4(CLBLM_L_X12Y146_SLICE_X16Y146_CO6),
.I5(1'b1),
.O5(CLBLM_L_X12Y145_SLICE_X16Y145_CO5),
.O6(CLBLM_L_X12Y145_SLICE_X16Y145_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfefefafafc54fcfc)
  ) CLBLM_L_X12Y145_SLICE_X16Y145_BLUT (
.I0(CLBLM_R_X7Y149_SLICE_X8Y149_AQ),
.I1(CLBLL_L_X4Y148_SLICE_X4Y148_CQ),
.I2(CLBLM_L_X12Y145_SLICE_X17Y145_DO6),
.I3(CLBLM_R_X7Y146_SLICE_X9Y146_CO6),
.I4(CLBLM_R_X7Y144_SLICE_X9Y144_B5Q),
.I5(CLBLM_R_X7Y153_SLICE_X8Y153_A5Q),
.O5(CLBLM_L_X12Y145_SLICE_X16Y145_BO5),
.O6(CLBLM_L_X12Y145_SLICE_X16Y145_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h03000202fcfcffff)
  ) CLBLM_L_X12Y145_SLICE_X16Y145_ALUT (
.I0(RIOB33_X105Y141_IOB_X1Y142_I),
.I1(CLBLM_R_X7Y144_SLICE_X9Y144_B5Q),
.I2(CLBLM_L_X12Y145_SLICE_X17Y145_CO6),
.I3(CLBLM_L_X12Y146_SLICE_X16Y146_CQ),
.I4(CLBLM_R_X7Y153_SLICE_X8Y153_A5Q),
.I5(1'b1),
.O5(CLBLM_L_X12Y145_SLICE_X16Y145_AO5),
.O6(CLBLM_L_X12Y145_SLICE_X16Y145_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h7fff7fff7fff7fff)
  ) CLBLM_L_X12Y145_SLICE_X17Y145_DLUT (
.I0(CLBLM_R_X5Y142_SLICE_X6Y142_D5Q),
.I1(CLBLL_L_X4Y147_SLICE_X4Y147_CQ),
.I2(CLBLM_L_X10Y146_SLICE_X12Y146_DQ),
.I3(CLBLM_R_X7Y151_SLICE_X8Y151_D5Q),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X12Y145_SLICE_X17Y145_DO5),
.O6(CLBLM_L_X12Y145_SLICE_X17Y145_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffffff7ffffff)
  ) CLBLM_L_X12Y145_SLICE_X17Y145_CLUT (
.I0(CLBLM_R_X5Y142_SLICE_X6Y142_D5Q),
.I1(CLBLL_L_X4Y147_SLICE_X4Y147_CQ),
.I2(CLBLM_R_X7Y149_SLICE_X8Y149_AQ),
.I3(CLBLM_R_X7Y151_SLICE_X8Y151_D5Q),
.I4(CLBLM_L_X10Y146_SLICE_X12Y146_DQ),
.I5(CLBLL_L_X4Y148_SLICE_X4Y148_CQ),
.O5(CLBLM_L_X12Y145_SLICE_X17Y145_CO5),
.O6(CLBLM_L_X12Y145_SLICE_X17Y145_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfff8ff88f8f88888)
  ) CLBLM_L_X12Y145_SLICE_X17Y145_BLUT (
.I0(RIOB33_X105Y141_IOB_X1Y142_I),
.I1(CLBLM_L_X12Y146_SLICE_X16Y146_CQ),
.I2(RIOB33_X105Y143_IOB_X1Y144_I),
.I3(RIOB33_X105Y143_IOB_X1Y143_I),
.I4(CLBLM_R_X5Y148_SLICE_X6Y148_CQ),
.I5(CLBLM_L_X12Y146_SLICE_X16Y146_AQ),
.O5(CLBLM_L_X12Y145_SLICE_X17Y145_BO5),
.O6(CLBLM_L_X12Y145_SLICE_X17Y145_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffdffffffbff)
  ) CLBLM_L_X12Y145_SLICE_X17Y145_ALUT (
.I0(CLBLM_R_X7Y149_SLICE_X8Y149_AQ),
.I1(CLBLM_R_X7Y153_SLICE_X8Y153_A5Q),
.I2(CLBLM_R_X7Y144_SLICE_X9Y144_B5Q),
.I3(CLBLL_L_X4Y148_SLICE_X4Y148_CQ),
.I4(CLBLM_L_X12Y145_SLICE_X17Y145_DO6),
.I5(1'b1),
.O5(CLBLM_L_X12Y145_SLICE_X17Y145_AO5),
.O6(CLBLM_L_X12Y145_SLICE_X17Y145_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y146_SLICE_X16Y146_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(LIOB33_X0Y61_IOB_X0Y62_I),
.D(CLBLM_R_X5Y144_SLICE_X6Y144_CQ),
.Q(CLBLM_L_X12Y146_SLICE_X16Y146_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y146_SLICE_X16Y146_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(LIOB33_X0Y61_IOB_X0Y62_I),
.D(CLBLM_L_X12Y146_SLICE_X16Y146_AQ),
.Q(CLBLM_L_X12Y146_SLICE_X16Y146_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y146_SLICE_X16Y146_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(LIOB33_X0Y61_IOB_X0Y62_I),
.D(CLBLM_L_X8Y152_SLICE_X11Y152_D5Q),
.Q(CLBLM_L_X12Y146_SLICE_X16Y146_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y146_SLICE_X16Y146_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(LIOB33_X0Y61_IOB_X0Y62_I),
.D(CLBLM_L_X12Y146_SLICE_X16Y146_CQ),
.Q(CLBLM_L_X12Y146_SLICE_X16Y146_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h000b0000000b000b)
  ) CLBLM_L_X12Y146_SLICE_X16Y146_DLUT (
.I0(CLBLM_L_X12Y145_SLICE_X17Y145_AO5),
.I1(RIOB33_X105Y147_IOB_X1Y147_I),
.I2(CLBLM_R_X11Y146_SLICE_X15Y146_CO6),
.I3(CLBLM_L_X12Y146_SLICE_X16Y146_AO5),
.I4(CLBLM_R_X11Y146_SLICE_X14Y146_DO6),
.I5(CLBLM_L_X12Y145_SLICE_X16Y145_BO6),
.O5(CLBLM_L_X12Y146_SLICE_X16Y146_DO5),
.O6(CLBLM_L_X12Y146_SLICE_X16Y146_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffffffffdffff)
  ) CLBLM_L_X12Y146_SLICE_X16Y146_CLUT (
.I0(CLBLM_R_X5Y142_SLICE_X6Y142_D5Q),
.I1(CLBLL_L_X4Y147_SLICE_X4Y147_CQ),
.I2(CLBLM_L_X10Y147_SLICE_X12Y147_BO6),
.I3(CLBLM_L_X10Y146_SLICE_X12Y146_DQ),
.I4(CLBLM_R_X7Y149_SLICE_X8Y149_AQ),
.I5(CLBLM_R_X7Y151_SLICE_X8Y151_D5Q),
.O5(CLBLM_L_X12Y146_SLICE_X16Y146_CO5),
.O6(CLBLM_L_X12Y146_SLICE_X16Y146_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'haabaaaaaaabababa)
  ) CLBLM_L_X12Y146_SLICE_X16Y146_BLUT (
.I0(CLBLM_R_X11Y144_SLICE_X14Y144_DO6),
.I1(CLBLM_L_X12Y145_SLICE_X16Y145_CO6),
.I2(CLBLM_L_X12Y146_SLICE_X17Y146_CO6),
.I3(CLBLM_L_X12Y145_SLICE_X16Y145_BO6),
.I4(CLBLM_R_X13Y146_SLICE_X18Y146_BO6),
.I5(CLBLM_L_X10Y146_SLICE_X13Y146_CQ),
.O5(CLBLM_L_X12Y146_SLICE_X16Y146_BO5),
.O6(CLBLM_L_X12Y146_SLICE_X16Y146_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0011001105000000)
  ) CLBLM_L_X12Y146_SLICE_X16Y146_ALUT (
.I0(CLBLM_R_X7Y153_SLICE_X8Y153_A5Q),
.I1(CLBLM_L_X10Y146_SLICE_X13Y146_DO6),
.I2(CLBLM_L_X12Y145_SLICE_X17Y145_CO6),
.I3(CLBLM_R_X7Y144_SLICE_X9Y144_B5Q),
.I4(RIOB33_X105Y141_IOB_X1Y141_I),
.I5(1'b1),
.O5(CLBLM_L_X12Y146_SLICE_X16Y146_AO5),
.O6(CLBLM_L_X12Y146_SLICE_X16Y146_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y146_SLICE_X17Y146_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X12Y146_SLICE_X17Y146_AO6),
.Q(CLBLM_L_X12Y146_SLICE_X17Y146_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hc4f5c4f50000c4f5)
  ) CLBLM_L_X12Y146_SLICE_X17Y146_DLUT (
.I0(CLBLM_L_X10Y147_SLICE_X13Y147_AQ),
.I1(CLBLM_L_X12Y147_SLICE_X17Y147_AO6),
.I2(CLBLM_L_X12Y145_SLICE_X17Y145_AO6),
.I3(CLBLM_R_X11Y150_SLICE_X14Y150_AQ),
.I4(RIOB33_X105Y139_IOB_X1Y139_I),
.I5(CLBLM_R_X13Y146_SLICE_X18Y146_AO6),
.O5(CLBLM_L_X12Y146_SLICE_X17Y146_DO5),
.O6(CLBLM_L_X12Y146_SLICE_X17Y146_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h88aaccff080a0c0f)
  ) CLBLM_L_X12Y146_SLICE_X17Y146_CLUT (
.I0(CLBLM_R_X13Y146_SLICE_X18Y146_AO6),
.I1(CLBLM_L_X12Y147_SLICE_X17Y147_AO6),
.I2(CLBLM_R_X11Y146_SLICE_X14Y146_AQ),
.I3(CLBLM_L_X10Y147_SLICE_X12Y147_AQ),
.I4(RIOB33_X105Y139_IOB_X1Y140_I),
.I5(CLBLM_L_X12Y145_SLICE_X17Y145_AO6),
.O5(CLBLM_L_X12Y146_SLICE_X17Y146_CO5),
.O6(CLBLM_L_X12Y146_SLICE_X17Y146_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffffffffefffc)
  ) CLBLM_L_X12Y146_SLICE_X17Y146_BLUT (
.I0(CLBLM_L_X12Y146_SLICE_X16Y146_DQ),
.I1(CLBLM_L_X12Y145_SLICE_X16Y145_DO6),
.I2(CLBLM_L_X12Y145_SLICE_X17Y145_BO6),
.I3(CLBLM_R_X11Y146_SLICE_X15Y146_AO5),
.I4(RIOB33_X105Y145_IOB_X1Y146_I),
.I5(CLBLM_L_X12Y147_SLICE_X17Y147_CO6),
.O5(CLBLM_L_X12Y146_SLICE_X17Y146_BO5),
.O6(CLBLM_L_X12Y146_SLICE_X17Y146_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffe0f0efffc0f0c)
  ) CLBLM_L_X12Y146_SLICE_X17Y146_ALUT (
.I0(CLBLM_R_X11Y150_SLICE_X14Y150_AQ),
.I1(CLBLM_R_X13Y146_SLICE_X18Y146_CO6),
.I2(LIOB33_X0Y61_IOB_X0Y62_I),
.I3(CLBLM_L_X12Y146_SLICE_X17Y146_BO6),
.I4(CLBLM_R_X7Y145_SLICE_X8Y145_DQ),
.I5(RIOB33_X105Y139_IOB_X1Y139_I),
.O5(CLBLM_L_X12Y146_SLICE_X17Y146_AO5),
.O6(CLBLM_L_X12Y146_SLICE_X17Y146_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffffffffcfffc)
  ) CLBLM_L_X12Y147_SLICE_X16Y147_DLUT (
.I0(1'b1),
.I1(CLBLM_R_X7Y151_SLICE_X8Y151_D5Q),
.I2(CLBLM_L_X10Y146_SLICE_X12Y146_DQ),
.I3(CLBLL_L_X4Y147_SLICE_X4Y147_CQ),
.I4(1'b1),
.I5(CLBLM_R_X5Y142_SLICE_X6Y142_D5Q),
.O5(CLBLM_L_X12Y147_SLICE_X16Y147_DO5),
.O6(CLBLM_L_X12Y147_SLICE_X16Y147_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hcceecceefcfefcfe)
  ) CLBLM_L_X12Y147_SLICE_X16Y147_CLUT (
.I0(CLBLM_L_X8Y147_SLICE_X11Y147_AQ),
.I1(CLBLM_L_X12Y147_SLICE_X17Y147_AO5),
.I2(RIOB33_X105Y145_IOB_X1Y145_I),
.I3(CLBLM_L_X12Y146_SLICE_X16Y146_CO6),
.I4(1'b1),
.I5(CLBLM_L_X12Y148_SLICE_X16Y148_AO6),
.O5(CLBLM_L_X12Y147_SLICE_X16Y147_CO5),
.O6(CLBLM_L_X12Y147_SLICE_X16Y147_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0030aaba00300030)
  ) CLBLM_L_X12Y147_SLICE_X16Y147_BLUT (
.I0(RIOB33_X105Y145_IOB_X1Y145_I),
.I1(CLBLM_R_X11Y147_SLICE_X14Y147_AO5),
.I2(CLBLM_L_X8Y147_SLICE_X11Y147_AQ),
.I3(CLBLM_R_X7Y146_SLICE_X9Y146_CO6),
.I4(CLBLM_L_X12Y145_SLICE_X17Y145_CO6),
.I5(CLBLM_L_X12Y147_SLICE_X16Y147_AO5),
.O5(CLBLM_L_X12Y147_SLICE_X16Y147_BO5),
.O6(CLBLM_L_X12Y147_SLICE_X16Y147_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0d00080000550055)
  ) CLBLM_L_X12Y147_SLICE_X16Y147_ALUT (
.I0(CLBLM_R_X7Y153_SLICE_X8Y153_A5Q),
.I1(CLBLM_L_X8Y149_SLICE_X10Y149_AQ),
.I2(CLBLM_L_X12Y145_SLICE_X17Y145_CO6),
.I3(CLBLM_R_X7Y144_SLICE_X9Y144_B5Q),
.I4(RIOB33_X105Y135_IOB_X1Y135_I),
.I5(1'b1),
.O5(CLBLM_L_X12Y147_SLICE_X16Y147_AO5),
.O6(CLBLM_L_X12Y147_SLICE_X16Y147_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'ha0a0f0f0aaaaffff)
  ) CLBLM_L_X12Y147_SLICE_X17Y147_DLUT (
.I0(CLBLM_L_X12Y145_SLICE_X17Y145_AO5),
.I1(1'b1),
.I2(CLBLM_R_X13Y146_SLICE_X18Y146_AO6),
.I3(1'b1),
.I4(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.I5(RIOB33_X105Y137_IOB_X1Y138_I),
.O5(CLBLM_L_X12Y147_SLICE_X17Y147_DO5),
.O6(CLBLM_L_X12Y147_SLICE_X17Y147_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hfafaf0f0aaaa0000)
  ) CLBLM_L_X12Y147_SLICE_X17Y147_CLUT (
.I0(CLBLM_L_X8Y149_SLICE_X10Y149_AQ),
.I1(1'b1),
.I2(CLBLM_R_X7Y148_SLICE_X8Y148_AQ),
.I3(1'b1),
.I4(RIOB33_X105Y135_IOB_X1Y135_I),
.I5(RIOB33_X105Y137_IOB_X1Y138_I),
.O5(CLBLM_L_X12Y147_SLICE_X17Y147_CO5),
.O6(CLBLM_L_X12Y147_SLICE_X17Y147_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000020223033)
  ) CLBLM_L_X12Y147_SLICE_X17Y147_BLUT (
.I0(CLBLM_R_X13Y146_SLICE_X18Y146_AO6),
.I1(CLBLM_L_X12Y147_SLICE_X16Y147_BO6),
.I2(CLBLM_L_X12Y145_SLICE_X17Y145_AO5),
.I3(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.I4(RIOB33_X105Y137_IOB_X1Y138_I),
.I5(CLBLM_L_X12Y147_SLICE_X17Y147_AO5),
.O5(CLBLM_L_X12Y147_SLICE_X17Y147_BO5),
.O6(CLBLM_L_X12Y147_SLICE_X17Y147_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff3f3f00008c80)
  ) CLBLM_L_X12Y147_SLICE_X17Y147_ALUT (
.I0(CLBLM_R_X7Y148_SLICE_X8Y148_AQ),
.I1(CLBLM_R_X7Y153_SLICE_X8Y153_A5Q),
.I2(CLBLM_R_X7Y144_SLICE_X9Y144_B5Q),
.I3(CLBLM_L_X12Y146_SLICE_X16Y146_BQ),
.I4(CLBLM_L_X12Y145_SLICE_X17Y145_CO6),
.I5(1'b1),
.O5(CLBLM_L_X12Y147_SLICE_X17Y147_AO5),
.O6(CLBLM_L_X12Y147_SLICE_X17Y147_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hff77ff55ff33ff00)
  ) CLBLM_L_X12Y148_SLICE_X16Y148_DLUT (
.I0(CLBLM_R_X13Y146_SLICE_X18Y146_AO6),
.I1(CLBLM_L_X12Y146_SLICE_X16Y146_CO6),
.I2(1'b1),
.I3(CLBLM_L_X12Y148_SLICE_X16Y148_AO5),
.I4(CLBLM_R_X5Y144_SLICE_X7Y144_AQ),
.I5(RIOB33_X105Y137_IOB_X1Y137_I),
.O5(CLBLM_L_X12Y148_SLICE_X16Y148_DO5),
.O6(CLBLM_L_X12Y148_SLICE_X16Y148_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h1100313011001100)
  ) CLBLM_L_X12Y148_SLICE_X16Y148_CLUT (
.I0(CLBLM_L_X12Y145_SLICE_X17Y145_CO6),
.I1(CLBLM_L_X10Y147_SLICE_X12Y147_BO6),
.I2(CLBLM_R_X7Y149_SLICE_X8Y149_AQ),
.I3(RIOB33_X105Y137_IOB_X1Y137_I),
.I4(CLBLM_R_X7Y146_SLICE_X9Y146_CO6),
.I5(CLBLM_R_X5Y144_SLICE_X7Y144_AQ),
.O5(CLBLM_L_X12Y148_SLICE_X16Y148_CO5),
.O6(CLBLM_L_X12Y148_SLICE_X16Y148_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000055051101)
  ) CLBLM_L_X12Y148_SLICE_X16Y148_BLUT (
.I0(CLBLM_L_X12Y148_SLICE_X16Y148_CO6),
.I1(RIOB33_X105Y145_IOB_X1Y146_I),
.I2(RIOB33_X105Y147_IOB_X1Y148_I),
.I3(CLBLM_L_X12Y145_SLICE_X17Y145_AO5),
.I4(CLBLM_L_X12Y148_SLICE_X16Y148_AO6),
.I5(CLBLM_L_X12Y148_SLICE_X16Y148_AO5),
.O5(CLBLM_L_X12Y148_SLICE_X16Y148_BO5),
.O6(CLBLM_L_X12Y148_SLICE_X16Y148_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffcfffc0c080008)
  ) CLBLM_L_X12Y148_SLICE_X16Y148_ALUT (
.I0(CLBLM_L_X12Y146_SLICE_X16Y146_DQ),
.I1(CLBLM_R_X7Y153_SLICE_X8Y153_A5Q),
.I2(CLBLM_L_X12Y145_SLICE_X17Y145_CO6),
.I3(CLBLM_R_X7Y144_SLICE_X9Y144_B5Q),
.I4(CLBLM_R_X7Y147_SLICE_X8Y147_AQ),
.I5(1'b1),
.O5(CLBLM_L_X12Y148_SLICE_X16Y148_AO5),
.O6(CLBLM_L_X12Y148_SLICE_X16Y148_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X12Y148_SLICE_X17Y148_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X12Y148_SLICE_X17Y148_DO5),
.O6(CLBLM_L_X12Y148_SLICE_X17Y148_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X12Y148_SLICE_X17Y148_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X12Y148_SLICE_X17Y148_CO5),
.O6(CLBLM_L_X12Y148_SLICE_X17Y148_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X12Y148_SLICE_X17Y148_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X12Y148_SLICE_X17Y148_BO5),
.O6(CLBLM_L_X12Y148_SLICE_X17Y148_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'haaffaaffaaffa2f3)
  ) CLBLM_L_X12Y148_SLICE_X17Y148_ALUT (
.I0(CLBLM_L_X12Y145_SLICE_X17Y145_AO5),
.I1(RIOB33_X105Y145_IOB_X1Y146_I),
.I2(CLBLM_R_X7Y144_SLICE_X9Y144_B5Q),
.I3(RIOB33_X105Y147_IOB_X1Y148_I),
.I4(CLBLM_L_X12Y145_SLICE_X17Y145_CO6),
.I5(CLBLM_R_X7Y153_SLICE_X8Y153_A5Q),
.O5(CLBLM_L_X12Y148_SLICE_X17Y148_AO5),
.O6(CLBLM_L_X12Y148_SLICE_X17Y148_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0f000000000a000a)
  ) CLBLM_L_X12Y149_SLICE_X16Y149_DLUT (
.I0(CLBLM_R_X7Y149_SLICE_X9Y149_BQ),
.I1(1'b1),
.I2(CLBLM_R_X11Y144_SLICE_X14Y144_AO6),
.I3(CLBLM_R_X7Y153_SLICE_X8Y153_A5Q),
.I4(CLBLL_L_X4Y144_SLICE_X4Y144_D5Q),
.I5(CLBLM_R_X7Y144_SLICE_X9Y144_B5Q),
.O5(CLBLM_L_X12Y149_SLICE_X16Y149_DO5),
.O6(CLBLM_L_X12Y149_SLICE_X16Y149_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0f3c03300fb403b8)
  ) CLBLM_L_X12Y149_SLICE_X16Y149_CLUT (
.I0(CLBLM_L_X12Y146_SLICE_X16Y146_BO6),
.I1(CLBLM_L_X12Y147_SLICE_X16Y147_DO6),
.I2(CLBLM_R_X11Y149_SLICE_X14Y149_DO6),
.I3(CLBLM_R_X11Y149_SLICE_X15Y149_DO6),
.I4(CLBLM_R_X11Y147_SLICE_X14Y147_DO6),
.I5(CLBLM_L_X8Y145_SLICE_X10Y145_BO6),
.O5(CLBLM_L_X12Y149_SLICE_X16Y149_CO5),
.O6(CLBLM_L_X12Y149_SLICE_X16Y149_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hff00ff00ff88ff30)
  ) CLBLM_L_X12Y149_SLICE_X16Y149_BLUT (
.I0(CLBLL_L_X4Y144_SLICE_X4Y144_D5Q),
.I1(CLBLM_R_X7Y144_SLICE_X9Y144_B5Q),
.I2(CLBLM_R_X7Y149_SLICE_X9Y149_BQ),
.I3(CLBLM_L_X8Y149_SLICE_X10Y149_AO6),
.I4(CLBLM_R_X7Y153_SLICE_X8Y153_A5Q),
.I5(CLBLM_R_X11Y144_SLICE_X14Y144_AO6),
.O5(CLBLM_L_X12Y149_SLICE_X16Y149_BO5),
.O6(CLBLM_L_X12Y149_SLICE_X16Y149_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000110031)
  ) CLBLM_L_X12Y149_SLICE_X16Y149_ALUT (
.I0(CLBLM_L_X12Y147_SLICE_X16Y147_DO6),
.I1(CLBLM_R_X11Y150_SLICE_X14Y150_BO6),
.I2(CLBLM_L_X12Y146_SLICE_X16Y146_BO6),
.I3(CLBLM_L_X12Y149_SLICE_X16Y149_BO6),
.I4(CLBLM_L_X8Y145_SLICE_X10Y145_BO6),
.I5(CLBLM_R_X7Y148_SLICE_X8Y148_CO6),
.O5(CLBLM_L_X12Y149_SLICE_X16Y149_AO5),
.O6(CLBLM_L_X12Y149_SLICE_X16Y149_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hff00ffaafff0fffa)
  ) CLBLM_L_X12Y149_SLICE_X17Y149_DLUT (
.I0(CLBLM_L_X8Y152_SLICE_X11Y152_CQ),
.I1(1'b1),
.I2(CLBLM_L_X10Y146_SLICE_X12Y146_AQ),
.I3(CLBLM_L_X10Y146_SLICE_X13Y146_DO6),
.I4(CLBLM_L_X12Y149_SLICE_X17Y149_BO5),
.I5(CLBLM_L_X12Y149_SLICE_X17Y149_BO6),
.O5(CLBLM_L_X12Y149_SLICE_X17Y149_DO5),
.O6(CLBLM_L_X12Y149_SLICE_X17Y149_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffffffffffffb)
  ) CLBLM_L_X12Y149_SLICE_X17Y149_CLUT (
.I0(CLBLM_L_X12Y147_SLICE_X16Y147_DO6),
.I1(CLBLL_L_X4Y148_SLICE_X4Y148_CQ),
.I2(CLBLM_R_X7Y149_SLICE_X8Y149_AQ),
.I3(CLBLM_R_X7Y153_SLICE_X8Y153_A5Q),
.I4(CLBLM_L_X10Y146_SLICE_X13Y146_DO6),
.I5(CLBLM_R_X7Y144_SLICE_X9Y144_B5Q),
.O5(CLBLM_L_X12Y149_SLICE_X17Y149_CO5),
.O6(CLBLM_L_X12Y149_SLICE_X17Y149_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffbffffbffff)
  ) CLBLM_L_X12Y149_SLICE_X17Y149_BLUT (
.I0(CLBLM_R_X7Y149_SLICE_X8Y149_AQ),
.I1(CLBLL_L_X4Y148_SLICE_X4Y148_CQ),
.I2(CLBLM_R_X7Y153_SLICE_X8Y153_A5Q),
.I3(CLBLM_L_X12Y147_SLICE_X16Y147_DO6),
.I4(CLBLM_R_X7Y144_SLICE_X9Y144_B5Q),
.I5(1'b1),
.O5(CLBLM_L_X12Y149_SLICE_X17Y149_BO5),
.O6(CLBLM_L_X12Y149_SLICE_X17Y149_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hbbbb11113f3f3f3f)
  ) CLBLM_L_X12Y149_SLICE_X17Y149_ALUT (
.I0(LIOB33_X0Y61_IOB_X0Y62_I),
.I1(CLBLM_R_X11Y149_SLICE_X15Y149_AO6),
.I2(CLBLM_L_X10Y148_SLICE_X12Y148_AQ),
.I3(1'b1),
.I4(CLBLM_L_X10Y148_SLICE_X13Y148_BQ),
.I5(1'b1),
.O5(CLBLM_L_X12Y149_SLICE_X17Y149_AO5),
.O6(CLBLM_L_X12Y149_SLICE_X17Y149_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X12Y150_SLICE_X16Y150_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X12Y150_SLICE_X16Y150_DO5),
.O6(CLBLM_L_X12Y150_SLICE_X16Y150_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000400000)
  ) CLBLM_L_X12Y150_SLICE_X16Y150_CLUT (
.I0(CLBLM_R_X7Y149_SLICE_X8Y149_AQ),
.I1(CLBLM_L_X10Y146_SLICE_X12Y146_AQ),
.I2(CLBLL_L_X4Y148_SLICE_X4Y148_CQ),
.I3(CLBLM_R_X7Y144_SLICE_X9Y144_B5Q),
.I4(CLBLM_R_X7Y153_SLICE_X8Y153_A5Q),
.I5(CLBLM_L_X12Y147_SLICE_X16Y147_DO6),
.O5(CLBLM_L_X12Y150_SLICE_X16Y150_CO5),
.O6(CLBLM_L_X12Y150_SLICE_X16Y150_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaaa2a2ffaaffa2)
  ) CLBLM_L_X12Y150_SLICE_X16Y150_BLUT (
.I0(CLBLM_L_X8Y152_SLICE_X10Y152_DQ),
.I1(CLBLM_L_X12Y147_SLICE_X16Y147_AO5),
.I2(CLBLM_R_X11Y144_SLICE_X14Y144_CO6),
.I3(CLBLL_L_X4Y150_SLICE_X4Y150_CQ),
.I4(CLBLM_L_X10Y146_SLICE_X13Y146_DO6),
.I5(CLBLM_R_X7Y148_SLICE_X8Y148_AO5),
.O5(CLBLM_L_X12Y150_SLICE_X16Y150_BO5),
.O6(CLBLM_L_X12Y150_SLICE_X16Y150_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0fff0fffffff00ff)
  ) CLBLM_L_X12Y150_SLICE_X16Y150_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(CLBLM_L_X8Y149_SLICE_X11Y149_BO6),
.I3(CLBLM_L_X10Y148_SLICE_X12Y148_AQ),
.I4(CLBLM_R_X11Y149_SLICE_X15Y149_CO6),
.I5(1'b1),
.O5(CLBLM_L_X12Y150_SLICE_X16Y150_AO5),
.O6(CLBLM_L_X12Y150_SLICE_X16Y150_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X12Y150_SLICE_X17Y150_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X12Y150_SLICE_X17Y150_DO5),
.O6(CLBLM_L_X12Y150_SLICE_X17Y150_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X12Y150_SLICE_X17Y150_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X12Y150_SLICE_X17Y150_CO5),
.O6(CLBLM_L_X12Y150_SLICE_X17Y150_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X12Y150_SLICE_X17Y150_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X12Y150_SLICE_X17Y150_BO5),
.O6(CLBLM_L_X12Y150_SLICE_X17Y150_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X12Y150_SLICE_X17Y150_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X12Y150_SLICE_X17Y150_AO5),
.O6(CLBLM_L_X12Y150_SLICE_X17Y150_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y151_SLICE_X16Y151_A_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_L_X12Y151_SLICE_X16Y151_AO6),
.Q(CLBLM_L_X12Y151_SLICE_X16Y151_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X12Y151_SLICE_X16Y151_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X12Y151_SLICE_X16Y151_DO5),
.O6(CLBLM_L_X12Y151_SLICE_X16Y151_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X12Y151_SLICE_X16Y151_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X12Y151_SLICE_X16Y151_CO5),
.O6(CLBLM_L_X12Y151_SLICE_X16Y151_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hff00fffff0f0ffff)
  ) CLBLM_L_X12Y151_SLICE_X16Y151_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(CLBLM_L_X10Y149_SLICE_X12Y149_CO6),
.I3(CLBLM_R_X11Y148_SLICE_X14Y148_AO6),
.I4(CLBLM_L_X10Y148_SLICE_X12Y148_AQ),
.I5(1'b1),
.O5(CLBLM_L_X12Y151_SLICE_X16Y151_BO5),
.O6(CLBLM_L_X12Y151_SLICE_X16Y151_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'haf05af050f0fffff)
  ) CLBLM_L_X12Y151_SLICE_X16Y151_ALUT (
.I0(LIOB33_X0Y61_IOB_X0Y62_I),
.I1(1'b1),
.I2(CLBLM_L_X12Y149_SLICE_X16Y149_AO6),
.I3(CLBLM_R_X11Y151_SLICE_X15Y151_A5Q),
.I4(CLBLM_L_X10Y148_SLICE_X12Y148_AQ),
.I5(1'b1),
.O5(CLBLM_L_X12Y151_SLICE_X16Y151_AO5),
.O6(CLBLM_L_X12Y151_SLICE_X16Y151_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X12Y151_SLICE_X17Y151_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X12Y151_SLICE_X17Y151_DO5),
.O6(CLBLM_L_X12Y151_SLICE_X17Y151_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X12Y151_SLICE_X17Y151_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X12Y151_SLICE_X17Y151_CO5),
.O6(CLBLM_L_X12Y151_SLICE_X17Y151_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X12Y151_SLICE_X17Y151_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X12Y151_SLICE_X17Y151_BO5),
.O6(CLBLM_L_X12Y151_SLICE_X17Y151_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X12Y151_SLICE_X17Y151_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X12Y151_SLICE_X17Y151_AO5),
.O6(CLBLM_L_X12Y151_SLICE_X17Y151_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X12Y152_SLICE_X16Y152_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X12Y152_SLICE_X16Y152_DO5),
.O6(CLBLM_L_X12Y152_SLICE_X16Y152_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X12Y152_SLICE_X16Y152_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X12Y152_SLICE_X16Y152_CO5),
.O6(CLBLM_L_X12Y152_SLICE_X16Y152_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X12Y152_SLICE_X16Y152_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X12Y152_SLICE_X16Y152_BO5),
.O6(CLBLM_L_X12Y152_SLICE_X16Y152_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'haaafaaaf0f0fffff)
  ) CLBLM_L_X12Y152_SLICE_X16Y152_ALUT (
.I0(RIOB33_X105Y133_IOB_X1Y133_I),
.I1(1'b1),
.I2(CLBLM_L_X10Y148_SLICE_X12Y148_AQ),
.I3(CLBLM_L_X8Y144_SLICE_X10Y144_BQ),
.I4(CLBLM_R_X11Y148_SLICE_X14Y148_BO6),
.I5(1'b1),
.O5(CLBLM_L_X12Y152_SLICE_X16Y152_AO5),
.O6(CLBLM_L_X12Y152_SLICE_X16Y152_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X12Y152_SLICE_X17Y152_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X12Y152_SLICE_X17Y152_DO5),
.O6(CLBLM_L_X12Y152_SLICE_X17Y152_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X12Y152_SLICE_X17Y152_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X12Y152_SLICE_X17Y152_CO5),
.O6(CLBLM_L_X12Y152_SLICE_X17Y152_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X12Y152_SLICE_X17Y152_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X12Y152_SLICE_X17Y152_BO5),
.O6(CLBLM_L_X12Y152_SLICE_X17Y152_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X12Y152_SLICE_X17Y152_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X12Y152_SLICE_X17Y152_AO5),
.O6(CLBLM_L_X12Y152_SLICE_X17Y152_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X12Y153_SLICE_X16Y153_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X12Y153_SLICE_X16Y153_DO5),
.O6(CLBLM_L_X12Y153_SLICE_X16Y153_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X12Y153_SLICE_X16Y153_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X12Y153_SLICE_X16Y153_CO5),
.O6(CLBLM_L_X12Y153_SLICE_X16Y153_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X12Y153_SLICE_X16Y153_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X12Y153_SLICE_X16Y153_BO5),
.O6(CLBLM_L_X12Y153_SLICE_X16Y153_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h3333ffffb1b1b1b1)
  ) CLBLM_L_X12Y153_SLICE_X16Y153_ALUT (
.I0(LIOB33_X0Y61_IOB_X0Y62_I),
.I1(CLBLM_R_X11Y149_SLICE_X14Y149_AO6),
.I2(CLBLM_R_X7Y153_SLICE_X9Y153_D5Q),
.I3(1'b1),
.I4(CLBLM_L_X10Y148_SLICE_X12Y148_AQ),
.I5(1'b1),
.O5(CLBLM_L_X12Y153_SLICE_X16Y153_AO5),
.O6(CLBLM_L_X12Y153_SLICE_X16Y153_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X12Y153_SLICE_X17Y153_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X12Y153_SLICE_X17Y153_DO5),
.O6(CLBLM_L_X12Y153_SLICE_X17Y153_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X12Y153_SLICE_X17Y153_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X12Y153_SLICE_X17Y153_CO5),
.O6(CLBLM_L_X12Y153_SLICE_X17Y153_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X12Y153_SLICE_X17Y153_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X12Y153_SLICE_X17Y153_BO5),
.O6(CLBLM_L_X12Y153_SLICE_X17Y153_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X12Y153_SLICE_X17Y153_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X12Y153_SLICE_X17Y153_AO5),
.O6(CLBLM_L_X12Y153_SLICE_X17Y153_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y142_SLICE_X2Y142_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y142_SLICE_X2Y142_AO6),
.Q(CLBLM_R_X3Y142_SLICE_X2Y142_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y142_SLICE_X2Y142_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y142_SLICE_X2Y142_DO5),
.O6(CLBLM_R_X3Y142_SLICE_X2Y142_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y142_SLICE_X2Y142_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y142_SLICE_X2Y142_CO5),
.O6(CLBLM_R_X3Y142_SLICE_X2Y142_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff77ffffff7fff)
  ) CLBLM_R_X3Y142_SLICE_X2Y142_BLUT (
.I0(CLBLL_L_X4Y142_SLICE_X4Y142_BQ),
.I1(CLBLM_R_X3Y142_SLICE_X3Y142_AQ),
.I2(CLBLM_R_X3Y142_SLICE_X2Y142_AQ),
.I3(CLBLM_R_X3Y143_SLICE_X2Y143_AQ),
.I4(CLBLM_R_X5Y147_SLICE_X6Y147_AQ),
.I5(1'b1),
.O5(CLBLM_R_X3Y142_SLICE_X2Y142_BO5),
.O6(CLBLM_R_X3Y142_SLICE_X2Y142_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hcccca0aacccc0000)
  ) CLBLM_R_X3Y142_SLICE_X2Y142_ALUT (
.I0(CLBLM_R_X3Y142_SLICE_X2Y142_BO5),
.I1(CLBLM_R_X3Y143_SLICE_X3Y143_AQ),
.I2(CLBLM_R_X3Y142_SLICE_X2Y142_AQ),
.I3(CLBLM_R_X3Y142_SLICE_X2Y142_BO6),
.I4(LIOB33_X0Y61_IOB_X0Y62_I),
.I5(CLBLM_L_X10Y144_SLICE_X12Y144_AO6),
.O5(CLBLM_R_X3Y142_SLICE_X2Y142_AO5),
.O6(CLBLM_R_X3Y142_SLICE_X2Y142_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y142_SLICE_X3Y142_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y142_SLICE_X3Y142_AO6),
.Q(CLBLM_R_X3Y142_SLICE_X3Y142_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y142_SLICE_X3Y142_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y142_SLICE_X3Y142_DO5),
.O6(CLBLM_R_X3Y142_SLICE_X3Y142_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffffffffffcfc)
  ) CLBLM_R_X3Y142_SLICE_X3Y142_CLUT (
.I0(1'b1),
.I1(CLBLM_R_X5Y145_SLICE_X7Y145_AQ),
.I2(CLBLL_L_X4Y143_SLICE_X4Y143_DQ),
.I3(1'b1),
.I4(CLBLM_R_X3Y145_SLICE_X2Y145_B5Q),
.I5(CLBLL_L_X4Y146_SLICE_X4Y146_C5Q),
.O5(CLBLM_R_X3Y142_SLICE_X3Y142_CO5),
.O6(CLBLM_R_X3Y142_SLICE_X3Y142_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000005)
  ) CLBLM_R_X3Y142_SLICE_X3Y142_BLUT (
.I0(CLBLM_R_X7Y146_SLICE_X8Y146_DQ),
.I1(1'b1),
.I2(CLBLM_R_X3Y147_SLICE_X3Y147_C5Q),
.I3(CLBLL_L_X4Y142_SLICE_X5Y142_CQ),
.I4(CLBLM_R_X5Y141_SLICE_X6Y141_BQ),
.I5(CLBLM_R_X3Y142_SLICE_X3Y142_CO6),
.O5(CLBLM_R_X3Y142_SLICE_X3Y142_BO5),
.O6(CLBLM_R_X3Y142_SLICE_X3Y142_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hafa0a0afa0a0a0a0)
  ) CLBLM_R_X3Y142_SLICE_X3Y142_ALUT (
.I0(CLBLM_R_X7Y142_SLICE_X9Y142_BQ),
.I1(1'b1),
.I2(LIOB33_X0Y61_IOB_X0Y62_I),
.I3(CLBLM_R_X3Y142_SLICE_X3Y142_AQ),
.I4(CLBLM_R_X5Y147_SLICE_X6Y147_AQ),
.I5(CLBLM_L_X10Y144_SLICE_X12Y144_AO6),
.O5(CLBLM_R_X3Y142_SLICE_X3Y142_AO5),
.O6(CLBLM_R_X3Y142_SLICE_X3Y142_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y143_SLICE_X2Y143_A5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y143_SLICE_X2Y143_BO6),
.Q(CLBLM_R_X3Y143_SLICE_X2Y143_A5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y143_SLICE_X2Y143_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y143_SLICE_X2Y143_AO6),
.Q(CLBLM_R_X3Y143_SLICE_X2Y143_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y143_SLICE_X2Y143_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y143_SLICE_X2Y143_DO5),
.O6(CLBLM_R_X3Y143_SLICE_X2Y143_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hff0ff00000008888)
  ) CLBLM_R_X3Y143_SLICE_X2Y143_CLUT (
.I0(CLBLL_L_X4Y142_SLICE_X4Y142_BQ),
.I1(CLBLM_R_X3Y142_SLICE_X3Y142_AQ),
.I2(LIOB33_X0Y61_IOB_X0Y62_I),
.I3(CLBLM_R_X5Y144_SLICE_X6Y144_AQ),
.I4(CLBLM_R_X5Y147_SLICE_X6Y147_AQ),
.I5(1'b1),
.O5(CLBLM_R_X3Y143_SLICE_X2Y143_CO5),
.O6(CLBLM_R_X3Y143_SLICE_X2Y143_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hb1f5e4a033333333)
  ) CLBLM_R_X3Y143_SLICE_X2Y143_BLUT (
.I0(LIOB33_X0Y61_IOB_X0Y62_I),
.I1(LIOB33_X0Y57_IOB_X0Y58_I),
.I2(CLBLL_L_X4Y145_SLICE_X4Y145_AQ),
.I3(CLBLM_R_X3Y143_SLICE_X3Y143_CQ),
.I4(CLBLM_R_X3Y143_SLICE_X2Y143_A5Q),
.I5(1'b1),
.O5(CLBLM_R_X3Y143_SLICE_X2Y143_BO5),
.O6(CLBLM_R_X3Y143_SLICE_X2Y143_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h8d88d8888d88d888)
  ) CLBLM_R_X3Y143_SLICE_X2Y143_ALUT (
.I0(LIOB33_X0Y61_IOB_X0Y62_I),
.I1(CLBLM_L_X8Y144_SLICE_X11Y144_B5Q),
.I2(CLBLM_R_X3Y143_SLICE_X2Y143_AQ),
.I3(CLBLM_L_X10Y144_SLICE_X12Y144_AO6),
.I4(CLBLM_R_X3Y143_SLICE_X2Y143_CO5),
.I5(1'b1),
.O5(CLBLM_R_X3Y143_SLICE_X2Y143_AO5),
.O6(CLBLM_R_X3Y143_SLICE_X2Y143_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y143_SLICE_X3Y143_C5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y143_SLICE_X3Y143_CO5),
.Q(CLBLM_R_X3Y143_SLICE_X3Y143_C5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y143_SLICE_X3Y143_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y143_SLICE_X3Y143_AO6),
.Q(CLBLM_R_X3Y143_SLICE_X3Y143_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y143_SLICE_X3Y143_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y143_SLICE_X3Y143_BO6),
.Q(CLBLM_R_X3Y143_SLICE_X3Y143_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y143_SLICE_X3Y143_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y143_SLICE_X3Y143_CO6),
.Q(CLBLM_R_X3Y143_SLICE_X3Y143_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h2222222222222222)
  ) CLBLM_R_X3Y143_SLICE_X3Y143_DLUT (
.I0(CLBLL_L_X4Y143_SLICE_X4Y143_C5Q),
.I1(CLBLL_L_X4Y144_SLICE_X4Y144_CQ),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y143_SLICE_X3Y143_DO5),
.O6(CLBLM_R_X3Y143_SLICE_X3Y143_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f033ccff00aaaa)
  ) CLBLM_R_X3Y143_SLICE_X3Y143_CLUT (
.I0(CLBLM_R_X3Y151_SLICE_X3Y151_AQ),
.I1(LIOB33_X0Y57_IOB_X0Y58_I),
.I2(CLBLM_R_X5Y146_SLICE_X6Y146_AQ),
.I3(CLBLM_R_X3Y143_SLICE_X3Y143_CQ),
.I4(LIOB33_X0Y61_IOB_X0Y62_I),
.I5(1'b1),
.O5(CLBLM_R_X3Y143_SLICE_X3Y143_CO5),
.O6(CLBLM_R_X3Y143_SLICE_X3Y143_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'he4e4f5f5a0a0a0a0)
  ) CLBLM_R_X3Y143_SLICE_X3Y143_BLUT (
.I0(LIOB33_X0Y61_IOB_X0Y62_I),
.I1(CLBLM_R_X3Y143_SLICE_X3Y143_BQ),
.I2(CLBLM_R_X5Y141_SLICE_X6Y141_BQ),
.I3(1'b1),
.I4(CLBLL_L_X4Y142_SLICE_X4Y142_AQ),
.I5(CLBLL_L_X4Y143_SLICE_X5Y143_B5Q),
.O5(CLBLM_R_X3Y143_SLICE_X3Y143_BO5),
.O6(CLBLM_R_X3Y143_SLICE_X3Y143_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfeaafefe54005454)
  ) CLBLM_R_X3Y143_SLICE_X3Y143_ALUT (
.I0(LIOB33_X0Y61_IOB_X0Y62_I),
.I1(CLBLM_R_X3Y147_SLICE_X3Y147_BQ),
.I2(CLBLM_R_X3Y143_SLICE_X3Y143_AQ),
.I3(CLBLL_L_X4Y151_SLICE_X4Y151_BQ),
.I4(CLBLM_R_X3Y145_SLICE_X3Y145_D5Q),
.I5(CLBLL_L_X4Y143_SLICE_X4Y143_D5Q),
.O5(CLBLM_R_X3Y143_SLICE_X3Y143_AO5),
.O6(CLBLM_R_X3Y143_SLICE_X3Y143_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y144_SLICE_X2Y144_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y144_SLICE_X2Y144_BO5),
.Q(CLBLM_R_X3Y144_SLICE_X2Y144_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0305000003050000)
  ) CLBLM_R_X3Y144_SLICE_X2Y144_DLUT (
.I0(CLBLM_R_X5Y153_SLICE_X6Y153_B5Q),
.I1(CLBLL_L_X2Y146_SLICE_X0Y146_DQ),
.I2(CLBLM_R_X3Y144_SLICE_X3Y144_AQ),
.I3(CLBLL_L_X2Y146_SLICE_X1Y146_B5Q),
.I4(CLBLM_R_X3Y145_SLICE_X3Y145_CQ),
.I5(1'b1),
.O5(CLBLM_R_X3Y144_SLICE_X2Y144_DO5),
.O6(CLBLM_R_X3Y144_SLICE_X2Y144_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff1000ffff9080)
  ) CLBLM_R_X3Y144_SLICE_X2Y144_CLUT (
.I0(CLBLL_L_X2Y146_SLICE_X1Y146_B5Q),
.I1(CLBLM_R_X3Y145_SLICE_X3Y145_CQ),
.I2(CLBLM_R_X3Y144_SLICE_X3Y144_AQ),
.I3(CLBLM_R_X5Y143_SLICE_X6Y143_D5Q),
.I4(CLBLM_R_X3Y144_SLICE_X2Y144_DO6),
.I5(CLBLM_R_X3Y144_SLICE_X2Y144_BO6),
.O5(CLBLM_R_X3Y144_SLICE_X2Y144_CO5),
.O6(CLBLM_R_X3Y144_SLICE_X2Y144_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h88880000f808f000)
  ) CLBLM_R_X3Y144_SLICE_X2Y144_BLUT (
.I0(CLBLM_R_X3Y143_SLICE_X2Y143_A5Q),
.I1(LIOB33_X0Y57_IOB_X0Y58_I),
.I2(LIOB33_X0Y61_IOB_X0Y62_I),
.I3(CLBLM_R_X3Y150_SLICE_X2Y150_AQ),
.I4(CLBLM_R_X3Y143_SLICE_X3Y143_CQ),
.I5(1'b1),
.O5(CLBLM_R_X3Y144_SLICE_X2Y144_BO5),
.O6(CLBLM_R_X3Y144_SLICE_X2Y144_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h20a8000088880000)
  ) CLBLM_R_X3Y144_SLICE_X2Y144_ALUT (
.I0(CLBLM_R_X3Y145_SLICE_X3Y145_CQ),
.I1(CLBLL_L_X2Y146_SLICE_X1Y146_B5Q),
.I2(CLBLM_R_X3Y144_SLICE_X2Y144_AQ),
.I3(CLBLM_R_X3Y144_SLICE_X2Y144_BO6),
.I4(CLBLM_R_X3Y144_SLICE_X3Y144_AQ),
.I5(1'b1),
.O5(CLBLM_R_X3Y144_SLICE_X2Y144_AO5),
.O6(CLBLM_R_X3Y144_SLICE_X2Y144_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y144_SLICE_X3Y144_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y144_SLICE_X3Y144_AO6),
.Q(CLBLM_R_X3Y144_SLICE_X3Y144_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0055000500550004)
  ) CLBLM_R_X3Y144_SLICE_X3Y144_DLUT (
.I0(CLBLL_L_X2Y146_SLICE_X1Y146_B5Q),
.I1(CLBLM_R_X5Y143_SLICE_X6Y143_D5Q),
.I2(CLBLM_R_X3Y144_SLICE_X2Y144_BO6),
.I3(CLBLM_R_X3Y145_SLICE_X3Y145_CQ),
.I4(CLBLM_R_X3Y144_SLICE_X3Y144_AQ),
.I5(CLBLM_R_X3Y142_SLICE_X3Y142_BO6),
.O5(CLBLM_R_X3Y144_SLICE_X3Y144_DO5),
.O6(CLBLM_R_X3Y144_SLICE_X3Y144_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hb333333300000000)
  ) CLBLM_R_X3Y144_SLICE_X3Y144_CLUT (
.I0(CLBLM_R_X3Y143_SLICE_X3Y143_CQ),
.I1(CLBLM_R_X3Y145_SLICE_X3Y145_CQ),
.I2(LIOB33_X0Y57_IOB_X0Y58_I),
.I3(CLBLM_R_X3Y143_SLICE_X2Y143_A5Q),
.I4(CLBLM_R_X3Y144_SLICE_X3Y144_AQ),
.I5(CLBLL_L_X2Y146_SLICE_X1Y146_B5Q),
.O5(CLBLM_R_X3Y144_SLICE_X3Y144_CO5),
.O6(CLBLM_R_X3Y144_SLICE_X3Y144_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffffa2a3a2a2)
  ) CLBLM_R_X3Y144_SLICE_X3Y144_BLUT (
.I0(CLBLM_R_X5Y147_SLICE_X6Y147_B5Q),
.I1(CLBLM_R_X3Y144_SLICE_X2Y144_BO6),
.I2(CLBLM_R_X3Y144_SLICE_X3Y144_AQ),
.I3(CLBLM_R_X3Y142_SLICE_X3Y142_BO6),
.I4(CLBLM_R_X5Y143_SLICE_X6Y143_D5Q),
.I5(CLBLM_R_X3Y145_SLICE_X3Y145_CQ),
.O5(CLBLM_R_X3Y144_SLICE_X3Y144_BO5),
.O6(CLBLM_R_X3Y144_SLICE_X3Y144_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hff00f0f0ff00fbfb)
  ) CLBLM_R_X3Y144_SLICE_X3Y144_ALUT (
.I0(CLBLM_R_X3Y144_SLICE_X3Y144_DO6),
.I1(CLBLL_L_X2Y144_SLICE_X1Y144_AO6),
.I2(CLBLM_R_X3Y144_SLICE_X2Y144_AO6),
.I3(CLBLL_L_X4Y153_SLICE_X4Y153_BQ),
.I4(LIOB33_X0Y61_IOB_X0Y62_I),
.I5(CLBLM_R_X5Y147_SLICE_X6Y147_B5Q),
.O5(CLBLM_R_X3Y144_SLICE_X3Y144_AO5),
.O6(CLBLM_R_X3Y144_SLICE_X3Y144_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y145_SLICE_X2Y145_B5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y145_SLICE_X2Y145_BO5),
.Q(CLBLM_R_X3Y145_SLICE_X2Y145_B5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "C5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y145_SLICE_X2Y145_C5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y145_SLICE_X2Y145_CO5),
.Q(CLBLM_R_X3Y145_SLICE_X2Y145_C5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y145_SLICE_X2Y145_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y145_SLICE_X2Y145_AO6),
.Q(CLBLM_R_X3Y145_SLICE_X2Y145_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y145_SLICE_X2Y145_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y145_SLICE_X2Y145_BO6),
.Q(CLBLM_R_X3Y145_SLICE_X2Y145_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y145_SLICE_X2Y145_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y145_SLICE_X2Y145_CO6),
.Q(CLBLM_R_X3Y145_SLICE_X2Y145_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffffffffffffe)
  ) CLBLM_R_X3Y145_SLICE_X2Y145_DLUT (
.I0(CLBLM_R_X3Y148_SLICE_X2Y148_A5Q),
.I1(CLBLL_L_X4Y145_SLICE_X4Y145_C5Q),
.I2(CLBLM_R_X3Y147_SLICE_X2Y147_DQ),
.I3(CLBLM_L_X10Y153_SLICE_X13Y153_CQ),
.I4(CLBLM_R_X5Y145_SLICE_X6Y145_B5Q),
.I5(CLBLL_L_X4Y145_SLICE_X5Y145_CQ),
.O5(CLBLM_R_X3Y145_SLICE_X2Y145_DO5),
.O6(CLBLM_R_X3Y145_SLICE_X2Y145_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hccf0ccf0ffaa00aa)
  ) CLBLM_R_X3Y145_SLICE_X2Y145_CLUT (
.I0(CLBLM_R_X5Y143_SLICE_X6Y143_C5Q),
.I1(CLBLL_L_X4Y147_SLICE_X5Y147_BQ),
.I2(CLBLL_L_X4Y147_SLICE_X5Y147_C5Q),
.I3(LIOB33_X0Y61_IOB_X0Y62_I),
.I4(CLBLM_R_X7Y144_SLICE_X9Y144_A5Q),
.I5(1'b1),
.O5(CLBLM_R_X3Y145_SLICE_X2Y145_CO5),
.O6(CLBLM_R_X3Y145_SLICE_X2Y145_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0fff000ccaaccaa)
  ) CLBLM_R_X3Y145_SLICE_X2Y145_BLUT (
.I0(CLBLL_L_X4Y146_SLICE_X4Y146_C5Q),
.I1(CLBLM_R_X3Y145_SLICE_X2Y145_BQ),
.I2(CLBLL_L_X4Y145_SLICE_X4Y145_B5Q),
.I3(LIOB33_X0Y61_IOB_X0Y62_I),
.I4(CLBLM_R_X3Y151_SLICE_X3Y151_BQ),
.I5(1'b1),
.O5(CLBLM_R_X3Y145_SLICE_X2Y145_BO5),
.O6(CLBLM_R_X3Y145_SLICE_X2Y145_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffa800a8fffc00fc)
  ) CLBLM_R_X3Y145_SLICE_X2Y145_ALUT (
.I0(CLBLM_L_X10Y145_SLICE_X12Y145_AQ),
.I1(CLBLM_R_X3Y145_SLICE_X2Y145_BQ),
.I2(CLBLM_R_X3Y145_SLICE_X2Y145_AQ),
.I3(LIOB33_X0Y61_IOB_X0Y62_I),
.I4(CLBLM_R_X3Y143_SLICE_X2Y143_AQ),
.I5(CLBLM_R_X5Y142_SLICE_X7Y142_BQ),
.O5(CLBLM_R_X3Y145_SLICE_X2Y145_AO5),
.O6(CLBLM_R_X3Y145_SLICE_X2Y145_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y145_SLICE_X3Y145_C5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y145_SLICE_X3Y145_CO5),
.Q(CLBLM_R_X3Y145_SLICE_X3Y145_C5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y145_SLICE_X3Y145_D5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y145_SLICE_X3Y145_DO5),
.Q(CLBLM_R_X3Y145_SLICE_X3Y145_D5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y145_SLICE_X3Y145_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y145_SLICE_X3Y145_AO6),
.Q(CLBLM_R_X3Y145_SLICE_X3Y145_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y145_SLICE_X3Y145_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y145_SLICE_X3Y145_BO6),
.Q(CLBLM_R_X3Y145_SLICE_X3Y145_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y145_SLICE_X3Y145_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y145_SLICE_X3Y145_CO6),
.Q(CLBLM_R_X3Y145_SLICE_X3Y145_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y145_SLICE_X3Y145_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y145_SLICE_X3Y145_DO6),
.Q(CLBLM_R_X3Y145_SLICE_X3Y145_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hffcc3300ee22ee22)
  ) CLBLM_R_X3Y145_SLICE_X3Y145_DLUT (
.I0(CLBLL_L_X4Y151_SLICE_X4Y151_BQ),
.I1(LIOB33_X0Y61_IOB_X0Y62_I),
.I2(1'b1),
.I3(CLBLM_R_X3Y146_SLICE_X2Y146_BQ),
.I4(CLBLM_R_X7Y146_SLICE_X8Y146_CQ),
.I5(1'b1),
.O5(CLBLM_R_X3Y145_SLICE_X3Y145_DO5),
.O6(CLBLM_R_X3Y145_SLICE_X3Y145_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hccfc0030bbbb8888)
  ) CLBLM_R_X3Y145_SLICE_X3Y145_CLUT (
.I0(CLBLM_R_X3Y143_SLICE_X2Y143_A5Q),
.I1(LIOB33_X0Y61_IOB_X0Y62_I),
.I2(CLBLM_R_X3Y144_SLICE_X3Y144_BO6),
.I3(CLBLM_R_X3Y144_SLICE_X3Y144_CO6),
.I4(CLBLM_L_X10Y151_SLICE_X13Y151_A5Q),
.I5(1'b1),
.O5(CLBLM_R_X3Y145_SLICE_X3Y145_CO5),
.O6(CLBLM_R_X3Y145_SLICE_X3Y145_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf3f3f3f3e2e2d1d1)
  ) CLBLM_R_X3Y145_SLICE_X3Y145_BLUT (
.I0(CLBLL_L_X4Y145_SLICE_X4Y145_DO6),
.I1(LIOB33_X0Y61_IOB_X0Y62_I),
.I2(CLBLM_R_X3Y146_SLICE_X2Y146_C5Q),
.I3(1'b1),
.I4(CLBLM_R_X3Y145_SLICE_X3Y145_BQ),
.I5(CLBLM_R_X3Y145_SLICE_X2Y145_CQ),
.O5(CLBLM_R_X3Y145_SLICE_X3Y145_BO5),
.O6(CLBLM_R_X3Y145_SLICE_X3Y145_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hbbb8bbb88888bbb8)
  ) CLBLM_R_X3Y145_SLICE_X3Y145_ALUT (
.I0(CLBLL_L_X4Y152_SLICE_X4Y152_DQ),
.I1(LIOB33_X0Y61_IOB_X0Y62_I),
.I2(CLBLL_L_X4Y145_SLICE_X4Y145_B5Q),
.I3(CLBLM_R_X3Y145_SLICE_X3Y145_AQ),
.I4(CLBLL_L_X4Y142_SLICE_X5Y142_DQ),
.I5(CLBLL_L_X4Y147_SLICE_X5Y147_CQ),
.O5(CLBLM_R_X3Y145_SLICE_X3Y145_AO5),
.O6(CLBLM_R_X3Y145_SLICE_X3Y145_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y146_SLICE_X2Y146_C5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y146_SLICE_X2Y146_CO5),
.Q(CLBLM_R_X3Y146_SLICE_X2Y146_C5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y146_SLICE_X2Y146_D5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y146_SLICE_X2Y146_DO5),
.Q(CLBLM_R_X3Y146_SLICE_X2Y146_D5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y146_SLICE_X2Y146_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y146_SLICE_X2Y146_AO6),
.Q(CLBLM_R_X3Y146_SLICE_X2Y146_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y146_SLICE_X2Y146_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y146_SLICE_X2Y146_BO6),
.Q(CLBLM_R_X3Y146_SLICE_X2Y146_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y146_SLICE_X2Y146_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y146_SLICE_X2Y146_CO6),
.Q(CLBLM_R_X3Y146_SLICE_X2Y146_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y146_SLICE_X2Y146_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y146_SLICE_X2Y146_DO6),
.Q(CLBLM_R_X3Y146_SLICE_X2Y146_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'haaf0aaf0f0ccf0cc)
  ) CLBLM_R_X3Y146_SLICE_X2Y146_DLUT (
.I0(CLBLL_L_X4Y147_SLICE_X4Y147_AQ),
.I1(CLBLM_R_X11Y148_SLICE_X14Y148_AO6),
.I2(CLBLL_L_X2Y145_SLICE_X1Y145_BQ),
.I3(LIOB33_X0Y61_IOB_X0Y62_I),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y146_SLICE_X2Y146_DO5),
.O6(CLBLM_R_X3Y146_SLICE_X2Y146_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hdd11dd11fcfc3030)
  ) CLBLM_R_X3Y146_SLICE_X2Y146_CLUT (
.I0(CLBLM_R_X5Y150_SLICE_X6Y150_C5Q),
.I1(LIOB33_X0Y61_IOB_X0Y62_I),
.I2(CLBLM_R_X3Y147_SLICE_X2Y147_D5Q),
.I3(CLBLM_R_X7Y142_SLICE_X9Y142_CQ),
.I4(CLBLL_L_X4Y149_SLICE_X5Y149_CQ),
.I5(1'b1),
.O5(CLBLM_R_X3Y146_SLICE_X2Y146_CO5),
.O6(CLBLM_R_X3Y146_SLICE_X2Y146_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaaaaaa03030c0c)
  ) CLBLM_R_X3Y146_SLICE_X2Y146_BLUT (
.I0(CLBLM_R_X5Y149_SLICE_X6Y149_B5Q),
.I1(CLBLM_R_X3Y146_SLICE_X2Y146_BQ),
.I2(CLBLL_L_X4Y143_SLICE_X4Y143_D5Q),
.I3(1'b1),
.I4(CLBLL_L_X2Y146_SLICE_X1Y146_DO6),
.I5(LIOB33_X0Y61_IOB_X0Y62_I),
.O5(CLBLM_R_X3Y146_SLICE_X2Y146_BO5),
.O6(CLBLM_R_X3Y146_SLICE_X2Y146_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffddfcdc33113010)
  ) CLBLM_R_X3Y146_SLICE_X2Y146_ALUT (
.I0(CLBLM_R_X5Y142_SLICE_X7Y142_BQ),
.I1(LIOB33_X0Y61_IOB_X0Y62_I),
.I2(CLBLM_R_X3Y146_SLICE_X2Y146_AQ),
.I3(CLBLM_L_X10Y145_SLICE_X12Y145_AQ),
.I4(CLBLM_R_X3Y143_SLICE_X3Y143_C5Q),
.I5(CLBLM_R_X3Y145_SLICE_X2Y145_C5Q),
.O5(CLBLM_R_X3Y146_SLICE_X2Y146_AO5),
.O6(CLBLM_R_X3Y146_SLICE_X2Y146_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y146_SLICE_X3Y146_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y146_SLICE_X3Y146_AO6),
.Q(CLBLM_R_X3Y146_SLICE_X3Y146_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y146_SLICE_X3Y146_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y146_SLICE_X3Y146_BO6),
.Q(CLBLM_R_X3Y146_SLICE_X3Y146_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h9009900990099009)
  ) CLBLM_R_X3Y146_SLICE_X3Y146_DLUT (
.I0(CLBLL_L_X2Y145_SLICE_X1Y145_BQ),
.I1(CLBLM_R_X3Y148_SLICE_X3Y148_C5Q),
.I2(CLBLL_L_X4Y149_SLICE_X4Y149_AQ),
.I3(CLBLM_R_X5Y150_SLICE_X7Y150_A5Q),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y146_SLICE_X3Y146_DO5),
.O6(CLBLM_R_X3Y146_SLICE_X3Y146_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hffbeffffffbeffff)
  ) CLBLM_R_X3Y146_SLICE_X3Y146_CLUT (
.I0(CLBLL_L_X4Y146_SLICE_X4Y146_DO5),
.I1(CLBLL_L_X2Y145_SLICE_X1Y145_CQ),
.I2(CLBLM_R_X3Y149_SLICE_X3Y149_DQ),
.I3(CLBLM_R_X5Y146_SLICE_X6Y146_CO6),
.I4(CLBLM_R_X3Y146_SLICE_X3Y146_DO6),
.I5(1'b1),
.O5(CLBLM_R_X3Y146_SLICE_X3Y146_CO5),
.O6(CLBLM_R_X3Y146_SLICE_X3Y146_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hacaca0afacacafaf)
  ) CLBLM_R_X3Y146_SLICE_X3Y146_BLUT (
.I0(CLBLM_R_X3Y146_SLICE_X2Y146_DQ),
.I1(CLBLM_R_X3Y146_SLICE_X3Y146_BQ),
.I2(LIOB33_X0Y61_IOB_X0Y62_I),
.I3(CLBLL_L_X4Y152_SLICE_X4Y152_DQ),
.I4(CLBLL_L_X4Y146_SLICE_X5Y146_AQ),
.I5(CLBLM_R_X3Y149_SLICE_X3Y149_CQ),
.O5(CLBLM_R_X3Y146_SLICE_X3Y146_BO5),
.O6(CLBLM_R_X3Y146_SLICE_X3Y146_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff3333cffc0330)
  ) CLBLM_R_X3Y146_SLICE_X3Y146_ALUT (
.I0(1'b1),
.I1(LIOB33_X0Y61_IOB_X0Y62_I),
.I2(CLBLM_R_X7Y146_SLICE_X8Y146_BQ),
.I3(CLBLM_R_X3Y146_SLICE_X2Y146_BQ),
.I4(CLBLM_R_X3Y145_SLICE_X3Y145_AQ),
.I5(CLBLM_R_X3Y146_SLICE_X3Y146_CO6),
.O5(CLBLM_R_X3Y146_SLICE_X3Y146_AO5),
.O6(CLBLM_R_X3Y146_SLICE_X3Y146_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y147_SLICE_X2Y147_D5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y147_SLICE_X2Y147_DO5),
.Q(CLBLM_R_X3Y147_SLICE_X2Y147_D5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y147_SLICE_X2Y147_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y147_SLICE_X2Y147_AO6),
.Q(CLBLM_R_X3Y147_SLICE_X2Y147_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y147_SLICE_X2Y147_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y147_SLICE_X2Y147_BO6),
.Q(CLBLM_R_X3Y147_SLICE_X2Y147_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y147_SLICE_X2Y147_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y147_SLICE_X2Y147_CO6),
.Q(CLBLM_R_X3Y147_SLICE_X2Y147_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y147_SLICE_X2Y147_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y147_SLICE_X2Y147_DO6),
.Q(CLBLM_R_X3Y147_SLICE_X2Y147_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hfc30fc30bbbb8888)
  ) CLBLM_R_X3Y147_SLICE_X2Y147_DLUT (
.I0(CLBLM_R_X7Y152_SLICE_X8Y152_CQ),
.I1(LIOB33_X0Y61_IOB_X0Y62_I),
.I2(CLBLM_L_X10Y153_SLICE_X13Y153_CQ),
.I3(CLBLM_L_X8Y147_SLICE_X10Y147_BQ),
.I4(CLBLL_L_X4Y142_SLICE_X5Y142_D5Q),
.I5(1'b1),
.O5(CLBLM_R_X3Y147_SLICE_X2Y147_DO5),
.O6(CLBLM_R_X3Y147_SLICE_X2Y147_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff0000060c060c)
  ) CLBLM_R_X3Y147_SLICE_X2Y147_CLUT (
.I0(CLBLL_L_X2Y146_SLICE_X1Y146_AQ),
.I1(CLBLM_R_X3Y147_SLICE_X2Y147_CQ),
.I2(CLBLL_L_X4Y143_SLICE_X4Y143_D5Q),
.I3(CLBLL_L_X4Y149_SLICE_X5Y149_CQ),
.I4(CLBLM_R_X3Y149_SLICE_X3Y149_DQ),
.I5(LIOB33_X0Y61_IOB_X0Y62_I),
.O5(CLBLM_R_X3Y147_SLICE_X2Y147_CO5),
.O6(CLBLM_R_X3Y147_SLICE_X2Y147_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaaaaaa3c00cc00)
  ) CLBLM_R_X3Y147_SLICE_X2Y147_BLUT (
.I0(CLBLM_R_X3Y148_SLICE_X2Y148_A5Q),
.I1(CLBLM_R_X3Y147_SLICE_X2Y147_BQ),
.I2(CLBLM_R_X3Y147_SLICE_X2Y147_AQ),
.I3(CLBLL_L_X2Y150_SLICE_X1Y150_AQ),
.I4(CLBLM_R_X3Y152_SLICE_X2Y152_AO6),
.I5(LIOB33_X0Y61_IOB_X0Y62_I),
.O5(CLBLM_R_X3Y147_SLICE_X2Y147_BO5),
.O6(CLBLM_R_X3Y147_SLICE_X2Y147_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hff00ff0028282828)
  ) CLBLM_R_X3Y147_SLICE_X2Y147_ALUT (
.I0(CLBLL_L_X2Y150_SLICE_X1Y150_AQ),
.I1(CLBLM_R_X3Y152_SLICE_X2Y152_AO6),
.I2(CLBLM_R_X3Y147_SLICE_X2Y147_AQ),
.I3(CLBLM_R_X3Y147_SLICE_X2Y147_D5Q),
.I4(1'b1),
.I5(LIOB33_X0Y61_IOB_X0Y62_I),
.O5(CLBLM_R_X3Y147_SLICE_X2Y147_AO5),
.O6(CLBLM_R_X3Y147_SLICE_X2Y147_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y147_SLICE_X3Y147_B5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y147_SLICE_X3Y147_BO5),
.Q(CLBLM_R_X3Y147_SLICE_X3Y147_B5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "C5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y147_SLICE_X3Y147_C5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y147_SLICE_X3Y147_CO5),
.Q(CLBLM_R_X3Y147_SLICE_X3Y147_C5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y147_SLICE_X3Y147_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y147_SLICE_X3Y147_AO6),
.Q(CLBLM_R_X3Y147_SLICE_X3Y147_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y147_SLICE_X3Y147_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y147_SLICE_X3Y147_BO6),
.Q(CLBLM_R_X3Y147_SLICE_X3Y147_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y147_SLICE_X3Y147_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y147_SLICE_X3Y147_CO6),
.Q(CLBLM_R_X3Y147_SLICE_X3Y147_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f00000f3f30000)
  ) CLBLM_R_X3Y147_SLICE_X3Y147_DLUT (
.I0(1'b1),
.I1(CLBLM_R_X5Y146_SLICE_X7Y146_BQ),
.I2(CLBLL_L_X4Y150_SLICE_X4Y150_DO6),
.I3(1'b1),
.I4(CLBLL_L_X2Y150_SLICE_X1Y150_AQ),
.I5(CLBLL_L_X4Y146_SLICE_X5Y146_BQ),
.O5(CLBLM_R_X3Y147_SLICE_X3Y147_DO5),
.O6(CLBLM_R_X3Y147_SLICE_X3Y147_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hccccaaaaaaaaff00)
  ) CLBLM_R_X3Y147_SLICE_X3Y147_CLUT (
.I0(CLBLL_L_X4Y147_SLICE_X5Y147_C5Q),
.I1(CLBLM_R_X5Y147_SLICE_X6Y147_CQ),
.I2(1'b1),
.I3(CLBLM_R_X7Y146_SLICE_X8Y146_DQ),
.I4(LIOB33_X0Y61_IOB_X0Y62_I),
.I5(1'b1),
.O5(CLBLM_R_X3Y147_SLICE_X3Y147_CO5),
.O6(CLBLM_R_X3Y147_SLICE_X3Y147_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hffaa5500d8d8d8d8)
  ) CLBLM_R_X3Y147_SLICE_X3Y147_BLUT (
.I0(LIOB33_X0Y61_IOB_X0Y62_I),
.I1(CLBLM_R_X3Y147_SLICE_X3Y147_BQ),
.I2(RIOB33_X105Y119_IOB_X1Y119_I),
.I3(CLBLM_R_X3Y145_SLICE_X3Y145_BQ),
.I4(CLBLM_R_X5Y151_SLICE_X6Y151_C5Q),
.I5(1'b1),
.O5(CLBLM_R_X3Y147_SLICE_X3Y147_BO5),
.O6(CLBLM_R_X3Y147_SLICE_X3Y147_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0eef022f0eef022)
  ) CLBLM_R_X3Y147_SLICE_X3Y147_ALUT (
.I0(CLBLM_R_X3Y147_SLICE_X3Y147_AQ),
.I1(CLBLM_R_X11Y148_SLICE_X15Y148_AO6),
.I2(CLBLM_R_X3Y143_SLICE_X3Y143_C5Q),
.I3(LIOB33_X0Y61_IOB_X0Y62_I),
.I4(CLBLM_R_X3Y145_SLICE_X3Y145_AQ),
.I5(1'b1),
.O5(CLBLM_R_X3Y147_SLICE_X3Y147_AO5),
.O6(CLBLM_R_X3Y147_SLICE_X3Y147_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y148_SLICE_X2Y148_A5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y148_SLICE_X2Y148_AO5),
.Q(CLBLM_R_X3Y148_SLICE_X2Y148_A5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y148_SLICE_X2Y148_B5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y148_SLICE_X2Y148_BO5),
.Q(CLBLM_R_X3Y148_SLICE_X2Y148_B5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y148_SLICE_X2Y148_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y148_SLICE_X2Y148_AO6),
.Q(CLBLM_R_X3Y148_SLICE_X2Y148_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y148_SLICE_X2Y148_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y148_SLICE_X2Y148_BO6),
.Q(CLBLM_R_X3Y148_SLICE_X2Y148_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffffffefefefe)
  ) CLBLM_R_X3Y148_SLICE_X2Y148_DLUT (
.I0(CLBLM_R_X5Y147_SLICE_X6Y147_CQ),
.I1(CLBLL_L_X4Y146_SLICE_X4Y146_B5Q),
.I2(CLBLM_R_X3Y150_SLICE_X3Y150_B5Q),
.I3(1'b1),
.I4(1'b1),
.I5(CLBLM_R_X3Y148_SLICE_X2Y148_AQ),
.O5(CLBLM_R_X3Y148_SLICE_X2Y148_DO5),
.O6(CLBLM_R_X3Y148_SLICE_X2Y148_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0fffffffa0000000)
  ) CLBLM_R_X3Y148_SLICE_X2Y148_CLUT (
.I0(CLBLM_R_X3Y149_SLICE_X2Y149_DQ),
.I1(1'b1),
.I2(CLBLL_L_X2Y146_SLICE_X1Y146_BQ),
.I3(CLBLL_L_X4Y149_SLICE_X4Y149_D5Q),
.I4(CLBLL_L_X4Y149_SLICE_X4Y149_DQ),
.I5(1'b1),
.O5(CLBLM_R_X3Y148_SLICE_X2Y148_CO5),
.O6(CLBLM_R_X3Y148_SLICE_X2Y148_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hc5c5cacafc0cfc0c)
  ) CLBLM_R_X3Y148_SLICE_X2Y148_BLUT (
.I0(CLBLM_R_X3Y148_SLICE_X2Y148_BQ),
.I1(CLBLM_R_X3Y148_SLICE_X3Y148_B5Q),
.I2(LIOB33_X0Y61_IOB_X0Y62_I),
.I3(CLBLM_L_X10Y154_SLICE_X12Y154_B5Q),
.I4(CLBLM_R_X3Y148_SLICE_X2Y148_CO5),
.I5(1'b1),
.O5(CLBLM_R_X3Y148_SLICE_X2Y148_BO5),
.O6(CLBLM_R_X3Y148_SLICE_X2Y148_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'ha3aca3acfafa0a0a)
  ) CLBLM_R_X3Y148_SLICE_X2Y148_ALUT (
.I0(CLBLM_R_X3Y147_SLICE_X2Y147_DQ),
.I1(CLBLM_R_X7Y148_SLICE_X9Y148_AQ),
.I2(LIOB33_X0Y61_IOB_X0Y62_I),
.I3(CLBLM_R_X3Y151_SLICE_X3Y151_CQ),
.I4(CLBLM_R_X3Y145_SLICE_X2Y145_AQ),
.I5(1'b1),
.O5(CLBLM_R_X3Y148_SLICE_X2Y148_AO5),
.O6(CLBLM_R_X3Y148_SLICE_X2Y148_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y148_SLICE_X3Y148_B5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y148_SLICE_X3Y148_BO5),
.Q(CLBLM_R_X3Y148_SLICE_X3Y148_B5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "C5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y148_SLICE_X3Y148_C5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y148_SLICE_X3Y148_CO5),
.Q(CLBLM_R_X3Y148_SLICE_X3Y148_C5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y148_SLICE_X3Y148_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y148_SLICE_X3Y148_AO6),
.Q(CLBLM_R_X3Y148_SLICE_X3Y148_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y148_SLICE_X3Y148_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y148_SLICE_X3Y148_BO6),
.Q(CLBLM_R_X3Y148_SLICE_X3Y148_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y148_SLICE_X3Y148_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y148_SLICE_X3Y148_CO6),
.Q(CLBLM_R_X3Y148_SLICE_X3Y148_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0f000f003333ffff)
  ) CLBLM_R_X3Y148_SLICE_X3Y148_DLUT (
.I0(1'b1),
.I1(CLBLM_R_X3Y149_SLICE_X3Y149_CQ),
.I2(CLBLL_L_X4Y148_SLICE_X4Y148_C5Q),
.I3(CLBLM_R_X3Y149_SLICE_X2Y149_CQ),
.I4(CLBLL_L_X4Y152_SLICE_X4Y152_DQ),
.I5(1'b1),
.O5(CLBLM_R_X3Y148_SLICE_X3Y148_DO5),
.O6(CLBLM_R_X3Y148_SLICE_X3Y148_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hccffcc00aaf0aaf0)
  ) CLBLM_R_X3Y148_SLICE_X3Y148_CLUT (
.I0(CLBLL_L_X4Y153_SLICE_X4Y153_AQ),
.I1(CLBLM_L_X12Y146_SLICE_X17Y146_AQ),
.I2(CLBLM_L_X10Y151_SLICE_X13Y151_A5Q),
.I3(LIOB33_X0Y61_IOB_X0Y62_I),
.I4(RIOB33_X105Y101_IOB_X1Y101_I),
.I5(1'b1),
.O5(CLBLM_R_X3Y148_SLICE_X3Y148_CO5),
.O6(CLBLM_R_X3Y148_SLICE_X3Y148_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfc30fc30eeee2222)
  ) CLBLM_R_X3Y148_SLICE_X3Y148_BLUT (
.I0(CLBLL_L_X4Y148_SLICE_X5Y148_A5Q),
.I1(LIOB33_X0Y61_IOB_X0Y62_I),
.I2(CLBLL_L_X4Y146_SLICE_X4Y146_C5Q),
.I3(CLBLM_R_X5Y145_SLICE_X6Y145_C5Q),
.I4(CLBLM_R_X7Y148_SLICE_X9Y148_AQ),
.I5(1'b1),
.O5(CLBLM_R_X3Y148_SLICE_X3Y148_BO5),
.O6(CLBLM_R_X3Y148_SLICE_X3Y148_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffddffd000dd00d0)
  ) CLBLM_R_X3Y148_SLICE_X3Y148_ALUT (
.I0(CLBLM_R_X5Y142_SLICE_X7Y142_BQ),
.I1(CLBLM_L_X10Y145_SLICE_X12Y145_AQ),
.I2(CLBLM_R_X3Y148_SLICE_X3Y148_AQ),
.I3(LIOB33_X0Y61_IOB_X0Y62_I),
.I4(CLBLM_R_X3Y150_SLICE_X3Y150_A5Q),
.I5(CLBLM_R_X3Y149_SLICE_X2Y149_CQ),
.O5(CLBLM_R_X3Y148_SLICE_X3Y148_AO5),
.O6(CLBLM_R_X3Y148_SLICE_X3Y148_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y149_SLICE_X2Y149_C5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y149_SLICE_X2Y149_CO5),
.Q(CLBLM_R_X3Y149_SLICE_X2Y149_C5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y149_SLICE_X2Y149_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y149_SLICE_X2Y149_AO6),
.Q(CLBLM_R_X3Y149_SLICE_X2Y149_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y149_SLICE_X2Y149_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y149_SLICE_X2Y149_BO6),
.Q(CLBLM_R_X3Y149_SLICE_X2Y149_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y149_SLICE_X2Y149_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y149_SLICE_X2Y149_CO6),
.Q(CLBLM_R_X3Y149_SLICE_X2Y149_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y149_SLICE_X2Y149_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y149_SLICE_X2Y149_DO6),
.Q(CLBLM_R_X3Y149_SLICE_X2Y149_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff0000f08ff08f)
  ) CLBLM_R_X3Y149_SLICE_X2Y149_DLUT (
.I0(CLBLM_R_X3Y148_SLICE_X2Y148_BQ),
.I1(LIOB33_X0Y55_IOB_X0Y55_I),
.I2(CLBLM_R_X3Y149_SLICE_X2Y149_DQ),
.I3(CLBLM_R_X3Y148_SLICE_X2Y148_CO6),
.I4(CLBLM_R_X3Y150_SLICE_X3Y150_DQ),
.I5(LIOB33_X0Y61_IOB_X0Y62_I),
.O5(CLBLM_R_X3Y149_SLICE_X2Y149_DO5),
.O6(CLBLM_R_X3Y149_SLICE_X2Y149_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'haaffaa00f0ccf0cc)
  ) CLBLM_R_X3Y149_SLICE_X2Y149_CLUT (
.I0(CLBLM_R_X3Y148_SLICE_X2Y148_BQ),
.I1(CLBLM_R_X3Y150_SLICE_X2Y150_DQ),
.I2(CLBLM_R_X3Y148_SLICE_X3Y148_AQ),
.I3(LIOB33_X0Y61_IOB_X0Y62_I),
.I4(RIOB33_X105Y121_IOB_X1Y121_I),
.I5(1'b1),
.O5(CLBLM_R_X3Y149_SLICE_X2Y149_CO5),
.O6(CLBLM_R_X3Y149_SLICE_X2Y149_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hff06ff0c0006000c)
  ) CLBLM_R_X3Y149_SLICE_X2Y149_BLUT (
.I0(CLBLL_L_X4Y149_SLICE_X4Y149_AQ),
.I1(CLBLM_R_X3Y149_SLICE_X2Y149_BQ),
.I2(CLBLL_L_X4Y143_SLICE_X4Y143_D5Q),
.I3(LIOB33_X0Y61_IOB_X0Y62_I),
.I4(CLBLL_L_X4Y146_SLICE_X4Y146_DO6),
.I5(CLBLM_R_X3Y150_SLICE_X2Y150_DQ),
.O5(CLBLM_R_X3Y149_SLICE_X2Y149_BO5),
.O6(CLBLM_R_X3Y149_SLICE_X2Y149_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hcc0acca0cc0acca0)
  ) CLBLM_R_X3Y149_SLICE_X2Y149_ALUT (
.I0(CLBLL_L_X2Y150_SLICE_X1Y150_AQ),
.I1(CLBLM_R_X3Y149_SLICE_X2Y149_DQ),
.I2(CLBLM_R_X3Y149_SLICE_X2Y149_AQ),
.I3(LIOB33_X0Y61_IOB_X0Y62_I),
.I4(CLBLM_R_X7Y153_SLICE_X9Y153_AQ),
.I5(1'b1),
.O5(CLBLM_R_X3Y149_SLICE_X2Y149_AO5),
.O6(CLBLM_R_X3Y149_SLICE_X2Y149_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y149_SLICE_X3Y149_D5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y149_SLICE_X3Y149_DO5),
.Q(CLBLM_R_X3Y149_SLICE_X3Y149_D5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y149_SLICE_X3Y149_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y149_SLICE_X3Y149_AO6),
.Q(CLBLM_R_X3Y149_SLICE_X3Y149_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y149_SLICE_X3Y149_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y149_SLICE_X3Y149_BO6),
.Q(CLBLM_R_X3Y149_SLICE_X3Y149_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y149_SLICE_X3Y149_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y149_SLICE_X3Y149_CO6),
.Q(CLBLM_R_X3Y149_SLICE_X3Y149_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y149_SLICE_X3Y149_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y149_SLICE_X3Y149_DO6),
.Q(CLBLM_R_X3Y149_SLICE_X3Y149_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'heeee2222d1d1d1d1)
  ) CLBLM_R_X3Y149_SLICE_X3Y149_DLUT (
.I0(CLBLM_R_X3Y146_SLICE_X2Y146_D5Q),
.I1(LIOB33_X0Y61_IOB_X0Y62_I),
.I2(CLBLM_R_X3Y150_SLICE_X3Y150_A5Q),
.I3(1'b1),
.I4(CLBLM_R_X3Y150_SLICE_X2Y150_CQ),
.I5(1'b1),
.O5(CLBLM_R_X3Y149_SLICE_X3Y149_DO5),
.O6(CLBLM_R_X3Y149_SLICE_X3Y149_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff000000070007)
  ) CLBLM_R_X3Y149_SLICE_X3Y149_CLUT (
.I0(CLBLM_R_X3Y149_SLICE_X3Y149_BQ),
.I1(CLBLM_R_X3Y149_SLICE_X3Y149_CQ),
.I2(CLBLM_R_X7Y146_SLICE_X8Y146_CQ),
.I3(CLBLM_R_X3Y147_SLICE_X3Y147_CQ),
.I4(CLBLM_R_X5Y153_SLICE_X6Y153_A5Q),
.I5(LIOB33_X0Y61_IOB_X0Y62_I),
.O5(CLBLM_R_X3Y149_SLICE_X3Y149_CO5),
.O6(CLBLM_R_X3Y149_SLICE_X3Y149_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf3f3f3f3f3e2f3e2)
  ) CLBLM_R_X3Y149_SLICE_X3Y149_BLUT (
.I0(CLBLM_R_X3Y149_SLICE_X3Y149_CQ),
.I1(LIOB33_X0Y61_IOB_X0Y62_I),
.I2(CLBLL_L_X4Y142_SLICE_X5Y142_C5Q),
.I3(CLBLM_R_X7Y146_SLICE_X8Y146_CQ),
.I4(1'b1),
.I5(CLBLM_R_X3Y147_SLICE_X3Y147_CQ),
.O5(CLBLM_R_X3Y149_SLICE_X3Y149_BO5),
.O6(CLBLM_R_X3Y149_SLICE_X3Y149_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hcccccccc0aa0a0a0)
  ) CLBLM_R_X3Y149_SLICE_X3Y149_ALUT (
.I0(CLBLL_L_X2Y150_SLICE_X1Y150_AQ),
.I1(CLBLM_R_X3Y149_SLICE_X3Y149_BQ),
.I2(CLBLM_R_X3Y149_SLICE_X3Y149_AQ),
.I3(CLBLM_R_X7Y153_SLICE_X9Y153_AQ),
.I4(CLBLM_R_X3Y149_SLICE_X2Y149_AQ),
.I5(LIOB33_X0Y61_IOB_X0Y62_I),
.O5(CLBLM_R_X3Y149_SLICE_X3Y149_AO5),
.O6(CLBLM_R_X3Y149_SLICE_X3Y149_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y150_SLICE_X2Y150_D5_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_R_X3Y150_SLICE_X2Y150_DO5),
.Q(CLBLM_R_X3Y150_SLICE_X2Y150_D5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y150_SLICE_X2Y150_A_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_R_X3Y150_SLICE_X2Y150_AO6),
.Q(CLBLM_R_X3Y150_SLICE_X2Y150_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y150_SLICE_X2Y150_B_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_R_X3Y150_SLICE_X2Y150_BO6),
.Q(CLBLM_R_X3Y150_SLICE_X2Y150_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y150_SLICE_X2Y150_C_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_R_X3Y150_SLICE_X2Y150_CO6),
.Q(CLBLM_R_X3Y150_SLICE_X2Y150_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y150_SLICE_X2Y150_D_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_R_X3Y150_SLICE_X2Y150_DO6),
.Q(CLBLM_R_X3Y150_SLICE_X2Y150_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hf033f033aa33aa33)
  ) CLBLM_R_X3Y150_SLICE_X2Y150_DLUT (
.I0(CLBLM_R_X3Y152_SLICE_X3Y152_AQ),
.I1(CLBLM_L_X10Y151_SLICE_X13Y151_AQ),
.I2(CLBLM_R_X3Y150_SLICE_X3Y150_B5Q),
.I3(LIOB33_X0Y61_IOB_X0Y62_I),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y150_SLICE_X2Y150_DO5),
.O6(CLBLM_R_X3Y150_SLICE_X2Y150_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hcccccccc0000550a)
  ) CLBLM_R_X3Y150_SLICE_X2Y150_CLUT (
.I0(CLBLM_R_X3Y150_SLICE_X2Y150_CQ),
.I1(CLBLL_L_X4Y144_SLICE_X5Y144_CQ),
.I2(CLBLM_R_X3Y150_SLICE_X2Y150_BQ),
.I3(CLBLM_R_X3Y150_SLICE_X3Y150_CQ),
.I4(CLBLM_R_X5Y153_SLICE_X6Y153_D5Q),
.I5(LIOB33_X0Y61_IOB_X0Y62_I),
.O5(CLBLM_R_X3Y150_SLICE_X2Y150_CO5),
.O6(CLBLM_R_X3Y150_SLICE_X2Y150_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hc0d1c0d1d1c0c0c0)
  ) CLBLM_R_X3Y150_SLICE_X2Y150_BLUT (
.I0(CLBLM_R_X5Y153_SLICE_X6Y153_D5Q),
.I1(LIOB33_X0Y61_IOB_X0Y62_I),
.I2(CLBLM_R_X3Y148_SLICE_X2Y148_AQ),
.I3(CLBLM_R_X3Y150_SLICE_X2Y150_CQ),
.I4(CLBLM_R_X3Y150_SLICE_X3Y150_CQ),
.I5(CLBLM_R_X3Y150_SLICE_X2Y150_BQ),
.O5(CLBLM_R_X3Y150_SLICE_X2Y150_BO5),
.O6(CLBLM_R_X3Y150_SLICE_X2Y150_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hccccfff0cccc5550)
  ) CLBLM_R_X3Y150_SLICE_X2Y150_ALUT (
.I0(CLBLM_R_X5Y142_SLICE_X7Y142_BQ),
.I1(CLBLL_L_X4Y152_SLICE_X5Y152_AQ),
.I2(CLBLM_R_X3Y150_SLICE_X2Y150_AQ),
.I3(CLBLM_R_X3Y150_SLICE_X3Y150_BQ),
.I4(LIOB33_X0Y61_IOB_X0Y62_I),
.I5(CLBLM_L_X10Y145_SLICE_X12Y145_AQ),
.O5(CLBLM_R_X3Y150_SLICE_X2Y150_AO5),
.O6(CLBLM_R_X3Y150_SLICE_X2Y150_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y150_SLICE_X3Y150_A5_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_R_X3Y150_SLICE_X3Y150_AO5),
.Q(CLBLM_R_X3Y150_SLICE_X3Y150_A5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y150_SLICE_X3Y150_B5_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_R_X3Y150_SLICE_X3Y150_BO5),
.Q(CLBLM_R_X3Y150_SLICE_X3Y150_B5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y150_SLICE_X3Y150_D5_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_R_X3Y150_SLICE_X3Y150_DO5),
.Q(CLBLM_R_X3Y150_SLICE_X3Y150_D5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y150_SLICE_X3Y150_A_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_R_X3Y150_SLICE_X3Y150_AO6),
.Q(CLBLM_R_X3Y150_SLICE_X3Y150_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y150_SLICE_X3Y150_B_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_R_X3Y150_SLICE_X3Y150_BO6),
.Q(CLBLM_R_X3Y150_SLICE_X3Y150_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y150_SLICE_X3Y150_C_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_R_X3Y150_SLICE_X3Y150_CO6),
.Q(CLBLM_R_X3Y150_SLICE_X3Y150_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y150_SLICE_X3Y150_D_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_R_X3Y150_SLICE_X3Y150_DO6),
.Q(CLBLM_R_X3Y150_SLICE_X3Y150_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'haffa0550dddd8888)
  ) CLBLM_R_X3Y150_SLICE_X3Y150_DLUT (
.I0(LIOB33_X0Y61_IOB_X0Y62_I),
.I1(CLBLL_L_X4Y152_SLICE_X4Y152_AQ),
.I2(CLBLM_R_X3Y150_SLICE_X2Y150_D5Q),
.I3(CLBLM_R_X3Y151_SLICE_X3Y151_BQ),
.I4(CLBLM_R_X3Y150_SLICE_X3Y150_AQ),
.I5(1'b1),
.O5(CLBLM_R_X3Y150_SLICE_X3Y150_DO5),
.O6(CLBLM_R_X3Y150_SLICE_X3Y150_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffbfbfb55515151)
  ) CLBLM_R_X3Y150_SLICE_X3Y150_CLUT (
.I0(LIOB33_X0Y61_IOB_X0Y62_I),
.I1(CLBLM_R_X3Y150_SLICE_X3Y150_CQ),
.I2(CLBLM_R_X5Y153_SLICE_X6Y153_D5Q),
.I3(CLBLM_R_X3Y150_SLICE_X2Y150_CQ),
.I4(CLBLM_R_X3Y150_SLICE_X2Y150_BQ),
.I5(CLBLL_L_X4Y150_SLICE_X4Y150_CQ),
.O5(CLBLM_R_X3Y150_SLICE_X3Y150_CO5),
.O6(CLBLM_R_X3Y150_SLICE_X3Y150_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0aaf0aaff660066)
  ) CLBLM_R_X3Y150_SLICE_X3Y150_BLUT (
.I0(CLBLL_L_X4Y151_SLICE_X5Y151_CQ),
.I1(CLBLM_R_X3Y149_SLICE_X3Y149_D5Q),
.I2(CLBLM_R_X3Y150_SLICE_X3Y150_CQ),
.I3(LIOB33_X0Y61_IOB_X0Y62_I),
.I4(CLBLM_R_X7Y151_SLICE_X9Y151_AQ),
.I5(1'b1),
.O5(CLBLM_R_X3Y150_SLICE_X3Y150_BO5),
.O6(CLBLM_R_X3Y150_SLICE_X3Y150_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hff0f000faaffaa00)
  ) CLBLM_R_X3Y150_SLICE_X3Y150_ALUT (
.I0(CLBLM_R_X3Y143_SLICE_X3Y143_BQ),
.I1(1'b1),
.I2(CLBLM_L_X10Y149_SLICE_X12Y149_BQ),
.I3(LIOB33_X0Y61_IOB_X0Y62_I),
.I4(CLBLL_L_X4Y151_SLICE_X4Y151_AQ),
.I5(1'b1),
.O5(CLBLM_R_X3Y150_SLICE_X3Y150_AO5),
.O6(CLBLM_R_X3Y150_SLICE_X3Y150_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y151_SLICE_X2Y151_A_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(LIOB33_X0Y61_IOB_X0Y62_I),
.D(CLBLL_L_X4Y151_SLICE_X4Y151_DQ),
.Q(CLBLM_R_X3Y151_SLICE_X2Y151_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y151_SLICE_X2Y151_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y151_SLICE_X2Y151_DO5),
.O6(CLBLM_R_X3Y151_SLICE_X2Y151_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hdf200000ff000000)
  ) CLBLM_R_X3Y151_SLICE_X2Y151_CLUT (
.I0(CLBLM_R_X3Y151_SLICE_X3Y151_AQ),
.I1(CLBLL_L_X4Y147_SLICE_X5Y147_DO6),
.I2(CLBLM_R_X3Y151_SLICE_X3Y151_CQ),
.I3(CLBLL_L_X4Y150_SLICE_X4Y150_B5Q),
.I4(CLBLL_L_X4Y147_SLICE_X4Y147_AQ),
.I5(CLBLM_R_X3Y151_SLICE_X3Y151_BQ),
.O5(CLBLM_R_X3Y151_SLICE_X2Y151_CO5),
.O6(CLBLM_R_X3Y151_SLICE_X2Y151_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hbbae110433cc33cc)
  ) CLBLM_R_X3Y151_SLICE_X2Y151_BLUT (
.I0(LIOB33_X0Y61_IOB_X0Y62_I),
.I1(CLBLL_L_X4Y142_SLICE_X4Y142_AQ),
.I2(CLBLL_L_X4Y151_SLICE_X4Y151_DQ),
.I3(CLBLM_R_X3Y143_SLICE_X3Y143_BQ),
.I4(CLBLM_R_X3Y149_SLICE_X2Y149_C5Q),
.I5(1'b1),
.O5(CLBLM_R_X3Y151_SLICE_X2Y151_BO5),
.O6(CLBLM_R_X3Y151_SLICE_X2Y151_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hcfc5cfc5ff55ff55)
  ) CLBLM_R_X3Y151_SLICE_X2Y151_ALUT (
.I0(CLBLM_R_X3Y151_SLICE_X3Y151_A5Q),
.I1(CLBLL_L_X4Y144_SLICE_X4Y144_B5Q),
.I2(LIOB33_X0Y61_IOB_X0Y62_I),
.I3(CLBLM_R_X5Y148_SLICE_X6Y148_BQ),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y151_SLICE_X2Y151_AO5),
.O6(CLBLM_R_X3Y151_SLICE_X2Y151_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y151_SLICE_X3Y151_A5_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_R_X3Y151_SLICE_X2Y151_BO6),
.Q(CLBLM_R_X3Y151_SLICE_X3Y151_A5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y151_SLICE_X3Y151_A_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_R_X3Y151_SLICE_X3Y151_AO6),
.Q(CLBLM_R_X3Y151_SLICE_X3Y151_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y151_SLICE_X3Y151_B_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_R_X3Y151_SLICE_X3Y151_BO6),
.Q(CLBLM_R_X3Y151_SLICE_X3Y151_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y151_SLICE_X3Y151_C_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_R_X3Y151_SLICE_X3Y151_CO6),
.Q(CLBLM_R_X3Y151_SLICE_X3Y151_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'heeee444400c000c0)
  ) CLBLM_R_X3Y151_SLICE_X3Y151_DLUT (
.I0(LIOB33_X0Y61_IOB_X0Y62_I),
.I1(CLBLM_R_X3Y151_SLICE_X3Y151_CQ),
.I2(CLBLM_R_X3Y151_SLICE_X3Y151_AQ),
.I3(CLBLL_L_X4Y147_SLICE_X5Y147_DO6),
.I4(CLBLM_L_X10Y150_SLICE_X12Y150_AQ),
.I5(1'b1),
.O5(CLBLM_R_X3Y151_SLICE_X3Y151_DO5),
.O6(CLBLM_R_X3Y151_SLICE_X3Y151_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hff55ff55eb41eb41)
  ) CLBLM_R_X3Y151_SLICE_X3Y151_CLUT (
.I0(LIOB33_X0Y61_IOB_X0Y62_I),
.I1(CLBLM_R_X3Y151_SLICE_X3Y151_CQ),
.I2(CLBLL_L_X4Y147_SLICE_X5Y147_DO6),
.I3(CLBLL_L_X4Y152_SLICE_X4Y152_CQ),
.I4(1'b1),
.I5(CLBLM_R_X3Y145_SLICE_X2Y145_CQ),
.O5(CLBLM_R_X3Y151_SLICE_X3Y151_CO5),
.O6(CLBLM_R_X3Y151_SLICE_X3Y151_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f01144f0f00000)
  ) CLBLM_R_X3Y151_SLICE_X3Y151_BLUT (
.I0(CLBLM_R_X3Y145_SLICE_X2Y145_CQ),
.I1(CLBLM_R_X3Y151_SLICE_X3Y151_BQ),
.I2(CLBLM_R_X5Y146_SLICE_X6Y146_BQ),
.I3(CLBLM_R_X3Y151_SLICE_X3Y151_DO5),
.I4(LIOB33_X0Y61_IOB_X0Y62_I),
.I5(CLBLL_L_X4Y147_SLICE_X4Y147_AQ),
.O5(CLBLM_R_X3Y151_SLICE_X3Y151_BO5),
.O6(CLBLM_R_X3Y151_SLICE_X3Y151_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffcffde00fc00de)
  ) CLBLM_R_X3Y151_SLICE_X3Y151_ALUT (
.I0(CLBLM_R_X3Y151_SLICE_X3Y151_CQ),
.I1(CLBLM_R_X3Y145_SLICE_X2Y145_CQ),
.I2(CLBLM_R_X3Y151_SLICE_X3Y151_AQ),
.I3(LIOB33_X0Y61_IOB_X0Y62_I),
.I4(CLBLL_L_X4Y147_SLICE_X5Y147_DO6),
.I5(CLBLM_L_X8Y154_SLICE_X10Y154_AQ),
.O5(CLBLM_R_X3Y151_SLICE_X3Y151_AO5),
.O6(CLBLM_R_X3Y151_SLICE_X3Y151_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y152_SLICE_X2Y152_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y152_SLICE_X2Y152_DO5),
.O6(CLBLM_R_X3Y152_SLICE_X2Y152_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y152_SLICE_X2Y152_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y152_SLICE_X2Y152_CO5),
.O6(CLBLM_R_X3Y152_SLICE_X2Y152_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y152_SLICE_X2Y152_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y152_SLICE_X2Y152_BO5),
.O6(CLBLM_R_X3Y152_SLICE_X2Y152_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'haa00000000000000)
  ) CLBLM_R_X3Y152_SLICE_X2Y152_ALUT (
.I0(CLBLL_L_X4Y152_SLICE_X5Y152_AQ),
.I1(1'b1),
.I2(1'b1),
.I3(CLBLL_L_X4Y152_SLICE_X5Y152_DO6),
.I4(CLBLM_R_X3Y152_SLICE_X3Y152_AQ),
.I5(CLBLL_L_X4Y152_SLICE_X5Y152_A5Q),
.O5(CLBLM_R_X3Y152_SLICE_X2Y152_AO5),
.O6(CLBLM_R_X3Y152_SLICE_X2Y152_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y152_SLICE_X3Y152_A_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_R_X3Y152_SLICE_X3Y152_AO6),
.Q(CLBLM_R_X3Y152_SLICE_X3Y152_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y152_SLICE_X3Y152_B_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_R_X3Y152_SLICE_X3Y152_BO6),
.Q(CLBLM_R_X3Y152_SLICE_X3Y152_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y152_SLICE_X3Y152_C_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_R_X3Y152_SLICE_X3Y152_CO6),
.Q(CLBLM_R_X3Y152_SLICE_X3Y152_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h8888888888888888)
  ) CLBLM_R_X3Y152_SLICE_X3Y152_DLUT (
.I0(CLBLM_R_X3Y150_SLICE_X2Y150_BQ),
.I1(CLBLM_R_X3Y150_SLICE_X2Y150_CQ),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y152_SLICE_X3Y152_DO5),
.O6(CLBLM_R_X3Y152_SLICE_X3Y152_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hfbfe5154fefe5454)
  ) CLBLM_R_X3Y152_SLICE_X3Y152_CLUT (
.I0(LIOB33_X0Y61_IOB_X0Y62_I),
.I1(CLBLM_R_X3Y152_SLICE_X3Y152_CQ),
.I2(CLBLM_R_X5Y153_SLICE_X6Y153_D5Q),
.I3(CLBLM_R_X3Y150_SLICE_X2Y150_CQ),
.I4(CLBLM_R_X5Y152_SLICE_X7Y152_CQ),
.I5(CLBLM_R_X3Y150_SLICE_X2Y150_BQ),
.O5(CLBLM_R_X3Y152_SLICE_X3Y152_CO5),
.O6(CLBLM_R_X3Y152_SLICE_X3Y152_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffc60000ffc6)
  ) CLBLM_R_X3Y152_SLICE_X3Y152_BLUT (
.I0(CLBLM_R_X3Y152_SLICE_X3Y152_DO6),
.I1(CLBLM_R_X3Y152_SLICE_X3Y152_BQ),
.I2(CLBLM_R_X3Y152_SLICE_X3Y152_CQ),
.I3(CLBLM_R_X5Y153_SLICE_X6Y153_D5Q),
.I4(LIOB33_X0Y61_IOB_X0Y62_I),
.I5(CLBLL_L_X4Y150_SLICE_X4Y150_AQ),
.O5(CLBLM_R_X3Y152_SLICE_X3Y152_BO5),
.O6(CLBLM_R_X3Y152_SLICE_X3Y152_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hbe14aa00fa50aa00)
  ) CLBLM_R_X3Y152_SLICE_X3Y152_ALUT (
.I0(LIOB33_X0Y61_IOB_X0Y62_I),
.I1(CLBLL_L_X4Y152_SLICE_X5Y152_A5Q),
.I2(CLBLM_R_X3Y152_SLICE_X3Y152_AQ),
.I3(CLBLL_L_X4Y151_SLICE_X5Y151_AQ),
.I4(CLBLL_L_X2Y150_SLICE_X1Y150_AQ),
.I5(CLBLL_L_X4Y152_SLICE_X5Y152_DO6),
.O5(CLBLM_R_X3Y152_SLICE_X3Y152_AO5),
.O6(CLBLM_R_X3Y152_SLICE_X3Y152_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y153_SLICE_X2Y153_A_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_R_X3Y151_SLICE_X2Y151_AO6),
.Q(CLBLM_R_X3Y153_SLICE_X2Y153_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y153_SLICE_X2Y153_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y153_SLICE_X2Y153_DO5),
.O6(CLBLM_R_X3Y153_SLICE_X2Y153_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y153_SLICE_X2Y153_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y153_SLICE_X2Y153_CO5),
.O6(CLBLM_R_X3Y153_SLICE_X2Y153_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y153_SLICE_X2Y153_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y153_SLICE_X2Y153_BO5),
.O6(CLBLM_R_X3Y153_SLICE_X2Y153_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y153_SLICE_X2Y153_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y153_SLICE_X2Y153_AO5),
.O6(CLBLM_R_X3Y153_SLICE_X2Y153_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y153_SLICE_X3Y153_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y153_SLICE_X3Y153_DO5),
.O6(CLBLM_R_X3Y153_SLICE_X3Y153_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y153_SLICE_X3Y153_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y153_SLICE_X3Y153_CO5),
.O6(CLBLM_R_X3Y153_SLICE_X3Y153_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y153_SLICE_X3Y153_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y153_SLICE_X3Y153_BO5),
.O6(CLBLM_R_X3Y153_SLICE_X3Y153_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y153_SLICE_X3Y153_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y153_SLICE_X3Y153_AO5),
.O6(CLBLM_R_X3Y153_SLICE_X3Y153_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y140_SLICE_X6Y140_A5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y140_SLICE_X6Y140_DO6),
.Q(CLBLM_R_X5Y140_SLICE_X6Y140_A5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y140_SLICE_X6Y140_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y140_SLICE_X6Y140_AO6),
.Q(CLBLM_R_X5Y140_SLICE_X6Y140_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y140_SLICE_X6Y140_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y140_SLICE_X6Y140_BO6),
.Q(CLBLM_R_X5Y140_SLICE_X6Y140_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y140_SLICE_X6Y140_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y140_SLICE_X6Y140_CO6),
.Q(CLBLM_R_X5Y140_SLICE_X6Y140_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0ccf0cca0a00000)
  ) CLBLM_R_X5Y140_SLICE_X6Y140_DLUT (
.I0(CLBLL_L_X4Y140_SLICE_X4Y140_AQ),
.I1(CLBLM_R_X5Y141_SLICE_X6Y141_BQ),
.I2(CLBLM_R_X5Y140_SLICE_X6Y140_AQ),
.I3(LIOB33_X0Y61_IOB_X0Y62_I),
.I4(CLBLM_R_X5Y140_SLICE_X6Y140_CQ),
.I5(1'b1),
.O5(CLBLM_R_X5Y140_SLICE_X6Y140_DO5),
.O6(CLBLM_R_X5Y140_SLICE_X6Y140_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hf066f000f066f000)
  ) CLBLM_R_X5Y140_SLICE_X6Y140_CLUT (
.I0(CLBLL_L_X4Y140_SLICE_X4Y140_AQ),
.I1(CLBLM_R_X5Y140_SLICE_X6Y140_CQ),
.I2(CLBLM_R_X7Y147_SLICE_X9Y147_DQ),
.I3(LIOB33_X0Y61_IOB_X0Y62_I),
.I4(CLBLL_L_X4Y140_SLICE_X4Y140_CO6),
.I5(1'b1),
.O5(CLBLM_R_X5Y140_SLICE_X6Y140_CO5),
.O6(CLBLM_R_X5Y140_SLICE_X6Y140_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf7fdf7fd070d070d)
  ) CLBLM_R_X5Y140_SLICE_X6Y140_BLUT (
.I0(CLBLL_L_X4Y140_SLICE_X4Y140_CO6),
.I1(CLBLM_R_X5Y140_SLICE_X6Y140_BQ),
.I2(LIOB33_X0Y61_IOB_X0Y62_I),
.I3(CLBLM_R_X5Y140_SLICE_X6Y140_DO5),
.I4(1'b1),
.I5(CLBLM_R_X5Y142_SLICE_X6Y142_CQ),
.O5(CLBLM_R_X5Y140_SLICE_X6Y140_BO5),
.O6(CLBLM_R_X5Y140_SLICE_X6Y140_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff00007bf37bf3)
  ) CLBLM_R_X5Y140_SLICE_X6Y140_ALUT (
.I0(CLBLM_R_X5Y140_SLICE_X6Y140_CQ),
.I1(CLBLL_L_X4Y140_SLICE_X4Y140_CO6),
.I2(CLBLM_R_X5Y140_SLICE_X6Y140_AQ),
.I3(CLBLL_L_X4Y140_SLICE_X4Y140_AQ),
.I4(CLBLM_R_X5Y144_SLICE_X6Y144_DQ),
.I5(LIOB33_X0Y61_IOB_X0Y62_I),
.O5(CLBLM_R_X5Y140_SLICE_X6Y140_AO5),
.O6(CLBLM_R_X5Y140_SLICE_X6Y140_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X5Y140_SLICE_X7Y140_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y140_SLICE_X7Y140_DO5),
.O6(CLBLM_R_X5Y140_SLICE_X7Y140_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X5Y140_SLICE_X7Y140_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y140_SLICE_X7Y140_CO5),
.O6(CLBLM_R_X5Y140_SLICE_X7Y140_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X5Y140_SLICE_X7Y140_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y140_SLICE_X7Y140_BO5),
.O6(CLBLM_R_X5Y140_SLICE_X7Y140_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X5Y140_SLICE_X7Y140_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y140_SLICE_X7Y140_AO5),
.O6(CLBLM_R_X5Y140_SLICE_X7Y140_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y141_SLICE_X6Y141_B5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y141_SLICE_X6Y141_BO5),
.Q(CLBLM_R_X5Y141_SLICE_X6Y141_B5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y141_SLICE_X6Y141_D5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y141_SLICE_X6Y141_DO5),
.Q(CLBLM_R_X5Y141_SLICE_X6Y141_D5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y141_SLICE_X6Y141_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y141_SLICE_X6Y141_AO6),
.Q(CLBLM_R_X5Y141_SLICE_X6Y141_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y141_SLICE_X6Y141_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y141_SLICE_X6Y141_BO6),
.Q(CLBLM_R_X5Y141_SLICE_X6Y141_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y141_SLICE_X6Y141_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y141_SLICE_X6Y141_DO6),
.Q(CLBLM_R_X5Y141_SLICE_X6Y141_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0aaf0aaccffcc00)
  ) CLBLM_R_X5Y141_SLICE_X6Y141_DLUT (
.I0(RIOB33_X105Y107_IOB_X1Y108_I),
.I1(CLBLM_R_X5Y141_SLICE_X6Y141_AQ),
.I2(CLBLM_L_X8Y146_SLICE_X11Y146_DQ),
.I3(LIOB33_X0Y61_IOB_X0Y62_I),
.I4(RIOB33_X105Y123_IOB_X1Y123_I),
.I5(1'b1),
.O5(CLBLM_R_X5Y141_SLICE_X6Y141_DO5),
.O6(CLBLM_R_X5Y141_SLICE_X6Y141_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hcfcfc0c000cc00cc)
  ) CLBLM_R_X5Y141_SLICE_X6Y141_CLUT (
.I0(1'b1),
.I1(CLBLM_R_X5Y141_SLICE_X6Y141_D5Q),
.I2(LIOB33_X0Y61_IOB_X0Y62_I),
.I3(CLBLM_L_X8Y151_SLICE_X10Y151_B5Q),
.I4(CLBLM_L_X10Y145_SLICE_X12Y145_AQ),
.I5(1'b1),
.O5(CLBLM_R_X5Y141_SLICE_X6Y141_CO5),
.O6(CLBLM_R_X5Y141_SLICE_X6Y141_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hee44ee44e4e4e4e4)
  ) CLBLM_R_X5Y141_SLICE_X6Y141_BLUT (
.I0(LIOB33_X0Y61_IOB_X0Y62_I),
.I1(CLBLM_R_X5Y145_SLICE_X7Y145_AQ),
.I2(CLBLM_R_X5Y140_SLICE_X6Y140_CQ),
.I3(CLBLM_L_X8Y144_SLICE_X10Y144_BQ),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y141_SLICE_X6Y141_BO5),
.O6(CLBLM_R_X5Y141_SLICE_X6Y141_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hdddd8888d8d8d8d8)
  ) CLBLM_R_X5Y141_SLICE_X6Y141_ALUT (
.I0(LIOB33_X0Y61_IOB_X0Y62_I),
.I1(CLBLM_R_X5Y141_SLICE_X6Y141_DQ),
.I2(CLBLM_R_X5Y141_SLICE_X6Y141_AQ),
.I3(1'b1),
.I4(CLBLM_R_X5Y142_SLICE_X6Y142_AQ),
.I5(CLBLM_R_X11Y146_SLICE_X14Y146_DO6),
.O5(CLBLM_R_X5Y141_SLICE_X6Y141_AO5),
.O6(CLBLM_R_X5Y141_SLICE_X6Y141_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X5Y141_SLICE_X7Y141_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y141_SLICE_X7Y141_DO5),
.O6(CLBLM_R_X5Y141_SLICE_X7Y141_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X5Y141_SLICE_X7Y141_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y141_SLICE_X7Y141_CO5),
.O6(CLBLM_R_X5Y141_SLICE_X7Y141_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X5Y141_SLICE_X7Y141_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y141_SLICE_X7Y141_BO5),
.O6(CLBLM_R_X5Y141_SLICE_X7Y141_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X5Y141_SLICE_X7Y141_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y141_SLICE_X7Y141_AO5),
.O6(CLBLM_R_X5Y141_SLICE_X7Y141_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y142_SLICE_X6Y142_D5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y142_SLICE_X6Y142_DO5),
.Q(CLBLM_R_X5Y142_SLICE_X6Y142_D5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y142_SLICE_X6Y142_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y142_SLICE_X6Y142_AO6),
.Q(CLBLM_R_X5Y142_SLICE_X6Y142_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y142_SLICE_X6Y142_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y142_SLICE_X6Y142_BO6),
.Q(CLBLM_R_X5Y142_SLICE_X6Y142_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y142_SLICE_X6Y142_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y142_SLICE_X6Y142_CO6),
.Q(CLBLM_R_X5Y142_SLICE_X6Y142_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y142_SLICE_X6Y142_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y142_SLICE_X6Y142_DO6),
.Q(CLBLM_R_X5Y142_SLICE_X6Y142_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hf000f0ffaa00aaff)
  ) CLBLM_R_X5Y142_SLICE_X6Y142_DLUT (
.I0(CLBLM_R_X3Y142_SLICE_X2Y142_AQ),
.I1(1'b1),
.I2(CLBLM_L_X8Y143_SLICE_X11Y143_DQ),
.I3(LIOB33_X0Y61_IOB_X0Y62_I),
.I4(CLBLM_R_X3Y146_SLICE_X2Y146_D5Q),
.I5(1'b1),
.O5(CLBLM_R_X5Y142_SLICE_X6Y142_DO5),
.O6(CLBLM_R_X5Y142_SLICE_X6Y142_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hff00e0e0ff00e0e0)
  ) CLBLM_R_X5Y142_SLICE_X6Y142_CLUT (
.I0(CLBLM_R_X5Y143_SLICE_X6Y143_AQ),
.I1(CLBLM_R_X5Y142_SLICE_X6Y142_CQ),
.I2(CLBLM_R_X13Y149_SLICE_X18Y149_AO6),
.I3(CLBLM_R_X7Y151_SLICE_X8Y151_C5Q),
.I4(LIOB33_X0Y61_IOB_X0Y62_I),
.I5(1'b1),
.O5(CLBLM_R_X5Y142_SLICE_X6Y142_CO5),
.O6(CLBLM_R_X5Y142_SLICE_X6Y142_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'haaffaa00aaccaacc)
  ) CLBLM_R_X5Y142_SLICE_X6Y142_BLUT (
.I0(CLBLL_L_X2Y146_SLICE_X0Y146_CQ),
.I1(CLBLM_R_X5Y142_SLICE_X6Y142_BQ),
.I2(1'b1),
.I3(LIOB33_X0Y61_IOB_X0Y62_I),
.I4(CLBLL_L_X4Y142_SLICE_X5Y142_BQ),
.I5(CLBLM_R_X13Y149_SLICE_X18Y149_AO6),
.O5(CLBLM_R_X5Y142_SLICE_X6Y142_BO5),
.O6(CLBLM_R_X5Y142_SLICE_X6Y142_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hccccccccfafa00fa)
  ) CLBLM_R_X5Y142_SLICE_X6Y142_ALUT (
.I0(CLBLM_L_X8Y143_SLICE_X11Y143_DQ),
.I1(CLBLM_R_X3Y151_SLICE_X3Y151_AQ),
.I2(CLBLM_R_X5Y142_SLICE_X6Y142_AQ),
.I3(CLBLM_R_X5Y142_SLICE_X7Y142_BQ),
.I4(CLBLM_L_X10Y145_SLICE_X12Y145_AQ),
.I5(LIOB33_X0Y61_IOB_X0Y62_I),
.O5(CLBLM_R_X5Y142_SLICE_X6Y142_AO5),
.O6(CLBLM_R_X5Y142_SLICE_X6Y142_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y142_SLICE_X7Y142_A5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y142_SLICE_X7Y142_AO5),
.Q(CLBLM_R_X5Y142_SLICE_X7Y142_A5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y142_SLICE_X7Y142_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y142_SLICE_X7Y142_AO6),
.Q(CLBLM_R_X5Y142_SLICE_X7Y142_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y142_SLICE_X7Y142_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y141_SLICE_X6Y141_CO6),
.Q(CLBLM_R_X5Y142_SLICE_X7Y142_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X5Y142_SLICE_X7Y142_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y142_SLICE_X7Y142_DO5),
.O6(CLBLM_R_X5Y142_SLICE_X7Y142_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000001100000011)
  ) CLBLM_R_X5Y142_SLICE_X7Y142_CLUT (
.I0(CLBLM_R_X5Y147_SLICE_X6Y147_C5Q),
.I1(CLBLM_R_X5Y144_SLICE_X7Y144_DO6),
.I2(1'b1),
.I3(LIOB33_X0Y61_IOB_X0Y61_I),
.I4(CLBLM_R_X5Y142_SLICE_X7Y142_AQ),
.I5(1'b1),
.O5(CLBLM_R_X5Y142_SLICE_X7Y142_CO5),
.O6(CLBLM_R_X5Y142_SLICE_X7Y142_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h77bb77bbddeeddee)
  ) CLBLM_R_X5Y142_SLICE_X7Y142_BLUT (
.I0(CLBLL_L_X4Y143_SLICE_X4Y143_DQ),
.I1(CLBLM_R_X5Y141_SLICE_X6Y141_BQ),
.I2(1'b1),
.I3(CLBLL_L_X4Y142_SLICE_X5Y142_C5Q),
.I4(1'b1),
.I5(CLBLM_R_X5Y140_SLICE_X6Y140_A5Q),
.O5(CLBLM_R_X5Y142_SLICE_X7Y142_BO5),
.O6(CLBLM_R_X5Y142_SLICE_X7Y142_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hccffcc00aaf0aaf0)
  ) CLBLM_R_X5Y142_SLICE_X7Y142_ALUT (
.I0(CLBLM_R_X5Y142_SLICE_X7Y142_AQ),
.I1(CLBLM_R_X7Y143_SLICE_X9Y143_CQ),
.I2(CLBLL_L_X4Y149_SLICE_X5Y149_C5Q),
.I3(LIOB33_X0Y61_IOB_X0Y62_I),
.I4(CLBLM_R_X5Y147_SLICE_X6Y147_C5Q),
.I5(1'b1),
.O5(CLBLM_R_X5Y142_SLICE_X7Y142_AO5),
.O6(CLBLM_R_X5Y142_SLICE_X7Y142_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y143_SLICE_X6Y143_C5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y143_SLICE_X6Y143_CO5),
.Q(CLBLM_R_X5Y143_SLICE_X6Y143_C5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y143_SLICE_X6Y143_D5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y143_SLICE_X6Y143_DO5),
.Q(CLBLM_R_X5Y143_SLICE_X6Y143_D5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y143_SLICE_X6Y143_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y143_SLICE_X6Y143_AO6),
.Q(CLBLM_R_X5Y143_SLICE_X6Y143_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y143_SLICE_X6Y143_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y143_SLICE_X6Y143_BO6),
.Q(CLBLM_R_X5Y143_SLICE_X6Y143_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y143_SLICE_X6Y143_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y143_SLICE_X6Y143_CO6),
.Q(CLBLM_R_X5Y143_SLICE_X6Y143_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y143_SLICE_X6Y143_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y143_SLICE_X6Y143_DO6),
.Q(CLBLM_R_X5Y143_SLICE_X6Y143_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f0ff00cccc5050)
  ) CLBLM_R_X5Y143_SLICE_X6Y143_DLUT (
.I0(CLBLM_R_X5Y153_SLICE_X6Y153_B5Q),
.I1(CLBLM_R_X5Y143_SLICE_X6Y143_AQ),
.I2(CLBLM_R_X3Y144_SLICE_X2Y144_AQ),
.I3(CLBLM_R_X7Y142_SLICE_X8Y142_D5Q),
.I4(LIOB33_X0Y61_IOB_X0Y62_I),
.I5(1'b1),
.O5(CLBLM_R_X5Y143_SLICE_X6Y143_DO5),
.O6(CLBLM_R_X5Y143_SLICE_X6Y143_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hff00fcfcf0f0aaaa)
  ) CLBLM_R_X5Y143_SLICE_X6Y143_CLUT (
.I0(RIOB33_X105Y111_IOB_X1Y111_I),
.I1(CLBLM_R_X5Y143_SLICE_X6Y143_CQ),
.I2(CLBLM_R_X5Y143_SLICE_X6Y143_D5Q),
.I3(CLBLM_L_X8Y143_SLICE_X10Y143_BQ),
.I4(LIOB33_X0Y61_IOB_X0Y62_I),
.I5(1'b1),
.O5(CLBLM_R_X5Y143_SLICE_X6Y143_CO5),
.O6(CLBLM_R_X5Y143_SLICE_X6Y143_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'ha0a0e4e4a0a0e4e4)
  ) CLBLM_R_X5Y143_SLICE_X6Y143_BLUT (
.I0(LIOB33_X0Y61_IOB_X0Y62_I),
.I1(CLBLL_L_X2Y145_SLICE_X1Y145_DO5),
.I2(CLBLM_R_X7Y143_SLICE_X8Y143_AQ),
.I3(1'b1),
.I4(CLBLL_L_X2Y146_SLICE_X1Y146_CO5),
.I5(1'b1),
.O5(CLBLM_R_X5Y143_SLICE_X6Y143_BO5),
.O6(CLBLM_R_X5Y143_SLICE_X6Y143_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaaff33aaaaf030)
  ) CLBLM_R_X5Y143_SLICE_X6Y143_ALUT (
.I0(CLBLM_R_X3Y151_SLICE_X2Y151_AQ),
.I1(CLBLM_R_X7Y142_SLICE_X8Y142_C5Q),
.I2(CLBLM_R_X5Y143_SLICE_X6Y143_AQ),
.I3(CLBLM_R_X7Y152_SLICE_X8Y152_D5Q),
.I4(LIOB33_X0Y61_IOB_X0Y62_I),
.I5(CLBLL_L_X4Y143_SLICE_X5Y143_DQ),
.O5(CLBLM_R_X5Y143_SLICE_X6Y143_AO5),
.O6(CLBLM_R_X5Y143_SLICE_X6Y143_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y143_SLICE_X7Y143_C5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y143_SLICE_X7Y143_CO5),
.Q(CLBLM_R_X5Y143_SLICE_X7Y143_C5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y143_SLICE_X7Y143_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y143_SLICE_X7Y143_AO6),
.Q(CLBLM_R_X5Y143_SLICE_X7Y143_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y143_SLICE_X7Y143_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y143_SLICE_X7Y143_BO6),
.Q(CLBLM_R_X5Y143_SLICE_X7Y143_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y143_SLICE_X7Y143_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y143_SLICE_X7Y143_CO6),
.Q(CLBLM_R_X5Y143_SLICE_X7Y143_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffff77bbddee)
  ) CLBLM_R_X5Y143_SLICE_X7Y143_DLUT (
.I0(CLBLM_R_X5Y145_SLICE_X7Y145_AQ),
.I1(CLBLL_L_X4Y142_SLICE_X5Y142_CQ),
.I2(1'b1),
.I3(CLBLM_R_X5Y141_SLICE_X6Y141_B5Q),
.I4(CLBLM_R_X7Y144_SLICE_X8Y144_CQ),
.I5(CLBLM_R_X5Y142_SLICE_X7Y142_BO6),
.O5(CLBLM_R_X5Y143_SLICE_X7Y143_DO5),
.O6(CLBLM_R_X5Y143_SLICE_X7Y143_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f0aaaaccccff00)
  ) CLBLM_R_X5Y143_SLICE_X7Y143_CLUT (
.I0(CLBLM_R_X3Y151_SLICE_X3Y151_BQ),
.I1(CLBLM_R_X5Y143_SLICE_X7Y143_CQ),
.I2(CLBLM_R_X5Y151_SLICE_X7Y151_AQ),
.I3(CLBLL_L_X4Y144_SLICE_X5Y144_CQ),
.I4(LIOB33_X0Y61_IOB_X0Y62_I),
.I5(1'b1),
.O5(CLBLM_R_X5Y143_SLICE_X7Y143_CO5),
.O6(CLBLM_R_X5Y143_SLICE_X7Y143_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hffee5544afae0504)
  ) CLBLM_R_X5Y143_SLICE_X7Y143_BLUT (
.I0(LIOB33_X0Y61_IOB_X0Y62_I),
.I1(CLBLM_R_X5Y143_SLICE_X7Y143_BQ),
.I2(CLBLM_R_X3Y145_SLICE_X3Y145_D5Q),
.I3(CLBLM_R_X7Y145_SLICE_X8Y145_C5Q),
.I4(CLBLM_R_X3Y151_SLICE_X3Y151_BQ),
.I5(CLBLL_L_X4Y151_SLICE_X4Y151_BQ),
.O5(CLBLM_R_X5Y143_SLICE_X7Y143_BO5),
.O6(CLBLM_R_X5Y143_SLICE_X7Y143_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffb800b8ff8b008b)
  ) CLBLM_R_X5Y143_SLICE_X7Y143_ALUT (
.I0(CLBLM_R_X5Y143_SLICE_X6Y143_DQ),
.I1(CLBLM_L_X8Y149_SLICE_X11Y149_AQ),
.I2(CLBLM_R_X5Y143_SLICE_X7Y143_AQ),
.I3(LIOB33_X0Y61_IOB_X0Y62_I),
.I4(CLBLM_R_X5Y142_SLICE_X6Y142_AQ),
.I5(CLBLM_R_X7Y143_SLICE_X8Y143_DO6),
.O5(CLBLM_R_X5Y143_SLICE_X7Y143_AO5),
.O6(CLBLM_R_X5Y143_SLICE_X7Y143_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y144_SLICE_X6Y144_D5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y144_SLICE_X6Y144_DO5),
.Q(CLBLM_R_X5Y144_SLICE_X6Y144_D5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y144_SLICE_X6Y144_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y144_SLICE_X6Y144_AO6),
.Q(CLBLM_R_X5Y144_SLICE_X6Y144_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y144_SLICE_X6Y144_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y144_SLICE_X6Y144_BO6),
.Q(CLBLM_R_X5Y144_SLICE_X6Y144_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y144_SLICE_X6Y144_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y144_SLICE_X6Y144_CO6),
.Q(CLBLM_R_X5Y144_SLICE_X6Y144_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y144_SLICE_X6Y144_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y144_SLICE_X6Y144_DO6),
.Q(CLBLM_R_X5Y144_SLICE_X6Y144_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaa0ff0ccccf0f0)
  ) CLBLM_R_X5Y144_SLICE_X6Y144_DLUT (
.I0(CLBLM_R_X5Y144_SLICE_X6Y144_BQ),
.I1(CLBLL_L_X4Y144_SLICE_X4Y144_BQ),
.I2(CLBLM_R_X5Y145_SLICE_X6Y145_D5Q),
.I3(CLBLL_L_X4Y144_SLICE_X4Y144_D5Q),
.I4(LIOB33_X0Y61_IOB_X0Y62_I),
.I5(1'b1),
.O5(CLBLM_R_X5Y144_SLICE_X6Y144_DO5),
.O6(CLBLM_R_X5Y144_SLICE_X6Y144_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff000300000003)
  ) CLBLM_R_X5Y144_SLICE_X6Y144_CLUT (
.I0(1'b1),
.I1(CLBLM_R_X5Y145_SLICE_X6Y145_D5Q),
.I2(CLBLL_L_X4Y143_SLICE_X4Y143_BQ),
.I3(CLBLL_L_X4Y145_SLICE_X4Y145_DO5),
.I4(LIOB33_X0Y61_IOB_X0Y62_I),
.I5(CLBLM_R_X5Y144_SLICE_X6Y144_D5Q),
.O5(CLBLM_R_X5Y144_SLICE_X6Y144_CO5),
.O6(CLBLM_R_X5Y144_SLICE_X6Y144_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hff00ff00e4e4e4e4)
  ) CLBLM_R_X5Y144_SLICE_X6Y144_BLUT (
.I0(CLBLM_R_X13Y149_SLICE_X18Y149_AO6),
.I1(CLBLM_R_X5Y144_SLICE_X6Y144_BQ),
.I2(CLBLL_L_X4Y145_SLICE_X4Y145_AQ),
.I3(CLBLM_L_X8Y150_SLICE_X11Y150_AQ),
.I4(1'b1),
.I5(LIOB33_X0Y61_IOB_X0Y62_I),
.O5(CLBLM_R_X5Y144_SLICE_X6Y144_BO5),
.O6(CLBLM_R_X5Y144_SLICE_X6Y144_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hee44ee44fa50fa50)
  ) CLBLM_R_X5Y144_SLICE_X6Y144_ALUT (
.I0(LIOB33_X0Y61_IOB_X0Y62_I),
.I1(CLBLM_R_X5Y152_SLICE_X6Y152_AQ),
.I2(CLBLM_R_X5Y144_SLICE_X6Y144_AQ),
.I3(CLBLM_R_X7Y144_SLICE_X8Y144_D5Q),
.I4(1'b1),
.I5(CLBLM_R_X11Y146_SLICE_X14Y146_DO6),
.O5(CLBLM_R_X5Y144_SLICE_X6Y144_AO5),
.O6(CLBLM_R_X5Y144_SLICE_X6Y144_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y144_SLICE_X7Y144_B5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y144_SLICE_X7Y144_BO5),
.Q(CLBLM_R_X5Y144_SLICE_X7Y144_B5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "C5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y144_SLICE_X7Y144_C5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y144_SLICE_X7Y144_CO5),
.Q(CLBLM_R_X5Y144_SLICE_X7Y144_C5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y144_SLICE_X7Y144_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y144_SLICE_X7Y144_AO6),
.Q(CLBLM_R_X5Y144_SLICE_X7Y144_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y144_SLICE_X7Y144_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y144_SLICE_X7Y144_BO6),
.Q(CLBLM_R_X5Y144_SLICE_X7Y144_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y144_SLICE_X7Y144_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y144_SLICE_X7Y144_CO6),
.Q(CLBLM_R_X5Y144_SLICE_X7Y144_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffefefffffefe)
  ) CLBLM_R_X5Y144_SLICE_X7Y144_DLUT (
.I0(CLBLM_R_X5Y144_SLICE_X7Y144_C5Q),
.I1(CLBLL_L_X4Y148_SLICE_X5Y148_B5Q),
.I2(CLBLM_L_X8Y142_SLICE_X10Y142_A5Q),
.I3(1'b1),
.I4(CLBLM_L_X8Y152_SLICE_X10Y152_C5Q),
.I5(1'b1),
.O5(CLBLM_R_X5Y144_SLICE_X7Y144_DO5),
.O6(CLBLM_R_X5Y144_SLICE_X7Y144_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hfafa0a0af000ff0f)
  ) CLBLM_R_X5Y144_SLICE_X7Y144_CLUT (
.I0(CLBLM_R_X5Y143_SLICE_X7Y143_C5Q),
.I1(1'b1),
.I2(LIOB33_X0Y61_IOB_X0Y62_I),
.I3(CLBLM_R_X7Y144_SLICE_X8Y144_C5Q),
.I4(CLBLM_L_X8Y145_SLICE_X11Y145_DQ),
.I5(1'b1),
.O5(CLBLM_R_X5Y144_SLICE_X7Y144_CO5),
.O6(CLBLM_R_X5Y144_SLICE_X7Y144_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hff330033f0ccf0cc)
  ) CLBLM_R_X5Y144_SLICE_X7Y144_BLUT (
.I0(1'b1),
.I1(CLBLM_R_X3Y146_SLICE_X2Y146_D5Q),
.I2(CLBLM_R_X5Y151_SLICE_X7Y151_B5Q),
.I3(LIOB33_X0Y61_IOB_X0Y62_I),
.I4(CLBLM_R_X5Y144_SLICE_X7Y144_C5Q),
.I5(1'b1),
.O5(CLBLM_R_X5Y144_SLICE_X7Y144_BO5),
.O6(CLBLM_R_X5Y144_SLICE_X7Y144_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hccccccccfff000f0)
  ) CLBLM_R_X5Y144_SLICE_X7Y144_ALUT (
.I0(1'b1),
.I1(CLBLL_L_X4Y150_SLICE_X4Y150_C5Q),
.I2(CLBLM_R_X5Y144_SLICE_X7Y144_AQ),
.I3(CLBLM_R_X11Y146_SLICE_X14Y146_DO6),
.I4(CLBLM_R_X3Y150_SLICE_X2Y150_AQ),
.I5(LIOB33_X0Y61_IOB_X0Y62_I),
.O5(CLBLM_R_X5Y144_SLICE_X7Y144_AO5),
.O6(CLBLM_R_X5Y144_SLICE_X7Y144_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y145_SLICE_X6Y145_B5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y145_SLICE_X6Y145_BO5),
.Q(CLBLM_R_X5Y145_SLICE_X6Y145_B5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "C5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y145_SLICE_X6Y145_C5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y145_SLICE_X6Y145_CO5),
.Q(CLBLM_R_X5Y145_SLICE_X6Y145_C5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y145_SLICE_X6Y145_D5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y145_SLICE_X6Y145_DO5),
.Q(CLBLM_R_X5Y145_SLICE_X6Y145_D5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y145_SLICE_X6Y145_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y145_SLICE_X6Y145_AO6),
.Q(CLBLM_R_X5Y145_SLICE_X6Y145_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y145_SLICE_X6Y145_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y145_SLICE_X6Y145_BO6),
.Q(CLBLM_R_X5Y145_SLICE_X6Y145_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y145_SLICE_X6Y145_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y145_SLICE_X6Y145_CO6),
.Q(CLBLM_R_X5Y145_SLICE_X6Y145_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y145_SLICE_X6Y145_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y145_SLICE_X6Y145_DO6),
.Q(CLBLM_R_X5Y145_SLICE_X6Y145_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hb8b8b8b8ee22ff33)
  ) CLBLM_R_X5Y145_SLICE_X6Y145_DLUT (
.I0(CLBLM_R_X3Y145_SLICE_X2Y145_CQ),
.I1(LIOB33_X0Y61_IOB_X0Y62_I),
.I2(CLBLM_R_X3Y151_SLICE_X3Y151_AQ),
.I3(CLBLM_R_X5Y149_SLICE_X7Y149_CQ),
.I4(CLBLM_R_X5Y145_SLICE_X6Y145_D5Q),
.I5(1'b1),
.O5(CLBLM_R_X5Y145_SLICE_X6Y145_DO5),
.O6(CLBLM_R_X5Y145_SLICE_X6Y145_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hf303f303afa0afa0)
  ) CLBLM_R_X5Y145_SLICE_X6Y145_CLUT (
.I0(CLBLM_L_X8Y142_SLICE_X10Y142_A5Q),
.I1(CLBLM_R_X3Y146_SLICE_X2Y146_D5Q),
.I2(LIOB33_X0Y61_IOB_X0Y62_I),
.I3(CLBLM_R_X5Y142_SLICE_X6Y142_DQ),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y145_SLICE_X6Y145_CO5),
.O6(CLBLM_R_X5Y145_SLICE_X6Y145_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'haa33aaccf0aaf0aa)
  ) CLBLM_R_X5Y145_SLICE_X6Y145_BLUT (
.I0(CLBLL_L_X4Y145_SLICE_X5Y145_CQ),
.I1(CLBLL_L_X4Y151_SLICE_X4Y151_AQ),
.I2(CLBLM_R_X5Y145_SLICE_X6Y145_AQ),
.I3(LIOB33_X0Y61_IOB_X0Y62_I),
.I4(CLBLM_R_X7Y149_SLICE_X8Y149_A5Q),
.I5(1'b1),
.O5(CLBLM_R_X5Y145_SLICE_X6Y145_BO5),
.O6(CLBLM_R_X5Y145_SLICE_X6Y145_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hff00ff00f6f60000)
  ) CLBLM_R_X5Y145_SLICE_X6Y145_ALUT (
.I0(RIOB33_X105Y109_IOB_X1Y109_I),
.I1(CLBLM_R_X5Y147_SLICE_X7Y147_C5Q),
.I2(CLBLM_R_X5Y145_SLICE_X6Y145_AQ),
.I3(CLBLL_L_X2Y146_SLICE_X0Y146_BQ),
.I4(CLBLM_R_X7Y151_SLICE_X9Y151_A5Q),
.I5(LIOB33_X0Y61_IOB_X0Y62_I),
.O5(CLBLM_R_X5Y145_SLICE_X6Y145_AO5),
.O6(CLBLM_R_X5Y145_SLICE_X6Y145_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y145_SLICE_X7Y145_A5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y145_SLICE_X7Y145_AO5),
.Q(CLBLM_R_X5Y145_SLICE_X7Y145_A5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y145_SLICE_X7Y145_B5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y145_SLICE_X7Y145_BO5),
.Q(CLBLM_R_X5Y145_SLICE_X7Y145_B5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y145_SLICE_X7Y145_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y145_SLICE_X7Y145_AO6),
.Q(CLBLM_R_X5Y145_SLICE_X7Y145_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y145_SLICE_X7Y145_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y145_SLICE_X7Y145_BO6),
.Q(CLBLM_R_X5Y145_SLICE_X7Y145_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h3cffff3c3cffff3c)
  ) CLBLM_R_X5Y145_SLICE_X7Y145_DLUT (
.I0(1'b1),
.I1(CLBLM_R_X7Y145_SLICE_X8Y145_BQ),
.I2(CLBLM_R_X7Y146_SLICE_X8Y146_DQ),
.I3(CLBLM_R_X5Y146_SLICE_X7Y146_D5Q),
.I4(CLBLM_R_X3Y145_SLICE_X2Y145_B5Q),
.I5(1'b1),
.O5(CLBLM_R_X5Y145_SLICE_X7Y145_DO5),
.O6(CLBLM_R_X5Y145_SLICE_X7Y145_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffff7dffffffbe)
  ) CLBLM_R_X5Y145_SLICE_X7Y145_CLUT (
.I0(CLBLM_R_X3Y147_SLICE_X3Y147_C5Q),
.I1(CLBLM_R_X3Y148_SLICE_X3Y148_BQ),
.I2(CLBLL_L_X4Y146_SLICE_X4Y146_C5Q),
.I3(CLBLM_R_X5Y143_SLICE_X7Y143_DO6),
.I4(CLBLM_R_X5Y145_SLICE_X7Y145_DO6),
.I5(CLBLM_R_X5Y147_SLICE_X7Y147_B5Q),
.O5(CLBLM_R_X5Y145_SLICE_X7Y145_CO5),
.O6(CLBLM_R_X5Y145_SLICE_X7Y145_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfcfc0c0cc5c0c5c0)
  ) CLBLM_R_X5Y145_SLICE_X7Y145_BLUT (
.I0(CLBLM_L_X8Y144_SLICE_X10Y144_AO5),
.I1(CLBLL_L_X4Y147_SLICE_X4Y147_D5Q),
.I2(LIOB33_X0Y61_IOB_X0Y62_I),
.I3(CLBLM_L_X10Y144_SLICE_X12Y144_AO6),
.I4(CLBLM_L_X10Y151_SLICE_X12Y151_CQ),
.I5(1'b1),
.O5(CLBLM_R_X5Y145_SLICE_X7Y145_BO5),
.O6(CLBLM_R_X5Y145_SLICE_X7Y145_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hacacacacc0c0cfcf)
  ) CLBLM_R_X5Y145_SLICE_X7Y145_ALUT (
.I0(CLBLM_R_X5Y147_SLICE_X7Y147_CQ),
.I1(CLBLM_R_X3Y145_SLICE_X2Y145_B5Q),
.I2(LIOB33_X0Y61_IOB_X0Y62_I),
.I3(1'b1),
.I4(CLBLM_L_X10Y153_SLICE_X13Y153_A5Q),
.I5(1'b1),
.O5(CLBLM_R_X5Y145_SLICE_X7Y145_AO5),
.O6(CLBLM_R_X5Y145_SLICE_X7Y145_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y146_SLICE_X6Y146_B5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y146_SLICE_X6Y146_BO5),
.Q(CLBLM_R_X5Y146_SLICE_X6Y146_B5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y146_SLICE_X6Y146_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y146_SLICE_X6Y146_AO6),
.Q(CLBLM_R_X5Y146_SLICE_X6Y146_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y146_SLICE_X6Y146_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y146_SLICE_X6Y146_BO6),
.Q(CLBLM_R_X5Y146_SLICE_X6Y146_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0ff0ffffffff0ff0)
  ) CLBLM_R_X5Y146_SLICE_X6Y146_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(CLBLM_R_X3Y147_SLICE_X2Y147_BQ),
.I3(CLBLL_L_X4Y144_SLICE_X4Y144_DQ),
.I4(CLBLM_R_X3Y145_SLICE_X3Y145_C5Q),
.I5(CLBLM_R_X3Y147_SLICE_X2Y147_AQ),
.O5(CLBLM_R_X5Y146_SLICE_X6Y146_DO5),
.O6(CLBLM_R_X5Y146_SLICE_X6Y146_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h7777ddddbbbbeeee)
  ) CLBLM_R_X5Y146_SLICE_X6Y146_CLUT (
.I0(CLBLL_L_X2Y145_SLICE_X1Y145_AQ),
.I1(CLBLM_R_X3Y149_SLICE_X2Y149_BQ),
.I2(1'b1),
.I3(1'b1),
.I4(CLBLM_R_X7Y147_SLICE_X9Y147_DQ),
.I5(CLBLM_R_X5Y142_SLICE_X7Y142_A5Q),
.O5(CLBLM_R_X5Y146_SLICE_X6Y146_CO5),
.O6(CLBLM_R_X5Y146_SLICE_X6Y146_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hcfcfc0c0ff0ff000)
  ) CLBLM_R_X5Y146_SLICE_X6Y146_BLUT (
.I0(1'b1),
.I1(CLBLM_R_X3Y146_SLICE_X3Y146_BQ),
.I2(LIOB33_X0Y61_IOB_X0Y62_I),
.I3(CLBLM_R_X7Y149_SLICE_X8Y149_A5Q),
.I4(CLBLL_L_X4Y149_SLICE_X5Y149_C5Q),
.I5(1'b1),
.O5(CLBLM_R_X5Y146_SLICE_X6Y146_BO5),
.O6(CLBLM_R_X5Y146_SLICE_X6Y146_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hff33cc00fc30fc30)
  ) CLBLM_R_X5Y146_SLICE_X6Y146_ALUT (
.I0(1'b1),
.I1(LIOB33_X0Y61_IOB_X0Y62_I),
.I2(CLBLM_R_X5Y146_SLICE_X6Y146_AQ),
.I3(CLBLM_R_X5Y147_SLICE_X6Y147_BQ),
.I4(CLBLL_L_X4Y144_SLICE_X5Y144_AQ),
.I5(CLBLM_R_X11Y148_SLICE_X15Y148_AO6),
.O5(CLBLM_R_X5Y146_SLICE_X6Y146_AO5),
.O6(CLBLM_R_X5Y146_SLICE_X6Y146_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y146_SLICE_X7Y146_C5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y146_SLICE_X7Y146_CO5),
.Q(CLBLM_R_X5Y146_SLICE_X7Y146_C5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y146_SLICE_X7Y146_D5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y146_SLICE_X7Y146_DO5),
.Q(CLBLM_R_X5Y146_SLICE_X7Y146_D5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y146_SLICE_X7Y146_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y146_SLICE_X7Y146_AO6),
.Q(CLBLM_R_X5Y146_SLICE_X7Y146_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y146_SLICE_X7Y146_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y146_SLICE_X7Y146_BO6),
.Q(CLBLM_R_X5Y146_SLICE_X7Y146_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y146_SLICE_X7Y146_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y146_SLICE_X7Y146_CO6),
.Q(CLBLM_R_X5Y146_SLICE_X7Y146_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y146_SLICE_X7Y146_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y146_SLICE_X7Y146_DO6),
.Q(CLBLM_R_X5Y146_SLICE_X7Y146_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'haaffaa00ccf0ccf0)
  ) CLBLM_R_X5Y146_SLICE_X7Y146_DLUT (
.I0(CLBLM_L_X8Y154_SLICE_X11Y154_AQ),
.I1(CLBLM_L_X8Y152_SLICE_X10Y152_DQ),
.I2(CLBLM_R_X3Y145_SLICE_X2Y145_B5Q),
.I3(LIOB33_X0Y61_IOB_X0Y62_I),
.I4(CLBLM_R_X5Y149_SLICE_X6Y149_B5Q),
.I5(1'b1),
.O5(CLBLM_R_X5Y146_SLICE_X7Y146_DO5),
.O6(CLBLM_R_X5Y146_SLICE_X7Y146_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hbbbb1111b1b1b1b1)
  ) CLBLM_R_X5Y146_SLICE_X7Y146_CLUT (
.I0(LIOB33_X0Y61_IOB_X0Y62_I),
.I1(CLBLM_L_X12Y151_SLICE_X16Y151_AQ),
.I2(CLBLM_R_X3Y146_SLICE_X2Y146_AQ),
.I3(1'b1),
.I4(CLBLM_R_X5Y145_SLICE_X7Y145_BQ),
.I5(1'b1),
.O5(CLBLM_R_X5Y146_SLICE_X7Y146_CO5),
.O6(CLBLM_R_X5Y146_SLICE_X7Y146_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hff00ff0000000c0c)
  ) CLBLM_R_X5Y146_SLICE_X7Y146_BLUT (
.I0(1'b1),
.I1(CLBLM_R_X5Y145_SLICE_X6Y145_D5Q),
.I2(CLBLL_L_X4Y145_SLICE_X4Y145_DO5),
.I3(CLBLM_L_X8Y148_SLICE_X11Y148_BQ),
.I4(CLBLL_L_X4Y143_SLICE_X4Y143_BQ),
.I5(LIOB33_X0Y61_IOB_X0Y62_I),
.O5(CLBLM_R_X5Y146_SLICE_X7Y146_BO5),
.O6(CLBLM_R_X5Y146_SLICE_X7Y146_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffb800b8ffaa00aa)
  ) CLBLM_R_X5Y146_SLICE_X7Y146_ALUT (
.I0(CLBLL_L_X4Y146_SLICE_X4Y146_BQ),
.I1(CLBLM_R_X7Y152_SLICE_X8Y152_D5Q),
.I2(CLBLM_R_X5Y146_SLICE_X7Y146_AQ),
.I3(LIOB33_X0Y61_IOB_X0Y62_I),
.I4(CLBLL_L_X2Y145_SLICE_X1Y145_AQ),
.I5(CLBLM_R_X7Y142_SLICE_X8Y142_C5Q),
.O5(CLBLM_R_X5Y146_SLICE_X7Y146_AO5),
.O6(CLBLM_R_X5Y146_SLICE_X7Y146_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y147_SLICE_X6Y147_B5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y147_SLICE_X6Y147_BO5),
.Q(CLBLM_R_X5Y147_SLICE_X6Y147_B5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "C5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y147_SLICE_X6Y147_C5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y147_SLICE_X6Y147_CO5),
.Q(CLBLM_R_X5Y147_SLICE_X6Y147_C5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y147_SLICE_X6Y147_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y147_SLICE_X6Y147_AO6),
.Q(CLBLM_R_X5Y147_SLICE_X6Y147_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y147_SLICE_X6Y147_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y147_SLICE_X6Y147_BO6),
.Q(CLBLM_R_X5Y147_SLICE_X6Y147_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y147_SLICE_X6Y147_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y147_SLICE_X6Y147_CO6),
.Q(CLBLM_R_X5Y147_SLICE_X6Y147_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h66ff66ffff66ff66)
  ) CLBLM_R_X5Y147_SLICE_X6Y147_DLUT (
.I0(CLBLM_R_X3Y147_SLICE_X2Y147_AQ),
.I1(CLBLM_R_X7Y144_SLICE_X8Y144_D5Q),
.I2(1'b1),
.I3(CLBLM_R_X5Y145_SLICE_X7Y145_A5Q),
.I4(1'b1),
.I5(CLBLM_R_X3Y147_SLICE_X2Y147_BQ),
.O5(CLBLM_R_X5Y147_SLICE_X6Y147_DO5),
.O6(CLBLM_R_X5Y147_SLICE_X6Y147_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hde12de12bbbb8888)
  ) CLBLM_R_X5Y147_SLICE_X6Y147_CLUT (
.I0(CLBLL_L_X4Y143_SLICE_X4Y143_BQ),
.I1(LIOB33_X0Y61_IOB_X0Y62_I),
.I2(CLBLM_R_X7Y153_SLICE_X8Y153_AQ),
.I3(CLBLL_L_X4Y151_SLICE_X4Y151_CQ),
.I4(CLBLM_L_X8Y154_SLICE_X10Y154_BO5),
.I5(1'b1),
.O5(CLBLM_R_X5Y147_SLICE_X6Y147_CO5),
.O6(CLBLM_R_X5Y147_SLICE_X6Y147_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hcfcfc0c0fa0afa0a)
  ) CLBLM_R_X5Y147_SLICE_X6Y147_BLUT (
.I0(CLBLM_R_X5Y153_SLICE_X6Y153_B5Q),
.I1(CLBLM_R_X7Y144_SLICE_X8Y144_B5Q),
.I2(LIOB33_X0Y61_IOB_X0Y62_I),
.I3(CLBLM_R_X3Y150_SLICE_X3Y150_BQ),
.I4(CLBLL_L_X4Y151_SLICE_X4Y151_AQ),
.I5(1'b1),
.O5(CLBLM_R_X5Y147_SLICE_X6Y147_BO5),
.O6(CLBLM_R_X5Y147_SLICE_X6Y147_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfaf0fbf00a000b00)
  ) CLBLM_R_X5Y147_SLICE_X6Y147_ALUT (
.I0(CLBLL_L_X4Y150_SLICE_X4Y150_DO6),
.I1(CLBLL_L_X4Y146_SLICE_X5Y146_BQ),
.I2(LIOB33_X0Y61_IOB_X0Y62_I),
.I3(CLBLL_L_X2Y150_SLICE_X1Y150_AQ),
.I4(CLBLM_R_X5Y146_SLICE_X7Y146_BQ),
.I5(CLBLM_L_X8Y147_SLICE_X11Y147_CQ),
.O5(CLBLM_R_X5Y147_SLICE_X6Y147_AO5),
.O6(CLBLM_R_X5Y147_SLICE_X6Y147_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y147_SLICE_X7Y147_B5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y147_SLICE_X7Y147_BO5),
.Q(CLBLM_R_X5Y147_SLICE_X7Y147_B5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "C5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y147_SLICE_X7Y147_C5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y147_SLICE_X7Y147_CO5),
.Q(CLBLM_R_X5Y147_SLICE_X7Y147_C5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y147_SLICE_X7Y147_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y147_SLICE_X7Y147_AO6),
.Q(CLBLM_R_X5Y147_SLICE_X7Y147_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y147_SLICE_X7Y147_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y147_SLICE_X7Y147_BO6),
.Q(CLBLM_R_X5Y147_SLICE_X7Y147_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y147_SLICE_X7Y147_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y147_SLICE_X7Y147_CO6),
.Q(CLBLM_R_X5Y147_SLICE_X7Y147_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000040004)
  ) CLBLM_R_X5Y147_SLICE_X7Y147_DLUT (
.I0(CLBLM_R_X7Y151_SLICE_X9Y151_DQ),
.I1(CLBLM_R_X7Y147_SLICE_X8Y147_AO6),
.I2(CLBLM_R_X7Y153_SLICE_X9Y153_CQ),
.I3(CLBLM_R_X3Y148_SLICE_X2Y148_DO6),
.I4(1'b1),
.I5(CLBLM_L_X8Y148_SLICE_X10Y148_BQ),
.O5(CLBLM_R_X5Y147_SLICE_X7Y147_DO5),
.O6(CLBLM_R_X5Y147_SLICE_X7Y147_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hffcc00ccaaf0aaf0)
  ) CLBLM_R_X5Y147_SLICE_X7Y147_CLUT (
.I0(CLBLM_R_X7Y151_SLICE_X9Y151_DQ),
.I1(CLBLM_R_X5Y145_SLICE_X6Y145_D5Q),
.I2(RIOB33_X105Y109_IOB_X1Y109_I),
.I3(LIOB33_X0Y61_IOB_X0Y62_I),
.I4(CLBLM_L_X10Y153_SLICE_X12Y153_A5Q),
.I5(1'b1),
.O5(CLBLM_R_X5Y147_SLICE_X7Y147_CO5),
.O6(CLBLM_R_X5Y147_SLICE_X7Y147_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hd8d8d8d8ff55aa00)
  ) CLBLM_R_X5Y147_SLICE_X7Y147_BLUT (
.I0(LIOB33_X0Y61_IOB_X0Y62_I),
.I1(CLBLM_R_X7Y154_SLICE_X8Y154_BQ),
.I2(RIOB33_X105Y123_IOB_X1Y124_I),
.I3(CLBLM_R_X7Y147_SLICE_X9Y147_CQ),
.I4(CLBLM_R_X3Y147_SLICE_X3Y147_C5Q),
.I5(1'b1),
.O5(CLBLM_R_X5Y147_SLICE_X7Y147_BO5),
.O6(CLBLM_R_X5Y147_SLICE_X7Y147_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff0000e2f0e2f0)
  ) CLBLM_R_X5Y147_SLICE_X7Y147_ALUT (
.I0(CLBLM_R_X5Y149_SLICE_X7Y149_DQ),
.I1(CLBLM_L_X8Y147_SLICE_X10Y147_C5Q),
.I2(CLBLM_R_X5Y147_SLICE_X7Y147_AQ),
.I3(CLBLM_L_X10Y144_SLICE_X13Y144_CQ),
.I4(CLBLM_R_X5Y148_SLICE_X7Y148_C5Q),
.I5(LIOB33_X0Y61_IOB_X0Y62_I),
.O5(CLBLM_R_X5Y147_SLICE_X7Y147_AO5),
.O6(CLBLM_R_X5Y147_SLICE_X7Y147_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y148_SLICE_X6Y148_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(LIOB33_X0Y61_IOB_X0Y62_I),
.D(CLBLL_L_X4Y151_SLICE_X5Y151_CQ),
.Q(CLBLM_R_X5Y148_SLICE_X6Y148_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y148_SLICE_X6Y148_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(LIOB33_X0Y61_IOB_X0Y62_I),
.D(CLBLL_L_X4Y147_SLICE_X5Y147_CQ),
.Q(CLBLM_R_X5Y148_SLICE_X6Y148_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y148_SLICE_X6Y148_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(LIOB33_X0Y61_IOB_X0Y62_I),
.D(CLBLM_R_X5Y149_SLICE_X7Y149_C5Q),
.Q(CLBLM_R_X5Y148_SLICE_X6Y148_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hffcfffffffffffff)
  ) CLBLM_R_X5Y148_SLICE_X6Y148_DLUT (
.I0(1'b1),
.I1(CLBLM_R_X7Y153_SLICE_X8Y153_CQ),
.I2(CLBLM_R_X3Y150_SLICE_X3Y150_A5Q),
.I3(CLBLM_R_X3Y144_SLICE_X3Y144_AQ),
.I4(CLBLM_L_X10Y148_SLICE_X13Y148_C5Q),
.I5(CLBLL_L_X4Y146_SLICE_X5Y146_AO5),
.O5(CLBLM_R_X5Y148_SLICE_X6Y148_DO5),
.O6(CLBLM_R_X5Y148_SLICE_X6Y148_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hff7fffffffffffff)
  ) CLBLM_R_X5Y148_SLICE_X6Y148_CLUT (
.I0(CLBLM_R_X7Y151_SLICE_X9Y151_BQ),
.I1(CLBLM_R_X5Y149_SLICE_X6Y149_AQ),
.I2(CLBLM_R_X5Y143_SLICE_X7Y143_AQ),
.I3(CLBLM_R_X7Y143_SLICE_X8Y143_DO6),
.I4(CLBLM_R_X7Y150_SLICE_X8Y150_AQ),
.I5(CLBLL_L_X4Y147_SLICE_X5Y147_AQ),
.O5(CLBLM_R_X5Y148_SLICE_X6Y148_CO5),
.O6(CLBLM_R_X5Y148_SLICE_X6Y148_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffffffeffffe)
  ) CLBLM_R_X5Y148_SLICE_X6Y148_BLUT (
.I0(CLBLM_R_X5Y146_SLICE_X6Y146_DO6),
.I1(CLBLM_R_X5Y148_SLICE_X7Y148_DO6),
.I2(CLBLM_R_X7Y142_SLICE_X8Y142_DQ),
.I3(CLBLM_R_X7Y148_SLICE_X8Y148_DO6),
.I4(CLBLL_L_X4Y152_SLICE_X5Y152_AQ),
.I5(CLBLM_R_X5Y149_SLICE_X6Y149_DO6),
.O5(CLBLM_R_X5Y148_SLICE_X6Y148_BO5),
.O6(CLBLM_R_X5Y148_SLICE_X6Y148_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hf7fffffff7f7ffff)
  ) CLBLM_R_X5Y148_SLICE_X6Y148_ALUT (
.I0(CLBLM_R_X7Y150_SLICE_X8Y150_AQ),
.I1(CLBLM_R_X7Y151_SLICE_X9Y151_BQ),
.I2(CLBLM_R_X7Y143_SLICE_X8Y143_DO6),
.I3(CLBLM_R_X5Y149_SLICE_X6Y149_AQ),
.I4(CLBLM_R_X5Y143_SLICE_X7Y143_AQ),
.I5(1'b1),
.O5(CLBLM_R_X5Y148_SLICE_X6Y148_AO5),
.O6(CLBLM_R_X5Y148_SLICE_X6Y148_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y148_SLICE_X7Y148_C5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y148_SLICE_X7Y148_CO5),
.Q(CLBLM_R_X5Y148_SLICE_X7Y148_C5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y148_SLICE_X7Y148_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y148_SLICE_X7Y148_AO6),
.Q(CLBLM_R_X5Y148_SLICE_X7Y148_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y148_SLICE_X7Y148_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y148_SLICE_X7Y148_BO6),
.Q(CLBLM_R_X5Y148_SLICE_X7Y148_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y148_SLICE_X7Y148_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y148_SLICE_X7Y148_CO6),
.Q(CLBLM_R_X5Y148_SLICE_X7Y148_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h77dd77ddbbeebbee)
  ) CLBLM_R_X5Y148_SLICE_X7Y148_DLUT (
.I0(CLBLM_R_X5Y154_SLICE_X6Y154_AQ),
.I1(CLBLM_R_X5Y154_SLICE_X6Y154_BQ),
.I2(1'b1),
.I3(CLBLM_R_X7Y148_SLICE_X9Y148_A5Q),
.I4(1'b1),
.I5(CLBLM_L_X8Y147_SLICE_X11Y147_CQ),
.O5(CLBLM_R_X5Y148_SLICE_X7Y148_DO5),
.O6(CLBLM_R_X5Y148_SLICE_X7Y148_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hcccc5a5aff00aaaa)
  ) CLBLM_R_X5Y148_SLICE_X7Y148_CLUT (
.I0(CLBLL_L_X4Y143_SLICE_X4Y143_BQ),
.I1(CLBLM_R_X5Y148_SLICE_X7Y148_AQ),
.I2(CLBLL_L_X4Y150_SLICE_X4Y150_CQ),
.I3(CLBLM_R_X7Y143_SLICE_X8Y143_BQ),
.I4(LIOB33_X0Y61_IOB_X0Y62_I),
.I5(1'b1),
.O5(CLBLM_R_X5Y148_SLICE_X7Y148_CO5),
.O6(CLBLM_R_X5Y148_SLICE_X7Y148_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff0000ee44ee44)
  ) CLBLM_R_X5Y148_SLICE_X7Y148_BLUT (
.I0(CLBLM_R_X11Y148_SLICE_X15Y148_AO6),
.I1(CLBLM_R_X5Y148_SLICE_X7Y148_BQ),
.I2(1'b1),
.I3(CLBLM_R_X5Y148_SLICE_X7Y148_AQ),
.I4(CLBLM_R_X5Y146_SLICE_X7Y146_D5Q),
.I5(LIOB33_X0Y61_IOB_X0Y62_I),
.O5(CLBLM_R_X5Y148_SLICE_X7Y148_BO5),
.O6(CLBLM_R_X5Y148_SLICE_X7Y148_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff0000fa32fa32)
  ) CLBLM_R_X5Y148_SLICE_X7Y148_ALUT (
.I0(CLBLM_R_X5Y147_SLICE_X7Y147_CQ),
.I1(CLBLL_L_X4Y142_SLICE_X5Y142_DQ),
.I2(CLBLM_R_X5Y148_SLICE_X7Y148_AQ),
.I3(CLBLL_L_X4Y147_SLICE_X5Y147_CQ),
.I4(CLBLM_R_X3Y148_SLICE_X3Y148_CQ),
.I5(LIOB33_X0Y61_IOB_X0Y62_I),
.O5(CLBLM_R_X5Y148_SLICE_X7Y148_AO5),
.O6(CLBLM_R_X5Y148_SLICE_X7Y148_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y149_SLICE_X6Y149_B5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y149_SLICE_X6Y149_BO5),
.Q(CLBLM_R_X5Y149_SLICE_X6Y149_B5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "C5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y149_SLICE_X6Y149_C5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y149_SLICE_X6Y149_CO5),
.Q(CLBLM_R_X5Y149_SLICE_X6Y149_C5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y149_SLICE_X6Y149_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y149_SLICE_X6Y149_AO6),
.Q(CLBLM_R_X5Y149_SLICE_X6Y149_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y149_SLICE_X6Y149_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y149_SLICE_X6Y149_BO6),
.Q(CLBLM_R_X5Y149_SLICE_X6Y149_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y149_SLICE_X6Y149_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y149_SLICE_X6Y149_CO6),
.Q(CLBLM_R_X5Y149_SLICE_X6Y149_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hbbeeffffffffbbee)
  ) CLBLM_R_X5Y149_SLICE_X6Y149_DLUT (
.I0(CLBLM_R_X3Y149_SLICE_X2Y149_AQ),
.I1(CLBLL_L_X4Y153_SLICE_X5Y153_AQ),
.I2(1'b1),
.I3(CLBLM_L_X8Y152_SLICE_X11Y152_D5Q),
.I4(CLBLM_L_X8Y144_SLICE_X11Y144_BQ),
.I5(CLBLM_R_X3Y152_SLICE_X3Y152_AQ),
.O5(CLBLM_R_X5Y149_SLICE_X6Y149_DO5),
.O6(CLBLM_R_X5Y149_SLICE_X6Y149_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hf000fc0cafafa0a0)
  ) CLBLM_R_X5Y149_SLICE_X6Y149_CLUT (
.I0(CLBLL_L_X4Y148_SLICE_X4Y148_C5Q),
.I1(CLBLM_L_X8Y151_SLICE_X10Y151_AQ),
.I2(LIOB33_X0Y61_IOB_X0Y62_I),
.I3(CLBLL_L_X4Y143_SLICE_X5Y143_DQ),
.I4(CLBLM_L_X8Y145_SLICE_X11Y145_DQ),
.I5(1'b1),
.O5(CLBLM_R_X5Y149_SLICE_X6Y149_CO5),
.O6(CLBLM_R_X5Y149_SLICE_X6Y149_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hffaa00aacc00ccff)
  ) CLBLM_R_X5Y149_SLICE_X6Y149_BLUT (
.I0(CLBLM_L_X10Y149_SLICE_X13Y149_AQ),
.I1(CLBLL_L_X4Y148_SLICE_X5Y148_BQ),
.I2(1'b1),
.I3(LIOB33_X0Y61_IOB_X0Y62_I),
.I4(CLBLM_R_X5Y148_SLICE_X6Y148_AQ),
.I5(1'b1),
.O5(CLBLM_R_X5Y149_SLICE_X6Y149_BO5),
.O6(CLBLM_R_X5Y149_SLICE_X6Y149_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hff00d8d8ff008d8d)
  ) CLBLM_R_X5Y149_SLICE_X6Y149_ALUT (
.I0(CLBLM_L_X8Y149_SLICE_X11Y149_AQ),
.I1(CLBLM_R_X7Y151_SLICE_X9Y151_C5Q),
.I2(CLBLM_R_X5Y149_SLICE_X6Y149_AQ),
.I3(CLBLL_L_X4Y145_SLICE_X5Y145_C5Q),
.I4(LIOB33_X0Y61_IOB_X0Y62_I),
.I5(CLBLM_R_X5Y148_SLICE_X6Y148_AO5),
.O5(CLBLM_R_X5Y149_SLICE_X6Y149_AO5),
.O6(CLBLM_R_X5Y149_SLICE_X6Y149_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y149_SLICE_X7Y149_C5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y149_SLICE_X7Y149_CO5),
.Q(CLBLM_R_X5Y149_SLICE_X7Y149_C5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y149_SLICE_X7Y149_D5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y149_SLICE_X7Y149_DO5),
.Q(CLBLM_R_X5Y149_SLICE_X7Y149_D5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y149_SLICE_X7Y149_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y149_SLICE_X7Y149_AO6),
.Q(CLBLM_R_X5Y149_SLICE_X7Y149_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y149_SLICE_X7Y149_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y149_SLICE_X7Y149_BO6),
.Q(CLBLM_R_X5Y149_SLICE_X7Y149_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y149_SLICE_X7Y149_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y149_SLICE_X7Y149_CO6),
.Q(CLBLM_R_X5Y149_SLICE_X7Y149_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y149_SLICE_X7Y149_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y149_SLICE_X7Y149_DO6),
.Q(CLBLM_R_X5Y149_SLICE_X7Y149_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hffcc3300bbbb8888)
  ) CLBLM_R_X5Y149_SLICE_X7Y149_DLUT (
.I0(CLBLM_R_X5Y150_SLICE_X6Y150_A5Q),
.I1(LIOB33_X0Y61_IOB_X0Y62_I),
.I2(1'b1),
.I3(CLBLL_L_X4Y149_SLICE_X4Y149_AQ),
.I4(CLBLM_R_X5Y149_SLICE_X7Y149_AQ),
.I5(1'b1),
.O5(CLBLM_R_X5Y149_SLICE_X7Y149_DO5),
.O6(CLBLM_R_X5Y149_SLICE_X7Y149_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hee22ee22cffc0330)
  ) CLBLM_R_X5Y149_SLICE_X7Y149_CLUT (
.I0(CLBLM_L_X10Y153_SLICE_X13Y153_A5Q),
.I1(LIOB33_X0Y61_IOB_X0Y62_I),
.I2(CLBLM_R_X3Y151_SLICE_X3Y151_BQ),
.I3(CLBLM_R_X7Y149_SLICE_X9Y149_CQ),
.I4(CLBLM_R_X7Y144_SLICE_X9Y144_AQ),
.I5(1'b1),
.O5(CLBLM_R_X5Y149_SLICE_X7Y149_CO5),
.O6(CLBLM_R_X5Y149_SLICE_X7Y149_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hafa0afafaca0acac)
  ) CLBLM_R_X5Y149_SLICE_X7Y149_BLUT (
.I0(CLBLM_R_X3Y144_SLICE_X3Y144_AQ),
.I1(CLBLM_R_X5Y149_SLICE_X7Y149_BQ),
.I2(LIOB33_X0Y61_IOB_X0Y62_I),
.I3(CLBLM_R_X7Y152_SLICE_X8Y152_D5Q),
.I4(CLBLM_R_X7Y142_SLICE_X8Y142_C5Q),
.I5(CLBLM_R_X5Y152_SLICE_X7Y152_B5Q),
.O5(CLBLM_R_X5Y149_SLICE_X7Y149_BO5),
.O6(CLBLM_R_X5Y149_SLICE_X7Y149_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfc30fc30dc10ec20)
  ) CLBLM_R_X5Y149_SLICE_X7Y149_ALUT (
.I0(CLBLL_L_X4Y151_SLICE_X4Y151_B5Q),
.I1(LIOB33_X0Y61_IOB_X0Y62_I),
.I2(CLBLM_R_X7Y151_SLICE_X9Y151_A5Q),
.I3(CLBLM_L_X10Y149_SLICE_X12Y149_A5Q),
.I4(RIOB33_X105Y107_IOB_X1Y107_I),
.I5(CLBLM_R_X5Y149_SLICE_X7Y149_AQ),
.O5(CLBLM_R_X5Y149_SLICE_X7Y149_AO5),
.O6(CLBLM_R_X5Y149_SLICE_X7Y149_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y150_SLICE_X6Y150_A5_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_R_X5Y150_SLICE_X6Y150_AO5),
.Q(CLBLM_R_X5Y150_SLICE_X6Y150_A5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y150_SLICE_X6Y150_B5_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_R_X5Y150_SLICE_X6Y150_BO5),
.Q(CLBLM_R_X5Y150_SLICE_X6Y150_B5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "C5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y150_SLICE_X6Y150_C5_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_R_X5Y150_SLICE_X6Y150_CO5),
.Q(CLBLM_R_X5Y150_SLICE_X6Y150_C5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y150_SLICE_X6Y150_A_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_R_X5Y150_SLICE_X6Y150_AO6),
.Q(CLBLM_R_X5Y150_SLICE_X6Y150_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y150_SLICE_X6Y150_B_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_R_X5Y150_SLICE_X6Y150_BO6),
.Q(CLBLM_R_X5Y150_SLICE_X6Y150_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y150_SLICE_X6Y150_C_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_R_X5Y150_SLICE_X6Y150_CO6),
.Q(CLBLM_R_X5Y150_SLICE_X6Y150_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000001)
  ) CLBLM_R_X5Y150_SLICE_X6Y150_DLUT (
.I0(CLBLM_R_X5Y150_SLICE_X6Y150_BQ),
.I1(CLBLM_R_X5Y151_SLICE_X7Y151_B5Q),
.I2(CLBLM_R_X5Y151_SLICE_X6Y151_DO6),
.I3(CLBLM_R_X5Y150_SLICE_X6Y150_A5Q),
.I4(CLBLM_R_X5Y145_SLICE_X6Y145_BQ),
.I5(CLBLM_L_X8Y146_SLICE_X11Y146_DQ),
.O5(CLBLM_R_X5Y150_SLICE_X6Y150_DO5),
.O6(CLBLM_R_X5Y150_SLICE_X6Y150_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hf5f5a0a0ffbb5511)
  ) CLBLM_R_X5Y150_SLICE_X6Y150_CLUT (
.I0(LIOB33_X0Y61_IOB_X0Y62_I),
.I1(CLBLM_R_X5Y144_SLICE_X6Y144_CQ),
.I2(CLBLM_L_X10Y144_SLICE_X13Y144_A5Q),
.I3(CLBLL_L_X4Y150_SLICE_X4Y150_DO6),
.I4(CLBLM_R_X5Y152_SLICE_X6Y152_B5Q),
.I5(1'b1),
.O5(CLBLM_R_X5Y150_SLICE_X6Y150_CO5),
.O6(CLBLM_R_X5Y150_SLICE_X6Y150_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'ha3aca3acfafa0a0a)
  ) CLBLM_R_X5Y150_SLICE_X6Y150_BLUT (
.I0(CLBLM_R_X5Y150_SLICE_X6Y150_CQ),
.I1(CLBLM_L_X8Y153_SLICE_X10Y153_BQ),
.I2(LIOB33_X0Y61_IOB_X0Y62_I),
.I3(CLBLL_L_X4Y143_SLICE_X4Y143_AQ),
.I4(CLBLM_R_X3Y142_SLICE_X3Y142_AQ),
.I5(1'b1),
.O5(CLBLM_R_X5Y150_SLICE_X6Y150_BO5),
.O6(CLBLM_R_X5Y150_SLICE_X6Y150_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hcfc0cfc0f505fa0a)
  ) CLBLM_R_X5Y150_SLICE_X6Y150_ALUT (
.I0(CLBLM_L_X8Y153_SLICE_X10Y153_DQ),
.I1(CLBLM_R_X5Y150_SLICE_X6Y150_BQ),
.I2(LIOB33_X0Y61_IOB_X0Y62_I),
.I3(CLBLL_L_X2Y145_SLICE_X1Y145_CQ),
.I4(CLBLM_R_X5Y152_SLICE_X6Y152_DQ),
.I5(1'b1),
.O5(CLBLM_R_X5Y150_SLICE_X6Y150_AO5),
.O6(CLBLM_R_X5Y150_SLICE_X6Y150_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y150_SLICE_X7Y150_A5_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_R_X5Y150_SLICE_X7Y150_AO5),
.Q(CLBLM_R_X5Y150_SLICE_X7Y150_A5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y150_SLICE_X7Y150_A_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_R_X5Y150_SLICE_X7Y150_AO6),
.Q(CLBLM_R_X5Y150_SLICE_X7Y150_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h3ff3cffc3ff3cffc)
  ) CLBLM_R_X5Y150_SLICE_X7Y150_DLUT (
.I0(1'b1),
.I1(CLBLM_R_X7Y153_SLICE_X9Y153_AQ),
.I2(CLBLM_R_X3Y149_SLICE_X3Y149_AQ),
.I3(CLBLM_R_X5Y149_SLICE_X7Y149_CQ),
.I4(CLBLM_R_X7Y152_SLICE_X8Y152_DQ),
.I5(1'b1),
.O5(CLBLM_R_X5Y150_SLICE_X7Y150_DO5),
.O6(CLBLM_R_X5Y150_SLICE_X7Y150_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h8400210000840021)
  ) CLBLM_R_X5Y150_SLICE_X7Y150_CLUT (
.I0(CLBLM_R_X5Y154_SLICE_X6Y154_AQ),
.I1(CLBLM_R_X5Y154_SLICE_X6Y154_BQ),
.I2(CLBLM_R_X7Y151_SLICE_X8Y151_CQ),
.I3(CLBLL_L_X4Y153_SLICE_X5Y153_AQ),
.I4(CLBLM_R_X7Y147_SLICE_X9Y147_D5Q),
.I5(CLBLM_R_X5Y149_SLICE_X6Y149_BQ),
.O5(CLBLM_R_X5Y150_SLICE_X7Y150_CO5),
.O6(CLBLM_R_X5Y150_SLICE_X7Y150_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffdfffeffffffff)
  ) CLBLM_R_X5Y150_SLICE_X7Y150_BLUT (
.I0(CLBLL_L_X4Y152_SLICE_X5Y152_A5Q),
.I1(CLBLM_R_X5Y151_SLICE_X7Y151_DO6),
.I2(CLBLM_R_X5Y147_SLICE_X6Y147_DO6),
.I3(CLBLM_R_X5Y150_SLICE_X7Y150_DO6),
.I4(CLBLM_R_X5Y146_SLICE_X6Y146_BQ),
.I5(CLBLM_R_X5Y150_SLICE_X7Y150_CO6),
.O5(CLBLM_R_X5Y150_SLICE_X7Y150_BO5),
.O6(CLBLM_R_X5Y150_SLICE_X7Y150_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hccaaccaaf0fff000)
  ) CLBLM_R_X5Y150_SLICE_X7Y150_ALUT (
.I0(CLBLL_L_X4Y150_SLICE_X4Y150_B5Q),
.I1(CLBLM_R_X5Y149_SLICE_X7Y149_DQ),
.I2(CLBLM_R_X5Y150_SLICE_X7Y150_AQ),
.I3(LIOB33_X0Y61_IOB_X0Y62_I),
.I4(CLBLM_L_X10Y153_SLICE_X13Y153_A5Q),
.I5(1'b1),
.O5(CLBLM_R_X5Y150_SLICE_X7Y150_AO5),
.O6(CLBLM_R_X5Y150_SLICE_X7Y150_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y151_SLICE_X6Y151_C5_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_R_X5Y151_SLICE_X6Y151_CO5),
.Q(CLBLM_R_X5Y151_SLICE_X6Y151_C5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y151_SLICE_X6Y151_A_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_R_X5Y151_SLICE_X6Y151_AO6),
.Q(CLBLM_R_X5Y151_SLICE_X6Y151_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y151_SLICE_X6Y151_B_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_R_X5Y151_SLICE_X6Y151_BO6),
.Q(CLBLM_R_X5Y151_SLICE_X6Y151_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y151_SLICE_X6Y151_C_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_R_X5Y151_SLICE_X6Y151_CO6),
.Q(CLBLM_R_X5Y151_SLICE_X6Y151_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffffffefefefe)
  ) CLBLM_R_X5Y151_SLICE_X6Y151_DLUT (
.I0(CLBLM_R_X5Y149_SLICE_X7Y149_C5Q),
.I1(CLBLM_R_X5Y151_SLICE_X6Y151_CQ),
.I2(CLBLL_L_X4Y144_SLICE_X4Y144_B5Q),
.I3(1'b1),
.I4(1'b1),
.I5(CLBLM_R_X7Y152_SLICE_X8Y152_BQ),
.O5(CLBLM_R_X5Y151_SLICE_X6Y151_DO5),
.O6(CLBLM_R_X5Y151_SLICE_X6Y151_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'haffa0550dd88dd88)
  ) CLBLM_R_X5Y151_SLICE_X6Y151_CLUT (
.I0(LIOB33_X0Y61_IOB_X0Y62_I),
.I1(CLBLM_R_X5Y146_SLICE_X6Y146_B5Q),
.I2(CLBLL_L_X4Y153_SLICE_X4Y153_B5Q),
.I3(CLBLM_R_X3Y151_SLICE_X3Y151_AQ),
.I4(CLBLM_L_X10Y152_SLICE_X12Y152_CQ),
.I5(1'b1),
.O5(CLBLM_R_X5Y151_SLICE_X6Y151_CO5),
.O6(CLBLM_R_X5Y151_SLICE_X6Y151_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hffa800a8ffa800a8)
  ) CLBLM_R_X5Y151_SLICE_X6Y151_BLUT (
.I0(CLBLM_R_X13Y149_SLICE_X18Y149_AO6),
.I1(CLBLM_R_X5Y151_SLICE_X6Y151_BQ),
.I2(CLBLM_R_X7Y147_SLICE_X9Y147_BQ),
.I3(LIOB33_X0Y61_IOB_X0Y62_I),
.I4(CLBLL_L_X2Y146_SLICE_X1Y146_B5Q),
.I5(1'b1),
.O5(CLBLM_R_X5Y151_SLICE_X6Y151_BO5),
.O6(CLBLM_R_X5Y151_SLICE_X6Y151_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f0aaaaf0f0aa00)
  ) CLBLM_R_X5Y151_SLICE_X6Y151_ALUT (
.I0(CLBLM_R_X13Y149_SLICE_X18Y149_AO6),
.I1(1'b1),
.I2(CLBLL_L_X4Y151_SLICE_X5Y151_D5Q),
.I3(CLBLM_R_X5Y151_SLICE_X6Y151_AQ),
.I4(LIOB33_X0Y61_IOB_X0Y62_I),
.I5(CLBLL_L_X4Y145_SLICE_X5Y145_AQ),
.O5(CLBLM_R_X5Y151_SLICE_X6Y151_AO5),
.O6(CLBLM_R_X5Y151_SLICE_X6Y151_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y151_SLICE_X7Y151_B5_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_R_X5Y151_SLICE_X7Y151_BO5),
.Q(CLBLM_R_X5Y151_SLICE_X7Y151_B5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y151_SLICE_X7Y151_A_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_R_X5Y151_SLICE_X7Y151_AO6),
.Q(CLBLM_R_X5Y151_SLICE_X7Y151_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y151_SLICE_X7Y151_B_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_R_X5Y151_SLICE_X7Y151_BO6),
.Q(CLBLM_R_X5Y151_SLICE_X7Y151_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h3f3fcfcff3f3fcfc)
  ) CLBLM_R_X5Y151_SLICE_X7Y151_DLUT (
.I0(1'b1),
.I1(CLBLM_R_X11Y151_SLICE_X15Y151_A5Q),
.I2(CLBLM_R_X7Y151_SLICE_X8Y151_DQ),
.I3(1'b1),
.I4(CLBLL_L_X4Y152_SLICE_X5Y152_AQ),
.I5(CLBLM_R_X3Y152_SLICE_X3Y152_AQ),
.O5(CLBLM_R_X5Y151_SLICE_X7Y151_DO5),
.O6(CLBLM_R_X5Y151_SLICE_X7Y151_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffefefffffefe)
  ) CLBLM_R_X5Y151_SLICE_X7Y151_CLUT (
.I0(CLBLM_R_X5Y148_SLICE_X7Y148_CQ),
.I1(CLBLM_R_X5Y144_SLICE_X6Y144_DQ),
.I2(CLBLL_L_X4Y151_SLICE_X5Y151_B5Q),
.I3(1'b1),
.I4(CLBLM_R_X7Y147_SLICE_X9Y147_AQ),
.I5(1'b1),
.O5(CLBLM_R_X5Y151_SLICE_X7Y151_CO5),
.O6(CLBLM_R_X5Y151_SLICE_X7Y151_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'he4e4e4e4bbee1144)
  ) CLBLM_R_X5Y151_SLICE_X7Y151_BLUT (
.I0(LIOB33_X0Y61_IOB_X0Y62_I),
.I1(CLBLL_L_X4Y151_SLICE_X5Y151_CQ),
.I2(CLBLL_L_X4Y151_SLICE_X4Y151_A5Q),
.I3(CLBLM_R_X7Y144_SLICE_X8Y144_B5Q),
.I4(CLBLM_L_X10Y154_SLICE_X12Y154_AQ),
.I5(1'b1),
.O5(CLBLM_R_X5Y151_SLICE_X7Y151_BO5),
.O6(CLBLM_R_X5Y151_SLICE_X7Y151_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hccfaccafcc50cc05)
  ) CLBLM_R_X5Y151_SLICE_X7Y151_ALUT (
.I0(CLBLM_L_X8Y149_SLICE_X11Y149_AQ),
.I1(CLBLM_R_X7Y145_SLICE_X8Y145_BQ),
.I2(CLBLM_R_X5Y151_SLICE_X7Y151_AQ),
.I3(LIOB33_X0Y61_IOB_X0Y62_I),
.I4(CLBLM_R_X5Y148_SLICE_X6Y148_CO6),
.I5(CLBLL_L_X4Y151_SLICE_X5Y151_D5Q),
.O5(CLBLM_R_X5Y151_SLICE_X7Y151_AO5),
.O6(CLBLM_R_X5Y151_SLICE_X7Y151_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y152_SLICE_X6Y152_B5_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_R_X5Y152_SLICE_X6Y152_BO5),
.Q(CLBLM_R_X5Y152_SLICE_X6Y152_B5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y152_SLICE_X6Y152_A_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_R_X5Y152_SLICE_X6Y152_AO6),
.Q(CLBLM_R_X5Y152_SLICE_X6Y152_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y152_SLICE_X6Y152_B_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_R_X5Y152_SLICE_X6Y152_BO6),
.Q(CLBLM_R_X5Y152_SLICE_X6Y152_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y152_SLICE_X6Y152_C_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_R_X5Y152_SLICE_X6Y152_CO6),
.Q(CLBLM_R_X5Y152_SLICE_X6Y152_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y152_SLICE_X6Y152_D_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_R_X5Y152_SLICE_X6Y152_DO6),
.Q(CLBLM_R_X5Y152_SLICE_X6Y152_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaaaaaaff3cfff0)
  ) CLBLM_R_X5Y152_SLICE_X6Y152_DLUT (
.I0(CLBLM_R_X5Y152_SLICE_X7Y152_AQ),
.I1(CLBLM_R_X5Y152_SLICE_X6Y152_CQ),
.I2(CLBLM_R_X5Y152_SLICE_X6Y152_DQ),
.I3(CLBLM_R_X3Y145_SLICE_X2Y145_CQ),
.I4(CLBLL_L_X4Y148_SLICE_X4Y148_DO6),
.I5(LIOB33_X0Y61_IOB_X0Y62_I),
.O5(CLBLM_R_X5Y152_SLICE_X6Y152_DO5),
.O6(CLBLM_R_X5Y152_SLICE_X6Y152_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaaaaaaff33ffcc)
  ) CLBLM_R_X5Y152_SLICE_X6Y152_CLUT (
.I0(CLBLM_R_X7Y147_SLICE_X9Y147_BQ),
.I1(CLBLM_R_X5Y152_SLICE_X6Y152_CQ),
.I2(1'b1),
.I3(CLBLM_R_X3Y145_SLICE_X2Y145_CQ),
.I4(CLBLL_L_X4Y148_SLICE_X4Y148_DO6),
.I5(LIOB33_X0Y61_IOB_X0Y62_I),
.O5(CLBLM_R_X5Y152_SLICE_X6Y152_CO5),
.O6(CLBLM_R_X5Y152_SLICE_X6Y152_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f0ff00aaaacccc)
  ) CLBLM_R_X5Y152_SLICE_X6Y152_BLUT (
.I0(CLBLL_L_X4Y152_SLICE_X5Y152_A5Q),
.I1(CLBLL_L_X4Y144_SLICE_X4Y144_C5Q),
.I2(CLBLM_R_X7Y153_SLICE_X8Y153_DQ),
.I3(CLBLM_R_X5Y144_SLICE_X7Y144_CQ),
.I4(LIOB33_X0Y61_IOB_X0Y62_I),
.I5(1'b1),
.O5(CLBLM_R_X5Y152_SLICE_X6Y152_BO5),
.O6(CLBLM_R_X5Y152_SLICE_X6Y152_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaaccffaaaac0f0)
  ) CLBLM_R_X5Y152_SLICE_X6Y152_ALUT (
.I0(CLBLM_L_X8Y153_SLICE_X11Y153_AQ),
.I1(CLBLM_L_X10Y145_SLICE_X12Y145_AQ),
.I2(CLBLM_R_X5Y152_SLICE_X6Y152_AQ),
.I3(CLBLM_R_X5Y142_SLICE_X7Y142_BQ),
.I4(LIOB33_X0Y61_IOB_X0Y62_I),
.I5(CLBLM_R_X5Y152_SLICE_X7Y152_CQ),
.O5(CLBLM_R_X5Y152_SLICE_X6Y152_AO5),
.O6(CLBLM_R_X5Y152_SLICE_X6Y152_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y152_SLICE_X7Y152_A5_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_R_X5Y152_SLICE_X7Y152_AO5),
.Q(CLBLM_R_X5Y152_SLICE_X7Y152_A5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y152_SLICE_X7Y152_B5_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_R_X5Y152_SLICE_X7Y152_BO5),
.Q(CLBLM_R_X5Y152_SLICE_X7Y152_B5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "C5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y152_SLICE_X7Y152_C5_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_R_X5Y152_SLICE_X7Y152_CO5),
.Q(CLBLM_R_X5Y152_SLICE_X7Y152_C5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y152_SLICE_X7Y152_A_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_R_X5Y152_SLICE_X7Y152_AO6),
.Q(CLBLM_R_X5Y152_SLICE_X7Y152_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y152_SLICE_X7Y152_B_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_R_X5Y152_SLICE_X7Y152_BO6),
.Q(CLBLM_R_X5Y152_SLICE_X7Y152_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y152_SLICE_X7Y152_C_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_R_X5Y152_SLICE_X7Y152_CO6),
.Q(CLBLM_R_X5Y152_SLICE_X7Y152_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y152_SLICE_X7Y152_D_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_R_X5Y152_SLICE_X7Y152_DO5),
.Q(CLBLM_R_X5Y152_SLICE_X7Y152_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hffaaffaaa3a3a0a0)
  ) CLBLM_R_X5Y152_SLICE_X7Y152_DLUT (
.I0(CLBLM_R_X3Y146_SLICE_X3Y146_AQ),
.I1(CLBLM_R_X5Y151_SLICE_X7Y151_CO6),
.I2(LIOB33_X0Y61_IOB_X0Y62_I),
.I3(CLBLM_R_X7Y153_SLICE_X9Y153_DQ),
.I4(CLBLM_R_X5Y150_SLICE_X6Y150_DO6),
.I5(1'b1),
.O5(CLBLM_R_X5Y152_SLICE_X7Y152_DO5),
.O6(CLBLM_R_X5Y152_SLICE_X7Y152_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaaf0f0ccccff00)
  ) CLBLM_R_X5Y152_SLICE_X7Y152_CLUT (
.I0(CLBLM_L_X8Y152_SLICE_X10Y152_BQ),
.I1(CLBLM_R_X5Y151_SLICE_X7Y151_BQ),
.I2(CLBLM_R_X5Y152_SLICE_X6Y152_CQ),
.I3(CLBLM_R_X5Y152_SLICE_X7Y152_A5Q),
.I4(LIOB33_X0Y61_IOB_X0Y62_I),
.I5(1'b1),
.O5(CLBLM_R_X5Y152_SLICE_X7Y152_CO5),
.O6(CLBLM_R_X5Y152_SLICE_X7Y152_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hffcc3300bb88bb88)
  ) CLBLM_R_X5Y152_SLICE_X7Y152_BLUT (
.I0(CLBLM_R_X5Y151_SLICE_X6Y151_CQ),
.I1(LIOB33_X0Y61_IOB_X0Y62_I),
.I2(1'b1),
.I3(CLBLL_L_X4Y145_SLICE_X5Y145_BQ),
.I4(CLBLM_R_X7Y155_SLICE_X8Y155_A5Q),
.I5(1'b1),
.O5(CLBLM_R_X5Y152_SLICE_X7Y152_BO5),
.O6(CLBLM_R_X5Y152_SLICE_X7Y152_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hbb88bb88c0c0f3f3)
  ) CLBLM_R_X5Y152_SLICE_X7Y152_ALUT (
.I0(CLBLL_L_X4Y146_SLICE_X4Y146_C5Q),
.I1(LIOB33_X0Y61_IOB_X0Y62_I),
.I2(CLBLM_R_X7Y151_SLICE_X8Y151_D5Q),
.I3(CLBLM_R_X5Y149_SLICE_X6Y149_CQ),
.I4(CLBLM_R_X7Y146_SLICE_X8Y146_A5Q),
.I5(1'b1),
.O5(CLBLM_R_X5Y152_SLICE_X7Y152_AO5),
.O6(CLBLM_R_X5Y152_SLICE_X7Y152_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y153_SLICE_X6Y153_A5_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_R_X5Y153_SLICE_X6Y153_AO5),
.Q(CLBLM_R_X5Y153_SLICE_X6Y153_A5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y153_SLICE_X6Y153_B5_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_R_X5Y153_SLICE_X6Y153_BO5),
.Q(CLBLM_R_X5Y153_SLICE_X6Y153_B5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y153_SLICE_X6Y153_D5_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_R_X5Y153_SLICE_X6Y153_DO5),
.Q(CLBLM_R_X5Y153_SLICE_X6Y153_D5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y153_SLICE_X6Y153_A_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_R_X5Y153_SLICE_X6Y153_AO6),
.Q(CLBLM_R_X5Y153_SLICE_X6Y153_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y153_SLICE_X6Y153_B_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_R_X5Y153_SLICE_X6Y153_BO6),
.Q(CLBLM_R_X5Y153_SLICE_X6Y153_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y153_SLICE_X6Y153_C_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_R_X5Y153_SLICE_X6Y153_CO6),
.Q(CLBLM_R_X5Y153_SLICE_X6Y153_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y153_SLICE_X6Y153_D_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_R_X5Y153_SLICE_X6Y153_DO6),
.Q(CLBLM_R_X5Y153_SLICE_X6Y153_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'ha0a0f5f5aa00ff55)
  ) CLBLM_R_X5Y153_SLICE_X6Y153_DLUT (
.I0(LIOB33_X0Y61_IOB_X0Y62_I),
.I1(1'b1),
.I2(CLBLM_L_X8Y153_SLICE_X10Y153_DQ),
.I3(CLBLM_L_X8Y144_SLICE_X11Y144_AQ),
.I4(CLBLL_L_X4Y153_SLICE_X4Y153_A5Q),
.I5(1'b1),
.O5(CLBLM_R_X5Y153_SLICE_X6Y153_DO5),
.O6(CLBLM_R_X5Y153_SLICE_X6Y153_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hccccccccafa0afa0)
  ) CLBLM_R_X5Y153_SLICE_X6Y153_CLUT (
.I0(CLBLM_R_X3Y153_SLICE_X2Y153_AQ),
.I1(CLBLM_R_X3Y147_SLICE_X2Y147_CQ),
.I2(CLBLM_L_X8Y144_SLICE_X10Y144_AQ),
.I3(RIOB33_X105Y105_IOB_X1Y106_I),
.I4(1'b1),
.I5(LIOB33_X0Y61_IOB_X0Y62_I),
.O5(CLBLM_R_X5Y153_SLICE_X6Y153_CO5),
.O6(CLBLM_R_X5Y153_SLICE_X6Y153_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'ha0a0afa0cacacaca)
  ) CLBLM_R_X5Y153_SLICE_X6Y153_BLUT (
.I0(CLBLM_R_X5Y153_SLICE_X6Y153_CQ),
.I1(CLBLM_R_X5Y153_SLICE_X7Y153_CQ),
.I2(LIOB33_X0Y61_IOB_X0Y62_I),
.I3(RIOB33_X105Y131_IOB_X1Y131_I),
.I4(CLBLM_R_X3Y151_SLICE_X2Y151_AQ),
.I5(1'b1),
.O5(CLBLM_R_X5Y153_SLICE_X6Y153_BO5),
.O6(CLBLM_R_X5Y153_SLICE_X6Y153_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hcfc0cfc0fcfc0c0c)
  ) CLBLM_R_X5Y153_SLICE_X6Y153_ALUT (
.I0(1'b1),
.I1(CLBLM_R_X5Y153_SLICE_X6Y153_BQ),
.I2(LIOB33_X0Y61_IOB_X0Y62_I),
.I3(CLBLL_L_X4Y148_SLICE_X5Y148_AQ),
.I4(CLBLM_R_X7Y152_SLICE_X8Y152_BQ),
.I5(1'b1),
.O5(CLBLM_R_X5Y153_SLICE_X6Y153_AO5),
.O6(CLBLM_R_X5Y153_SLICE_X6Y153_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y153_SLICE_X7Y153_A_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_R_X5Y153_SLICE_X7Y153_AO6),
.Q(CLBLM_R_X5Y153_SLICE_X7Y153_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y153_SLICE_X7Y153_B_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_R_X5Y153_SLICE_X7Y153_BO6),
.Q(CLBLM_R_X5Y153_SLICE_X7Y153_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y153_SLICE_X7Y153_C_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_R_X5Y153_SLICE_X7Y153_CO6),
.Q(CLBLM_R_X5Y153_SLICE_X7Y153_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h00dc00cc50505050)
  ) CLBLM_R_X5Y153_SLICE_X7Y153_DLUT (
.I0(CLBLM_R_X5Y148_SLICE_X6Y148_CO6),
.I1(CLBLM_L_X8Y153_SLICE_X10Y153_A5Q),
.I2(CLBLM_R_X5Y151_SLICE_X7Y151_AQ),
.I3(CLBLM_L_X8Y149_SLICE_X11Y149_AQ),
.I4(CLBLM_R_X5Y153_SLICE_X7Y153_AQ),
.I5(1'b1),
.O5(CLBLM_R_X5Y153_SLICE_X7Y153_DO5),
.O6(CLBLM_R_X5Y153_SLICE_X7Y153_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaaff33aaaacc00)
  ) CLBLM_R_X5Y153_SLICE_X7Y153_CLUT (
.I0(CLBLM_L_X12Y151_SLICE_X16Y151_AQ),
.I1(CLBLM_R_X11Y148_SLICE_X15Y148_AO6),
.I2(1'b1),
.I3(CLBLM_R_X5Y153_SLICE_X7Y153_BQ),
.I4(LIOB33_X0Y61_IOB_X0Y62_I),
.I5(CLBLM_R_X5Y153_SLICE_X7Y153_CQ),
.O5(CLBLM_R_X5Y153_SLICE_X7Y153_CO5),
.O6(CLBLM_R_X5Y153_SLICE_X7Y153_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfef00e00fefe0e0e)
  ) CLBLM_R_X5Y153_SLICE_X7Y153_BLUT (
.I0(CLBLM_R_X7Y152_SLICE_X9Y152_CQ),
.I1(CLBLM_R_X5Y153_SLICE_X7Y153_BQ),
.I2(LIOB33_X0Y61_IOB_X0Y62_I),
.I3(CLBLL_L_X4Y147_SLICE_X5Y147_CQ),
.I4(CLBLL_L_X4Y153_SLICE_X4Y153_A5Q),
.I5(CLBLL_L_X4Y142_SLICE_X5Y142_DQ),
.O5(CLBLM_R_X5Y153_SLICE_X7Y153_BO5),
.O6(CLBLM_R_X5Y153_SLICE_X7Y153_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfcfc0c0cf5fa050a)
  ) CLBLM_R_X5Y153_SLICE_X7Y153_ALUT (
.I0(CLBLM_R_X5Y153_SLICE_X7Y153_AQ),
.I1(CLBLM_R_X7Y153_SLICE_X9Y153_D5Q),
.I2(LIOB33_X0Y61_IOB_X0Y62_I),
.I3(CLBLM_R_X5Y153_SLICE_X7Y153_DO5),
.I4(CLBLL_L_X4Y147_SLICE_X4Y147_B5Q),
.I5(CLBLM_L_X8Y149_SLICE_X11Y149_AQ),
.O5(CLBLM_R_X5Y153_SLICE_X7Y153_AO5),
.O6(CLBLM_R_X5Y153_SLICE_X7Y153_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y154_SLICE_X6Y154_A_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_R_X5Y154_SLICE_X6Y154_AO6),
.Q(CLBLM_R_X5Y154_SLICE_X6Y154_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y154_SLICE_X6Y154_B_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_R_X5Y154_SLICE_X6Y154_BO6),
.Q(CLBLM_R_X5Y154_SLICE_X6Y154_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X5Y154_SLICE_X6Y154_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y154_SLICE_X6Y154_DO5),
.O6(CLBLM_R_X5Y154_SLICE_X6Y154_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X5Y154_SLICE_X6Y154_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y154_SLICE_X6Y154_CO5),
.O6(CLBLM_R_X5Y154_SLICE_X6Y154_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf202f808f202f808)
  ) CLBLM_R_X5Y154_SLICE_X6Y154_BLUT (
.I0(CLBLL_L_X2Y150_SLICE_X1Y150_AQ),
.I1(CLBLM_R_X5Y154_SLICE_X6Y154_BQ),
.I2(LIOB33_X0Y61_IOB_X0Y62_I),
.I3(CLBLM_R_X5Y148_SLICE_X7Y148_CQ),
.I4(CLBLL_L_X4Y153_SLICE_X5Y153_BO5),
.I5(1'b1),
.O5(CLBLM_R_X5Y154_SLICE_X6Y154_BO5),
.O6(CLBLM_R_X5Y154_SLICE_X6Y154_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff2a8000002a80)
  ) CLBLM_R_X5Y154_SLICE_X6Y154_ALUT (
.I0(CLBLL_L_X2Y150_SLICE_X1Y150_AQ),
.I1(CLBLM_R_X5Y154_SLICE_X6Y154_BQ),
.I2(CLBLL_L_X4Y153_SLICE_X5Y153_BO5),
.I3(CLBLM_R_X5Y154_SLICE_X6Y154_AQ),
.I4(LIOB33_X0Y61_IOB_X0Y62_I),
.I5(CLBLM_L_X10Y153_SLICE_X12Y153_BQ),
.O5(CLBLM_R_X5Y154_SLICE_X6Y154_AO5),
.O6(CLBLM_R_X5Y154_SLICE_X6Y154_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y154_SLICE_X7Y154_A_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_R_X5Y154_SLICE_X7Y154_AO6),
.Q(CLBLM_R_X5Y154_SLICE_X7Y154_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X5Y154_SLICE_X7Y154_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y154_SLICE_X7Y154_DO5),
.O6(CLBLM_R_X5Y154_SLICE_X7Y154_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X5Y154_SLICE_X7Y154_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y154_SLICE_X7Y154_CO5),
.O6(CLBLM_R_X5Y154_SLICE_X7Y154_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X5Y154_SLICE_X7Y154_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y154_SLICE_X7Y154_BO5),
.O6(CLBLM_R_X5Y154_SLICE_X7Y154_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfd0dfd0dfe0efe0e)
  ) CLBLM_R_X5Y154_SLICE_X7Y154_ALUT (
.I0(CLBLL_L_X4Y150_SLICE_X4Y150_A5Q),
.I1(CLBLM_R_X5Y150_SLICE_X7Y150_BO6),
.I2(LIOB33_X0Y61_IOB_X0Y62_I),
.I3(CLBLM_R_X5Y154_SLICE_X6Y154_BQ),
.I4(1'b1),
.I5(CLBLM_R_X3Y149_SLICE_X2Y149_AQ),
.O5(CLBLM_R_X5Y154_SLICE_X7Y154_AO5),
.O6(CLBLM_R_X5Y154_SLICE_X7Y154_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X7Y141_SLICE_X8Y141_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y141_SLICE_X8Y141_DO5),
.O6(CLBLM_R_X7Y141_SLICE_X8Y141_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X7Y141_SLICE_X8Y141_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y141_SLICE_X8Y141_CO5),
.O6(CLBLM_R_X7Y141_SLICE_X8Y141_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hc000c00000000000)
  ) CLBLM_R_X7Y141_SLICE_X8Y141_BLUT (
.I0(1'b1),
.I1(CLBLM_R_X7Y145_SLICE_X8Y145_AQ),
.I2(CLBLM_R_X3Y151_SLICE_X2Y151_AQ),
.I3(CLBLM_L_X10Y147_SLICE_X12Y147_CO6),
.I4(1'b1),
.I5(RIOB33_SING_X105Y100_IOB_X1Y100_I),
.O5(CLBLM_R_X7Y141_SLICE_X8Y141_BO5),
.O6(CLBLM_R_X7Y141_SLICE_X8Y141_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h777777770c000000)
  ) CLBLM_R_X7Y141_SLICE_X8Y141_ALUT (
.I0(CLBLM_L_X8Y145_SLICE_X11Y145_DQ),
.I1(RIOB33_X105Y131_IOB_X1Y131_I),
.I2(RIOB33_X105Y101_IOB_X1Y102_I),
.I3(CLBLM_L_X10Y147_SLICE_X12Y147_CO6),
.I4(CLBLM_R_X3Y151_SLICE_X2Y151_AQ),
.I5(1'b1),
.O5(CLBLM_R_X7Y141_SLICE_X8Y141_AO5),
.O6(CLBLM_R_X7Y141_SLICE_X8Y141_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y141_SLICE_X9Y141_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y141_SLICE_X9Y141_AO6),
.Q(CLBLM_R_X7Y141_SLICE_X9Y141_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X7Y141_SLICE_X9Y141_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y141_SLICE_X9Y141_DO5),
.O6(CLBLM_R_X7Y141_SLICE_X9Y141_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X7Y141_SLICE_X9Y141_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y141_SLICE_X9Y141_CO5),
.O6(CLBLM_R_X7Y141_SLICE_X9Y141_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X7Y141_SLICE_X9Y141_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y141_SLICE_X9Y141_BO5),
.O6(CLBLM_R_X7Y141_SLICE_X9Y141_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hdf13cf03dd11cc00)
  ) CLBLM_R_X7Y141_SLICE_X9Y141_ALUT (
.I0(CLBLM_R_X7Y141_SLICE_X9Y141_AQ),
.I1(LIOB33_X0Y61_IOB_X0Y62_I),
.I2(CLBLM_R_X7Y141_SLICE_X8Y141_AO6),
.I3(CLBLM_R_X7Y144_SLICE_X9Y144_BQ),
.I4(CLBLM_L_X8Y142_SLICE_X10Y142_DO6),
.I5(CLBLL_L_X4Y151_SLICE_X4Y151_CQ),
.O5(CLBLM_R_X7Y141_SLICE_X9Y141_AO5),
.O6(CLBLM_R_X7Y141_SLICE_X9Y141_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y142_SLICE_X8Y142_C5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y142_SLICE_X8Y142_CO5),
.Q(CLBLM_R_X7Y142_SLICE_X8Y142_C5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y142_SLICE_X8Y142_D5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y142_SLICE_X8Y142_DO5),
.Q(CLBLM_R_X7Y142_SLICE_X8Y142_D5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y142_SLICE_X8Y142_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y142_SLICE_X8Y142_AO6),
.Q(CLBLM_R_X7Y142_SLICE_X8Y142_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y142_SLICE_X8Y142_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y142_SLICE_X8Y142_BO6),
.Q(CLBLM_R_X7Y142_SLICE_X8Y142_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y142_SLICE_X8Y142_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y142_SLICE_X8Y142_CO6),
.Q(CLBLM_R_X7Y142_SLICE_X8Y142_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y142_SLICE_X8Y142_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y142_SLICE_X8Y142_DO6),
.Q(CLBLM_R_X7Y142_SLICE_X8Y142_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hafa0afa0cfc0cfc0)
  ) CLBLM_R_X7Y142_SLICE_X8Y142_DLUT (
.I0(CLBLM_R_X5Y147_SLICE_X7Y147_C5Q),
.I1(CLBLM_R_X7Y142_SLICE_X8Y142_CQ),
.I2(LIOB33_X0Y61_IOB_X0Y62_I),
.I3(CLBLL_L_X4Y149_SLICE_X5Y149_C5Q),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y142_SLICE_X8Y142_DO5),
.O6(CLBLM_R_X7Y142_SLICE_X8Y142_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hdd88dd88eeee4444)
  ) CLBLM_R_X7Y142_SLICE_X8Y142_CLUT (
.I0(LIOB33_X0Y61_IOB_X0Y62_I),
.I1(CLBLM_R_X7Y152_SLICE_X8Y152_D5Q),
.I2(1'b1),
.I3(CLBLM_R_X5Y145_SLICE_X6Y145_D5Q),
.I4(CLBLL_L_X4Y142_SLICE_X4Y142_A5Q),
.I5(1'b1),
.O5(CLBLM_R_X7Y142_SLICE_X8Y142_CO5),
.O6(CLBLM_R_X7Y142_SLICE_X8Y142_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffc000000fc00)
  ) CLBLM_R_X7Y142_SLICE_X8Y142_BLUT (
.I0(1'b1),
.I1(CLBLM_R_X7Y142_SLICE_X8Y142_BQ),
.I2(CLBLM_R_X7Y142_SLICE_X8Y142_AQ),
.I3(CLBLM_R_X13Y149_SLICE_X18Y149_AO6),
.I4(LIOB33_X0Y61_IOB_X0Y62_I),
.I5(CLBLM_R_X5Y143_SLICE_X6Y143_DQ),
.O5(CLBLM_R_X7Y142_SLICE_X8Y142_BO5),
.O6(CLBLM_R_X7Y142_SLICE_X8Y142_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfdfcecfc31302030)
  ) CLBLM_R_X7Y142_SLICE_X8Y142_ALUT (
.I0(CLBLM_L_X8Y147_SLICE_X10Y147_C5Q),
.I1(LIOB33_X0Y61_IOB_X0Y62_I),
.I2(CLBLM_R_X7Y142_SLICE_X8Y142_AQ),
.I3(CLBLM_L_X10Y144_SLICE_X13Y144_CQ),
.I4(CLBLM_R_X5Y150_SLICE_X6Y150_AQ),
.I5(CLBLM_L_X8Y142_SLICE_X10Y142_BQ),
.O5(CLBLM_R_X7Y142_SLICE_X8Y142_AO5),
.O6(CLBLM_R_X7Y142_SLICE_X8Y142_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y142_SLICE_X9Y142_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y142_SLICE_X9Y142_AO6),
.Q(CLBLM_R_X7Y142_SLICE_X9Y142_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y142_SLICE_X9Y142_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y142_SLICE_X9Y142_BO6),
.Q(CLBLM_R_X7Y142_SLICE_X9Y142_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y142_SLICE_X9Y142_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y142_SLICE_X9Y142_CO6),
.Q(CLBLM_R_X7Y142_SLICE_X9Y142_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hbfffbfffffffffff)
  ) CLBLM_R_X7Y142_SLICE_X9Y142_DLUT (
.I0(CLBLM_R_X3Y151_SLICE_X2Y151_AQ),
.I1(CLBLM_R_X7Y145_SLICE_X8Y145_AQ),
.I2(RIOB33_SING_X105Y100_IOB_X1Y100_I),
.I3(RIOB33_X105Y131_IOB_X1Y131_I),
.I4(1'b1),
.I5(RIOB33_X105Y101_IOB_X1Y101_I),
.O5(CLBLM_R_X7Y142_SLICE_X9Y142_DO5),
.O6(CLBLM_R_X7Y142_SLICE_X9Y142_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f0f0f00000aaaa)
  ) CLBLM_R_X7Y142_SLICE_X9Y142_CLUT (
.I0(CLBLM_L_X10Y147_SLICE_X12Y147_CO6),
.I1(1'b1),
.I2(CLBLM_R_X7Y145_SLICE_X8Y145_CQ),
.I3(1'b1),
.I4(CLBLM_R_X7Y142_SLICE_X9Y142_DO6),
.I5(LIOB33_X0Y61_IOB_X0Y62_I),
.O5(CLBLM_R_X7Y142_SLICE_X9Y142_CO5),
.O6(CLBLM_R_X7Y142_SLICE_X9Y142_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf202f202fe0efe0e)
  ) CLBLM_R_X7Y142_SLICE_X9Y142_BLUT (
.I0(RIOB33_X105Y105_IOB_X1Y105_I),
.I1(CLBLM_R_X7Y142_SLICE_X9Y142_BQ),
.I2(LIOB33_X0Y61_IOB_X0Y62_I),
.I3(CLBLM_R_X7Y146_SLICE_X8Y146_BQ),
.I4(1'b1),
.I5(CLBLL_L_X4Y152_SLICE_X4Y152_B5Q),
.O5(CLBLM_R_X7Y142_SLICE_X9Y142_BO5),
.O6(CLBLM_R_X7Y142_SLICE_X9Y142_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'heeecfffc22203330)
  ) CLBLM_R_X7Y142_SLICE_X9Y142_ALUT (
.I0(CLBLL_L_X4Y151_SLICE_X4Y151_BQ),
.I1(LIOB33_X0Y61_IOB_X0Y62_I),
.I2(CLBLM_R_X7Y142_SLICE_X9Y142_AQ),
.I3(CLBLL_L_X4Y143_SLICE_X5Y143_D5Q),
.I4(CLBLM_R_X3Y145_SLICE_X3Y145_D5Q),
.I5(CLBLM_R_X5Y145_SLICE_X6Y145_D5Q),
.O5(CLBLM_R_X7Y142_SLICE_X9Y142_AO5),
.O6(CLBLM_R_X7Y142_SLICE_X9Y142_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y143_SLICE_X8Y143_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y143_SLICE_X8Y143_AO6),
.Q(CLBLM_R_X7Y143_SLICE_X8Y143_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y143_SLICE_X8Y143_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y143_SLICE_X8Y143_BO6),
.Q(CLBLM_R_X7Y143_SLICE_X8Y143_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h7fffffffffffffff)
  ) CLBLM_R_X7Y143_SLICE_X8Y143_DLUT (
.I0(CLBLM_R_X7Y143_SLICE_X9Y143_AQ),
.I1(CLBLM_R_X7Y143_SLICE_X8Y143_AQ),
.I2(CLBLM_L_X10Y144_SLICE_X13Y144_DQ),
.I3(CLBLM_R_X7Y144_SLICE_X8Y144_AQ),
.I4(CLBLM_L_X10Y143_SLICE_X12Y143_BQ),
.I5(CLBLM_L_X8Y143_SLICE_X10Y143_BQ),
.O5(CLBLM_R_X7Y143_SLICE_X8Y143_DO5),
.O6(CLBLM_R_X7Y143_SLICE_X8Y143_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h7fffffff7fff7fff)
  ) CLBLM_R_X7Y143_SLICE_X8Y143_CLUT (
.I0(CLBLM_R_X7Y143_SLICE_X9Y143_AQ),
.I1(CLBLM_L_X10Y143_SLICE_X12Y143_BQ),
.I2(CLBLM_L_X10Y144_SLICE_X13Y144_DQ),
.I3(CLBLM_L_X8Y143_SLICE_X10Y143_BQ),
.I4(CLBLM_R_X7Y144_SLICE_X8Y144_AQ),
.I5(1'b1),
.O5(CLBLM_R_X7Y143_SLICE_X8Y143_CO5),
.O6(CLBLM_R_X7Y143_SLICE_X8Y143_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfaeefaee50445044)
  ) CLBLM_R_X7Y143_SLICE_X8Y143_BLUT (
.I0(LIOB33_X0Y61_IOB_X0Y62_I),
.I1(CLBLM_R_X7Y143_SLICE_X8Y143_BQ),
.I2(CLBLM_R_X3Y143_SLICE_X3Y143_AQ),
.I3(CLBLM_L_X12Y149_SLICE_X17Y149_CO6),
.I4(1'b1),
.I5(CLBLM_R_X7Y144_SLICE_X8Y144_CQ),
.O5(CLBLM_R_X7Y143_SLICE_X8Y143_BO5),
.O6(CLBLM_R_X7Y143_SLICE_X8Y143_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfeba5410efab4501)
  ) CLBLM_R_X7Y143_SLICE_X8Y143_ALUT (
.I0(LIOB33_X0Y61_IOB_X0Y62_I),
.I1(CLBLM_L_X8Y149_SLICE_X11Y149_AQ),
.I2(CLBLM_R_X7Y143_SLICE_X8Y143_AQ),
.I3(CLBLM_L_X10Y146_SLICE_X12Y146_D5Q),
.I4(CLBLL_L_X4Y147_SLICE_X5Y147_B5Q),
.I5(CLBLM_R_X7Y143_SLICE_X8Y143_CO6),
.O5(CLBLM_R_X7Y143_SLICE_X8Y143_AO5),
.O6(CLBLM_R_X7Y143_SLICE_X8Y143_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y143_SLICE_X9Y143_B5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y143_SLICE_X9Y143_BO5),
.Q(CLBLM_R_X7Y143_SLICE_X9Y143_B5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y143_SLICE_X9Y143_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y143_SLICE_X9Y143_AO6),
.Q(CLBLM_R_X7Y143_SLICE_X9Y143_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y143_SLICE_X9Y143_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y143_SLICE_X9Y143_BO6),
.Q(CLBLM_R_X7Y143_SLICE_X9Y143_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y143_SLICE_X9Y143_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y143_SLICE_X9Y143_CO6),
.Q(CLBLM_R_X7Y143_SLICE_X9Y143_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0033003300330033)
  ) CLBLM_R_X7Y143_SLICE_X9Y143_DLUT (
.I0(1'b1),
.I1(CLBLM_L_X8Y142_SLICE_X10Y142_CQ),
.I2(1'b1),
.I3(CLBLM_R_X7Y141_SLICE_X9Y141_AQ),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y143_SLICE_X9Y143_DO5),
.O6(CLBLM_R_X7Y143_SLICE_X9Y143_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hf5f0f5f405000504)
  ) CLBLM_R_X7Y143_SLICE_X9Y143_CLUT (
.I0(CLBLM_R_X11Y146_SLICE_X14Y146_BO6),
.I1(CLBLM_R_X7Y143_SLICE_X9Y143_CQ),
.I2(LIOB33_X0Y61_IOB_X0Y62_I),
.I3(CLBLL_L_X4Y151_SLICE_X4Y151_CQ),
.I4(CLBLM_R_X7Y143_SLICE_X9Y143_DO6),
.I5(CLBLL_L_X2Y146_SLICE_X1Y146_BQ),
.O5(CLBLM_R_X7Y143_SLICE_X9Y143_CO5),
.O6(CLBLM_R_X7Y143_SLICE_X9Y143_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0aaf0aaffcc00cc)
  ) CLBLM_R_X7Y143_SLICE_X9Y143_BLUT (
.I0(CLBLM_R_X7Y144_SLICE_X8Y144_BQ),
.I1(RIOB33_X105Y113_IOB_X1Y113_I),
.I2(CLBLM_R_X5Y143_SLICE_X7Y143_C5Q),
.I3(LIOB33_X0Y61_IOB_X0Y62_I),
.I4(CLBLM_L_X8Y144_SLICE_X10Y144_AQ),
.I5(1'b1),
.O5(CLBLM_R_X7Y143_SLICE_X9Y143_BO5),
.O6(CLBLM_R_X7Y143_SLICE_X9Y143_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'haaccaa0faaccaa0f)
  ) CLBLM_R_X7Y143_SLICE_X9Y143_ALUT (
.I0(CLBLM_R_X7Y151_SLICE_X9Y151_A5Q),
.I1(CLBLM_R_X7Y151_SLICE_X9Y151_CQ),
.I2(CLBLM_R_X7Y143_SLICE_X9Y143_AQ),
.I3(LIOB33_X0Y61_IOB_X0Y62_I),
.I4(CLBLM_L_X8Y149_SLICE_X11Y149_AQ),
.I5(1'b1),
.O5(CLBLM_R_X7Y143_SLICE_X9Y143_AO5),
.O6(CLBLM_R_X7Y143_SLICE_X9Y143_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y144_SLICE_X8Y144_B5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y144_SLICE_X8Y144_BO5),
.Q(CLBLM_R_X7Y144_SLICE_X8Y144_B5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "C5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y144_SLICE_X8Y144_C5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y144_SLICE_X8Y144_CO5),
.Q(CLBLM_R_X7Y144_SLICE_X8Y144_C5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y144_SLICE_X8Y144_D5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y144_SLICE_X8Y144_DO5),
.Q(CLBLM_R_X7Y144_SLICE_X8Y144_D5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y144_SLICE_X8Y144_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y144_SLICE_X8Y144_AO6),
.Q(CLBLM_R_X7Y144_SLICE_X8Y144_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y144_SLICE_X8Y144_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y144_SLICE_X8Y144_BO6),
.Q(CLBLM_R_X7Y144_SLICE_X8Y144_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y144_SLICE_X8Y144_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y144_SLICE_X8Y144_CO6),
.Q(CLBLM_R_X7Y144_SLICE_X8Y144_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y144_SLICE_X8Y144_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y144_SLICE_X8Y144_DO6),
.Q(CLBLM_R_X7Y144_SLICE_X8Y144_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hff003333f0f03333)
  ) CLBLM_R_X7Y144_SLICE_X8Y144_DLUT (
.I0(1'b1),
.I1(CLBLM_L_X10Y149_SLICE_X12Y149_BQ),
.I2(CLBLM_R_X5Y142_SLICE_X6Y142_BQ),
.I3(CLBLM_L_X10Y147_SLICE_X12Y147_BQ),
.I4(LIOB33_X0Y61_IOB_X0Y62_I),
.I5(1'b1),
.O5(CLBLM_R_X7Y144_SLICE_X8Y144_DO5),
.O6(CLBLM_R_X7Y144_SLICE_X8Y144_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0ccf0ccccffcc00)
  ) CLBLM_R_X7Y144_SLICE_X8Y144_CLUT (
.I0(1'b1),
.I1(CLBLL_L_X4Y142_SLICE_X5Y142_CQ),
.I2(CLBLM_R_X7Y144_SLICE_X9Y144_B5Q),
.I3(LIOB33_X0Y61_IOB_X0Y62_I),
.I4(CLBLM_R_X11Y149_SLICE_X15Y149_CO6),
.I5(1'b1),
.O5(CLBLM_R_X7Y144_SLICE_X8Y144_CO5),
.O6(CLBLM_R_X7Y144_SLICE_X8Y144_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hff550055f055f055)
  ) CLBLM_R_X7Y144_SLICE_X8Y144_BLUT (
.I0(CLBLM_R_X3Y146_SLICE_X2Y146_D5Q),
.I1(1'b1),
.I2(CLBLM_R_X7Y144_SLICE_X8Y144_AQ),
.I3(LIOB33_X0Y61_IOB_X0Y62_I),
.I4(CLBLL_L_X4Y147_SLICE_X5Y147_AQ),
.I5(1'b1),
.O5(CLBLM_R_X7Y144_SLICE_X8Y144_BO5),
.O6(CLBLM_R_X7Y144_SLICE_X8Y144_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hff00ff00d8d88d8d)
  ) CLBLM_R_X7Y144_SLICE_X8Y144_ALUT (
.I0(CLBLM_L_X8Y149_SLICE_X11Y149_AQ),
.I1(CLBLM_R_X5Y145_SLICE_X6Y145_C5Q),
.I2(CLBLM_R_X7Y144_SLICE_X8Y144_AQ),
.I3(CLBLM_R_X5Y152_SLICE_X6Y152_CQ),
.I4(CLBLM_R_X7Y143_SLICE_X8Y143_CO5),
.I5(LIOB33_X0Y61_IOB_X0Y62_I),
.O5(CLBLM_R_X7Y144_SLICE_X8Y144_AO5),
.O6(CLBLM_R_X7Y144_SLICE_X8Y144_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y144_SLICE_X9Y144_A5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y144_SLICE_X10Y144_BO5),
.Q(CLBLM_R_X7Y144_SLICE_X9Y144_A5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y144_SLICE_X9Y144_B5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y144_SLICE_X9Y144_BO5),
.Q(CLBLM_R_X7Y144_SLICE_X9Y144_B5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y144_SLICE_X9Y144_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y144_SLICE_X9Y144_AO6),
.Q(CLBLM_R_X7Y144_SLICE_X9Y144_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y144_SLICE_X9Y144_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y144_SLICE_X9Y144_BO6),
.Q(CLBLM_R_X7Y144_SLICE_X9Y144_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h00ee000000220000)
  ) CLBLM_R_X7Y144_SLICE_X9Y144_DLUT (
.I0(CLBLM_R_X5Y146_SLICE_X7Y146_C5Q),
.I1(CLBLM_R_X7Y153_SLICE_X8Y153_A5Q),
.I2(1'b1),
.I3(CLBLM_R_X7Y144_SLICE_X9Y144_CO6),
.I4(CLBLM_R_X7Y144_SLICE_X9Y144_B5Q),
.I5(CLBLM_R_X5Y148_SLICE_X6Y148_BQ),
.O5(CLBLM_R_X7Y144_SLICE_X9Y144_DO5),
.O6(CLBLM_R_X7Y144_SLICE_X9Y144_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffffffffffff7)
  ) CLBLM_R_X7Y144_SLICE_X9Y144_CLUT (
.I0(CLBLM_R_X5Y142_SLICE_X6Y142_D5Q),
.I1(CLBLL_L_X4Y148_SLICE_X4Y148_CQ),
.I2(CLBLM_R_X7Y149_SLICE_X8Y149_AQ),
.I3(CLBLL_L_X4Y147_SLICE_X4Y147_CQ),
.I4(CLBLM_R_X7Y151_SLICE_X8Y151_D5Q),
.I5(CLBLM_L_X10Y146_SLICE_X12Y146_DQ),
.O5(CLBLM_R_X7Y144_SLICE_X9Y144_CO5),
.O6(CLBLM_R_X7Y144_SLICE_X9Y144_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf000f0ffaa00aaff)
  ) CLBLM_R_X7Y144_SLICE_X9Y144_BLUT (
.I0(CLBLL_L_X4Y146_SLICE_X4Y146_BQ),
.I1(1'b1),
.I2(CLBLM_L_X8Y143_SLICE_X10Y143_AQ),
.I3(LIOB33_X0Y61_IOB_X0Y62_I),
.I4(CLBLM_L_X12Y151_SLICE_X16Y151_AQ),
.I5(1'b1),
.O5(CLBLM_R_X7Y144_SLICE_X9Y144_BO5),
.O6(CLBLM_R_X7Y144_SLICE_X9Y144_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffee3322cfce0302)
  ) CLBLM_R_X7Y144_SLICE_X9Y144_ALUT (
.I0(CLBLM_R_X7Y144_SLICE_X9Y144_AQ),
.I1(LIOB33_X0Y61_IOB_X0Y62_I),
.I2(CLBLM_R_X3Y145_SLICE_X3Y145_D5Q),
.I3(CLBLM_R_X5Y144_SLICE_X6Y144_D5Q),
.I4(CLBLM_L_X10Y144_SLICE_X13Y144_C5Q),
.I5(CLBLL_L_X4Y151_SLICE_X4Y151_BQ),
.O5(CLBLM_R_X7Y144_SLICE_X9Y144_AO5),
.O6(CLBLM_R_X7Y144_SLICE_X9Y144_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y145_SLICE_X8Y145_A5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y145_SLICE_X8Y145_AO5),
.Q(CLBLM_R_X7Y145_SLICE_X8Y145_A5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y145_SLICE_X8Y145_B5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y145_SLICE_X8Y145_BO5),
.Q(CLBLM_R_X7Y145_SLICE_X8Y145_B5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "C5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y145_SLICE_X8Y145_C5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y145_SLICE_X8Y145_CO5),
.Q(CLBLM_R_X7Y145_SLICE_X8Y145_C5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y145_SLICE_X8Y145_D5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y145_SLICE_X8Y145_DO5),
.Q(CLBLM_R_X7Y145_SLICE_X8Y145_D5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y145_SLICE_X8Y145_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y145_SLICE_X8Y145_AO6),
.Q(CLBLM_R_X7Y145_SLICE_X8Y145_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y145_SLICE_X8Y145_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y145_SLICE_X8Y145_BO6),
.Q(CLBLM_R_X7Y145_SLICE_X8Y145_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y145_SLICE_X8Y145_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y145_SLICE_X8Y145_CO6),
.Q(CLBLM_R_X7Y145_SLICE_X8Y145_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y145_SLICE_X8Y145_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y145_SLICE_X8Y145_DO6),
.Q(CLBLM_R_X7Y145_SLICE_X8Y145_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hd1e2d1e2eeee2222)
  ) CLBLM_R_X7Y145_SLICE_X8Y145_DLUT (
.I0(CLBLM_R_X5Y145_SLICE_X6Y145_D5Q),
.I1(LIOB33_X0Y61_IOB_X0Y62_I),
.I2(CLBLM_R_X5Y150_SLICE_X7Y150_A5Q),
.I3(CLBLM_R_X7Y144_SLICE_X9Y144_A5Q),
.I4(CLBLM_R_X5Y153_SLICE_X6Y153_D5Q),
.I5(1'b1),
.O5(CLBLM_R_X7Y145_SLICE_X8Y145_DO5),
.O6(CLBLM_R_X7Y145_SLICE_X8Y145_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hc5cac5cafff00f00)
  ) CLBLM_R_X7Y145_SLICE_X8Y145_CLUT (
.I0(CLBLM_L_X8Y153_SLICE_X10Y153_D5Q),
.I1(CLBLL_L_X4Y142_SLICE_X4Y142_CQ),
.I2(LIOB33_X0Y61_IOB_X0Y62_I),
.I3(CLBLM_R_X5Y152_SLICE_X6Y152_DQ),
.I4(CLBLM_R_X5Y147_SLICE_X7Y147_B5Q),
.I5(1'b1),
.O5(CLBLM_R_X7Y145_SLICE_X8Y145_CO5),
.O6(CLBLM_R_X7Y145_SLICE_X8Y145_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0aaf0aaaaccaacc)
  ) CLBLM_R_X7Y145_SLICE_X8Y145_BLUT (
.I0(CLBLM_R_X7Y146_SLICE_X8Y146_DQ),
.I1(CLBLM_L_X8Y152_SLICE_X10Y152_A5Q),
.I2(CLBLM_R_X7Y149_SLICE_X8Y149_AQ),
.I3(LIOB33_X0Y61_IOB_X0Y62_I),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y145_SLICE_X8Y145_BO5),
.O6(CLBLM_R_X7Y145_SLICE_X8Y145_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'heeee22228b888b88)
  ) CLBLM_R_X7Y145_SLICE_X8Y145_ALUT (
.I0(CLBLM_R_X7Y145_SLICE_X8Y145_B5Q),
.I1(LIOB33_X0Y61_IOB_X0Y62_I),
.I2(CLBLL_L_X4Y153_SLICE_X5Y153_A5Q),
.I3(CLBLM_L_X8Y154_SLICE_X10Y154_BO5),
.I4(CLBLL_L_X4Y143_SLICE_X5Y143_D5Q),
.I5(1'b1),
.O5(CLBLM_R_X7Y145_SLICE_X8Y145_AO5),
.O6(CLBLM_R_X7Y145_SLICE_X8Y145_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h3050005030000000)
  ) CLBLM_R_X7Y145_SLICE_X9Y145_DLUT (
.I0(CLBLM_R_X7Y144_SLICE_X9Y144_CO6),
.I1(CLBLM_R_X7Y146_SLICE_X9Y146_CO5),
.I2(CLBLM_R_X7Y144_SLICE_X9Y144_B5Q),
.I3(CLBLM_R_X7Y153_SLICE_X8Y153_A5Q),
.I4(CLBLM_R_X7Y145_SLICE_X8Y145_BQ),
.I5(CLBLM_R_X3Y148_SLICE_X3Y148_C5Q),
.O5(CLBLM_R_X7Y145_SLICE_X9Y145_DO5),
.O6(CLBLM_R_X7Y145_SLICE_X9Y145_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h00400040f0400040)
  ) CLBLM_R_X7Y145_SLICE_X9Y145_CLUT (
.I0(CLBLM_R_X7Y144_SLICE_X9Y144_CO6),
.I1(CLBLM_R_X5Y142_SLICE_X7Y142_A5Q),
.I2(CLBLM_R_X7Y144_SLICE_X9Y144_B5Q),
.I3(CLBLM_R_X7Y153_SLICE_X8Y153_A5Q),
.I4(CLBLM_R_X5Y147_SLICE_X7Y147_B5Q),
.I5(CLBLM_R_X7Y146_SLICE_X9Y146_CO5),
.O5(CLBLM_R_X7Y145_SLICE_X9Y145_CO5),
.O6(CLBLM_R_X7Y145_SLICE_X9Y145_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h202020200000aa00)
  ) CLBLM_R_X7Y145_SLICE_X9Y145_BLUT (
.I0(CLBLM_R_X7Y144_SLICE_X9Y144_B5Q),
.I1(CLBLM_R_X7Y146_SLICE_X9Y146_CO5),
.I2(CLBLM_R_X3Y148_SLICE_X3Y148_BQ),
.I3(CLBLM_R_X7Y146_SLICE_X8Y146_BQ),
.I4(CLBLM_R_X7Y144_SLICE_X9Y144_CO6),
.I5(CLBLM_R_X7Y153_SLICE_X8Y153_A5Q),
.O5(CLBLM_R_X7Y145_SLICE_X9Y145_BO5),
.O6(CLBLM_R_X7Y145_SLICE_X9Y145_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h220022000000a0a0)
  ) CLBLM_R_X7Y145_SLICE_X9Y145_ALUT (
.I0(CLBLM_R_X7Y144_SLICE_X9Y144_B5Q),
.I1(CLBLM_R_X7Y146_SLICE_X9Y146_CO5),
.I2(CLBLM_R_X7Y147_SLICE_X9Y147_DQ),
.I3(CLBLM_R_X5Y141_SLICE_X6Y141_B5Q),
.I4(CLBLM_R_X7Y144_SLICE_X9Y144_CO6),
.I5(CLBLM_R_X7Y153_SLICE_X8Y153_A5Q),
.O5(CLBLM_R_X7Y145_SLICE_X9Y145_AO5),
.O6(CLBLM_R_X7Y145_SLICE_X9Y145_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y146_SLICE_X8Y146_A5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y146_SLICE_X8Y146_AO5),
.Q(CLBLM_R_X7Y146_SLICE_X8Y146_A5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y146_SLICE_X8Y146_B5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y146_SLICE_X8Y146_BO5),
.Q(CLBLM_R_X7Y146_SLICE_X8Y146_B5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "C5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y146_SLICE_X8Y146_C5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y146_SLICE_X8Y146_CO5),
.Q(CLBLM_R_X7Y146_SLICE_X8Y146_C5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y146_SLICE_X8Y146_D5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y146_SLICE_X8Y146_DO5),
.Q(CLBLM_R_X7Y146_SLICE_X8Y146_D5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y146_SLICE_X8Y146_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y146_SLICE_X8Y146_AO6),
.Q(CLBLM_R_X7Y146_SLICE_X8Y146_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y146_SLICE_X8Y146_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y146_SLICE_X8Y146_BO6),
.Q(CLBLM_R_X7Y146_SLICE_X8Y146_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y146_SLICE_X8Y146_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y146_SLICE_X8Y146_CO6),
.Q(CLBLM_R_X7Y146_SLICE_X8Y146_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y146_SLICE_X8Y146_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y146_SLICE_X8Y146_DO6),
.Q(CLBLM_R_X7Y146_SLICE_X8Y146_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hccccff00f0f0aaaa)
  ) CLBLM_R_X7Y146_SLICE_X8Y146_DLUT (
.I0(CLBLM_R_X7Y153_SLICE_X9Y153_A5Q),
.I1(CLBLM_R_X5Y145_SLICE_X7Y145_A5Q),
.I2(CLBLM_R_X7Y145_SLICE_X8Y145_A5Q),
.I3(CLBLM_R_X5Y147_SLICE_X6Y147_B5Q),
.I4(LIOB33_X0Y61_IOB_X0Y62_I),
.I5(1'b1),
.O5(CLBLM_R_X7Y146_SLICE_X8Y146_DO5),
.O6(CLBLM_R_X7Y146_SLICE_X8Y146_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hff00f0f0aaaacccc)
  ) CLBLM_R_X7Y146_SLICE_X8Y146_CLUT (
.I0(CLBLM_R_X7Y147_SLICE_X8Y147_AQ),
.I1(CLBLM_R_X5Y146_SLICE_X7Y146_CQ),
.I2(CLBLL_L_X4Y153_SLICE_X4Y153_AQ),
.I3(CLBLM_R_X5Y140_SLICE_X6Y140_A5Q),
.I4(LIOB33_X0Y61_IOB_X0Y62_I),
.I5(1'b1),
.O5(CLBLM_R_X7Y146_SLICE_X8Y146_CO5),
.O6(CLBLM_R_X7Y146_SLICE_X8Y146_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf5a0f5a0dd88dd88)
  ) CLBLM_R_X7Y146_SLICE_X8Y146_BLUT (
.I0(LIOB33_X0Y61_IOB_X0Y62_I),
.I1(CLBLM_R_X7Y142_SLICE_X8Y142_BQ),
.I2(CLBLM_R_X5Y154_SLICE_X6Y154_AQ),
.I3(CLBLM_L_X10Y149_SLICE_X13Y149_AQ),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y146_SLICE_X8Y146_BO5),
.O6(CLBLM_R_X7Y146_SLICE_X8Y146_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'heeee4444fa50fa50)
  ) CLBLM_R_X7Y146_SLICE_X8Y146_ALUT (
.I0(LIOB33_X0Y61_IOB_X0Y62_I),
.I1(CLBLM_R_X3Y147_SLICE_X2Y147_CQ),
.I2(CLBLM_R_X3Y146_SLICE_X2Y146_C5Q),
.I3(CLBLM_L_X8Y150_SLICE_X10Y150_AQ),
.I4(CLBLM_R_X7Y142_SLICE_X8Y142_AQ),
.I5(1'b1),
.O5(CLBLM_R_X7Y146_SLICE_X8Y146_AO5),
.O6(CLBLM_R_X7Y146_SLICE_X8Y146_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y146_SLICE_X9Y146_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y146_SLICE_X9Y146_AO6),
.Q(CLBLM_R_X7Y146_SLICE_X9Y146_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y146_SLICE_X9Y146_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y146_SLICE_X9Y146_BO6),
.Q(CLBLM_R_X7Y146_SLICE_X9Y146_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffffffffdffff)
  ) CLBLM_R_X7Y146_SLICE_X9Y146_DLUT (
.I0(CLBLM_R_X7Y149_SLICE_X8Y149_AQ),
.I1(CLBLM_L_X10Y146_SLICE_X12Y146_DQ),
.I2(CLBLM_R_X7Y151_SLICE_X8Y151_D5Q),
.I3(CLBLL_L_X4Y147_SLICE_X4Y147_CQ),
.I4(CLBLM_R_X5Y142_SLICE_X6Y142_D5Q),
.I5(CLBLM_R_X11Y146_SLICE_X15Y146_BO6),
.O5(CLBLM_R_X7Y146_SLICE_X9Y146_DO5),
.O6(CLBLM_R_X7Y146_SLICE_X9Y146_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffcfffffffdffff)
  ) CLBLM_R_X7Y146_SLICE_X9Y146_CLUT (
.I0(CLBLM_R_X7Y149_SLICE_X8Y149_AQ),
.I1(CLBLM_L_X10Y146_SLICE_X12Y146_DQ),
.I2(CLBLM_R_X7Y151_SLICE_X8Y151_D5Q),
.I3(CLBLL_L_X4Y147_SLICE_X4Y147_CQ),
.I4(CLBLM_R_X5Y142_SLICE_X6Y142_D5Q),
.I5(1'b1),
.O5(CLBLM_R_X7Y146_SLICE_X9Y146_CO5),
.O6(CLBLM_R_X7Y146_SLICE_X9Y146_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hffee5544afae0504)
  ) CLBLM_R_X7Y146_SLICE_X9Y146_BLUT (
.I0(LIOB33_X0Y61_IOB_X0Y62_I),
.I1(CLBLM_R_X7Y146_SLICE_X9Y146_BQ),
.I2(CLBLL_L_X4Y142_SLICE_X5Y142_DQ),
.I3(CLBLM_R_X5Y152_SLICE_X7Y152_BQ),
.I4(CLBLM_R_X7Y144_SLICE_X8Y144_BQ),
.I5(CLBLL_L_X4Y147_SLICE_X5Y147_CQ),
.O5(CLBLM_R_X7Y146_SLICE_X9Y146_BO5),
.O6(CLBLM_R_X7Y146_SLICE_X9Y146_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hbbb88888bbb8bbb8)
  ) CLBLM_R_X7Y146_SLICE_X9Y146_ALUT (
.I0(CLBLM_R_X7Y143_SLICE_X9Y143_B5Q),
.I1(LIOB33_X0Y61_IOB_X0Y62_I),
.I2(CLBLM_R_X7Y146_SLICE_X9Y146_AQ),
.I3(CLBLM_R_X5Y148_SLICE_X7Y148_C5Q),
.I4(CLBLM_L_X10Y145_SLICE_X12Y145_AQ),
.I5(CLBLM_R_X5Y142_SLICE_X7Y142_BQ),
.O5(CLBLM_R_X7Y146_SLICE_X9Y146_AO5),
.O6(CLBLM_R_X7Y146_SLICE_X9Y146_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y147_SLICE_X8Y147_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(LIOB33_X0Y61_IOB_X0Y62_I),
.D(CLBLL_L_X2Y150_SLICE_X1Y150_AQ),
.Q(CLBLM_R_X7Y147_SLICE_X8Y147_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hbfafbfafbbaabbaa)
  ) CLBLM_R_X7Y147_SLICE_X8Y147_DLUT (
.I0(CLBLM_R_X7Y147_SLICE_X8Y147_CO6),
.I1(CLBLM_R_X11Y147_SLICE_X14Y147_AO6),
.I2(CLBLM_L_X8Y150_SLICE_X11Y150_BO6),
.I3(CLBLM_R_X5Y145_SLICE_X6Y145_CQ),
.I4(1'b1),
.I5(CLBLM_R_X7Y142_SLICE_X8Y142_BQ),
.O5(CLBLM_R_X7Y147_SLICE_X8Y147_DO5),
.O6(CLBLM_R_X7Y147_SLICE_X8Y147_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000c4c400008080)
  ) CLBLM_R_X7Y147_SLICE_X8Y147_CLUT (
.I0(CLBLM_R_X7Y144_SLICE_X9Y144_B5Q),
.I1(CLBLM_R_X7Y153_SLICE_X8Y153_A5Q),
.I2(CLBLM_R_X7Y144_SLICE_X8Y144_B5Q),
.I3(1'b1),
.I4(CLBLM_R_X11Y144_SLICE_X14Y144_AO6),
.I5(CLBLM_R_X5Y144_SLICE_X7Y144_BQ),
.O5(CLBLM_R_X7Y147_SLICE_X8Y147_CO5),
.O6(CLBLM_R_X7Y147_SLICE_X8Y147_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000f00022)
  ) CLBLM_R_X7Y147_SLICE_X8Y147_BLUT (
.I0(CLBLL_L_X4Y144_SLICE_X4Y144_AQ),
.I1(CLBLM_L_X10Y146_SLICE_X13Y146_DO6),
.I2(CLBLM_R_X5Y144_SLICE_X6Y144_BQ),
.I3(CLBLM_R_X7Y153_SLICE_X8Y153_A5Q),
.I4(CLBLM_R_X7Y144_SLICE_X9Y144_B5Q),
.I5(CLBLM_R_X11Y144_SLICE_X14Y144_CO6),
.O5(CLBLM_R_X7Y147_SLICE_X8Y147_BO5),
.O6(CLBLM_R_X7Y147_SLICE_X8Y147_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000001)
  ) CLBLM_R_X7Y147_SLICE_X8Y147_ALUT (
.I0(CLBLM_R_X7Y145_SLICE_X8Y145_DQ),
.I1(CLBLM_L_X8Y145_SLICE_X10Y145_A5Q),
.I2(CLBLM_R_X7Y147_SLICE_X9Y147_C5Q),
.I3(CLBLM_L_X8Y153_SLICE_X10Y153_C5Q),
.I4(CLBLM_R_X7Y145_SLICE_X8Y145_CQ),
.I5(CLBLM_R_X3Y150_SLICE_X3Y150_DQ),
.O5(CLBLM_R_X7Y147_SLICE_X8Y147_AO5),
.O6(CLBLM_R_X7Y147_SLICE_X8Y147_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y147_SLICE_X9Y147_A5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y147_SLICE_X9Y147_AO5),
.Q(CLBLM_R_X7Y147_SLICE_X9Y147_A5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "C5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y147_SLICE_X9Y147_C5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y147_SLICE_X9Y147_CO5),
.Q(CLBLM_R_X7Y147_SLICE_X9Y147_C5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y147_SLICE_X9Y147_D5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y147_SLICE_X9Y147_DO5),
.Q(CLBLM_R_X7Y147_SLICE_X9Y147_D5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y147_SLICE_X9Y147_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y147_SLICE_X9Y147_AO6),
.Q(CLBLM_R_X7Y147_SLICE_X9Y147_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y147_SLICE_X9Y147_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y147_SLICE_X9Y147_BO6),
.Q(CLBLM_R_X7Y147_SLICE_X9Y147_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y147_SLICE_X9Y147_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y147_SLICE_X9Y147_CO6),
.Q(CLBLM_R_X7Y147_SLICE_X9Y147_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y147_SLICE_X9Y147_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y147_SLICE_X9Y147_DO6),
.Q(CLBLM_R_X7Y147_SLICE_X9Y147_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h8b8b8b8bcf03cf03)
  ) CLBLM_R_X7Y147_SLICE_X9Y147_DLUT (
.I0(CLBLM_L_X8Y147_SLICE_X10Y147_AQ),
.I1(LIOB33_X0Y61_IOB_X0Y62_I),
.I2(CLBLM_L_X10Y151_SLICE_X13Y151_AQ),
.I3(CLBLL_L_X4Y149_SLICE_X5Y149_AQ),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y147_SLICE_X9Y147_DO5),
.O6(CLBLM_R_X7Y147_SLICE_X9Y147_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hf5f5a0a0bb11ee44)
  ) CLBLM_R_X7Y147_SLICE_X9Y147_CLUT (
.I0(LIOB33_X0Y61_IOB_X0Y62_I),
.I1(CLBLM_R_X5Y145_SLICE_X6Y145_CQ),
.I2(CLBLM_R_X7Y146_SLICE_X9Y146_BQ),
.I3(CLBLM_L_X8Y146_SLICE_X11Y146_AQ),
.I4(CLBLL_L_X4Y150_SLICE_X4Y150_B5Q),
.I5(1'b1),
.O5(CLBLM_R_X7Y147_SLICE_X9Y147_CO5),
.O6(CLBLM_R_X7Y147_SLICE_X9Y147_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hacafacacaca0acac)
  ) CLBLM_R_X7Y147_SLICE_X9Y147_BLUT (
.I0(CLBLL_L_X4Y151_SLICE_X4Y151_BQ),
.I1(CLBLM_R_X7Y147_SLICE_X9Y147_BQ),
.I2(LIOB33_X0Y61_IOB_X0Y62_I),
.I3(CLBLM_L_X8Y147_SLICE_X10Y147_C5Q),
.I4(CLBLM_L_X10Y144_SLICE_X13Y144_CQ),
.I5(CLBLM_R_X7Y147_SLICE_X9Y147_A5Q),
.O5(CLBLM_R_X7Y147_SLICE_X9Y147_BO5),
.O6(CLBLM_R_X7Y147_SLICE_X9Y147_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hff006666f0f0ff00)
  ) CLBLM_R_X7Y147_SLICE_X9Y147_ALUT (
.I0(CLBLM_R_X3Y145_SLICE_X3Y145_BQ),
.I1(CLBLM_R_X7Y146_SLICE_X8Y146_B5Q),
.I2(CLBLM_R_X3Y146_SLICE_X2Y146_D5Q),
.I3(CLBLM_R_X3Y149_SLICE_X2Y149_BQ),
.I4(LIOB33_X0Y61_IOB_X0Y62_I),
.I5(1'b1),
.O5(CLBLM_R_X7Y147_SLICE_X9Y147_AO5),
.O6(CLBLM_R_X7Y147_SLICE_X9Y147_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y148_SLICE_X8Y148_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(LIOB33_X0Y61_IOB_X0Y62_I),
.D(CLBLM_R_X7Y147_SLICE_X9Y147_AQ),
.Q(CLBLM_R_X7Y148_SLICE_X8Y148_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h7d7d7d7dbebebebe)
  ) CLBLM_R_X7Y148_SLICE_X8Y148_DLUT (
.I0(CLBLM_R_X3Y149_SLICE_X3Y149_AQ),
.I1(CLBLM_R_X5Y144_SLICE_X7Y144_B5Q),
.I2(CLBLL_L_X4Y152_SLICE_X5Y152_A5Q),
.I3(1'b1),
.I4(1'b1),
.I5(CLBLM_R_X7Y144_SLICE_X9Y144_BQ),
.O5(CLBLM_R_X7Y148_SLICE_X8Y148_DO5),
.O6(CLBLM_R_X7Y148_SLICE_X8Y148_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffff4f4f4444)
  ) CLBLM_R_X7Y148_SLICE_X8Y148_CLUT (
.I0(CLBLM_R_X7Y148_SLICE_X8Y148_AO6),
.I1(CLBLM_R_X7Y144_SLICE_X9Y144_A5Q),
.I2(CLBLM_L_X8Y150_SLICE_X11Y150_BO6),
.I3(1'b1),
.I4(CLBLM_R_X5Y142_SLICE_X6Y142_BQ),
.I5(CLBLM_R_X7Y148_SLICE_X8Y148_BO6),
.O5(CLBLM_R_X7Y148_SLICE_X8Y148_CO5),
.O6(CLBLM_R_X7Y148_SLICE_X8Y148_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f2f0f0f0e2f0e0)
  ) CLBLM_R_X7Y148_SLICE_X8Y148_BLUT (
.I0(CLBLM_R_X7Y144_SLICE_X9Y144_B5Q),
.I1(CLBLM_R_X11Y144_SLICE_X14Y144_CO6),
.I2(CLBLM_R_X5Y149_SLICE_X7Y149_BQ),
.I3(CLBLM_R_X7Y153_SLICE_X8Y153_A5Q),
.I4(CLBLM_L_X8Y146_SLICE_X11Y146_C5Q),
.I5(CLBLM_L_X10Y146_SLICE_X13Y146_DO6),
.O5(CLBLM_R_X7Y148_SLICE_X8Y148_BO5),
.O6(CLBLM_R_X7Y148_SLICE_X8Y148_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfff7fffff7ffffff)
  ) CLBLM_R_X7Y148_SLICE_X8Y148_ALUT (
.I0(CLBLM_R_X7Y144_SLICE_X9Y144_B5Q),
.I1(CLBLL_L_X4Y148_SLICE_X4Y148_CQ),
.I2(CLBLM_L_X12Y147_SLICE_X16Y147_DO6),
.I3(CLBLM_R_X7Y153_SLICE_X8Y153_A5Q),
.I4(CLBLM_R_X7Y149_SLICE_X8Y149_AQ),
.I5(1'b1),
.O5(CLBLM_R_X7Y148_SLICE_X8Y148_AO5),
.O6(CLBLM_R_X7Y148_SLICE_X8Y148_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y148_SLICE_X9Y148_A5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y148_SLICE_X9Y148_AO5),
.Q(CLBLM_R_X7Y148_SLICE_X9Y148_A5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "C5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y148_SLICE_X9Y148_C5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y148_SLICE_X9Y148_CO5),
.Q(CLBLM_R_X7Y148_SLICE_X9Y148_C5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y148_SLICE_X9Y148_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y148_SLICE_X9Y148_AO6),
.Q(CLBLM_R_X7Y148_SLICE_X9Y148_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y148_SLICE_X9Y148_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y148_SLICE_X9Y148_BO6),
.Q(CLBLM_R_X7Y148_SLICE_X9Y148_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y148_SLICE_X9Y148_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y148_SLICE_X9Y148_CO6),
.Q(CLBLM_R_X7Y148_SLICE_X9Y148_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h1000100010111000)
  ) CLBLM_R_X7Y148_SLICE_X9Y148_DLUT (
.I0(CLBLM_R_X11Y146_SLICE_X15Y146_BO6),
.I1(CLBLM_R_X7Y146_SLICE_X9Y146_CO6),
.I2(CLBLM_R_X5Y146_SLICE_X7Y146_D5Q),
.I3(CLBLM_R_X7Y149_SLICE_X8Y149_AQ),
.I4(CLBLM_R_X5Y144_SLICE_X7Y144_B5Q),
.I5(CLBLL_L_X4Y148_SLICE_X4Y148_CQ),
.O5(CLBLM_R_X7Y148_SLICE_X9Y148_DO5),
.O6(CLBLM_R_X7Y148_SLICE_X9Y148_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hff00ccccaaaaf0f0)
  ) CLBLM_R_X7Y148_SLICE_X9Y148_CLUT (
.I0(CLBLM_L_X8Y148_SLICE_X10Y148_BQ),
.I1(CLBLM_R_X3Y151_SLICE_X3Y151_BQ),
.I2(CLBLM_R_X5Y152_SLICE_X6Y152_CQ),
.I3(CLBLM_R_X7Y151_SLICE_X9Y151_CQ),
.I4(LIOB33_X0Y61_IOB_X0Y62_I),
.I5(1'b1),
.O5(CLBLM_R_X7Y148_SLICE_X9Y148_CO5),
.O6(CLBLM_R_X7Y148_SLICE_X9Y148_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff0000f0ccf0cc)
  ) CLBLM_R_X7Y148_SLICE_X9Y148_BLUT (
.I0(1'b1),
.I1(CLBLM_R_X7Y148_SLICE_X9Y148_BQ),
.I2(CLBLM_R_X5Y143_SLICE_X7Y143_BQ),
.I3(CLBLM_L_X12Y149_SLICE_X17Y149_CO6),
.I4(CLBLM_L_X8Y148_SLICE_X10Y148_AQ),
.I5(LIOB33_X0Y61_IOB_X0Y62_I),
.O5(CLBLM_R_X7Y148_SLICE_X9Y148_BO5),
.O6(CLBLM_R_X7Y148_SLICE_X9Y148_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hcfcfc0c0ff0ff000)
  ) CLBLM_R_X7Y148_SLICE_X9Y148_ALUT (
.I0(1'b1),
.I1(CLBLM_R_X3Y148_SLICE_X3Y148_BQ),
.I2(LIOB33_X0Y61_IOB_X0Y62_I),
.I3(CLBLM_L_X8Y143_SLICE_X10Y143_CQ),
.I4(CLBLM_L_X10Y149_SLICE_X12Y149_BQ),
.I5(1'b1),
.O5(CLBLM_R_X7Y148_SLICE_X9Y148_AO5),
.O6(CLBLM_R_X7Y148_SLICE_X9Y148_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y149_SLICE_X8Y149_A5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y149_SLICE_X8Y149_AO5),
.Q(CLBLM_R_X7Y149_SLICE_X8Y149_A5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y149_SLICE_X8Y149_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y149_SLICE_X8Y149_AO6),
.Q(CLBLM_R_X7Y149_SLICE_X8Y149_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffff5d0c5d0c)
  ) CLBLM_R_X7Y149_SLICE_X8Y149_DLUT (
.I0(CLBLM_R_X7Y148_SLICE_X8Y148_AO5),
.I1(CLBLL_L_X4Y151_SLICE_X5Y151_AQ),
.I2(CLBLM_R_X13Y149_SLICE_X18Y149_AO6),
.I3(CLBLM_R_X7Y149_SLICE_X8Y149_A5Q),
.I4(1'b1),
.I5(CLBLM_R_X7Y149_SLICE_X8Y149_BO6),
.O5(CLBLM_R_X7Y149_SLICE_X8Y149_DO5),
.O6(CLBLM_R_X7Y149_SLICE_X8Y149_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hfafffefffafafefe)
  ) CLBLM_R_X7Y149_SLICE_X8Y149_CLUT (
.I0(CLBLM_L_X10Y146_SLICE_X13Y146_DO6),
.I1(CLBLM_R_X3Y149_SLICE_X3Y149_D5Q),
.I2(CLBLM_R_X7Y147_SLICE_X8Y147_BO6),
.I3(CLBLM_L_X10Y150_SLICE_X12Y150_BO6),
.I4(CLBLM_R_X7Y148_SLICE_X8Y148_AO6),
.I5(CLBLM_R_X5Y149_SLICE_X7Y149_D5Q),
.O5(CLBLM_R_X7Y149_SLICE_X8Y149_CO5),
.O6(CLBLM_R_X7Y149_SLICE_X8Y149_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h050500c0000000c0)
  ) CLBLM_R_X7Y149_SLICE_X8Y149_BLUT (
.I0(CLBLM_R_X11Y144_SLICE_X14Y144_AO6),
.I1(CLBLM_R_X5Y142_SLICE_X6Y142_CQ),
.I2(CLBLM_R_X7Y144_SLICE_X9Y144_B5Q),
.I3(CLBLM_R_X11Y144_SLICE_X14Y144_CO6),
.I4(CLBLM_R_X7Y153_SLICE_X8Y153_A5Q),
.I5(CLBLM_R_X7Y149_SLICE_X9Y149_CQ),
.O5(CLBLM_R_X7Y149_SLICE_X8Y149_BO5),
.O6(CLBLM_R_X7Y149_SLICE_X8Y149_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hcccc00ffaaaa00ff)
  ) CLBLM_R_X7Y149_SLICE_X8Y149_ALUT (
.I0(CLBLM_R_X5Y152_SLICE_X7Y152_B5Q),
.I1(CLBLM_L_X8Y149_SLICE_X10Y149_AQ),
.I2(1'b1),
.I3(CLBLM_L_X10Y151_SLICE_X13Y151_AQ),
.I4(LIOB33_X0Y61_IOB_X0Y62_I),
.I5(1'b1),
.O5(CLBLM_R_X7Y149_SLICE_X8Y149_AO5),
.O6(CLBLM_R_X7Y149_SLICE_X8Y149_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y149_SLICE_X9Y149_A5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y149_SLICE_X9Y149_AO5),
.Q(CLBLM_R_X7Y149_SLICE_X9Y149_A5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y149_SLICE_X9Y149_B5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y149_SLICE_X9Y149_BO5),
.Q(CLBLM_R_X7Y149_SLICE_X9Y149_B5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "C5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y149_SLICE_X9Y149_C5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y149_SLICE_X9Y149_CO5),
.Q(CLBLM_R_X7Y149_SLICE_X9Y149_C5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y149_SLICE_X9Y149_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y149_SLICE_X9Y149_AO6),
.Q(CLBLM_R_X7Y149_SLICE_X9Y149_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y149_SLICE_X9Y149_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y149_SLICE_X9Y149_BO6),
.Q(CLBLM_R_X7Y149_SLICE_X9Y149_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y149_SLICE_X9Y149_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y149_SLICE_X9Y149_CO6),
.Q(CLBLM_R_X7Y149_SLICE_X9Y149_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h000000000c0a0c0a)
  ) CLBLM_R_X7Y149_SLICE_X9Y149_DLUT (
.I0(CLBLM_R_X7Y148_SLICE_X9Y148_AQ),
.I1(CLBLM_R_X7Y153_SLICE_X8Y153_AQ),
.I2(CLBLM_R_X11Y144_SLICE_X14Y144_AO6),
.I3(CLBLM_R_X7Y144_SLICE_X9Y144_B5Q),
.I4(1'b1),
.I5(CLBLM_R_X7Y153_SLICE_X8Y153_A5Q),
.O5(CLBLM_R_X7Y149_SLICE_X9Y149_DO5),
.O6(CLBLM_R_X7Y149_SLICE_X9Y149_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'ha3a3a3a3f303f303)
  ) CLBLM_R_X7Y149_SLICE_X9Y149_CLUT (
.I0(CLBLM_R_X7Y151_SLICE_X9Y151_C5Q),
.I1(CLBLM_L_X10Y151_SLICE_X13Y151_AQ),
.I2(LIOB33_X0Y61_IOB_X0Y62_I),
.I3(CLBLM_R_X7Y149_SLICE_X9Y149_AQ),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y149_SLICE_X9Y149_CO5),
.O6(CLBLM_R_X7Y149_SLICE_X9Y149_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'haa00ff55888d888d)
  ) CLBLM_R_X7Y149_SLICE_X9Y149_BLUT (
.I0(LIOB33_X0Y61_IOB_X0Y62_I),
.I1(CLBLM_R_X7Y146_SLICE_X8Y146_B5Q),
.I2(CLBLL_L_X4Y150_SLICE_X5Y150_AQ),
.I3(CLBLL_L_X4Y149_SLICE_X5Y149_DQ),
.I4(CLBLM_L_X12Y151_SLICE_X16Y151_AQ),
.I5(1'b1),
.O5(CLBLM_R_X7Y149_SLICE_X9Y149_BO5),
.O6(CLBLM_R_X7Y149_SLICE_X9Y149_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hbb88bb88fcfc3030)
  ) CLBLM_R_X7Y149_SLICE_X9Y149_ALUT (
.I0(CLBLM_R_X7Y149_SLICE_X9Y149_B5Q),
.I1(LIOB33_X0Y61_IOB_X0Y62_I),
.I2(CLBLM_L_X8Y148_SLICE_X11Y148_AQ),
.I3(CLBLM_L_X8Y153_SLICE_X10Y153_AQ),
.I4(CLBLM_R_X7Y149_SLICE_X9Y149_C5Q),
.I5(1'b1),
.O5(CLBLM_R_X7Y149_SLICE_X9Y149_AO5),
.O6(CLBLM_R_X7Y149_SLICE_X9Y149_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y150_SLICE_X8Y150_A_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_R_X7Y150_SLICE_X8Y150_AO6),
.Q(CLBLM_R_X7Y150_SLICE_X8Y150_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0013001100030000)
  ) CLBLM_R_X7Y150_SLICE_X8Y150_DLUT (
.I0(CLBLM_R_X11Y147_SLICE_X15Y147_BO6),
.I1(CLBLM_R_X7Y153_SLICE_X8Y153_A5Q),
.I2(CLBLM_R_X11Y144_SLICE_X14Y144_BO6),
.I3(CLBLM_R_X7Y144_SLICE_X9Y144_B5Q),
.I4(CLBLM_R_X7Y144_SLICE_X8Y144_D5Q),
.I5(CLBLM_R_X3Y151_SLICE_X2Y151_AQ),
.O5(CLBLM_R_X7Y150_SLICE_X8Y150_DO5),
.O6(CLBLM_R_X7Y150_SLICE_X8Y150_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffcc88fffffcf8)
  ) CLBLM_R_X7Y150_SLICE_X8Y150_CLUT (
.I0(CLBLM_R_X7Y153_SLICE_X8Y153_CQ),
.I1(CLBLM_R_X11Y148_SLICE_X15Y148_AO6),
.I2(CLBLM_R_X7Y149_SLICE_X9Y149_A5Q),
.I3(CLBLM_L_X10Y146_SLICE_X13Y146_DO6),
.I4(CLBLM_R_X7Y150_SLICE_X8Y150_DO6),
.I5(CLBLM_L_X10Y150_SLICE_X12Y150_BO6),
.O5(CLBLM_R_X7Y150_SLICE_X8Y150_CO5),
.O6(CLBLM_R_X7Y150_SLICE_X8Y150_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff3f3fffff3333)
  ) CLBLM_R_X7Y150_SLICE_X8Y150_BLUT (
.I0(1'b1),
.I1(CLBLM_R_X5Y143_SLICE_X7Y143_AQ),
.I2(CLBLM_R_X7Y150_SLICE_X8Y150_AQ),
.I3(1'b1),
.I4(CLBLM_R_X7Y143_SLICE_X8Y143_DO6),
.I5(1'b1),
.O5(CLBLM_R_X7Y150_SLICE_X8Y150_BO5),
.O6(CLBLM_R_X7Y150_SLICE_X8Y150_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hccccccccff00a5a5)
  ) CLBLM_R_X7Y150_SLICE_X8Y150_ALUT (
.I0(CLBLM_R_X7Y150_SLICE_X8Y150_BO5),
.I1(CLBLM_L_X10Y151_SLICE_X12Y151_AQ),
.I2(CLBLM_R_X7Y150_SLICE_X8Y150_AQ),
.I3(CLBLM_R_X7Y146_SLICE_X8Y146_D5Q),
.I4(CLBLM_L_X8Y149_SLICE_X11Y149_AQ),
.I5(LIOB33_X0Y61_IOB_X0Y62_I),
.O5(CLBLM_R_X7Y150_SLICE_X8Y150_AO5),
.O6(CLBLM_R_X7Y150_SLICE_X8Y150_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h00cc00ccaaeeaaee)
  ) CLBLM_R_X7Y150_SLICE_X9Y150_DLUT (
.I0(CLBLM_R_X7Y151_SLICE_X8Y151_AQ),
.I1(CLBLL_L_X4Y153_SLICE_X4Y153_B5Q),
.I2(1'b1),
.I3(CLBLM_L_X8Y150_SLICE_X10Y150_BO5),
.I4(1'b1),
.I5(CLBLM_L_X8Y150_SLICE_X11Y150_BO6),
.O5(CLBLM_R_X7Y150_SLICE_X9Y150_DO5),
.O6(CLBLM_R_X7Y150_SLICE_X9Y150_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000540010)
  ) CLBLM_R_X7Y150_SLICE_X9Y150_CLUT (
.I0(CLBLM_R_X11Y146_SLICE_X15Y146_BO6),
.I1(CLBLL_L_X4Y148_SLICE_X4Y148_CQ),
.I2(CLBLM_R_X5Y142_SLICE_X6Y142_DQ),
.I3(CLBLM_L_X12Y147_SLICE_X16Y147_DO6),
.I4(CLBLM_R_X3Y147_SLICE_X3Y147_AQ),
.I5(CLBLM_R_X7Y149_SLICE_X8Y149_AQ),
.O5(CLBLM_R_X7Y150_SLICE_X9Y150_CO5),
.O6(CLBLM_R_X7Y150_SLICE_X9Y150_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffffffff2f22)
  ) CLBLM_R_X7Y150_SLICE_X9Y150_BLUT (
.I0(CLBLM_R_X3Y149_SLICE_X2Y149_C5Q),
.I1(CLBLM_L_X8Y150_SLICE_X10Y150_BO6),
.I2(CLBLM_R_X7Y148_SLICE_X8Y148_AO6),
.I3(CLBLM_R_X7Y149_SLICE_X9Y149_C5Q),
.I4(CLBLM_R_X7Y150_SLICE_X9Y150_AO6),
.I5(CLBLM_L_X10Y146_SLICE_X13Y146_DO6),
.O5(CLBLM_R_X7Y150_SLICE_X9Y150_BO5),
.O6(CLBLM_R_X7Y150_SLICE_X9Y150_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h00aa000004040404)
  ) CLBLM_R_X7Y150_SLICE_X9Y150_ALUT (
.I0(CLBLM_R_X7Y153_SLICE_X8Y153_A5Q),
.I1(CLBLM_R_X3Y150_SLICE_X2Y150_D5Q),
.I2(CLBLM_R_X11Y144_SLICE_X14Y144_AO6),
.I3(CLBLM_R_X11Y144_SLICE_X14Y144_CO6),
.I4(CLBLM_R_X5Y151_SLICE_X6Y151_BQ),
.I5(CLBLM_R_X7Y144_SLICE_X9Y144_B5Q),
.O5(CLBLM_R_X7Y150_SLICE_X9Y150_AO5),
.O6(CLBLM_R_X7Y150_SLICE_X9Y150_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y151_SLICE_X8Y151_C5_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_R_X7Y151_SLICE_X8Y151_CO5),
.Q(CLBLM_R_X7Y151_SLICE_X8Y151_C5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y151_SLICE_X8Y151_D5_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_R_X7Y151_SLICE_X8Y151_DO5),
.Q(CLBLM_R_X7Y151_SLICE_X8Y151_D5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y151_SLICE_X8Y151_A_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_R_X7Y151_SLICE_X8Y151_AO6),
.Q(CLBLM_R_X7Y151_SLICE_X8Y151_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y151_SLICE_X8Y151_B_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_R_X7Y151_SLICE_X8Y151_BO6),
.Q(CLBLM_R_X7Y151_SLICE_X8Y151_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y151_SLICE_X8Y151_C_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_R_X7Y151_SLICE_X8Y151_CO6),
.Q(CLBLM_R_X7Y151_SLICE_X8Y151_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y151_SLICE_X8Y151_D_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_R_X7Y151_SLICE_X8Y151_DO6),
.Q(CLBLM_R_X7Y151_SLICE_X8Y151_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hd8d8d8d8fa50fa50)
  ) CLBLM_R_X7Y151_SLICE_X8Y151_DLUT (
.I0(LIOB33_X0Y61_IOB_X0Y62_I),
.I1(CLBLM_R_X5Y149_SLICE_X7Y149_BQ),
.I2(CLBLM_L_X10Y151_SLICE_X13Y151_A5Q),
.I3(CLBLM_L_X8Y152_SLICE_X10Y152_A5Q),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y151_SLICE_X8Y151_DO5),
.O6(CLBLM_R_X7Y151_SLICE_X8Y151_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaa00fff0f0cccc)
  ) CLBLM_R_X7Y151_SLICE_X8Y151_CLUT (
.I0(CLBLM_R_X3Y147_SLICE_X3Y147_AQ),
.I1(CLBLL_L_X4Y151_SLICE_X5Y151_BQ),
.I2(CLBLM_R_X7Y155_SLICE_X8Y155_AQ),
.I3(CLBLM_R_X3Y146_SLICE_X2Y146_D5Q),
.I4(LIOB33_X0Y61_IOB_X0Y62_I),
.I5(1'b1),
.O5(CLBLM_R_X7Y151_SLICE_X8Y151_CO5),
.O6(CLBLM_R_X7Y151_SLICE_X8Y151_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfafa5050eefa4450)
  ) CLBLM_R_X7Y151_SLICE_X8Y151_BLUT (
.I0(LIOB33_X0Y61_IOB_X0Y62_I),
.I1(CLBLM_R_X7Y151_SLICE_X8Y151_BQ),
.I2(CLBLM_R_X5Y151_SLICE_X6Y151_C5Q),
.I3(CLBLM_R_X3Y145_SLICE_X3Y145_D5Q),
.I4(CLBLL_L_X4Y150_SLICE_X5Y150_AQ),
.I5(CLBLL_L_X4Y151_SLICE_X4Y151_BQ),
.O5(CLBLM_R_X7Y151_SLICE_X8Y151_BO5),
.O6(CLBLM_R_X7Y151_SLICE_X8Y151_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hff00ff00c8c8c8c8)
  ) CLBLM_R_X7Y151_SLICE_X8Y151_ALUT (
.I0(CLBLM_R_X5Y147_SLICE_X7Y147_AQ),
.I1(CLBLM_R_X13Y149_SLICE_X18Y149_AO6),
.I2(CLBLM_R_X7Y151_SLICE_X8Y151_AQ),
.I3(CLBLM_R_X5Y144_SLICE_X7Y144_AQ),
.I4(1'b1),
.I5(LIOB33_X0Y61_IOB_X0Y62_I),
.O5(CLBLM_R_X7Y151_SLICE_X8Y151_AO5),
.O6(CLBLM_R_X7Y151_SLICE_X8Y151_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y151_SLICE_X9Y151_A5_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_R_X7Y152_SLICE_X9Y152_DO5),
.Q(CLBLM_R_X7Y151_SLICE_X9Y151_A5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "C5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y151_SLICE_X9Y151_C5_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_R_X7Y151_SLICE_X9Y151_CO5),
.Q(CLBLM_R_X7Y151_SLICE_X9Y151_C5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y151_SLICE_X9Y151_D5_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_R_X7Y151_SLICE_X9Y151_DO5),
.Q(CLBLM_R_X7Y151_SLICE_X9Y151_D5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y151_SLICE_X9Y151_A_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_R_X7Y151_SLICE_X9Y151_AO6),
.Q(CLBLM_R_X7Y151_SLICE_X9Y151_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y151_SLICE_X9Y151_B_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_R_X7Y151_SLICE_X9Y151_BO6),
.Q(CLBLM_R_X7Y151_SLICE_X9Y151_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y151_SLICE_X9Y151_C_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_R_X7Y151_SLICE_X9Y151_CO6),
.Q(CLBLM_R_X7Y151_SLICE_X9Y151_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y151_SLICE_X9Y151_D_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_R_X7Y151_SLICE_X9Y151_DO6),
.Q(CLBLM_R_X7Y151_SLICE_X9Y151_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hb1b1e4e4fa50fa50)
  ) CLBLM_R_X7Y151_SLICE_X9Y151_DLUT (
.I0(LIOB33_X0Y61_IOB_X0Y62_I),
.I1(CLBLL_L_X4Y151_SLICE_X4Y151_AQ),
.I2(CLBLM_L_X10Y153_SLICE_X12Y153_AQ),
.I3(CLBLL_L_X2Y146_SLICE_X0Y146_DQ),
.I4(CLBLM_R_X7Y149_SLICE_X9Y149_C5Q),
.I5(1'b1),
.O5(CLBLM_R_X7Y151_SLICE_X9Y151_DO5),
.O6(CLBLM_R_X7Y151_SLICE_X9Y151_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hfc30fc30bb88bb88)
  ) CLBLM_R_X7Y151_SLICE_X9Y151_CLUT (
.I0(CLBLM_R_X7Y151_SLICE_X8Y151_AQ),
.I1(LIOB33_X0Y61_IOB_X0Y62_I),
.I2(CLBLM_R_X11Y151_SLICE_X15Y151_AQ),
.I3(CLBLM_R_X3Y150_SLICE_X3Y150_D5Q),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y151_SLICE_X9Y151_CO5),
.O6(CLBLM_R_X7Y151_SLICE_X9Y151_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfdf8f8fd0d08080d)
  ) CLBLM_R_X7Y151_SLICE_X9Y151_BLUT (
.I0(CLBLM_L_X8Y149_SLICE_X11Y149_AQ),
.I1(CLBLM_R_X7Y152_SLICE_X9Y152_C5Q),
.I2(LIOB33_X0Y61_IOB_X0Y62_I),
.I3(CLBLM_R_X7Y150_SLICE_X8Y150_BO6),
.I4(CLBLM_R_X7Y151_SLICE_X9Y151_BQ),
.I5(CLBLM_L_X10Y153_SLICE_X13Y153_CQ),
.O5(CLBLM_R_X7Y151_SLICE_X9Y151_BO5),
.O6(CLBLM_R_X7Y151_SLICE_X9Y151_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff0000ddd0ddd0)
  ) CLBLM_R_X7Y151_SLICE_X9Y151_ALUT (
.I0(CLBLM_R_X7Y142_SLICE_X8Y142_C5Q),
.I1(CLBLM_R_X7Y152_SLICE_X8Y152_D5Q),
.I2(CLBLM_R_X7Y151_SLICE_X9Y151_AQ),
.I3(CLBLL_L_X4Y151_SLICE_X4Y151_C5Q),
.I4(CLBLM_L_X8Y153_SLICE_X10Y153_AQ),
.I5(LIOB33_X0Y61_IOB_X0Y62_I),
.O5(CLBLM_R_X7Y151_SLICE_X9Y151_AO5),
.O6(CLBLM_R_X7Y151_SLICE_X9Y151_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y152_SLICE_X8Y152_B5_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_R_X7Y152_SLICE_X8Y152_BO5),
.Q(CLBLM_R_X7Y152_SLICE_X8Y152_B5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y152_SLICE_X8Y152_D5_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_R_X7Y152_SLICE_X8Y152_DO5),
.Q(CLBLM_R_X7Y152_SLICE_X8Y152_D5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y152_SLICE_X8Y152_A_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_R_X7Y152_SLICE_X8Y152_AO6),
.Q(CLBLM_R_X7Y152_SLICE_X8Y152_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y152_SLICE_X8Y152_B_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_R_X7Y152_SLICE_X8Y152_BO6),
.Q(CLBLM_R_X7Y152_SLICE_X8Y152_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y152_SLICE_X8Y152_C_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_R_X7Y152_SLICE_X8Y152_CO6),
.Q(CLBLM_R_X7Y152_SLICE_X8Y152_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y152_SLICE_X8Y152_D_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_R_X7Y152_SLICE_X8Y152_DO6),
.Q(CLBLM_R_X7Y152_SLICE_X8Y152_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f0aaaaff00cccc)
  ) CLBLM_R_X7Y152_SLICE_X8Y152_DLUT (
.I0(CLBLM_L_X12Y151_SLICE_X16Y151_AQ),
.I1(RIOB33_X105Y111_IOB_X1Y112_I),
.I2(CLBLM_R_X3Y152_SLICE_X3Y152_BQ),
.I3(CLBLM_R_X7Y152_SLICE_X8Y152_AQ),
.I4(LIOB33_X0Y61_IOB_X0Y62_I),
.I5(1'b1),
.O5(CLBLM_R_X7Y152_SLICE_X8Y152_DO5),
.O6(CLBLM_R_X7Y152_SLICE_X8Y152_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hf5a0f5a0e4a0e4a0)
  ) CLBLM_R_X7Y152_SLICE_X8Y152_CLUT (
.I0(LIOB33_X0Y61_IOB_X0Y62_I),
.I1(CLBLM_R_X7Y152_SLICE_X8Y152_CQ),
.I2(CLBLM_R_X7Y153_SLICE_X8Y153_BQ),
.I3(CLBLM_L_X12Y149_SLICE_X17Y149_CO6),
.I4(1'b1),
.I5(CLBLM_R_X7Y152_SLICE_X8Y152_AQ),
.O5(CLBLM_R_X7Y152_SLICE_X8Y152_CO5),
.O6(CLBLM_R_X7Y152_SLICE_X8Y152_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hbe14be14eeee4444)
  ) CLBLM_R_X7Y152_SLICE_X8Y152_BLUT (
.I0(LIOB33_X0Y61_IOB_X0Y62_I),
.I1(CLBLM_R_X3Y151_SLICE_X3Y151_CQ),
.I2(CLBLL_L_X4Y150_SLICE_X4Y150_AQ),
.I3(CLBLL_L_X4Y152_SLICE_X4Y152_B5Q),
.I4(CLBLM_L_X8Y146_SLICE_X10Y146_BQ),
.I5(1'b1),
.O5(CLBLM_R_X7Y152_SLICE_X8Y152_BO5),
.O6(CLBLM_R_X7Y152_SLICE_X8Y152_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hefefefaa45454500)
  ) CLBLM_R_X7Y152_SLICE_X8Y152_ALUT (
.I0(LIOB33_X0Y61_IOB_X0Y62_I),
.I1(CLBLL_L_X4Y151_SLICE_X4Y151_BQ),
.I2(CLBLM_R_X3Y145_SLICE_X3Y145_D5Q),
.I3(CLBLM_R_X7Y152_SLICE_X8Y152_AQ),
.I4(CLBLM_R_X5Y151_SLICE_X7Y151_BQ),
.I5(CLBLM_R_X3Y151_SLICE_X3Y151_CQ),
.O5(CLBLM_R_X7Y152_SLICE_X8Y152_AO5),
.O6(CLBLM_R_X7Y152_SLICE_X8Y152_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y152_SLICE_X9Y152_B5_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_R_X7Y152_SLICE_X9Y152_BO5),
.Q(CLBLM_R_X7Y152_SLICE_X9Y152_B5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "C5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y152_SLICE_X9Y152_C5_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_R_X7Y152_SLICE_X9Y152_CO5),
.Q(CLBLM_R_X7Y152_SLICE_X9Y152_C5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y152_SLICE_X9Y152_A_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_R_X7Y152_SLICE_X9Y152_AO6),
.Q(CLBLM_R_X7Y152_SLICE_X9Y152_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y152_SLICE_X9Y152_B_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_R_X7Y152_SLICE_X9Y152_BO6),
.Q(CLBLM_R_X7Y152_SLICE_X9Y152_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y152_SLICE_X9Y152_C_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_R_X7Y152_SLICE_X9Y152_CO6),
.Q(CLBLM_R_X7Y152_SLICE_X9Y152_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'heeeefffffff00f00)
  ) CLBLM_R_X7Y152_SLICE_X9Y152_DLUT (
.I0(CLBLM_L_X8Y152_SLICE_X10Y152_BQ),
.I1(CLBLM_R_X7Y152_SLICE_X9Y152_AQ),
.I2(LIOB33_X0Y61_IOB_X0Y62_I),
.I3(CLBLL_L_X4Y145_SLICE_X5Y145_C5Q),
.I4(CLBLM_L_X8Y152_SLICE_X10Y152_AQ),
.I5(1'b1),
.O5(CLBLM_R_X7Y152_SLICE_X9Y152_DO5),
.O6(CLBLM_R_X7Y152_SLICE_X9Y152_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hcacacacaff0ff000)
  ) CLBLM_R_X7Y152_SLICE_X9Y152_CLUT (
.I0(CLBLL_L_X4Y143_SLICE_X4Y143_BQ),
.I1(CLBLM_R_X7Y152_SLICE_X9Y152_AQ),
.I2(LIOB33_X0Y61_IOB_X0Y62_I),
.I3(CLBLM_L_X8Y153_SLICE_X10Y153_BQ),
.I4(CLBLM_R_X7Y146_SLICE_X8Y146_C5Q),
.I5(1'b1),
.O5(CLBLM_R_X7Y152_SLICE_X9Y152_CO5),
.O6(CLBLM_R_X7Y152_SLICE_X9Y152_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfa50fa50ffaa5500)
  ) CLBLM_R_X7Y152_SLICE_X9Y152_BLUT (
.I0(LIOB33_X0Y61_IOB_X0Y62_I),
.I1(1'b1),
.I2(CLBLM_R_X5Y152_SLICE_X7Y152_AQ),
.I3(CLBLM_L_X10Y149_SLICE_X12Y149_BQ),
.I4(CLBLM_R_X7Y142_SLICE_X8Y142_D5Q),
.I5(1'b1),
.O5(CLBLM_R_X7Y152_SLICE_X9Y152_BO5),
.O6(CLBLM_R_X7Y152_SLICE_X9Y152_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hcccccccc000f0005)
  ) CLBLM_R_X7Y152_SLICE_X9Y152_ALUT (
.I0(CLBLM_L_X8Y152_SLICE_X10Y152_AQ),
.I1(CLBLL_L_X4Y151_SLICE_X4Y151_C5Q),
.I2(CLBLM_R_X7Y152_SLICE_X9Y152_AQ),
.I3(RIOB33_X105Y131_IOB_X1Y131_I),
.I4(CLBLM_L_X8Y152_SLICE_X10Y152_BQ),
.I5(LIOB33_X0Y61_IOB_X0Y62_I),
.O5(CLBLM_R_X7Y152_SLICE_X9Y152_AO5),
.O6(CLBLM_R_X7Y152_SLICE_X9Y152_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y153_SLICE_X8Y153_A5_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_R_X7Y153_SLICE_X8Y153_AO5),
.Q(CLBLM_R_X7Y153_SLICE_X8Y153_A5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y153_SLICE_X8Y153_A_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_R_X7Y153_SLICE_X8Y153_AO6),
.Q(CLBLM_R_X7Y153_SLICE_X8Y153_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y153_SLICE_X8Y153_B_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_R_X7Y153_SLICE_X8Y153_BO6),
.Q(CLBLM_R_X7Y153_SLICE_X8Y153_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y153_SLICE_X8Y153_C_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_R_X7Y153_SLICE_X8Y153_CO6),
.Q(CLBLM_R_X7Y153_SLICE_X8Y153_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y153_SLICE_X8Y153_D_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_R_X7Y153_SLICE_X8Y153_DO6),
.Q(CLBLM_R_X7Y153_SLICE_X8Y153_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hccccff00ccccf0f0)
  ) CLBLM_R_X7Y153_SLICE_X8Y153_DLUT (
.I0(1'b1),
.I1(CLBLM_R_X7Y147_SLICE_X9Y147_C5Q),
.I2(CLBLM_R_X7Y153_SLICE_X8Y153_DQ),
.I3(CLBLM_R_X7Y153_SLICE_X8Y153_BQ),
.I4(LIOB33_X0Y61_IOB_X0Y62_I),
.I5(CLBLM_R_X11Y148_SLICE_X15Y148_AO6),
.O5(CLBLM_R_X7Y153_SLICE_X8Y153_DO5),
.O6(CLBLM_R_X7Y153_SLICE_X8Y153_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffc540000fc54)
  ) CLBLM_R_X7Y153_SLICE_X8Y153_CLUT (
.I0(CLBLL_L_X4Y142_SLICE_X5Y142_DQ),
.I1(CLBLM_R_X7Y153_SLICE_X8Y153_CQ),
.I2(CLBLM_L_X10Y148_SLICE_X13Y148_C5Q),
.I3(CLBLL_L_X4Y147_SLICE_X5Y147_CQ),
.I4(LIOB33_X0Y61_IOB_X0Y62_I),
.I5(CLBLM_R_X7Y153_SLICE_X8Y153_AQ),
.O5(CLBLM_R_X7Y153_SLICE_X8Y153_CO5),
.O6(CLBLM_R_X7Y153_SLICE_X8Y153_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'he4e4f5f5e4a0f5a0)
  ) CLBLM_R_X7Y153_SLICE_X8Y153_BLUT (
.I0(LIOB33_X0Y61_IOB_X0Y62_I),
.I1(CLBLL_L_X4Y147_SLICE_X5Y147_CQ),
.I2(CLBLM_L_X8Y153_SLICE_X11Y153_BQ),
.I3(CLBLM_R_X5Y147_SLICE_X6Y147_BQ),
.I4(CLBLL_L_X4Y142_SLICE_X5Y142_DQ),
.I5(CLBLM_R_X7Y153_SLICE_X8Y153_BQ),
.O5(CLBLM_R_X7Y153_SLICE_X8Y153_BO5),
.O6(CLBLM_R_X7Y153_SLICE_X8Y153_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hf033f033ff330033)
  ) CLBLM_R_X7Y153_SLICE_X8Y153_ALUT (
.I0(1'b1),
.I1(CLBLM_L_X10Y149_SLICE_X12Y149_BQ),
.I2(CLBLM_R_X7Y148_SLICE_X8Y148_AQ),
.I3(LIOB33_X0Y61_IOB_X0Y62_I),
.I4(CLBLM_R_X3Y153_SLICE_X2Y153_AQ),
.I5(1'b1),
.O5(CLBLM_R_X7Y153_SLICE_X8Y153_AO5),
.O6(CLBLM_R_X7Y153_SLICE_X8Y153_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y153_SLICE_X9Y153_A5_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_R_X7Y153_SLICE_X9Y153_AO5),
.Q(CLBLM_R_X7Y153_SLICE_X9Y153_A5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "C5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y153_SLICE_X9Y153_C5_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_R_X7Y153_SLICE_X9Y153_CO5),
.Q(CLBLM_R_X7Y153_SLICE_X9Y153_C5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y153_SLICE_X9Y153_D5_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_R_X7Y153_SLICE_X9Y153_DO5),
.Q(CLBLM_R_X7Y153_SLICE_X9Y153_D5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y153_SLICE_X9Y153_A_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_R_X7Y153_SLICE_X9Y153_AO6),
.Q(CLBLM_R_X7Y153_SLICE_X9Y153_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y153_SLICE_X9Y153_B_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_R_X7Y153_SLICE_X9Y153_BO6),
.Q(CLBLM_R_X7Y153_SLICE_X9Y153_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y153_SLICE_X9Y153_C_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_R_X7Y153_SLICE_X9Y153_CO6),
.Q(CLBLM_R_X7Y153_SLICE_X9Y153_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y153_SLICE_X9Y153_D_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_R_X7Y153_SLICE_X9Y153_DO6),
.Q(CLBLM_R_X7Y153_SLICE_X9Y153_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hccaaccaaaaf0aaf0)
  ) CLBLM_R_X7Y153_SLICE_X9Y153_DLUT (
.I0(CLBLM_R_X5Y153_SLICE_X6Y153_AQ),
.I1(CLBLM_R_X7Y152_SLICE_X9Y152_B5Q),
.I2(CLBLM_R_X7Y143_SLICE_X9Y143_BQ),
.I3(LIOB33_X0Y61_IOB_X0Y62_I),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y153_SLICE_X9Y153_DO5),
.O6(CLBLM_R_X7Y153_SLICE_X9Y153_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'ha0afafa0cacacaca)
  ) CLBLM_R_X7Y153_SLICE_X9Y153_CLUT (
.I0(CLBLM_R_X7Y151_SLICE_X9Y151_D5Q),
.I1(CLBLM_R_X7Y154_SLICE_X8Y154_AQ),
.I2(LIOB33_X0Y61_IOB_X0Y62_I),
.I3(CLBLL_L_X4Y145_SLICE_X5Y145_BQ),
.I4(CLBLM_R_X7Y149_SLICE_X9Y149_BQ),
.I5(1'b1),
.O5(CLBLM_R_X7Y153_SLICE_X9Y153_CO5),
.O6(CLBLM_R_X7Y153_SLICE_X9Y153_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfafa0a0afcfa0c0a)
  ) CLBLM_R_X7Y153_SLICE_X9Y153_BLUT (
.I0(CLBLM_R_X7Y147_SLICE_X9Y147_CQ),
.I1(CLBLM_R_X7Y153_SLICE_X9Y153_BQ),
.I2(LIOB33_X0Y61_IOB_X0Y62_I),
.I3(CLBLM_R_X3Y145_SLICE_X3Y145_D5Q),
.I4(CLBLM_R_X5Y147_SLICE_X6Y147_AQ),
.I5(CLBLL_L_X4Y151_SLICE_X4Y151_BQ),
.O5(CLBLM_R_X7Y153_SLICE_X9Y153_BO5),
.O6(CLBLM_R_X7Y153_SLICE_X9Y153_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hcc0fcc00f0aaf0aa)
  ) CLBLM_R_X7Y153_SLICE_X9Y153_ALUT (
.I0(CLBLM_L_X10Y151_SLICE_X13Y151_A5Q),
.I1(CLBLM_L_X8Y152_SLICE_X10Y152_CQ),
.I2(CLBLM_R_X7Y153_SLICE_X9Y153_AQ),
.I3(LIOB33_X0Y61_IOB_X0Y62_I),
.I4(CLBLL_L_X2Y150_SLICE_X1Y150_AQ),
.I5(1'b1),
.O5(CLBLM_R_X7Y153_SLICE_X9Y153_AO5),
.O6(CLBLM_R_X7Y153_SLICE_X9Y153_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y154_SLICE_X8Y154_A_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_R_X7Y154_SLICE_X8Y154_AO6),
.Q(CLBLM_R_X7Y154_SLICE_X8Y154_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y154_SLICE_X8Y154_B_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_R_X7Y154_SLICE_X8Y154_BO6),
.Q(CLBLM_R_X7Y154_SLICE_X8Y154_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hf7fff7ffffffffff)
  ) CLBLM_R_X7Y154_SLICE_X8Y154_DLUT (
.I0(CLBLM_R_X7Y155_SLICE_X8Y155_AQ),
.I1(CLBLM_L_X8Y154_SLICE_X10Y154_AQ),
.I2(CLBLM_R_X7Y154_SLICE_X9Y154_DO6),
.I3(CLBLM_R_X7Y154_SLICE_X8Y154_BQ),
.I4(1'b1),
.I5(CLBLM_R_X7Y154_SLICE_X8Y154_AQ),
.O5(CLBLM_R_X7Y154_SLICE_X8Y154_DO5),
.O6(CLBLM_R_X7Y154_SLICE_X8Y154_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h3fffffff0000aaaa)
  ) CLBLM_R_X7Y154_SLICE_X8Y154_CLUT (
.I0(CLBLM_R_X5Y152_SLICE_X6Y152_BQ),
.I1(CLBLM_R_X7Y154_SLICE_X8Y154_AQ),
.I2(CLBLM_L_X8Y154_SLICE_X10Y154_AQ),
.I3(CLBLM_R_X7Y155_SLICE_X8Y155_BO5),
.I4(CLBLM_R_X7Y154_SLICE_X8Y154_DO6),
.I5(1'b1),
.O5(CLBLM_R_X7Y154_SLICE_X8Y154_CO5),
.O6(CLBLM_R_X7Y154_SLICE_X8Y154_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'haaf0aafcaaffaaff)
  ) CLBLM_R_X7Y154_SLICE_X8Y154_BLUT (
.I0(CLBLM_R_X5Y152_SLICE_X7Y152_C5Q),
.I1(CLBLM_R_X7Y154_SLICE_X8Y154_BQ),
.I2(CLBLM_R_X5Y150_SLICE_X6Y150_B5Q),
.I3(LIOB33_X0Y61_IOB_X0Y62_I),
.I4(CLBLM_R_X7Y154_SLICE_X8Y154_CO5),
.I5(CLBLM_R_X7Y154_SLICE_X8Y154_CO6),
.O5(CLBLM_R_X7Y154_SLICE_X8Y154_BO5),
.O6(CLBLM_R_X7Y154_SLICE_X8Y154_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hacafacafafacafac)
  ) CLBLM_R_X7Y154_SLICE_X8Y154_ALUT (
.I0(CLBLM_R_X7Y148_SLICE_X9Y148_A5Q),
.I1(CLBLM_R_X5Y150_SLICE_X6Y150_B5Q),
.I2(LIOB33_X0Y61_IOB_X0Y62_I),
.I3(CLBLM_R_X7Y154_SLICE_X8Y154_AQ),
.I4(1'b1),
.I5(CLBLM_R_X7Y155_SLICE_X8Y155_BO5),
.O5(CLBLM_R_X7Y154_SLICE_X8Y154_AO5),
.O6(CLBLM_R_X7Y154_SLICE_X8Y154_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y154_SLICE_X9Y154_A_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_R_X7Y154_SLICE_X9Y154_AO6),
.Q(CLBLM_R_X7Y154_SLICE_X9Y154_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y154_SLICE_X9Y154_B_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_R_X7Y154_SLICE_X9Y154_BO6),
.Q(CLBLM_R_X7Y154_SLICE_X9Y154_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h7fff7fffffffffff)
  ) CLBLM_R_X7Y154_SLICE_X9Y154_DLUT (
.I0(CLBLM_L_X8Y154_SLICE_X11Y154_AQ),
.I1(CLBLM_R_X7Y154_SLICE_X9Y154_AQ),
.I2(CLBLM_R_X7Y154_SLICE_X9Y154_BQ),
.I3(CLBLM_L_X8Y153_SLICE_X11Y153_AQ),
.I4(1'b1),
.I5(CLBLM_L_X10Y153_SLICE_X12Y153_A5Q),
.O5(CLBLM_R_X7Y154_SLICE_X9Y154_DO5),
.O6(CLBLM_R_X7Y154_SLICE_X9Y154_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h8000000080800000)
  ) CLBLM_R_X7Y154_SLICE_X9Y154_CLUT (
.I0(CLBLM_R_X5Y152_SLICE_X6Y152_BQ),
.I1(CLBLM_L_X10Y153_SLICE_X12Y153_A5Q),
.I2(CLBLM_L_X8Y154_SLICE_X11Y154_AQ),
.I3(CLBLM_R_X7Y154_SLICE_X9Y154_BQ),
.I4(CLBLM_L_X8Y153_SLICE_X11Y153_AQ),
.I5(1'b1),
.O5(CLBLM_R_X7Y154_SLICE_X9Y154_CO5),
.O6(CLBLM_R_X7Y154_SLICE_X9Y154_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf3c0f3f3f3f3f3c0)
  ) CLBLM_R_X7Y154_SLICE_X9Y154_BLUT (
.I0(1'b1),
.I1(LIOB33_X0Y61_IOB_X0Y62_I),
.I2(CLBLL_L_X4Y149_SLICE_X4Y149_AQ),
.I3(CLBLM_R_X5Y150_SLICE_X6Y150_B5Q),
.I4(CLBLM_R_X7Y154_SLICE_X9Y154_CO5),
.I5(CLBLM_R_X7Y154_SLICE_X9Y154_BQ),
.O5(CLBLM_R_X7Y154_SLICE_X9Y154_BO5),
.O6(CLBLM_R_X7Y154_SLICE_X9Y154_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hafafa0afafafafa0)
  ) CLBLM_R_X7Y154_SLICE_X9Y154_ALUT (
.I0(CLBLL_L_X4Y143_SLICE_X4Y143_AQ),
.I1(1'b1),
.I2(LIOB33_X0Y61_IOB_X0Y62_I),
.I3(CLBLM_R_X7Y154_SLICE_X9Y154_AQ),
.I4(CLBLM_R_X5Y150_SLICE_X6Y150_B5Q),
.I5(CLBLM_R_X7Y154_SLICE_X9Y154_CO6),
.O5(CLBLM_R_X7Y154_SLICE_X9Y154_AO5),
.O6(CLBLM_R_X7Y154_SLICE_X9Y154_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y155_SLICE_X8Y155_A5_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_R_X7Y155_SLICE_X8Y155_BO6),
.Q(CLBLM_R_X7Y155_SLICE_X8Y155_A5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y155_SLICE_X8Y155_A_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_R_X7Y155_SLICE_X8Y155_AO6),
.Q(CLBLM_R_X7Y155_SLICE_X8Y155_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X7Y155_SLICE_X8Y155_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y155_SLICE_X8Y155_DO5),
.O6(CLBLM_R_X7Y155_SLICE_X8Y155_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X7Y155_SLICE_X8Y155_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y155_SLICE_X8Y155_CO5),
.O6(CLBLM_R_X7Y155_SLICE_X8Y155_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hffaa5500c0c00000)
  ) CLBLM_R_X7Y155_SLICE_X8Y155_BLUT (
.I0(LIOB33_X0Y61_IOB_X0Y62_I),
.I1(CLBLM_R_X7Y154_SLICE_X9Y154_CO6),
.I2(CLBLM_R_X7Y155_SLICE_X8Y155_AQ),
.I3(CLBLL_L_X4Y153_SLICE_X4Y153_BQ),
.I4(CLBLM_R_X7Y154_SLICE_X9Y154_AQ),
.I5(1'b1),
.O5(CLBLM_R_X7Y155_SLICE_X8Y155_BO5),
.O6(CLBLM_R_X7Y155_SLICE_X8Y155_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hff55ff55be14fa50)
  ) CLBLM_R_X7Y155_SLICE_X8Y155_ALUT (
.I0(LIOB33_X0Y61_IOB_X0Y62_I),
.I1(CLBLM_R_X7Y154_SLICE_X9Y154_CO6),
.I2(CLBLM_R_X7Y155_SLICE_X8Y155_AQ),
.I3(CLBLL_L_X4Y140_SLICE_X4Y140_A5Q),
.I4(CLBLM_R_X7Y154_SLICE_X9Y154_AQ),
.I5(CLBLM_R_X5Y150_SLICE_X6Y150_B5Q),
.O5(CLBLM_R_X7Y155_SLICE_X8Y155_AO5),
.O6(CLBLM_R_X7Y155_SLICE_X8Y155_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X7Y155_SLICE_X9Y155_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y155_SLICE_X9Y155_DO5),
.O6(CLBLM_R_X7Y155_SLICE_X9Y155_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X7Y155_SLICE_X9Y155_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y155_SLICE_X9Y155_CO5),
.O6(CLBLM_R_X7Y155_SLICE_X9Y155_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X7Y155_SLICE_X9Y155_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y155_SLICE_X9Y155_BO5),
.O6(CLBLM_R_X7Y155_SLICE_X9Y155_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X7Y155_SLICE_X9Y155_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y155_SLICE_X9Y155_AO5),
.O6(CLBLM_R_X7Y155_SLICE_X9Y155_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000200000022)
  ) CLBLM_R_X11Y144_SLICE_X14Y144_DLUT (
.I0(CLBLM_R_X5Y142_SLICE_X6Y142_D5Q),
.I1(CLBLL_L_X4Y147_SLICE_X4Y147_CQ),
.I2(CLBLM_R_X7Y149_SLICE_X8Y149_AQ),
.I3(CLBLM_R_X7Y151_SLICE_X8Y151_D5Q),
.I4(CLBLM_L_X10Y146_SLICE_X12Y146_DQ),
.I5(CLBLL_L_X4Y148_SLICE_X4Y148_CQ),
.O5(CLBLM_R_X11Y144_SLICE_X14Y144_DO5),
.O6(CLBLM_R_X11Y144_SLICE_X14Y144_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffffffffffef)
  ) CLBLM_R_X11Y144_SLICE_X14Y144_CLUT (
.I0(CLBLM_R_X5Y142_SLICE_X6Y142_D5Q),
.I1(CLBLL_L_X4Y147_SLICE_X4Y147_CQ),
.I2(CLBLM_R_X7Y149_SLICE_X8Y149_AQ),
.I3(CLBLM_R_X7Y151_SLICE_X8Y151_D5Q),
.I4(CLBLM_L_X10Y146_SLICE_X12Y146_DQ),
.I5(CLBLL_L_X4Y148_SLICE_X4Y148_CQ),
.O5(CLBLM_R_X11Y144_SLICE_X14Y144_CO5),
.O6(CLBLM_R_X11Y144_SLICE_X14Y144_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffffffffffef)
  ) CLBLM_R_X11Y144_SLICE_X14Y144_BLUT (
.I0(CLBLM_L_X10Y146_SLICE_X12Y146_DQ),
.I1(CLBLL_L_X4Y148_SLICE_X4Y148_CQ),
.I2(CLBLM_R_X5Y142_SLICE_X6Y142_D5Q),
.I3(CLBLM_R_X7Y151_SLICE_X8Y151_D5Q),
.I4(CLBLM_R_X7Y149_SLICE_X8Y149_AQ),
.I5(CLBLL_L_X4Y147_SLICE_X4Y147_CQ),
.O5(CLBLM_R_X11Y144_SLICE_X14Y144_BO5),
.O6(CLBLM_R_X11Y144_SLICE_X14Y144_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffffffffbffff)
  ) CLBLM_R_X11Y144_SLICE_X14Y144_ALUT (
.I0(CLBLM_L_X10Y146_SLICE_X12Y146_DQ),
.I1(CLBLM_R_X7Y149_SLICE_X8Y149_AQ),
.I2(CLBLM_R_X5Y142_SLICE_X6Y142_D5Q),
.I3(CLBLM_R_X7Y151_SLICE_X8Y151_D5Q),
.I4(CLBLL_L_X4Y148_SLICE_X4Y148_CQ),
.I5(CLBLL_L_X4Y147_SLICE_X4Y147_CQ),
.O5(CLBLM_R_X11Y144_SLICE_X14Y144_AO5),
.O6(CLBLM_R_X11Y144_SLICE_X14Y144_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X11Y144_SLICE_X15Y144_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X11Y144_SLICE_X15Y144_DO5),
.O6(CLBLM_R_X11Y144_SLICE_X15Y144_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X11Y144_SLICE_X15Y144_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X11Y144_SLICE_X15Y144_CO5),
.O6(CLBLM_R_X11Y144_SLICE_X15Y144_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X11Y144_SLICE_X15Y144_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X11Y144_SLICE_X15Y144_BO5),
.O6(CLBLM_R_X11Y144_SLICE_X15Y144_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X11Y144_SLICE_X15Y144_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X11Y144_SLICE_X15Y144_AO5),
.O6(CLBLM_R_X11Y144_SLICE_X15Y144_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff0000ffff0a0f)
  ) CLBLM_R_X11Y145_SLICE_X14Y145_DLUT (
.I0(CLBLM_R_X11Y146_SLICE_X14Y146_DO6),
.I1(1'b1),
.I2(CLBLM_R_X11Y145_SLICE_X15Y145_BO6),
.I3(CLBLM_L_X12Y145_SLICE_X16Y145_BO6),
.I4(CLBLM_R_X11Y144_SLICE_X14Y144_DO6),
.I5(CLBLM_R_X11Y145_SLICE_X14Y145_BO6),
.O5(CLBLM_R_X11Y145_SLICE_X14Y145_DO5),
.O6(CLBLM_R_X11Y145_SLICE_X14Y145_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h020202020202ff02)
  ) CLBLM_R_X11Y145_SLICE_X14Y145_CLUT (
.I0(CLBLM_R_X5Y144_SLICE_X6Y144_AQ),
.I1(CLBLM_R_X11Y147_SLICE_X14Y147_AO5),
.I2(CLBLM_R_X7Y146_SLICE_X9Y146_CO6),
.I3(LIOB33_X0Y51_IOB_X0Y51_I),
.I4(CLBLM_L_X12Y145_SLICE_X17Y145_DO6),
.I5(CLBLM_R_X11Y146_SLICE_X14Y146_CO5),
.O5(CLBLM_R_X11Y145_SLICE_X14Y145_CO5),
.O6(CLBLM_R_X11Y145_SLICE_X14Y145_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0500050037330500)
  ) CLBLM_R_X11Y145_SLICE_X14Y145_BLUT (
.I0(CLBLM_L_X12Y145_SLICE_X17Y145_CO6),
.I1(CLBLM_L_X12Y145_SLICE_X17Y145_DO6),
.I2(CLBLM_L_X10Y147_SLICE_X12Y147_BO6),
.I3(RIOB33_X105Y135_IOB_X1Y136_I),
.I4(LIOB33_SING_X0Y50_IOB_X0Y50_I),
.I5(CLBLM_R_X11Y146_SLICE_X14Y146_CO5),
.O5(CLBLM_R_X11Y145_SLICE_X14Y145_BO5),
.O6(CLBLM_R_X11Y145_SLICE_X14Y145_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffeeff0f0f0e0f)
  ) CLBLM_R_X11Y145_SLICE_X14Y145_ALUT (
.I0(CLBLM_R_X7Y153_SLICE_X8Y153_A5Q),
.I1(CLBLM_L_X12Y145_SLICE_X17Y145_CO6),
.I2(LIOB33_X0Y51_IOB_X0Y52_I),
.I3(RIOB33_X105Y143_IOB_X1Y144_I),
.I4(CLBLM_R_X7Y144_SLICE_X9Y144_B5Q),
.I5(CLBLM_L_X12Y145_SLICE_X17Y145_AO5),
.O5(CLBLM_R_X11Y145_SLICE_X14Y145_AO5),
.O6(CLBLM_R_X11Y145_SLICE_X14Y145_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y145_SLICE_X15Y145_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y145_SLICE_X15Y145_AO6),
.Q(CLBLM_R_X11Y145_SLICE_X15Y145_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X11Y145_SLICE_X15Y145_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X11Y145_SLICE_X15Y145_DO5),
.O6(CLBLM_R_X11Y145_SLICE_X15Y145_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0fafcfef0fafcfe)
  ) CLBLM_R_X11Y145_SLICE_X15Y145_CLUT (
.I0(CLBLM_R_X5Y141_SLICE_X6Y141_AQ),
.I1(CLBLM_R_X5Y148_SLICE_X6Y148_CQ),
.I2(CLBLM_R_X11Y146_SLICE_X15Y146_BO5),
.I3(CLBLM_L_X12Y146_SLICE_X16Y146_CO6),
.I4(CLBLM_L_X12Y145_SLICE_X16Y145_AO5),
.I5(1'b1),
.O5(CLBLM_R_X11Y145_SLICE_X15Y145_CO5),
.O6(CLBLM_R_X11Y145_SLICE_X15Y145_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000303055007530)
  ) CLBLM_R_X11Y145_SLICE_X15Y145_BLUT (
.I0(CLBLM_R_X7Y146_SLICE_X9Y146_CO6),
.I1(CLBLM_R_X11Y146_SLICE_X15Y146_BO6),
.I2(CLBLM_L_X12Y145_SLICE_X16Y145_AQ),
.I3(CLBLM_R_X11Y145_SLICE_X15Y145_AQ),
.I4(CLBLM_L_X12Y145_SLICE_X17Y145_CO6),
.I5(CLBLM_R_X11Y147_SLICE_X14Y147_AO5),
.O5(CLBLM_R_X11Y145_SLICE_X15Y145_BO5),
.O6(CLBLM_R_X11Y145_SLICE_X15Y145_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'haaccaaf0aaccaaf0)
  ) CLBLM_R_X11Y145_SLICE_X15Y145_ALUT (
.I0(CLBLM_L_X10Y144_SLICE_X13Y144_DQ),
.I1(CLBLM_L_X10Y146_SLICE_X13Y146_BQ),
.I2(CLBLM_R_X11Y145_SLICE_X15Y145_AQ),
.I3(LIOB33_X0Y61_IOB_X0Y62_I),
.I4(CLBLM_R_X11Y146_SLICE_X14Y146_DO6),
.I5(1'b1),
.O5(CLBLM_R_X11Y145_SLICE_X15Y145_AO5),
.O6(CLBLM_R_X11Y145_SLICE_X15Y145_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y146_SLICE_X14Y146_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y146_SLICE_X14Y146_AO6),
.Q(CLBLM_R_X11Y146_SLICE_X14Y146_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000001000)
  ) CLBLM_R_X11Y146_SLICE_X14Y146_DLUT (
.I0(CLBLM_L_X10Y146_SLICE_X13Y146_DO6),
.I1(CLBLM_R_X7Y153_SLICE_X8Y153_A5Q),
.I2(CLBLL_L_X4Y148_SLICE_X4Y148_CQ),
.I3(CLBLM_R_X7Y149_SLICE_X8Y149_AQ),
.I4(CLBLM_R_X7Y146_SLICE_X9Y146_CO6),
.I5(CLBLM_R_X7Y144_SLICE_X9Y144_B5Q),
.O5(CLBLM_R_X11Y146_SLICE_X14Y146_DO5),
.O6(CLBLM_R_X11Y146_SLICE_X14Y146_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffbfffefffefff)
  ) CLBLM_R_X11Y146_SLICE_X14Y146_CLUT (
.I0(CLBLM_R_X7Y149_SLICE_X8Y149_AQ),
.I1(CLBLM_R_X7Y144_SLICE_X9Y144_B5Q),
.I2(CLBLL_L_X4Y148_SLICE_X4Y148_CQ),
.I3(CLBLM_R_X7Y153_SLICE_X8Y153_A5Q),
.I4(CLBLM_R_X7Y146_SLICE_X9Y146_CO6),
.I5(1'b1),
.O5(CLBLM_R_X11Y146_SLICE_X14Y146_CO5),
.O6(CLBLM_R_X11Y146_SLICE_X14Y146_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h3f373f37ff77ff77)
  ) CLBLM_R_X11Y146_SLICE_X14Y146_BLUT (
.I0(CLBLM_L_X8Y142_SLICE_X11Y142_BQ),
.I1(RIOB33_X105Y131_IOB_X1Y131_I),
.I2(CLBLM_L_X8Y145_SLICE_X11Y145_DQ),
.I3(CLBLL_L_X4Y151_SLICE_X4Y151_CQ),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X11Y146_SLICE_X14Y146_BO5),
.O6(CLBLM_R_X11Y146_SLICE_X14Y146_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hd8d8ddddd8d8d8d8)
  ) CLBLM_R_X11Y146_SLICE_X14Y146_ALUT (
.I0(LIOB33_X0Y61_IOB_X0Y62_I),
.I1(CLBLM_L_X10Y147_SLICE_X12Y147_CQ),
.I2(CLBLM_R_X11Y146_SLICE_X14Y146_AQ),
.I3(1'b1),
.I4(CLBLM_L_X10Y146_SLICE_X13Y146_DO5),
.I5(CLBLM_L_X10Y144_SLICE_X13Y144_AQ),
.O5(CLBLM_R_X11Y146_SLICE_X14Y146_AO5),
.O6(CLBLM_R_X11Y146_SLICE_X14Y146_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hff77ff33ff55ff00)
  ) CLBLM_R_X11Y146_SLICE_X15Y146_DLUT (
.I0(CLBLM_L_X12Y145_SLICE_X17Y145_AO5),
.I1(CLBLM_L_X12Y146_SLICE_X16Y146_CO6),
.I2(1'b1),
.I3(CLBLM_R_X13Y146_SLICE_X18Y146_AO5),
.I4(LIOB33_X0Y53_IOB_X0Y53_I),
.I5(CLBLM_L_X8Y146_SLICE_X11Y146_AQ),
.O5(CLBLM_R_X11Y146_SLICE_X15Y146_DO5),
.O6(CLBLM_R_X11Y146_SLICE_X15Y146_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h00000c0c55005d0c)
  ) CLBLM_R_X11Y146_SLICE_X15Y146_CLUT (
.I0(CLBLM_L_X12Y145_SLICE_X17Y145_CO6),
.I1(CLBLM_L_X10Y146_SLICE_X13Y146_AQ),
.I2(CLBLM_R_X11Y147_SLICE_X14Y147_AO5),
.I3(CLBLM_L_X10Y147_SLICE_X12Y147_CQ),
.I4(CLBLM_R_X7Y146_SLICE_X9Y146_CO6),
.I5(CLBLM_R_X11Y146_SLICE_X15Y146_BO6),
.O5(CLBLM_R_X11Y146_SLICE_X15Y146_CO5),
.O6(CLBLM_R_X11Y146_SLICE_X15Y146_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h55ff55ff31002000)
  ) CLBLM_R_X11Y146_SLICE_X15Y146_BLUT (
.I0(CLBLM_R_X7Y153_SLICE_X8Y153_A5Q),
.I1(CLBLM_L_X12Y145_SLICE_X17Y145_CO6),
.I2(CLBLM_L_X8Y146_SLICE_X10Y146_BQ),
.I3(CLBLM_R_X7Y144_SLICE_X9Y144_B5Q),
.I4(CLBLM_R_X5Y152_SLICE_X7Y152_C5Q),
.I5(1'b1),
.O5(CLBLM_R_X11Y146_SLICE_X15Y146_BO5),
.O6(CLBLM_R_X11Y146_SLICE_X15Y146_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h55ff55fffcccf000)
  ) CLBLM_R_X11Y146_SLICE_X15Y146_ALUT (
.I0(CLBLM_R_X7Y146_SLICE_X8Y146_A5Q),
.I1(CLBLM_L_X12Y146_SLICE_X16Y146_BQ),
.I2(CLBLM_L_X8Y146_SLICE_X10Y146_BQ),
.I3(CLBLM_R_X5Y152_SLICE_X7Y152_C5Q),
.I4(RIOB33_X105Y145_IOB_X1Y145_I),
.I5(1'b1),
.O5(CLBLM_R_X11Y146_SLICE_X15Y146_AO5),
.O6(CLBLM_R_X11Y146_SLICE_X15Y146_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h000c000c000c000e)
  ) CLBLM_R_X11Y147_SLICE_X14Y147_DLUT (
.I0(CLBLM_R_X11Y145_SLICE_X14Y145_AO6),
.I1(CLBLM_R_X11Y144_SLICE_X14Y144_DO6),
.I2(CLBLM_L_X10Y148_SLICE_X12Y148_DO6),
.I3(CLBLM_L_X8Y146_SLICE_X10Y146_DO6),
.I4(CLBLM_R_X11Y147_SLICE_X14Y147_BO5),
.I5(CLBLM_R_X11Y145_SLICE_X15Y145_CO6),
.O5(CLBLM_R_X11Y147_SLICE_X14Y147_DO5),
.O6(CLBLM_R_X11Y147_SLICE_X14Y147_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hccccccceccecccee)
  ) CLBLM_R_X11Y147_SLICE_X14Y147_CLUT (
.I0(CLBLM_R_X11Y145_SLICE_X14Y145_AO6),
.I1(CLBLM_R_X11Y144_SLICE_X14Y144_DO6),
.I2(CLBLM_R_X13Y146_SLICE_X18Y146_BO6),
.I3(CLBLM_R_X11Y145_SLICE_X15Y145_CO6),
.I4(CLBLM_R_X3Y146_SLICE_X2Y146_AQ),
.I5(CLBLM_L_X12Y145_SLICE_X16Y145_BO6),
.O5(CLBLM_R_X11Y147_SLICE_X14Y147_CO5),
.O6(CLBLM_R_X11Y147_SLICE_X14Y147_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfa0afa0afc0cfc0c)
  ) CLBLM_R_X11Y147_SLICE_X14Y147_BLUT (
.I0(CLBLM_L_X10Y148_SLICE_X13Y148_AQ),
.I1(CLBLM_R_X3Y146_SLICE_X2Y146_AQ),
.I2(CLBLM_R_X13Y146_SLICE_X18Y146_BO6),
.I3(CLBLM_L_X12Y145_SLICE_X16Y145_BO6),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X11Y147_SLICE_X14Y147_BO5),
.O6(CLBLM_R_X11Y147_SLICE_X14Y147_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffefffafafffff)
  ) CLBLM_R_X11Y147_SLICE_X14Y147_ALUT (
.I0(CLBLM_R_X7Y153_SLICE_X8Y153_A5Q),
.I1(CLBLM_L_X12Y147_SLICE_X16Y147_DO6),
.I2(CLBLM_R_X7Y149_SLICE_X8Y149_AQ),
.I3(CLBLL_L_X4Y148_SLICE_X4Y148_CQ),
.I4(CLBLM_R_X7Y144_SLICE_X9Y144_B5Q),
.I5(1'b1),
.O5(CLBLM_R_X11Y147_SLICE_X14Y147_AO5),
.O6(CLBLM_R_X11Y147_SLICE_X14Y147_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff0000ffff5151)
  ) CLBLM_R_X11Y147_SLICE_X15Y147_DLUT (
.I0(CLBLM_L_X12Y147_SLICE_X16Y147_AO6),
.I1(CLBLM_L_X12Y145_SLICE_X16Y145_BO6),
.I2(CLBLM_R_X11Y146_SLICE_X14Y146_DO6),
.I3(1'b1),
.I4(CLBLM_R_X11Y144_SLICE_X14Y144_DO6),
.I5(CLBLM_R_X11Y145_SLICE_X14Y145_CO6),
.O5(CLBLM_R_X11Y147_SLICE_X15Y147_DO5),
.O6(CLBLM_R_X11Y147_SLICE_X15Y147_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h000000000f0f0100)
  ) CLBLM_R_X11Y147_SLICE_X15Y147_CLUT (
.I0(CLBLM_R_X11Y147_SLICE_X14Y147_BO6),
.I1(CLBLM_R_X11Y146_SLICE_X15Y146_DO6),
.I2(CLBLM_L_X8Y146_SLICE_X10Y146_BO5),
.I3(CLBLM_L_X12Y146_SLICE_X17Y146_DO6),
.I4(CLBLM_R_X11Y144_SLICE_X14Y144_DO6),
.I5(CLBLM_L_X8Y146_SLICE_X10Y146_CO6),
.O5(CLBLM_R_X11Y147_SLICE_X15Y147_CO5),
.O6(CLBLM_R_X11Y147_SLICE_X15Y147_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffffffffffffe)
  ) CLBLM_R_X11Y147_SLICE_X15Y147_BLUT (
.I0(CLBLL_L_X4Y147_SLICE_X4Y147_CQ),
.I1(CLBLM_R_X7Y151_SLICE_X8Y151_D5Q),
.I2(CLBLM_R_X5Y142_SLICE_X6Y142_D5Q),
.I3(CLBLL_L_X4Y148_SLICE_X4Y148_CQ),
.I4(CLBLM_R_X7Y149_SLICE_X8Y149_AQ),
.I5(CLBLM_L_X10Y146_SLICE_X12Y146_DQ),
.O5(CLBLM_R_X11Y147_SLICE_X15Y147_BO5),
.O6(CLBLM_R_X11Y147_SLICE_X15Y147_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f0f1f0f3f0f1f0)
  ) CLBLM_R_X11Y147_SLICE_X15Y147_ALUT (
.I0(CLBLM_L_X10Y148_SLICE_X13Y148_AQ),
.I1(CLBLM_R_X11Y146_SLICE_X15Y146_DO6),
.I2(CLBLM_R_X11Y144_SLICE_X14Y144_DO6),
.I3(CLBLM_L_X12Y146_SLICE_X17Y146_DO6),
.I4(CLBLM_R_X13Y146_SLICE_X18Y146_BO6),
.I5(CLBLM_L_X12Y145_SLICE_X16Y145_BO6),
.O5(CLBLM_R_X11Y147_SLICE_X15Y147_AO5),
.O6(CLBLM_R_X11Y147_SLICE_X15Y147_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000ffff0000028a)
  ) CLBLM_R_X11Y148_SLICE_X14Y148_DLUT (
.I0(CLBLM_L_X12Y148_SLICE_X16Y148_BO6),
.I1(CLBLM_R_X13Y146_SLICE_X18Y146_BO6),
.I2(CLBLM_L_X10Y151_SLICE_X12Y151_AQ),
.I3(CLBLM_L_X12Y145_SLICE_X16Y145_BO6),
.I4(CLBLM_L_X8Y148_SLICE_X10Y148_CO6),
.I5(CLBLM_R_X11Y144_SLICE_X14Y144_DO6),
.O5(CLBLM_R_X11Y148_SLICE_X14Y148_DO5),
.O6(CLBLM_R_X11Y148_SLICE_X14Y148_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000ffff00002700)
  ) CLBLM_R_X11Y148_SLICE_X14Y148_CLUT (
.I0(CLBLM_R_X13Y146_SLICE_X18Y146_BO6),
.I1(CLBLM_L_X12Y145_SLICE_X16Y145_BO6),
.I2(CLBLM_R_X3Y145_SLICE_X2Y145_AQ),
.I3(CLBLM_L_X12Y147_SLICE_X17Y147_BO6),
.I4(CLBLM_L_X10Y147_SLICE_X12Y147_DO6),
.I5(CLBLM_R_X11Y144_SLICE_X14Y144_DO6),
.O5(CLBLM_R_X11Y148_SLICE_X14Y148_CO5),
.O6(CLBLM_R_X11Y148_SLICE_X14Y148_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0111011101110011)
  ) CLBLM_R_X11Y148_SLICE_X14Y148_BLUT (
.I0(CLBLM_L_X10Y148_SLICE_X12Y148_CO6),
.I1(CLBLM_L_X8Y148_SLICE_X10Y148_DO6),
.I2(CLBLM_L_X10Y145_SLICE_X12Y145_DO6),
.I3(CLBLM_L_X12Y147_SLICE_X16Y147_DO6),
.I4(CLBLM_L_X12Y146_SLICE_X16Y146_DO6),
.I5(CLBLM_R_X11Y144_SLICE_X14Y144_DO6),
.O5(CLBLM_R_X11Y148_SLICE_X14Y148_BO5),
.O6(CLBLM_R_X11Y148_SLICE_X14Y148_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffffffefeeee)
  ) CLBLM_R_X11Y148_SLICE_X14Y148_ALUT (
.I0(CLBLM_R_X7Y147_SLICE_X8Y147_DO6),
.I1(CLBLM_R_X11Y150_SLICE_X15Y150_AO6),
.I2(CLBLM_R_X11Y148_SLICE_X15Y148_CO6),
.I3(CLBLM_L_X8Y148_SLICE_X10Y148_CO6),
.I4(CLBLM_L_X12Y147_SLICE_X16Y147_DO6),
.I5(CLBLM_R_X7Y149_SLICE_X8Y149_CO6),
.O5(CLBLM_R_X11Y148_SLICE_X14Y148_AO5),
.O6(CLBLM_R_X11Y148_SLICE_X14Y148_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hff44ff44ff440cb7)
  ) CLBLM_R_X11Y148_SLICE_X15Y148_DLUT (
.I0(CLBLM_R_X11Y147_SLICE_X15Y147_CO6),
.I1(CLBLM_L_X12Y147_SLICE_X16Y147_DO6),
.I2(CLBLM_R_X11Y148_SLICE_X14Y148_DO6),
.I3(CLBLM_R_X11Y150_SLICE_X15Y150_CO6),
.I4(CLBLM_R_X7Y147_SLICE_X8Y147_DO6),
.I5(CLBLM_R_X11Y150_SLICE_X15Y150_BO6),
.O5(CLBLM_R_X11Y148_SLICE_X15Y148_DO5),
.O6(CLBLM_R_X11Y148_SLICE_X15Y148_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hcccccceeccceccce)
  ) CLBLM_R_X11Y148_SLICE_X15Y148_CLUT (
.I0(CLBLM_L_X12Y148_SLICE_X17Y148_AO6),
.I1(CLBLM_R_X11Y144_SLICE_X14Y144_DO6),
.I2(CLBLM_L_X10Y151_SLICE_X12Y151_AQ),
.I3(CLBLM_L_X12Y148_SLICE_X16Y148_DO6),
.I4(CLBLM_L_X12Y145_SLICE_X16Y145_BO6),
.I5(CLBLM_R_X13Y146_SLICE_X18Y146_BO6),
.O5(CLBLM_R_X11Y148_SLICE_X15Y148_CO5),
.O6(CLBLM_R_X11Y148_SLICE_X15Y148_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hcccccccececccece)
  ) CLBLM_R_X11Y148_SLICE_X15Y148_BLUT (
.I0(CLBLM_L_X12Y147_SLICE_X17Y147_DO6),
.I1(CLBLM_R_X11Y144_SLICE_X14Y144_DO6),
.I2(CLBLM_L_X12Y147_SLICE_X16Y147_CO6),
.I3(CLBLM_R_X13Y146_SLICE_X18Y146_BO6),
.I4(CLBLM_R_X3Y145_SLICE_X2Y145_AQ),
.I5(CLBLM_L_X12Y145_SLICE_X16Y145_BO6),
.O5(CLBLM_R_X11Y148_SLICE_X15Y148_BO5),
.O6(CLBLM_R_X11Y148_SLICE_X15Y148_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffffffffffdff)
  ) CLBLM_R_X11Y148_SLICE_X15Y148_ALUT (
.I0(CLBLM_R_X7Y153_SLICE_X8Y153_A5Q),
.I1(CLBLM_R_X7Y149_SLICE_X8Y149_AQ),
.I2(CLBLM_R_X7Y144_SLICE_X9Y144_B5Q),
.I3(CLBLL_L_X4Y148_SLICE_X4Y148_CQ),
.I4(CLBLM_L_X12Y147_SLICE_X16Y147_DO6),
.I5(CLBLM_L_X10Y146_SLICE_X13Y146_DO6),
.O5(CLBLM_R_X11Y148_SLICE_X15Y148_AO5),
.O6(CLBLM_R_X11Y148_SLICE_X15Y148_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffffefffffffe)
  ) CLBLM_R_X11Y149_SLICE_X14Y149_DLUT (
.I0(CLBLM_L_X8Y149_SLICE_X11Y149_CO6),
.I1(CLBLM_R_X11Y150_SLICE_X14Y150_CO6),
.I2(CLBLM_R_X7Y150_SLICE_X9Y150_DO6),
.I3(CLBLM_L_X10Y149_SLICE_X13Y149_DO6),
.I4(CLBLM_L_X8Y150_SLICE_X10Y150_DO6),
.I5(1'b1),
.O5(CLBLM_R_X11Y149_SLICE_X14Y149_DO5),
.O6(CLBLM_R_X11Y149_SLICE_X14Y149_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h9969996666966699)
  ) CLBLM_R_X11Y149_SLICE_X14Y149_CLUT (
.I0(CLBLM_L_X8Y149_SLICE_X11Y149_BO6),
.I1(CLBLM_L_X10Y147_SLICE_X13Y147_CO6),
.I2(CLBLM_R_X11Y148_SLICE_X14Y148_CO6),
.I3(CLBLM_L_X10Y149_SLICE_X12Y149_DO6),
.I4(CLBLM_L_X12Y147_SLICE_X16Y147_DO6),
.I5(CLBLM_R_X11Y148_SLICE_X14Y148_BO6),
.O5(CLBLM_R_X11Y149_SLICE_X14Y149_CO5),
.O6(CLBLM_R_X11Y149_SLICE_X14Y149_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffefffffffee)
  ) CLBLM_R_X11Y149_SLICE_X14Y149_BLUT (
.I0(CLBLM_R_X7Y150_SLICE_X9Y150_DO6),
.I1(CLBLM_L_X8Y149_SLICE_X11Y149_CO6),
.I2(CLBLM_R_X13Y149_SLICE_X18Y149_AO6),
.I3(CLBLM_L_X10Y149_SLICE_X13Y149_DO6),
.I4(CLBLM_L_X12Y149_SLICE_X17Y149_DO6),
.I5(CLBLM_R_X5Y146_SLICE_X7Y146_AQ),
.O5(CLBLM_R_X11Y149_SLICE_X14Y149_BO5),
.O6(CLBLM_R_X11Y149_SLICE_X14Y149_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0011001500110011)
  ) CLBLM_R_X11Y149_SLICE_X14Y149_ALUT (
.I0(CLBLM_L_X8Y150_SLICE_X10Y150_DO6),
.I1(CLBLM_L_X12Y147_SLICE_X16Y147_DO6),
.I2(CLBLM_L_X10Y148_SLICE_X12Y148_DO6),
.I3(CLBLM_R_X11Y149_SLICE_X14Y149_BO6),
.I4(CLBLM_L_X8Y146_SLICE_X10Y146_DO6),
.I5(CLBLM_R_X11Y147_SLICE_X14Y147_CO6),
.O5(CLBLM_R_X11Y149_SLICE_X14Y149_AO5),
.O6(CLBLM_R_X11Y149_SLICE_X14Y149_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffffffffffee)
  ) CLBLM_R_X11Y149_SLICE_X15Y149_DLUT (
.I0(CLBLM_L_X10Y150_SLICE_X13Y150_BO5),
.I1(CLBLM_L_X12Y149_SLICE_X16Y149_DO6),
.I2(1'b1),
.I3(CLBLM_R_X7Y148_SLICE_X8Y148_CO6),
.I4(CLBLM_R_X11Y150_SLICE_X14Y150_AO6),
.I5(CLBLM_L_X8Y149_SLICE_X10Y149_AO6),
.O5(CLBLM_R_X11Y149_SLICE_X15Y149_DO5),
.O6(CLBLM_R_X11Y149_SLICE_X15Y149_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h3cc3aaaac33caaaa)
  ) CLBLM_R_X11Y149_SLICE_X15Y149_CLUT (
.I0(CLBLM_L_X10Y145_SLICE_X13Y145_BO6),
.I1(CLBLM_R_X11Y149_SLICE_X14Y149_CO6),
.I2(CLBLM_R_X11Y152_SLICE_X15Y152_AQ),
.I3(CLBLM_R_X11Y148_SLICE_X15Y148_DO6),
.I4(RIOB33_X105Y131_IOB_X1Y132_I),
.I5(CLBLM_L_X12Y149_SLICE_X16Y149_CO6),
.O5(CLBLM_R_X11Y149_SLICE_X15Y149_CO5),
.O6(CLBLM_R_X11Y149_SLICE_X15Y149_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffcf00ffffefaa)
  ) CLBLM_R_X11Y149_SLICE_X15Y149_BLUT (
.I0(CLBLL_L_X4Y150_SLICE_X4Y150_CQ),
.I1(CLBLM_R_X11Y144_SLICE_X14Y144_CO6),
.I2(CLBLM_L_X12Y146_SLICE_X16Y146_AO6),
.I3(CLBLM_L_X8Y152_SLICE_X10Y152_DQ),
.I4(CLBLM_L_X8Y151_SLICE_X11Y151_BO6),
.I5(CLBLM_R_X7Y148_SLICE_X8Y148_AO5),
.O5(CLBLM_R_X11Y149_SLICE_X15Y149_BO5),
.O6(CLBLM_R_X11Y149_SLICE_X15Y149_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000110051)
  ) CLBLM_R_X11Y149_SLICE_X15Y149_ALUT (
.I0(CLBLM_R_X11Y151_SLICE_X14Y151_CO6),
.I1(CLBLM_L_X12Y147_SLICE_X16Y147_DO6),
.I2(CLBLM_R_X11Y147_SLICE_X15Y147_AO6),
.I3(CLBLM_R_X11Y149_SLICE_X15Y149_BO6),
.I4(CLBLM_L_X8Y146_SLICE_X10Y146_BO6),
.I5(CLBLM_L_X8Y149_SLICE_X10Y149_DO6),
.O5(CLBLM_R_X11Y149_SLICE_X15Y149_AO5),
.O6(CLBLM_R_X11Y149_SLICE_X15Y149_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y150_SLICE_X14Y150_A_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(LIOB33_X0Y61_IOB_X0Y62_I),
.D(CLBLM_L_X10Y150_SLICE_X13Y150_AQ),
.Q(CLBLM_R_X11Y150_SLICE_X14Y150_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000222200f00000)
  ) CLBLM_R_X11Y150_SLICE_X14Y150_DLUT (
.I0(CLBLM_R_X7Y146_SLICE_X8Y146_C5Q),
.I1(CLBLM_R_X11Y147_SLICE_X15Y147_BO6),
.I2(CLBLM_R_X7Y152_SLICE_X8Y152_DQ),
.I3(CLBLM_R_X11Y144_SLICE_X14Y144_BO6),
.I4(CLBLM_R_X7Y144_SLICE_X9Y144_B5Q),
.I5(CLBLM_R_X7Y153_SLICE_X8Y153_A5Q),
.O5(CLBLM_R_X11Y150_SLICE_X14Y150_DO5),
.O6(CLBLM_R_X11Y150_SLICE_X14Y150_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffffff5fdf0fc)
  ) CLBLM_R_X11Y150_SLICE_X14Y150_CLUT (
.I0(CLBLM_L_X12Y149_SLICE_X17Y149_BO5),
.I1(CLBLM_R_X5Y146_SLICE_X7Y146_AQ),
.I2(CLBLM_L_X10Y146_SLICE_X13Y146_DO6),
.I3(CLBLM_R_X13Y149_SLICE_X18Y149_AO6),
.I4(CLBLM_L_X8Y152_SLICE_X11Y152_CQ),
.I5(CLBLM_L_X12Y150_SLICE_X16Y150_CO6),
.O5(CLBLM_R_X11Y150_SLICE_X14Y150_CO5),
.O6(CLBLM_R_X11Y150_SLICE_X14Y150_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffff0fcfffffafe)
  ) CLBLM_R_X11Y150_SLICE_X14Y150_BLUT (
.I0(CLBLM_R_X7Y152_SLICE_X8Y152_DQ),
.I1(CLBLM_R_X7Y146_SLICE_X8Y146_C5Q),
.I2(CLBLM_L_X10Y150_SLICE_X13Y150_BO6),
.I3(CLBLM_L_X8Y150_SLICE_X10Y150_BO6),
.I4(CLBLM_R_X11Y150_SLICE_X14Y150_AO6),
.I5(CLBLM_L_X10Y148_SLICE_X12Y148_AO6),
.O5(CLBLM_R_X11Y150_SLICE_X14Y150_BO5),
.O6(CLBLM_R_X11Y150_SLICE_X14Y150_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffefffeecfcfcccc)
  ) CLBLM_R_X11Y150_SLICE_X14Y150_ALUT (
.I0(CLBLM_L_X10Y146_SLICE_X13Y146_DO6),
.I1(CLBLM_R_X11Y151_SLICE_X14Y151_BO6),
.I2(CLBLM_L_X12Y149_SLICE_X17Y149_BO5),
.I3(CLBLM_R_X7Y146_SLICE_X9Y146_BQ),
.I4(CLBLM_R_X11Y151_SLICE_X14Y151_AQ),
.I5(CLBLM_R_X11Y148_SLICE_X15Y148_AO6),
.O5(CLBLM_R_X11Y150_SLICE_X14Y150_AO5),
.O6(CLBLM_R_X11Y150_SLICE_X14Y150_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0c0cff0c0c0cff0c)
  ) CLBLM_R_X11Y150_SLICE_X15Y150_DLUT (
.I0(1'b1),
.I1(CLBLM_R_X7Y151_SLICE_X8Y151_CQ),
.I2(CLBLM_L_X10Y148_SLICE_X12Y148_AO6),
.I3(CLBLM_R_X7Y152_SLICE_X8Y152_CQ),
.I4(CLBLM_L_X12Y149_SLICE_X17Y149_BO5),
.I5(1'b1),
.O5(CLBLM_R_X11Y150_SLICE_X15Y150_DO5),
.O6(CLBLM_R_X11Y150_SLICE_X15Y150_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffffffffffefe)
  ) CLBLM_R_X11Y150_SLICE_X15Y150_CLUT (
.I0(CLBLM_L_X12Y150_SLICE_X16Y150_BO6),
.I1(CLBLM_R_X7Y150_SLICE_X8Y150_CO6),
.I2(CLBLM_L_X8Y149_SLICE_X10Y149_DO6),
.I3(1'b1),
.I4(CLBLM_R_X11Y151_SLICE_X14Y151_DO6),
.I5(CLBLM_L_X8Y151_SLICE_X11Y151_BO6),
.O5(CLBLM_R_X11Y150_SLICE_X15Y150_CO5),
.O6(CLBLM_R_X11Y150_SLICE_X15Y150_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffffffffffba)
  ) CLBLM_R_X11Y150_SLICE_X15Y150_BLUT (
.I0(CLBLM_R_X11Y150_SLICE_X15Y150_DO6),
.I1(CLBLM_L_X12Y149_SLICE_X17Y149_CO6),
.I2(CLBLM_R_X7Y153_SLICE_X9Y153_BQ),
.I3(CLBLM_L_X8Y150_SLICE_X11Y150_DO6),
.I4(CLBLM_R_X7Y149_SLICE_X8Y149_CO6),
.I5(CLBLM_R_X11Y151_SLICE_X15Y151_BO6),
.O5(CLBLM_R_X11Y150_SLICE_X15Y150_BO5),
.O6(CLBLM_R_X11Y150_SLICE_X15Y150_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffbaffbaffffffba)
  ) CLBLM_R_X11Y150_SLICE_X15Y150_ALUT (
.I0(CLBLM_R_X11Y150_SLICE_X15Y150_DO6),
.I1(CLBLM_L_X12Y149_SLICE_X17Y149_CO6),
.I2(CLBLM_R_X7Y153_SLICE_X9Y153_BQ),
.I3(CLBLM_L_X8Y150_SLICE_X11Y150_DO6),
.I4(CLBLM_R_X7Y143_SLICE_X9Y143_BQ),
.I5(CLBLM_L_X8Y150_SLICE_X10Y150_BO6),
.O5(CLBLM_R_X11Y150_SLICE_X15Y150_AO5),
.O6(CLBLM_R_X11Y150_SLICE_X15Y150_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y151_SLICE_X14Y151_A_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_R_X11Y151_SLICE_X14Y151_AO6),
.Q(CLBLM_R_X11Y151_SLICE_X14Y151_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffff50dc50dc)
  ) CLBLM_R_X11Y151_SLICE_X14Y151_DLUT (
.I0(CLBLM_L_X10Y148_SLICE_X12Y148_AO6),
.I1(CLBLM_R_X3Y150_SLICE_X3Y150_D5Q),
.I2(CLBLL_L_X4Y150_SLICE_X4Y150_A5Q),
.I3(CLBLM_L_X8Y150_SLICE_X10Y150_BO6),
.I4(1'b1),
.I5(CLBLM_L_X10Y151_SLICE_X13Y151_DO6),
.O5(CLBLM_R_X11Y151_SLICE_X14Y151_DO5),
.O6(CLBLM_R_X11Y151_SLICE_X14Y151_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffffdfddcfcc)
  ) CLBLM_R_X11Y151_SLICE_X14Y151_CLUT (
.I0(CLBLM_L_X10Y148_SLICE_X12Y148_AO6),
.I1(CLBLM_R_X7Y150_SLICE_X8Y150_CO6),
.I2(CLBLM_L_X8Y150_SLICE_X10Y150_BO6),
.I3(CLBLM_R_X3Y150_SLICE_X3Y150_D5Q),
.I4(CLBLL_L_X4Y150_SLICE_X4Y150_A5Q),
.I5(CLBLM_L_X10Y151_SLICE_X13Y151_DO6),
.O5(CLBLM_R_X11Y151_SLICE_X14Y151_CO5),
.O6(CLBLM_R_X11Y151_SLICE_X14Y151_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h00cc000010101010)
  ) CLBLM_R_X11Y151_SLICE_X14Y151_BLUT (
.I0(CLBLM_R_X11Y144_SLICE_X14Y144_BO6),
.I1(CLBLM_R_X7Y153_SLICE_X8Y153_A5Q),
.I2(CLBLM_R_X11Y151_SLICE_X15Y151_A5Q),
.I3(CLBLM_R_X11Y147_SLICE_X15Y147_BO6),
.I4(CLBLM_R_X11Y151_SLICE_X15Y151_AQ),
.I5(CLBLM_R_X7Y144_SLICE_X9Y144_B5Q),
.O5(CLBLM_R_X11Y151_SLICE_X14Y151_BO5),
.O6(CLBLM_R_X11Y151_SLICE_X14Y151_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffb8b80000b8b8)
  ) CLBLM_R_X11Y151_SLICE_X14Y151_ALUT (
.I0(CLBLM_R_X7Y144_SLICE_X9Y144_AQ),
.I1(CLBLM_L_X12Y149_SLICE_X17Y149_CO6),
.I2(CLBLM_R_X11Y151_SLICE_X14Y151_AQ),
.I3(1'b1),
.I4(LIOB33_X0Y61_IOB_X0Y62_I),
.I5(CLBLM_R_X7Y153_SLICE_X9Y153_DQ),
.O5(CLBLM_R_X11Y151_SLICE_X14Y151_AO5),
.O6(CLBLM_R_X11Y151_SLICE_X14Y151_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y151_SLICE_X15Y151_A5_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_R_X11Y151_SLICE_X15Y151_AO5),
.Q(CLBLM_R_X11Y151_SLICE_X15Y151_A5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y151_SLICE_X15Y151_A_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_R_X11Y151_SLICE_X15Y151_AO6),
.Q(CLBLM_R_X11Y151_SLICE_X15Y151_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X11Y151_SLICE_X15Y151_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X11Y151_SLICE_X15Y151_DO5),
.O6(CLBLM_R_X11Y151_SLICE_X15Y151_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X11Y151_SLICE_X15Y151_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X11Y151_SLICE_X15Y151_CO5),
.O6(CLBLM_R_X11Y151_SLICE_X15Y151_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000400000000)
  ) CLBLM_R_X11Y151_SLICE_X15Y151_BLUT (
.I0(CLBLL_L_X4Y148_SLICE_X4Y148_CQ),
.I1(CLBLM_R_X7Y153_SLICE_X8Y153_A5Q),
.I2(CLBLM_L_X12Y147_SLICE_X16Y147_DO6),
.I3(CLBLM_R_X7Y144_SLICE_X9Y144_B5Q),
.I4(CLBLM_R_X7Y149_SLICE_X8Y149_AQ),
.I5(CLBLM_R_X7Y143_SLICE_X9Y143_BQ),
.O5(CLBLM_R_X11Y151_SLICE_X15Y151_BO5),
.O6(CLBLM_R_X11Y151_SLICE_X15Y151_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0ff000fc0cfc0cf)
  ) CLBLM_R_X11Y151_SLICE_X15Y151_ALUT (
.I0(1'b1),
.I1(CLBLM_R_X5Y149_SLICE_X7Y149_D5Q),
.I2(LIOB33_X0Y61_IOB_X0Y62_I),
.I3(CLBLM_L_X12Y151_SLICE_X16Y151_AQ),
.I4(CLBLM_R_X11Y151_SLICE_X14Y151_AQ),
.I5(1'b1),
.O5(CLBLM_R_X11Y151_SLICE_X15Y151_AO5),
.O6(CLBLM_R_X11Y151_SLICE_X15Y151_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X11Y152_SLICE_X14Y152_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X11Y152_SLICE_X14Y152_DO5),
.O6(CLBLM_R_X11Y152_SLICE_X14Y152_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X11Y152_SLICE_X14Y152_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X11Y152_SLICE_X14Y152_CO5),
.O6(CLBLM_R_X11Y152_SLICE_X14Y152_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X11Y152_SLICE_X14Y152_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X11Y152_SLICE_X14Y152_BO5),
.O6(CLBLM_R_X11Y152_SLICE_X14Y152_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000004000)
  ) CLBLM_R_X11Y152_SLICE_X14Y152_ALUT (
.I0(CLBLM_L_X10Y153_SLICE_X13Y153_CQ),
.I1(CLBLM_L_X8Y152_SLICE_X10Y152_CQ),
.I2(CLBLM_R_X7Y146_SLICE_X8Y146_A5Q),
.I3(CLBLM_L_X10Y152_SLICE_X12Y152_AQ),
.I4(CLBLM_R_X11Y153_SLICE_X14Y153_AQ),
.I5(CLBLM_R_X5Y147_SLICE_X6Y147_AQ),
.O5(CLBLM_R_X11Y152_SLICE_X14Y152_AO5),
.O6(CLBLM_R_X11Y152_SLICE_X14Y152_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y152_SLICE_X15Y152_A5_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_R_X11Y152_SLICE_X15Y152_AO5),
.Q(CLBLM_R_X11Y152_SLICE_X15Y152_A5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y152_SLICE_X15Y152_B5_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_R_X11Y152_SLICE_X15Y152_BO5),
.Q(CLBLM_R_X11Y152_SLICE_X15Y152_B5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y152_SLICE_X15Y152_A_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_R_X11Y152_SLICE_X15Y152_AO6),
.Q(CLBLM_R_X11Y152_SLICE_X15Y152_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y152_SLICE_X15Y152_B_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_R_X11Y152_SLICE_X15Y152_BO6),
.Q(CLBLM_R_X11Y152_SLICE_X15Y152_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y152_SLICE_X15Y152_C_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_R_X11Y152_SLICE_X15Y152_CO6),
.Q(CLBLM_R_X11Y152_SLICE_X15Y152_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X11Y152_SLICE_X15Y152_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X11Y152_SLICE_X15Y152_DO5),
.O6(CLBLM_R_X11Y152_SLICE_X15Y152_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hcc33cc33cc33cc33)
  ) CLBLM_R_X11Y152_SLICE_X15Y152_CLUT (
.I0(1'b1),
.I1(CLBLM_R_X11Y152_SLICE_X15Y152_CQ),
.I2(1'b1),
.I3(CLBLM_L_X10Y151_SLICE_X13Y151_CO6),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X11Y152_SLICE_X15Y152_CO5),
.O6(CLBLM_R_X11Y152_SLICE_X15Y152_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hcc9ccc9cff1000ef)
  ) CLBLM_R_X11Y152_SLICE_X15Y152_BLUT (
.I0(CLBLM_R_X11Y152_SLICE_X15Y152_CQ),
.I1(CLBLM_R_X11Y152_SLICE_X15Y152_BQ),
.I2(CLBLM_R_X11Y152_SLICE_X15Y152_A5Q),
.I3(CLBLM_L_X10Y151_SLICE_X13Y151_CO6),
.I4(CLBLM_R_X11Y152_SLICE_X15Y152_B5Q),
.I5(1'b1),
.O5(CLBLM_R_X11Y152_SLICE_X15Y152_BO5),
.O6(CLBLM_R_X11Y152_SLICE_X15Y152_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h00001010f05af05a)
  ) CLBLM_R_X11Y152_SLICE_X15Y152_ALUT (
.I0(CLBLM_R_X11Y152_SLICE_X15Y152_CQ),
.I1(CLBLM_R_X11Y152_SLICE_X15Y152_BQ),
.I2(CLBLM_R_X11Y152_SLICE_X15Y152_A5Q),
.I3(CLBLM_L_X10Y151_SLICE_X13Y151_CO6),
.I4(CLBLM_R_X11Y152_SLICE_X15Y152_B5Q),
.I5(1'b1),
.O5(CLBLM_R_X11Y152_SLICE_X15Y152_AO5),
.O6(CLBLM_R_X11Y152_SLICE_X15Y152_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y153_SLICE_X14Y153_A5_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_R_X11Y153_SLICE_X14Y153_AO5),
.Q(CLBLM_R_X11Y153_SLICE_X14Y153_A5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y153_SLICE_X14Y153_A_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_R_X11Y153_SLICE_X14Y153_AO6),
.Q(CLBLM_R_X11Y153_SLICE_X14Y153_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h7fff7fffffffffff)
  ) CLBLM_R_X11Y153_SLICE_X14Y153_DLUT (
.I0(CLBLM_L_X10Y152_SLICE_X13Y152_AQ),
.I1(CLBLM_L_X10Y152_SLICE_X13Y152_BQ),
.I2(CLBLM_R_X11Y153_SLICE_X14Y153_AQ),
.I3(CLBLM_L_X10Y152_SLICE_X12Y152_AQ),
.I4(1'b1),
.I5(CLBLM_L_X8Y152_SLICE_X10Y152_CQ),
.O5(CLBLM_R_X11Y153_SLICE_X14Y153_DO5),
.O6(CLBLM_R_X11Y153_SLICE_X14Y153_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h4444c6cc4444cccc)
  ) CLBLM_R_X11Y153_SLICE_X14Y153_CLUT (
.I0(CLBLM_R_X7Y146_SLICE_X8Y146_A5Q),
.I1(CLBLM_R_X11Y153_SLICE_X14Y153_AQ),
.I2(CLBLM_R_X5Y147_SLICE_X6Y147_AQ),
.I3(CLBLM_L_X10Y152_SLICE_X12Y152_AQ),
.I4(CLBLM_L_X10Y153_SLICE_X13Y153_CQ),
.I5(CLBLM_L_X8Y152_SLICE_X10Y152_CQ),
.O5(CLBLM_R_X11Y153_SLICE_X14Y153_CO5),
.O6(CLBLM_R_X11Y153_SLICE_X14Y153_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h8000000000000000)
  ) CLBLM_R_X11Y153_SLICE_X14Y153_BLUT (
.I0(CLBLM_L_X8Y152_SLICE_X10Y152_CQ),
.I1(CLBLM_L_X10Y152_SLICE_X13Y152_BQ),
.I2(CLBLM_R_X11Y153_SLICE_X14Y153_AQ),
.I3(CLBLM_L_X10Y152_SLICE_X12Y152_AQ),
.I4(CLBLM_L_X10Y152_SLICE_X13Y152_AQ),
.I5(CLBLM_R_X11Y153_SLICE_X15Y153_BO5),
.O5(CLBLM_R_X11Y153_SLICE_X14Y153_BO5),
.O6(CLBLM_R_X11Y153_SLICE_X14Y153_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hff0ff000acacacac)
  ) CLBLM_R_X11Y153_SLICE_X14Y153_ALUT (
.I0(CLBLM_L_X10Y148_SLICE_X13Y148_C5Q),
.I1(CLBLM_R_X11Y153_SLICE_X15Y153_BO6),
.I2(LIOB33_X0Y61_IOB_X0Y62_I),
.I3(CLBLM_L_X8Y152_SLICE_X10Y152_C5Q),
.I4(CLBLM_R_X11Y153_SLICE_X14Y153_CO6),
.I5(1'b1),
.O5(CLBLM_R_X11Y153_SLICE_X14Y153_AO5),
.O6(CLBLM_R_X11Y153_SLICE_X14Y153_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y153_SLICE_X15Y153_A_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_R_X11Y153_SLICE_X15Y153_AO6),
.Q(CLBLM_R_X11Y153_SLICE_X15Y153_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hf3f3f3f3ffffffff)
  ) CLBLM_R_X11Y153_SLICE_X15Y153_DLUT (
.I0(1'b1),
.I1(CLBLM_R_X11Y153_SLICE_X14Y153_A5Q),
.I2(CLBLM_R_X11Y153_SLICE_X14Y153_DO6),
.I3(1'b1),
.I4(1'b1),
.I5(CLBLM_R_X11Y153_SLICE_X15Y153_AQ),
.O5(CLBLM_R_X11Y153_SLICE_X15Y153_DO5),
.O6(CLBLM_R_X11Y153_SLICE_X15Y153_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h5555fff75555ffff)
  ) CLBLM_R_X11Y153_SLICE_X15Y153_CLUT (
.I0(CLBLM_R_X7Y146_SLICE_X8Y146_A5Q),
.I1(CLBLM_R_X11Y153_SLICE_X14Y153_A5Q),
.I2(CLBLM_R_X11Y153_SLICE_X14Y153_DO6),
.I3(CLBLM_R_X5Y147_SLICE_X6Y147_AQ),
.I4(CLBLM_L_X10Y153_SLICE_X13Y153_CQ),
.I5(CLBLM_R_X11Y153_SLICE_X15Y153_AQ),
.O5(CLBLM_R_X11Y153_SLICE_X15Y153_CO5),
.O6(CLBLM_R_X11Y153_SLICE_X15Y153_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0a09aaaa000f0000)
  ) CLBLM_R_X11Y153_SLICE_X15Y153_BLUT (
.I0(CLBLM_R_X11Y153_SLICE_X14Y153_A5Q),
.I1(CLBLM_R_X11Y153_SLICE_X14Y153_DO6),
.I2(CLBLM_L_X10Y153_SLICE_X13Y153_CQ),
.I3(CLBLM_R_X5Y147_SLICE_X6Y147_AQ),
.I4(CLBLM_R_X7Y146_SLICE_X8Y146_A5Q),
.I5(1'b1),
.O5(CLBLM_R_X11Y153_SLICE_X15Y153_BO5),
.O6(CLBLM_R_X11Y153_SLICE_X15Y153_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hff00f8f8ff000808)
  ) CLBLM_R_X11Y153_SLICE_X15Y153_ALUT (
.I0(CLBLM_R_X11Y153_SLICE_X14Y153_A5Q),
.I1(CLBLM_R_X11Y153_SLICE_X14Y153_BO6),
.I2(CLBLM_R_X11Y153_SLICE_X15Y153_AQ),
.I3(CLBLM_L_X8Y148_SLICE_X11Y148_B5Q),
.I4(LIOB33_X0Y61_IOB_X0Y62_I),
.I5(CLBLM_R_X11Y153_SLICE_X15Y153_CO6),
.O5(CLBLM_R_X11Y153_SLICE_X15Y153_AO5),
.O6(CLBLM_R_X11Y153_SLICE_X15Y153_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X13Y146_SLICE_X18Y146_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X13Y146_SLICE_X18Y146_DO5),
.O6(CLBLM_R_X13Y146_SLICE_X18Y146_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hfaf0faf0aa00aa00)
  ) CLBLM_R_X13Y146_SLICE_X18Y146_CLUT (
.I0(RIOB33_X105Y141_IOB_X1Y141_I),
.I1(1'b1),
.I2(CLBLM_L_X10Y147_SLICE_X12Y147_AQ),
.I3(CLBLM_L_X10Y147_SLICE_X12Y147_CQ),
.I4(1'b1),
.I5(RIOB33_X105Y139_IOB_X1Y140_I),
.O5(CLBLM_R_X13Y146_SLICE_X18Y146_CO5),
.O6(CLBLM_R_X13Y146_SLICE_X18Y146_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffffffffefff)
  ) CLBLM_R_X13Y146_SLICE_X18Y146_BLUT (
.I0(CLBLM_R_X7Y153_SLICE_X8Y153_A5Q),
.I1(CLBLM_R_X7Y144_SLICE_X9Y144_B5Q),
.I2(CLBLM_R_X7Y149_SLICE_X8Y149_AQ),
.I3(CLBLL_L_X4Y148_SLICE_X4Y148_CQ),
.I4(CLBLM_R_X7Y146_SLICE_X9Y146_CO6),
.I5(CLBLM_L_X10Y146_SLICE_X13Y146_DO6),
.O5(CLBLM_R_X13Y146_SLICE_X18Y146_BO5),
.O6(CLBLM_R_X13Y146_SLICE_X18Y146_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffbbbb00003210)
  ) CLBLM_R_X13Y146_SLICE_X18Y146_ALUT (
.I0(CLBLM_R_X7Y153_SLICE_X8Y153_A5Q),
.I1(CLBLM_R_X7Y144_SLICE_X9Y144_B5Q),
.I2(RIOB33_X105Y143_IOB_X1Y143_I),
.I3(CLBLM_L_X12Y146_SLICE_X16Y146_AQ),
.I4(CLBLM_L_X12Y145_SLICE_X17Y145_CO6),
.I5(1'b1),
.O5(CLBLM_R_X13Y146_SLICE_X18Y146_AO5),
.O6(CLBLM_R_X13Y146_SLICE_X18Y146_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X13Y146_SLICE_X19Y146_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X13Y146_SLICE_X19Y146_DO5),
.O6(CLBLM_R_X13Y146_SLICE_X19Y146_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X13Y146_SLICE_X19Y146_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X13Y146_SLICE_X19Y146_CO5),
.O6(CLBLM_R_X13Y146_SLICE_X19Y146_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X13Y146_SLICE_X19Y146_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X13Y146_SLICE_X19Y146_BO5),
.O6(CLBLM_R_X13Y146_SLICE_X19Y146_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X13Y146_SLICE_X19Y146_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X13Y146_SLICE_X19Y146_AO5),
.O6(CLBLM_R_X13Y146_SLICE_X19Y146_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X13Y149_SLICE_X18Y149_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X13Y149_SLICE_X18Y149_DO5),
.O6(CLBLM_R_X13Y149_SLICE_X18Y149_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X13Y149_SLICE_X18Y149_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X13Y149_SLICE_X18Y149_CO5),
.O6(CLBLM_R_X13Y149_SLICE_X18Y149_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X13Y149_SLICE_X18Y149_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X13Y149_SLICE_X18Y149_BO5),
.O6(CLBLM_R_X13Y149_SLICE_X18Y149_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffffffffffef)
  ) CLBLM_R_X13Y149_SLICE_X18Y149_ALUT (
.I0(CLBLM_R_X7Y144_SLICE_X9Y144_B5Q),
.I1(CLBLM_R_X7Y153_SLICE_X8Y153_A5Q),
.I2(CLBLM_R_X7Y149_SLICE_X8Y149_AQ),
.I3(CLBLL_L_X4Y148_SLICE_X4Y148_CQ),
.I4(CLBLM_L_X12Y147_SLICE_X16Y147_DO6),
.I5(CLBLM_L_X10Y146_SLICE_X13Y146_DO6),
.O5(CLBLM_R_X13Y149_SLICE_X18Y149_AO5),
.O6(CLBLM_R_X13Y149_SLICE_X18Y149_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X13Y149_SLICE_X19Y149_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X13Y149_SLICE_X19Y149_DO5),
.O6(CLBLM_R_X13Y149_SLICE_X19Y149_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X13Y149_SLICE_X19Y149_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X13Y149_SLICE_X19Y149_CO5),
.O6(CLBLM_R_X13Y149_SLICE_X19Y149_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X13Y149_SLICE_X19Y149_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X13Y149_SLICE_X19Y149_BO5),
.O6(CLBLM_R_X13Y149_SLICE_X19Y149_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X13Y149_SLICE_X19Y149_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X13Y149_SLICE_X19Y149_AO5),
.O6(CLBLM_R_X13Y149_SLICE_X19Y149_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y178_SLICE_X162Y178_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y178_SLICE_X162Y178_DO5),
.O6(CLBLM_R_X103Y178_SLICE_X162Y178_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y178_SLICE_X162Y178_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y178_SLICE_X162Y178_CO5),
.O6(CLBLM_R_X103Y178_SLICE_X162Y178_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y178_SLICE_X162Y178_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y178_SLICE_X162Y178_BO5),
.O6(CLBLM_R_X103Y178_SLICE_X162Y178_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y178_SLICE_X162Y178_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y178_SLICE_X162Y178_AO5),
.O6(CLBLM_R_X103Y178_SLICE_X162Y178_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y178_SLICE_X163Y178_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y178_SLICE_X163Y178_DO5),
.O6(CLBLM_R_X103Y178_SLICE_X163Y178_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y178_SLICE_X163Y178_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y178_SLICE_X163Y178_CO5),
.O6(CLBLM_R_X103Y178_SLICE_X163Y178_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y178_SLICE_X163Y178_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y178_SLICE_X163Y178_BO5),
.O6(CLBLM_R_X103Y178_SLICE_X163Y178_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hccccccccff00ff00)
  ) CLBLM_R_X103Y178_SLICE_X163Y178_ALUT (
.I0(1'b1),
.I1(RIOB33_X105Y125_IOB_X1Y125_I),
.I2(1'b1),
.I3(RIOB33_X105Y125_IOB_X1Y126_I),
.I4(1'b1),
.I5(RIOB33_X105Y127_IOB_X1Y127_I),
.O5(CLBLM_R_X103Y178_SLICE_X163Y178_AO5),
.O6(CLBLM_R_X103Y178_SLICE_X163Y178_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "BUFGCTRL" *)
  BUFGCTRL #(
    .INIT_OUT(0),
    .IS_CE0_INVERTED(0),
    .IS_CE1_INVERTED(1),
    .IS_IGNORE0_INVERTED(1),
    .IS_IGNORE1_INVERTED(0),
    .IS_S0_INVERTED(0),
    .IS_S1_INVERTED(1),
    .PRESELECT_I0("TRUE"),
    .PRESELECT_I1("FALSE")
  ) CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_BUFGCTRL (
.CE0(1'b1),
.CE1(1'b1),
.I0(LIOB33_X0Y77_IOB_X0Y78_I),
.I1(1'b1),
.IGNORE0(1'b1),
.IGNORE1(1'b1),
.O(CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_O),
.S0(1'b1),
.S1(1'b1)
  );


  (* KEEP, DONT_TOUCH, BEL = "BUFHCE" *)
  BUFHCE #(
    .CE_TYPE("SYNC"),
    .INIT_OUT(0),
    .IS_CE_INVERTED(0)
  ) CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_BUFHCE (
.CE(1'b1),
.I(CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_O),
.O(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O)
  );


  (* KEEP, DONT_TOUCH, BEL = "BUFHCE" *)
  BUFHCE #(
    .CE_TYPE("SYNC"),
    .INIT_OUT(0),
    .IS_CE_INVERTED(0)
  ) CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_BUFHCE (
.CE(1'b1),
.I(CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_O),
.O(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y51_IOB_X0Y51_IBUF (
.I(LIOB33_X0Y51_IOB_X0Y51_IPAD),
.O(LIOB33_X0Y51_IOB_X0Y51_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y51_IOB_X0Y52_IBUF (
.I(LIOB33_X0Y51_IOB_X0Y52_IPAD),
.O(LIOB33_X0Y51_IOB_X0Y52_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y53_IOB_X0Y53_IBUF (
.I(LIOB33_X0Y53_IOB_X0Y53_IPAD),
.O(LIOB33_X0Y53_IOB_X0Y53_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y53_IOB_X0Y54_IBUF (
.I(LIOB33_X0Y53_IOB_X0Y54_IPAD),
.O(LIOB33_X0Y53_IOB_X0Y54_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y55_IOB_X0Y55_IBUF (
.I(LIOB33_X0Y55_IOB_X0Y55_IPAD),
.O(LIOB33_X0Y55_IOB_X0Y55_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y55_IOB_X0Y56_IBUF (
.I(LIOB33_X0Y55_IOB_X0Y56_IPAD),
.O(LIOB33_X0Y55_IOB_X0Y56_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y57_IOB_X0Y57_IBUF (
.I(LIOB33_X0Y57_IOB_X0Y57_IPAD),
.O(LIOB33_X0Y57_IOB_X0Y57_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y57_IOB_X0Y58_IBUF (
.I(LIOB33_X0Y57_IOB_X0Y58_IPAD),
.O(LIOB33_X0Y57_IOB_X0Y58_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y59_IOB_X0Y59_IBUF (
.I(LIOB33_X0Y59_IOB_X0Y59_IPAD),
.O(LIOB33_X0Y59_IOB_X0Y59_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y59_IOB_X0Y60_IBUF (
.I(LIOB33_X0Y59_IOB_X0Y60_IPAD),
.O(LIOB33_X0Y59_IOB_X0Y60_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y61_IOB_X0Y61_IBUF (
.I(LIOB33_X0Y61_IOB_X0Y61_IPAD),
.O(LIOB33_X0Y61_IOB_X0Y61_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y61_IOB_X0Y62_IBUF (
.I(LIOB33_X0Y61_IOB_X0Y62_IPAD),
.O(LIOB33_X0Y61_IOB_X0Y62_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y63_IOB_X0Y63_IBUF (
.I(LIOB33_X0Y63_IOB_X0Y63_IPAD),
.O(LIOB33_X0Y63_IOB_X0Y63_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y63_IOB_X0Y64_OBUF (
.I(CLBLM_R_X7Y141_SLICE_X8Y141_AO5),
.O(LIOB33_X0Y63_IOB_X0Y64_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y65_IOB_X0Y65_OBUF (
.I(CLBLM_R_X7Y141_SLICE_X8Y141_BO6),
.O(LIOB33_X0Y65_IOB_X0Y65_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y65_IOB_X0Y66_OBUF (
.I(CLBLL_L_X4Y151_SLICE_X4Y151_CQ),
.O(LIOB33_X0Y65_IOB_X0Y66_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y77_IOB_X0Y78_IBUF (
.I(LIOB33_X0Y77_IOB_X0Y78_IPAD),
.O(LIOB33_X0Y77_IOB_X0Y78_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y101_IOB_X0Y101_OBUF (
.I(CLBLM_L_X8Y145_SLICE_X11Y145_C5Q),
.O(LIOB33_X0Y101_IOB_X0Y101_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y101_IOB_X0Y102_OBUF (
.I(CLBLM_R_X5Y141_SLICE_X6Y141_DQ),
.O(LIOB33_X0Y101_IOB_X0Y102_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y103_IOB_X0Y103_OBUF (
.I(CLBLM_R_X5Y145_SLICE_X7Y145_BQ),
.O(LIOB33_X0Y103_IOB_X0Y103_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y103_IOB_X0Y104_OBUF (
.I(CLBLM_R_X3Y145_SLICE_X2Y145_C5Q),
.O(LIOB33_X0Y103_IOB_X0Y104_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y105_IOB_X0Y105_OBUF (
.I(CLBLL_L_X4Y150_SLICE_X4Y150_C5Q),
.O(LIOB33_X0Y105_IOB_X0Y105_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y105_IOB_X0Y106_OBUF (
.I(CLBLM_R_X3Y146_SLICE_X3Y146_BQ),
.O(LIOB33_X0Y105_IOB_X0Y106_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y107_IOB_X0Y107_OBUF (
.I(CLBLM_R_X7Y146_SLICE_X8Y146_DQ),
.O(LIOB33_X0Y107_IOB_X0Y107_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y107_IOB_X0Y108_OBUF (
.I(CLBLL_L_X4Y143_SLICE_X4Y143_DQ),
.O(LIOB33_X0Y107_IOB_X0Y108_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y109_IOB_X0Y109_OBUF (
.I(CLBLM_R_X5Y141_SLICE_X6Y141_BQ),
.O(LIOB33_X0Y109_IOB_X0Y109_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y109_IOB_X0Y110_OBUF (
.I(CLBLM_R_X5Y145_SLICE_X7Y145_AQ),
.O(LIOB33_X0Y109_IOB_X0Y110_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y111_IOB_X0Y111_OBUF (
.I(CLBLM_R_X3Y145_SLICE_X2Y145_B5Q),
.O(LIOB33_X0Y111_IOB_X0Y111_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y111_IOB_X0Y112_OBUF (
.I(CLBLL_L_X4Y146_SLICE_X4Y146_C5Q),
.O(LIOB33_X0Y111_IOB_X0Y112_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y113_IOB_X0Y113_OBUF (
.I(CLBLM_R_X3Y147_SLICE_X3Y147_C5Q),
.O(LIOB33_X0Y113_IOB_X0Y113_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y113_IOB_X0Y114_OBUF (
.I(CLBLM_L_X8Y142_SLICE_X10Y142_A5Q),
.O(LIOB33_X0Y113_IOB_X0Y114_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y115_IOB_X0Y115_OBUF (
.I(CLBLM_R_X5Y147_SLICE_X6Y147_C5Q),
.O(LIOB33_X0Y115_IOB_X0Y115_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y115_IOB_X0Y116_OBUF (
.I(CLBLM_R_X7Y143_SLICE_X9Y143_B5Q),
.O(LIOB33_X0Y115_IOB_X0Y116_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y117_IOB_X0Y117_OBUF (
.I(CLBLM_L_X10Y143_SLICE_X13Y143_C5Q),
.O(LIOB33_X0Y117_IOB_X0Y117_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y117_IOB_X0Y118_OBUF (
.I(CLBLM_R_X7Y142_SLICE_X9Y142_BQ),
.O(LIOB33_X0Y117_IOB_X0Y118_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y119_IOB_X0Y119_OBUF (
.I(CLBLL_L_X2Y146_SLICE_X0Y146_CQ),
.O(LIOB33_X0Y119_IOB_X0Y119_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y119_IOB_X0Y120_OBUF (
.I(CLBLL_L_X4Y147_SLICE_X4Y147_AQ),
.O(LIOB33_X0Y119_IOB_X0Y120_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y121_IOB_X0Y121_OBUF (
.I(CLBLM_L_X8Y147_SLICE_X10Y147_C5Q),
.O(LIOB33_X0Y121_IOB_X0Y121_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y121_IOB_X0Y122_OBUF (
.I(CLBLL_L_X4Y144_SLICE_X5Y144_CQ),
.O(LIOB33_X0Y121_IOB_X0Y122_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y123_IOB_X0Y123_OBUF (
.I(CLBLL_L_X2Y146_SLICE_X0Y146_CQ),
.O(LIOB33_X0Y123_IOB_X0Y123_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y123_IOB_X0Y124_OBUF (
.I(CLBLL_L_X4Y151_SLICE_X4Y151_CQ),
.O(LIOB33_X0Y123_IOB_X0Y124_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y125_IOB_X0Y125_OBUF (
.I(CLBLL_L_X4Y151_SLICE_X4Y151_BQ),
.O(LIOB33_X0Y125_IOB_X0Y125_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y125_IOB_X0Y126_OBUF (
.I(CLBLL_L_X4Y147_SLICE_X5Y147_CQ),
.O(LIOB33_X0Y125_IOB_X0Y126_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y127_IOB_X0Y127_OBUF (
.I(CLBLM_R_X7Y152_SLICE_X8Y152_D5Q),
.O(LIOB33_X0Y127_IOB_X0Y127_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y127_IOB_X0Y128_OBUF (
.I(CLBLM_L_X10Y145_SLICE_X12Y145_AQ),
.O(LIOB33_X0Y127_IOB_X0Y128_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y129_IOB_X0Y129_OBUF (
.I(CLBLL_L_X2Y146_SLICE_X0Y146_CQ),
.O(LIOB33_X0Y129_IOB_X0Y129_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y129_IOB_X0Y130_OBUF (
.I(CLBLL_L_X2Y145_SLICE_X0Y145_BQ),
.O(LIOB33_X0Y129_IOB_X0Y130_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y131_IOB_X0Y131_OBUF (
.I(CLBLL_L_X2Y75_SLICE_X0Y75_AO6),
.O(LIOB33_X0Y131_IOB_X0Y131_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y131_IOB_X0Y132_OBUF (
.I(CLBLM_R_X3Y143_SLICE_X2Y143_BO5),
.O(LIOB33_X0Y131_IOB_X0Y132_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y133_IOB_X0Y133_OBUF (
.I(CLBLL_L_X4Y140_SLICE_X4Y140_BO5),
.O(LIOB33_X0Y133_IOB_X0Y133_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y133_IOB_X0Y134_OBUF (
.I(CLBLL_L_X2Y145_SLICE_X0Y145_BQ),
.O(LIOB33_X0Y133_IOB_X0Y134_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y135_IOB_X0Y135_OBUF (
.I(CLBLL_L_X2Y145_SLICE_X0Y145_BQ),
.O(LIOB33_X0Y135_IOB_X0Y135_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y135_IOB_X0Y136_OBUF (
.I(CLBLM_L_X10Y153_SLICE_X13Y153_CQ),
.O(LIOB33_X0Y135_IOB_X0Y136_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y137_IOB_X0Y137_OBUF (
.I(CLBLM_R_X5Y153_SLICE_X6Y153_B5Q),
.O(LIOB33_X0Y137_IOB_X0Y137_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y137_IOB_X0Y138_OBUF (
.I(CLBLM_R_X3Y148_SLICE_X2Y148_A5Q),
.O(LIOB33_X0Y137_IOB_X0Y138_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y139_IOB_X0Y139_OBUF (
.I(CLBLM_R_X3Y147_SLICE_X2Y147_DQ),
.O(LIOB33_X0Y139_IOB_X0Y139_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y139_IOB_X0Y140_OBUF (
.I(CLBLL_L_X4Y145_SLICE_X4Y145_C5Q),
.O(LIOB33_X0Y139_IOB_X0Y140_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y141_IOB_X0Y141_OBUF (
.I(CLBLL_L_X4Y145_SLICE_X5Y145_CQ),
.O(LIOB33_X0Y141_IOB_X0Y141_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y141_IOB_X0Y142_OBUF (
.I(CLBLL_L_X2Y146_SLICE_X0Y146_CQ),
.O(LIOB33_X0Y141_IOB_X0Y142_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y143_IOB_X0Y143_OBUF (
.I(CLBLM_R_X3Y151_SLICE_X2Y151_BO5),
.O(LIOB33_X0Y143_IOB_X0Y143_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y145_IOB_X0Y145_OBUF (
.I(CLBLM_R_X3Y148_SLICE_X3Y148_DO6),
.O(LIOB33_X0Y145_IOB_X0Y145_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y145_IOB_X0Y146_OBUF (
.I(CLBLM_R_X3Y143_SLICE_X3Y143_DO6),
.O(LIOB33_X0Y145_IOB_X0Y146_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y147_IOB_X0Y147_OBUF (
.I(CLBLM_R_X5Y141_SLICE_X6Y141_CO5),
.O(LIOB33_X0Y147_IOB_X0Y147_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y147_IOB_X0Y148_OBUF (
.I(CLBLL_L_X2Y147_SLICE_X1Y147_AO6),
.O(LIOB33_X0Y147_IOB_X0Y148_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y151_IOB_X0Y151_OBUF (
.I(CLBLL_L_X2Y146_SLICE_X0Y146_CQ),
.O(LIOB33_X0Y151_IOB_X0Y151_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y151_IOB_X0Y152_OBUF (
.I(CLBLL_L_X4Y147_SLICE_X5Y147_C5Q),
.O(LIOB33_X0Y151_IOB_X0Y152_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y153_IOB_X0Y153_OBUF (
.I(CLBLM_L_X8Y153_SLICE_X10Y153_A5Q),
.O(LIOB33_X0Y153_IOB_X0Y153_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y153_IOB_X0Y154_OBUF (
.I(CLBLM_R_X7Y153_SLICE_X9Y153_DQ),
.O(LIOB33_X0Y153_IOB_X0Y154_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y155_IOB_X0Y155_OBUF (
.I(CLBLM_R_X5Y154_SLICE_X7Y154_AQ),
.O(LIOB33_X0Y155_IOB_X0Y155_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y155_IOB_X0Y156_OBUF (
.I(CLBLM_R_X3Y152_SLICE_X3Y152_CQ),
.O(LIOB33_X0Y155_IOB_X0Y156_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y157_IOB_X0Y157_OBUF (
.I(CLBLM_R_X3Y152_SLICE_X3Y152_BQ),
.O(LIOB33_X0Y157_IOB_X0Y157_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y157_IOB_X0Y158_OBUF (
.I(RIOB33_X105Y133_IOB_X1Y134_I),
.O(LIOB33_X0Y157_IOB_X0Y158_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y159_IOB_X0Y159_OBUF (
.I(CLBLL_L_X2Y146_SLICE_X0Y146_CQ),
.O(LIOB33_X0Y159_IOB_X0Y159_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y159_IOB_X0Y160_OBUF (
.I(CLBLL_L_X2Y148_SLICE_X0Y148_AQ),
.O(LIOB33_X0Y159_IOB_X0Y160_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y161_IOB_X0Y161_OBUF (
.I(CLBLM_R_X5Y152_SLICE_X7Y152_DQ),
.O(LIOB33_X0Y161_IOB_X0Y161_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y161_IOB_X0Y162_OBUF (
.I(CLBLM_L_X10Y144_SLICE_X12Y144_BO6),
.O(LIOB33_X0Y161_IOB_X0Y162_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y163_IOB_X0Y163_OBUF (
.I(CLBLM_R_X5Y152_SLICE_X7Y152_DO6),
.O(LIOB33_X0Y163_IOB_X0Y163_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y163_IOB_X0Y164_OBUF (
.I(RIOB33_X105Y101_IOB_X1Y102_I),
.O(LIOB33_X0Y163_IOB_X0Y164_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y165_IOB_X0Y165_OBUF (
.I(LIOB33_X0Y57_IOB_X0Y57_I),
.O(LIOB33_X0Y165_IOB_X0Y165_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y165_IOB_X0Y166_OBUF (
.I(RIOB33_SING_X105Y100_IOB_X1Y100_I),
.O(LIOB33_X0Y165_IOB_X0Y166_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y167_IOB_X0Y167_OBUF (
.I(RIOB33_X105Y105_IOB_X1Y106_I),
.O(LIOB33_X0Y167_IOB_X0Y167_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y167_IOB_X0Y168_OBUF (
.I(RIOB33_X105Y101_IOB_X1Y101_I),
.O(LIOB33_X0Y167_IOB_X0Y168_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y169_IOB_X0Y169_OBUF (
.I(RIOB33_X105Y117_IOB_X1Y117_I),
.O(LIOB33_X0Y169_IOB_X0Y169_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y169_IOB_X0Y170_OBUF (
.I(RIOB33_X105Y117_IOB_X1Y118_I),
.O(LIOB33_X0Y169_IOB_X0Y170_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y171_IOB_X0Y171_OBUF (
.I(RIOB33_X105Y119_IOB_X1Y119_I),
.O(LIOB33_X0Y171_IOB_X0Y171_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y171_IOB_X0Y172_OBUF (
.I(RIOB33_X105Y119_IOB_X1Y120_I),
.O(LIOB33_X0Y171_IOB_X0Y172_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y173_IOB_X0Y173_OBUF (
.I(RIOB33_X105Y121_IOB_X1Y121_I),
.O(LIOB33_X0Y173_IOB_X0Y173_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y173_IOB_X0Y174_OBUF (
.I(RIOB33_X105Y121_IOB_X1Y122_I),
.O(LIOB33_X0Y173_IOB_X0Y174_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y175_IOB_X0Y175_OBUF (
.I(RIOB33_X105Y123_IOB_X1Y123_I),
.O(LIOB33_X0Y175_IOB_X0Y175_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y175_IOB_X0Y176_OBUF (
.I(RIOB33_X105Y115_IOB_X1Y116_I),
.O(LIOB33_X0Y175_IOB_X0Y176_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y177_IOB_X0Y177_OBUF (
.I(RIOB33_X105Y123_IOB_X1Y124_I),
.O(LIOB33_X0Y177_IOB_X0Y177_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y177_IOB_X0Y178_OBUF (
.I(RIOB33_X105Y125_IOB_X1Y125_I),
.O(LIOB33_X0Y177_IOB_X0Y178_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y179_IOB_X0Y179_OBUF (
.I(RIOB33_X105Y125_IOB_X1Y126_I),
.O(LIOB33_X0Y179_IOB_X0Y179_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y179_IOB_X0Y180_OBUF (
.I(RIOB33_X105Y127_IOB_X1Y127_I),
.O(LIOB33_X0Y179_IOB_X0Y180_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y181_IOB_X0Y181_OBUF (
.I(RIOB33_X105Y127_IOB_X1Y128_I),
.O(LIOB33_X0Y181_IOB_X0Y181_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y181_IOB_X0Y182_OBUF (
.I(RIOB33_X105Y129_IOB_X1Y129_I),
.O(LIOB33_X0Y181_IOB_X0Y182_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y183_IOB_X0Y183_OBUF (
.I(RIOB33_X105Y129_IOB_X1Y130_I),
.O(LIOB33_X0Y183_IOB_X0Y183_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y183_IOB_X0Y184_OBUF (
.I(RIOB33_X105Y131_IOB_X1Y132_I),
.O(LIOB33_X0Y183_IOB_X0Y184_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y185_IOB_X0Y185_OBUF (
.I(RIOB33_X105Y133_IOB_X1Y133_I),
.O(LIOB33_X0Y185_IOB_X0Y185_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y185_IOB_X0Y186_OBUF (
.I(RIOB33_X105Y119_IOB_X1Y120_I),
.O(LIOB33_X0Y185_IOB_X0Y186_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y187_IOB_X0Y187_OBUF (
.I(CLBLM_L_X8Y145_SLICE_X11Y145_DQ),
.O(LIOB33_X0Y187_IOB_X0Y187_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y187_IOB_X0Y188_OBUF (
.I(CLBLM_R_X5Y147_SLICE_X6Y147_AQ),
.O(LIOB33_X0Y187_IOB_X0Y188_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y189_IOB_X0Y189_OBUF (
.I(CLBLM_L_X8Y147_SLICE_X10Y147_BQ),
.O(LIOB33_X0Y189_IOB_X0Y189_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y189_IOB_X0Y190_OBUF (
.I(CLBLM_L_X10Y154_SLICE_X12Y154_CO5),
.O(LIOB33_X0Y189_IOB_X0Y190_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y191_IOB_X0Y191_OBUF (
.I(CLBLL_L_X2Y148_SLICE_X1Y148_CO6),
.O(LIOB33_X0Y191_IOB_X0Y191_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y191_IOB_X0Y192_OBUF (
.I(CLBLL_L_X4Y153_SLICE_X4Y153_DO5),
.O(LIOB33_X0Y191_IOB_X0Y192_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y193_IOB_X0Y193_OBUF (
.I(CLBLL_L_X2Y166_SLICE_X0Y166_AO6),
.O(LIOB33_X0Y193_IOB_X0Y193_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y193_IOB_X0Y194_OBUF (
.I(RIOB33_X105Y103_IOB_X1Y103_I),
.O(LIOB33_X0Y193_IOB_X0Y194_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y195_IOB_X0Y195_OBUF (
.I(CLBLM_R_X3Y151_SLICE_X2Y151_AO5),
.O(LIOB33_X0Y195_IOB_X0Y195_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y195_IOB_X0Y196_OBUF (
.I(CLBLM_R_X3Y148_SLICE_X3Y148_DO5),
.O(LIOB33_X0Y195_IOB_X0Y196_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y197_IOB_X0Y197_OBUF (
.I(CLBLL_L_X4Y153_SLICE_X4Y153_CO5),
.O(LIOB33_X0Y197_IOB_X0Y197_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y197_IOB_X0Y198_OBUF (
.I(1'b1),
.O(LIOB33_X0Y197_IOB_X0Y198_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_SING_X0Y50_IOB_X0Y50_IBUF (
.I(LIOB33_SING_X0Y50_IOB_X0Y50_IPAD),
.O(LIOB33_SING_X0Y50_IOB_X0Y50_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_SING_X0Y100_IOB_X0Y100_OBUF (
.I(CLBLM_R_X3Y148_SLICE_X2Y148_B5Q),
.O(LIOB33_SING_X0Y100_IOB_X0Y100_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_SING_X0Y149_IOB_X0Y149_OBUF (
.I(RIOB33_X105Y115_IOB_X1Y115_I),
.O(LIOB33_SING_X0Y149_IOB_X0Y149_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_SING_X0Y150_IOB_X0Y150_OBUF (
.I(CLBLM_R_X3Y144_SLICE_X2Y144_AO5),
.O(LIOB33_SING_X0Y150_IOB_X0Y150_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_SING_X0Y199_IOB_X0Y199_OBUF (
.I(1'b1),
.O(LIOB33_SING_X0Y199_IOB_X0Y199_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y101_IOB_X1Y101_IBUF (
.I(RIOB33_X105Y101_IOB_X1Y101_IPAD),
.O(RIOB33_X105Y101_IOB_X1Y101_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y101_IOB_X1Y102_IBUF (
.I(RIOB33_X105Y101_IOB_X1Y102_IPAD),
.O(RIOB33_X105Y101_IOB_X1Y102_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y103_IOB_X1Y103_IBUF (
.I(RIOB33_X105Y103_IOB_X1Y103_IPAD),
.O(RIOB33_X105Y103_IOB_X1Y103_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y103_IOB_X1Y104_IBUF (
.I(RIOB33_X105Y103_IOB_X1Y104_IPAD),
.O(RIOB33_X105Y103_IOB_X1Y104_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y105_IOB_X1Y105_IBUF (
.I(RIOB33_X105Y105_IOB_X1Y105_IPAD),
.O(RIOB33_X105Y105_IOB_X1Y105_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y105_IOB_X1Y106_IBUF (
.I(RIOB33_X105Y105_IOB_X1Y106_IPAD),
.O(RIOB33_X105Y105_IOB_X1Y106_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y107_IOB_X1Y107_IBUF (
.I(RIOB33_X105Y107_IOB_X1Y107_IPAD),
.O(RIOB33_X105Y107_IOB_X1Y107_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y107_IOB_X1Y108_IBUF (
.I(RIOB33_X105Y107_IOB_X1Y108_IPAD),
.O(RIOB33_X105Y107_IOB_X1Y108_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y109_IOB_X1Y109_IBUF (
.I(RIOB33_X105Y109_IOB_X1Y109_IPAD),
.O(RIOB33_X105Y109_IOB_X1Y109_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y109_IOB_X1Y110_IBUF (
.I(RIOB33_X105Y109_IOB_X1Y110_IPAD),
.O(RIOB33_X105Y109_IOB_X1Y110_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y111_IOB_X1Y111_IBUF (
.I(RIOB33_X105Y111_IOB_X1Y111_IPAD),
.O(RIOB33_X105Y111_IOB_X1Y111_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y111_IOB_X1Y112_IBUF (
.I(RIOB33_X105Y111_IOB_X1Y112_IPAD),
.O(RIOB33_X105Y111_IOB_X1Y112_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y113_IOB_X1Y113_IBUF (
.I(RIOB33_X105Y113_IOB_X1Y113_IPAD),
.O(RIOB33_X105Y113_IOB_X1Y113_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y113_IOB_X1Y114_IBUF (
.I(RIOB33_X105Y113_IOB_X1Y114_IPAD),
.O(RIOB33_X105Y113_IOB_X1Y114_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y115_IOB_X1Y115_IBUF (
.I(RIOB33_X105Y115_IOB_X1Y115_IPAD),
.O(RIOB33_X105Y115_IOB_X1Y115_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y115_IOB_X1Y116_IBUF (
.I(RIOB33_X105Y115_IOB_X1Y116_IPAD),
.O(RIOB33_X105Y115_IOB_X1Y116_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y117_IOB_X1Y117_IBUF (
.I(RIOB33_X105Y117_IOB_X1Y117_IPAD),
.O(RIOB33_X105Y117_IOB_X1Y117_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y117_IOB_X1Y118_IBUF (
.I(RIOB33_X105Y117_IOB_X1Y118_IPAD),
.O(RIOB33_X105Y117_IOB_X1Y118_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y119_IOB_X1Y119_IBUF (
.I(RIOB33_X105Y119_IOB_X1Y119_IPAD),
.O(RIOB33_X105Y119_IOB_X1Y119_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y119_IOB_X1Y120_IBUF (
.I(RIOB33_X105Y119_IOB_X1Y120_IPAD),
.O(RIOB33_X105Y119_IOB_X1Y120_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y121_IOB_X1Y121_IBUF (
.I(RIOB33_X105Y121_IOB_X1Y121_IPAD),
.O(RIOB33_X105Y121_IOB_X1Y121_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y121_IOB_X1Y122_IBUF (
.I(RIOB33_X105Y121_IOB_X1Y122_IPAD),
.O(RIOB33_X105Y121_IOB_X1Y122_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y123_IOB_X1Y123_IBUF (
.I(RIOB33_X105Y123_IOB_X1Y123_IPAD),
.O(RIOB33_X105Y123_IOB_X1Y123_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y123_IOB_X1Y124_IBUF (
.I(RIOB33_X105Y123_IOB_X1Y124_IPAD),
.O(RIOB33_X105Y123_IOB_X1Y124_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y125_IOB_X1Y125_IBUF (
.I(RIOB33_X105Y125_IOB_X1Y125_IPAD),
.O(RIOB33_X105Y125_IOB_X1Y125_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y125_IOB_X1Y126_IBUF (
.I(RIOB33_X105Y125_IOB_X1Y126_IPAD),
.O(RIOB33_X105Y125_IOB_X1Y126_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y127_IOB_X1Y127_IBUF (
.I(RIOB33_X105Y127_IOB_X1Y127_IPAD),
.O(RIOB33_X105Y127_IOB_X1Y127_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y127_IOB_X1Y128_IBUF (
.I(RIOB33_X105Y127_IOB_X1Y128_IPAD),
.O(RIOB33_X105Y127_IOB_X1Y128_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y129_IOB_X1Y129_IBUF (
.I(RIOB33_X105Y129_IOB_X1Y129_IPAD),
.O(RIOB33_X105Y129_IOB_X1Y129_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y129_IOB_X1Y130_IBUF (
.I(RIOB33_X105Y129_IOB_X1Y130_IPAD),
.O(RIOB33_X105Y129_IOB_X1Y130_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y131_IOB_X1Y131_IBUF (
.I(RIOB33_X105Y131_IOB_X1Y131_IPAD),
.O(RIOB33_X105Y131_IOB_X1Y131_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y131_IOB_X1Y132_IBUF (
.I(RIOB33_X105Y131_IOB_X1Y132_IPAD),
.O(RIOB33_X105Y131_IOB_X1Y132_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y133_IOB_X1Y133_IBUF (
.I(RIOB33_X105Y133_IOB_X1Y133_IPAD),
.O(RIOB33_X105Y133_IOB_X1Y133_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y133_IOB_X1Y134_IBUF (
.I(RIOB33_X105Y133_IOB_X1Y134_IPAD),
.O(RIOB33_X105Y133_IOB_X1Y134_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y135_IOB_X1Y135_IBUF (
.I(RIOB33_X105Y135_IOB_X1Y135_IPAD),
.O(RIOB33_X105Y135_IOB_X1Y135_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y135_IOB_X1Y136_IBUF (
.I(RIOB33_X105Y135_IOB_X1Y136_IPAD),
.O(RIOB33_X105Y135_IOB_X1Y136_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y137_IOB_X1Y137_IBUF (
.I(RIOB33_X105Y137_IOB_X1Y137_IPAD),
.O(RIOB33_X105Y137_IOB_X1Y137_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y137_IOB_X1Y138_IBUF (
.I(RIOB33_X105Y137_IOB_X1Y138_IPAD),
.O(RIOB33_X105Y137_IOB_X1Y138_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y139_IOB_X1Y139_IBUF (
.I(RIOB33_X105Y139_IOB_X1Y139_IPAD),
.O(RIOB33_X105Y139_IOB_X1Y139_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y139_IOB_X1Y140_IBUF (
.I(RIOB33_X105Y139_IOB_X1Y140_IPAD),
.O(RIOB33_X105Y139_IOB_X1Y140_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y141_IOB_X1Y141_IBUF (
.I(RIOB33_X105Y141_IOB_X1Y141_IPAD),
.O(RIOB33_X105Y141_IOB_X1Y141_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y141_IOB_X1Y142_IBUF (
.I(RIOB33_X105Y141_IOB_X1Y142_IPAD),
.O(RIOB33_X105Y141_IOB_X1Y142_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y143_IOB_X1Y143_IBUF (
.I(RIOB33_X105Y143_IOB_X1Y143_IPAD),
.O(RIOB33_X105Y143_IOB_X1Y143_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y143_IOB_X1Y144_IBUF (
.I(RIOB33_X105Y143_IOB_X1Y144_IPAD),
.O(RIOB33_X105Y143_IOB_X1Y144_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y145_IOB_X1Y145_IBUF (
.I(RIOB33_X105Y145_IOB_X1Y145_IPAD),
.O(RIOB33_X105Y145_IOB_X1Y145_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y145_IOB_X1Y146_IBUF (
.I(RIOB33_X105Y145_IOB_X1Y146_IPAD),
.O(RIOB33_X105Y145_IOB_X1Y146_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y147_IOB_X1Y147_IBUF (
.I(RIOB33_X105Y147_IOB_X1Y147_IPAD),
.O(RIOB33_X105Y147_IOB_X1Y147_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y147_IOB_X1Y148_IBUF (
.I(RIOB33_X105Y147_IOB_X1Y148_IPAD),
.O(RIOB33_X105Y147_IOB_X1Y148_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y151_IOB_X1Y151_OBUF (
.I(1'b1),
.O(RIOB33_X105Y151_IOB_X1Y151_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y151_IOB_X1Y152_OBUF (
.I(1'b1),
.O(RIOB33_X105Y151_IOB_X1Y152_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y153_IOB_X1Y153_OBUF (
.I(1'b1),
.O(RIOB33_X105Y153_IOB_X1Y153_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y153_IOB_X1Y154_OBUF (
.I(1'b1),
.O(RIOB33_X105Y153_IOB_X1Y154_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y155_IOB_X1Y155_OBUF (
.I(1'b1),
.O(RIOB33_X105Y155_IOB_X1Y155_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y155_IOB_X1Y156_OBUF (
.I(1'b1),
.O(RIOB33_X105Y155_IOB_X1Y156_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y157_IOB_X1Y157_OBUF (
.I(1'b1),
.O(RIOB33_X105Y157_IOB_X1Y157_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y157_IOB_X1Y158_OBUF (
.I(1'b1),
.O(RIOB33_X105Y157_IOB_X1Y158_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y159_IOB_X1Y159_OBUF (
.I(1'b1),
.O(RIOB33_X105Y159_IOB_X1Y159_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y159_IOB_X1Y160_OBUF (
.I(1'b1),
.O(RIOB33_X105Y159_IOB_X1Y160_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y161_IOB_X1Y161_OBUF (
.I(CLBLM_L_X10Y154_SLICE_X12Y154_DO5),
.O(RIOB33_X105Y161_IOB_X1Y161_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y161_IOB_X1Y162_OBUF (
.I(CLBLM_R_X7Y153_SLICE_X9Y153_C5Q),
.O(RIOB33_X105Y161_IOB_X1Y162_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y163_IOB_X1Y163_OBUF (
.I(CLBLM_R_X7Y151_SLICE_X9Y151_D5Q),
.O(RIOB33_X105Y163_IOB_X1Y163_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y163_IOB_X1Y164_OBUF (
.I(CLBLM_L_X10Y153_SLICE_X12Y153_AQ),
.O(RIOB33_X105Y163_IOB_X1Y164_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y165_IOB_X1Y165_OBUF (
.I(CLBLM_L_X12Y152_SLICE_X16Y152_AO6),
.O(RIOB33_X105Y165_IOB_X1Y165_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y165_IOB_X1Y166_OBUF (
.I(CLBLM_L_X8Y153_SLICE_X10Y153_A5Q),
.O(RIOB33_X105Y165_IOB_X1Y166_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y167_IOB_X1Y167_OBUF (
.I(CLBLM_R_X7Y153_SLICE_X9Y153_DQ),
.O(RIOB33_X105Y167_IOB_X1Y167_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y167_IOB_X1Y168_OBUF (
.I(CLBLM_R_X5Y154_SLICE_X7Y154_AQ),
.O(RIOB33_X105Y167_IOB_X1Y168_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y169_IOB_X1Y169_OBUF (
.I(CLBLM_R_X3Y152_SLICE_X3Y152_CQ),
.O(RIOB33_X105Y169_IOB_X1Y169_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y169_IOB_X1Y170_OBUF (
.I(CLBLM_R_X3Y152_SLICE_X3Y152_BQ),
.O(RIOB33_X105Y169_IOB_X1Y170_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y171_IOB_X1Y171_OBUF (
.I(CLBLM_L_X8Y153_SLICE_X11Y153_DO6),
.O(RIOB33_X105Y171_IOB_X1Y171_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y171_IOB_X1Y172_OBUF (
.I(CLBLL_L_X2Y148_SLICE_X0Y148_AQ),
.O(RIOB33_X105Y171_IOB_X1Y172_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y173_IOB_X1Y173_OBUF (
.I(CLBLM_R_X5Y152_SLICE_X7Y152_DQ),
.O(RIOB33_X105Y173_IOB_X1Y173_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y173_IOB_X1Y174_OBUF (
.I(CLBLM_R_X5Y152_SLICE_X7Y152_DO6),
.O(RIOB33_X105Y173_IOB_X1Y174_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y175_IOB_X1Y175_OBUF (
.I(CLBLM_L_X10Y144_SLICE_X12Y144_BO6),
.O(RIOB33_X105Y175_IOB_X1Y175_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y175_IOB_X1Y176_OBUF (
.I(CLBLL_L_X2Y148_SLICE_X1Y148_BO6),
.O(RIOB33_X105Y175_IOB_X1Y176_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y177_IOB_X1Y177_OBUF (
.I(CLBLL_L_X2Y146_SLICE_X1Y146_B5Q),
.O(RIOB33_X105Y177_IOB_X1Y177_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y177_IOB_X1Y178_OBUF (
.I(CLBLM_R_X5Y147_SLICE_X6Y147_AQ),
.O(RIOB33_X105Y177_IOB_X1Y178_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y179_IOB_X1Y179_OBUF (
.I(CLBLM_L_X8Y147_SLICE_X10Y147_BQ),
.O(RIOB33_X105Y179_IOB_X1Y179_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y179_IOB_X1Y180_OBUF (
.I(CLBLM_L_X8Y145_SLICE_X11Y145_DQ),
.O(RIOB33_X105Y179_IOB_X1Y180_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y181_IOB_X1Y181_OBUF (
.I(CLBLM_L_X10Y154_SLICE_X12Y154_CO5),
.O(RIOB33_X105Y181_IOB_X1Y181_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y181_IOB_X1Y182_OBUF (
.I(CLBLM_R_X11Y146_SLICE_X14Y146_BO5),
.O(RIOB33_X105Y181_IOB_X1Y182_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y183_IOB_X1Y183_OBUF (
.I(1'b0),
.O(RIOB33_X105Y183_IOB_X1Y183_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y183_IOB_X1Y184_OBUF (
.I(CLBLM_R_X3Y148_SLICE_X3Y148_DO5),
.O(RIOB33_X105Y183_IOB_X1Y184_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y185_IOB_X1Y185_OBUF (
.I(CLBLM_L_X10Y153_SLICE_X12Y153_DO6),
.O(RIOB33_X105Y185_IOB_X1Y185_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y185_IOB_X1Y186_OBUF (
.I(CLBLM_L_X10Y149_SLICE_X13Y149_BO6),
.O(RIOB33_X105Y185_IOB_X1Y186_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y187_IOB_X1Y187_OBUF (
.I(CLBLM_R_X103Y178_SLICE_X163Y178_AO6),
.O(RIOB33_X105Y187_IOB_X1Y187_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y187_IOB_X1Y188_OBUF (
.I(CLBLM_R_X11Y146_SLICE_X14Y146_BO5),
.O(RIOB33_X105Y187_IOB_X1Y188_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y189_IOB_X1Y189_OBUF (
.I(CLBLM_R_X103Y178_SLICE_X163Y178_AO6),
.O(RIOB33_X105Y189_IOB_X1Y189_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y189_IOB_X1Y190_OBUF (
.I(CLBLM_L_X12Y151_SLICE_X16Y151_AO5),
.O(RIOB33_X105Y189_IOB_X1Y190_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y191_IOB_X1Y191_OBUF (
.I(CLBLM_L_X12Y149_SLICE_X17Y149_AO5),
.O(RIOB33_X105Y191_IOB_X1Y191_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y191_IOB_X1Y192_OBUF (
.I(CLBLM_L_X12Y153_SLICE_X16Y153_AO6),
.O(RIOB33_X105Y191_IOB_X1Y192_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y193_IOB_X1Y193_OBUF (
.I(CLBLM_L_X12Y151_SLICE_X16Y151_BO5),
.O(RIOB33_X105Y193_IOB_X1Y193_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y193_IOB_X1Y194_OBUF (
.I(CLBLM_L_X12Y151_SLICE_X16Y151_BO6),
.O(RIOB33_X105Y193_IOB_X1Y194_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y195_IOB_X1Y195_OBUF (
.I(CLBLM_L_X10Y149_SLICE_X13Y149_AO5),
.O(RIOB33_X105Y195_IOB_X1Y195_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y195_IOB_X1Y196_OBUF (
.I(CLBLM_L_X12Y150_SLICE_X16Y150_AO6),
.O(RIOB33_X105Y195_IOB_X1Y196_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y197_IOB_X1Y197_OBUF (
.I(CLBLM_L_X12Y152_SLICE_X16Y152_AO5),
.O(RIOB33_X105Y197_IOB_X1Y197_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y197_IOB_X1Y198_OBUF (
.I(CLBLM_L_X12Y150_SLICE_X16Y150_AO5),
.O(RIOB33_X105Y197_IOB_X1Y198_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_SING_X105Y100_IOB_X1Y100_IBUF (
.I(RIOB33_SING_X105Y100_IOB_X1Y100_IPAD),
.O(RIOB33_SING_X105Y100_IOB_X1Y100_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_SING_X105Y149_IOB_X1Y149_IBUF (
.I(RIOB33_SING_X105Y149_IOB_X1Y149_IPAD),
.O(RIOB33_SING_X105Y149_IOB_X1Y149_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_SING_X105Y150_IOB_X1Y150_OBUF (
.I(1'b1),
.O(RIOB33_SING_X105Y150_IOB_X1Y150_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_SING_X105Y199_IOB_X1Y199_OBUF (
.I(CLBLM_R_X7Y153_SLICE_X8Y153_A5Q),
.O(RIOB33_SING_X105Y199_IOB_X1Y199_OPAD)
  );
  assign CLBLL_L_X2Y75_SLICE_X0Y75_A = CLBLL_L_X2Y75_SLICE_X0Y75_AO6;
  assign CLBLL_L_X2Y75_SLICE_X0Y75_B = CLBLL_L_X2Y75_SLICE_X0Y75_BO6;
  assign CLBLL_L_X2Y75_SLICE_X0Y75_C = CLBLL_L_X2Y75_SLICE_X0Y75_CO6;
  assign CLBLL_L_X2Y75_SLICE_X0Y75_D = CLBLL_L_X2Y75_SLICE_X0Y75_DO6;
  assign CLBLL_L_X2Y75_SLICE_X1Y75_A = CLBLL_L_X2Y75_SLICE_X1Y75_AO6;
  assign CLBLL_L_X2Y75_SLICE_X1Y75_B = CLBLL_L_X2Y75_SLICE_X1Y75_BO6;
  assign CLBLL_L_X2Y75_SLICE_X1Y75_C = CLBLL_L_X2Y75_SLICE_X1Y75_CO6;
  assign CLBLL_L_X2Y75_SLICE_X1Y75_D = CLBLL_L_X2Y75_SLICE_X1Y75_DO6;
  assign CLBLL_L_X2Y144_SLICE_X0Y144_A = CLBLL_L_X2Y144_SLICE_X0Y144_AO6;
  assign CLBLL_L_X2Y144_SLICE_X0Y144_B = CLBLL_L_X2Y144_SLICE_X0Y144_BO6;
  assign CLBLL_L_X2Y144_SLICE_X0Y144_C = CLBLL_L_X2Y144_SLICE_X0Y144_CO6;
  assign CLBLL_L_X2Y144_SLICE_X0Y144_D = CLBLL_L_X2Y144_SLICE_X0Y144_DO6;
  assign CLBLL_L_X2Y144_SLICE_X1Y144_A = CLBLL_L_X2Y144_SLICE_X1Y144_AO6;
  assign CLBLL_L_X2Y144_SLICE_X1Y144_B = CLBLL_L_X2Y144_SLICE_X1Y144_BO6;
  assign CLBLL_L_X2Y144_SLICE_X1Y144_C = CLBLL_L_X2Y144_SLICE_X1Y144_CO6;
  assign CLBLL_L_X2Y144_SLICE_X1Y144_D = CLBLL_L_X2Y144_SLICE_X1Y144_DO6;
  assign CLBLL_L_X2Y145_SLICE_X0Y145_A = CLBLL_L_X2Y145_SLICE_X0Y145_AO6;
  assign CLBLL_L_X2Y145_SLICE_X0Y145_B = CLBLL_L_X2Y145_SLICE_X0Y145_BO6;
  assign CLBLL_L_X2Y145_SLICE_X0Y145_C = CLBLL_L_X2Y145_SLICE_X0Y145_CO6;
  assign CLBLL_L_X2Y145_SLICE_X0Y145_D = CLBLL_L_X2Y145_SLICE_X0Y145_DO6;
  assign CLBLL_L_X2Y145_SLICE_X1Y145_A = CLBLL_L_X2Y145_SLICE_X1Y145_AO6;
  assign CLBLL_L_X2Y145_SLICE_X1Y145_B = CLBLL_L_X2Y145_SLICE_X1Y145_BO6;
  assign CLBLL_L_X2Y145_SLICE_X1Y145_C = CLBLL_L_X2Y145_SLICE_X1Y145_CO6;
  assign CLBLL_L_X2Y145_SLICE_X1Y145_D = CLBLL_L_X2Y145_SLICE_X1Y145_DO6;
  assign CLBLL_L_X2Y145_SLICE_X1Y145_DMUX = CLBLL_L_X2Y145_SLICE_X1Y145_DO5;
  assign CLBLL_L_X2Y146_SLICE_X0Y146_A = CLBLL_L_X2Y146_SLICE_X0Y146_AO6;
  assign CLBLL_L_X2Y146_SLICE_X0Y146_B = CLBLL_L_X2Y146_SLICE_X0Y146_BO6;
  assign CLBLL_L_X2Y146_SLICE_X0Y146_C = CLBLL_L_X2Y146_SLICE_X0Y146_CO6;
  assign CLBLL_L_X2Y146_SLICE_X0Y146_D = CLBLL_L_X2Y146_SLICE_X0Y146_DO6;
  assign CLBLL_L_X2Y146_SLICE_X1Y146_A = CLBLL_L_X2Y146_SLICE_X1Y146_AO6;
  assign CLBLL_L_X2Y146_SLICE_X1Y146_B = CLBLL_L_X2Y146_SLICE_X1Y146_BO6;
  assign CLBLL_L_X2Y146_SLICE_X1Y146_C = CLBLL_L_X2Y146_SLICE_X1Y146_CO6;
  assign CLBLL_L_X2Y146_SLICE_X1Y146_D = CLBLL_L_X2Y146_SLICE_X1Y146_DO6;
  assign CLBLL_L_X2Y146_SLICE_X1Y146_BMUX = CLBLL_L_X2Y146_SLICE_X1Y146_B5Q;
  assign CLBLL_L_X2Y146_SLICE_X1Y146_CMUX = CLBLL_L_X2Y146_SLICE_X1Y146_CO5;
  assign CLBLL_L_X2Y147_SLICE_X0Y147_A = CLBLL_L_X2Y147_SLICE_X0Y147_AO6;
  assign CLBLL_L_X2Y147_SLICE_X0Y147_B = CLBLL_L_X2Y147_SLICE_X0Y147_BO6;
  assign CLBLL_L_X2Y147_SLICE_X0Y147_C = CLBLL_L_X2Y147_SLICE_X0Y147_CO6;
  assign CLBLL_L_X2Y147_SLICE_X0Y147_D = CLBLL_L_X2Y147_SLICE_X0Y147_DO6;
  assign CLBLL_L_X2Y147_SLICE_X1Y147_A = CLBLL_L_X2Y147_SLICE_X1Y147_AO6;
  assign CLBLL_L_X2Y147_SLICE_X1Y147_B = CLBLL_L_X2Y147_SLICE_X1Y147_BO6;
  assign CLBLL_L_X2Y147_SLICE_X1Y147_C = CLBLL_L_X2Y147_SLICE_X1Y147_CO6;
  assign CLBLL_L_X2Y147_SLICE_X1Y147_D = CLBLL_L_X2Y147_SLICE_X1Y147_DO6;
  assign CLBLL_L_X2Y148_SLICE_X0Y148_A = CLBLL_L_X2Y148_SLICE_X0Y148_AO6;
  assign CLBLL_L_X2Y148_SLICE_X0Y148_B = CLBLL_L_X2Y148_SLICE_X0Y148_BO6;
  assign CLBLL_L_X2Y148_SLICE_X0Y148_C = CLBLL_L_X2Y148_SLICE_X0Y148_CO6;
  assign CLBLL_L_X2Y148_SLICE_X0Y148_D = CLBLL_L_X2Y148_SLICE_X0Y148_DO6;
  assign CLBLL_L_X2Y148_SLICE_X1Y148_A = CLBLL_L_X2Y148_SLICE_X1Y148_AO6;
  assign CLBLL_L_X2Y148_SLICE_X1Y148_B = CLBLL_L_X2Y148_SLICE_X1Y148_BO6;
  assign CLBLL_L_X2Y148_SLICE_X1Y148_C = CLBLL_L_X2Y148_SLICE_X1Y148_CO6;
  assign CLBLL_L_X2Y148_SLICE_X1Y148_D = CLBLL_L_X2Y148_SLICE_X1Y148_DO6;
  assign CLBLL_L_X2Y150_SLICE_X0Y150_A = CLBLL_L_X2Y150_SLICE_X0Y150_AO6;
  assign CLBLL_L_X2Y150_SLICE_X0Y150_B = CLBLL_L_X2Y150_SLICE_X0Y150_BO6;
  assign CLBLL_L_X2Y150_SLICE_X0Y150_C = CLBLL_L_X2Y150_SLICE_X0Y150_CO6;
  assign CLBLL_L_X2Y150_SLICE_X0Y150_D = CLBLL_L_X2Y150_SLICE_X0Y150_DO6;
  assign CLBLL_L_X2Y150_SLICE_X1Y150_A = CLBLL_L_X2Y150_SLICE_X1Y150_AO6;
  assign CLBLL_L_X2Y150_SLICE_X1Y150_B = CLBLL_L_X2Y150_SLICE_X1Y150_BO6;
  assign CLBLL_L_X2Y150_SLICE_X1Y150_C = CLBLL_L_X2Y150_SLICE_X1Y150_CO6;
  assign CLBLL_L_X2Y150_SLICE_X1Y150_D = CLBLL_L_X2Y150_SLICE_X1Y150_DO6;
  assign CLBLL_L_X2Y166_SLICE_X0Y166_A = CLBLL_L_X2Y166_SLICE_X0Y166_AO6;
  assign CLBLL_L_X2Y166_SLICE_X0Y166_B = CLBLL_L_X2Y166_SLICE_X0Y166_BO6;
  assign CLBLL_L_X2Y166_SLICE_X0Y166_C = CLBLL_L_X2Y166_SLICE_X0Y166_CO6;
  assign CLBLL_L_X2Y166_SLICE_X0Y166_D = CLBLL_L_X2Y166_SLICE_X0Y166_DO6;
  assign CLBLL_L_X2Y166_SLICE_X1Y166_A = CLBLL_L_X2Y166_SLICE_X1Y166_AO6;
  assign CLBLL_L_X2Y166_SLICE_X1Y166_B = CLBLL_L_X2Y166_SLICE_X1Y166_BO6;
  assign CLBLL_L_X2Y166_SLICE_X1Y166_C = CLBLL_L_X2Y166_SLICE_X1Y166_CO6;
  assign CLBLL_L_X2Y166_SLICE_X1Y166_D = CLBLL_L_X2Y166_SLICE_X1Y166_DO6;
  assign CLBLL_L_X4Y140_SLICE_X4Y140_A = CLBLL_L_X4Y140_SLICE_X4Y140_AO6;
  assign CLBLL_L_X4Y140_SLICE_X4Y140_B = CLBLL_L_X4Y140_SLICE_X4Y140_BO6;
  assign CLBLL_L_X4Y140_SLICE_X4Y140_C = CLBLL_L_X4Y140_SLICE_X4Y140_CO6;
  assign CLBLL_L_X4Y140_SLICE_X4Y140_D = CLBLL_L_X4Y140_SLICE_X4Y140_DO6;
  assign CLBLL_L_X4Y140_SLICE_X4Y140_AMUX = CLBLL_L_X4Y140_SLICE_X4Y140_A5Q;
  assign CLBLL_L_X4Y140_SLICE_X4Y140_BMUX = CLBLL_L_X4Y140_SLICE_X4Y140_BO5;
  assign CLBLL_L_X4Y140_SLICE_X5Y140_A = CLBLL_L_X4Y140_SLICE_X5Y140_AO6;
  assign CLBLL_L_X4Y140_SLICE_X5Y140_B = CLBLL_L_X4Y140_SLICE_X5Y140_BO6;
  assign CLBLL_L_X4Y140_SLICE_X5Y140_C = CLBLL_L_X4Y140_SLICE_X5Y140_CO6;
  assign CLBLL_L_X4Y140_SLICE_X5Y140_D = CLBLL_L_X4Y140_SLICE_X5Y140_DO6;
  assign CLBLL_L_X4Y140_SLICE_X5Y140_CMUX = CLBLL_L_X4Y140_SLICE_X5Y140_CO5;
  assign CLBLL_L_X4Y142_SLICE_X4Y142_A = CLBLL_L_X4Y142_SLICE_X4Y142_AO6;
  assign CLBLL_L_X4Y142_SLICE_X4Y142_B = CLBLL_L_X4Y142_SLICE_X4Y142_BO6;
  assign CLBLL_L_X4Y142_SLICE_X4Y142_C = CLBLL_L_X4Y142_SLICE_X4Y142_CO6;
  assign CLBLL_L_X4Y142_SLICE_X4Y142_D = CLBLL_L_X4Y142_SLICE_X4Y142_DO6;
  assign CLBLL_L_X4Y142_SLICE_X4Y142_AMUX = CLBLL_L_X4Y142_SLICE_X4Y142_A5Q;
  assign CLBLL_L_X4Y142_SLICE_X5Y142_A = CLBLL_L_X4Y142_SLICE_X5Y142_AO6;
  assign CLBLL_L_X4Y142_SLICE_X5Y142_B = CLBLL_L_X4Y142_SLICE_X5Y142_BO6;
  assign CLBLL_L_X4Y142_SLICE_X5Y142_C = CLBLL_L_X4Y142_SLICE_X5Y142_CO6;
  assign CLBLL_L_X4Y142_SLICE_X5Y142_D = CLBLL_L_X4Y142_SLICE_X5Y142_DO6;
  assign CLBLL_L_X4Y142_SLICE_X5Y142_CMUX = CLBLL_L_X4Y142_SLICE_X5Y142_C5Q;
  assign CLBLL_L_X4Y142_SLICE_X5Y142_DMUX = CLBLL_L_X4Y142_SLICE_X5Y142_D5Q;
  assign CLBLL_L_X4Y143_SLICE_X4Y143_A = CLBLL_L_X4Y143_SLICE_X4Y143_AO6;
  assign CLBLL_L_X4Y143_SLICE_X4Y143_B = CLBLL_L_X4Y143_SLICE_X4Y143_BO6;
  assign CLBLL_L_X4Y143_SLICE_X4Y143_C = CLBLL_L_X4Y143_SLICE_X4Y143_CO6;
  assign CLBLL_L_X4Y143_SLICE_X4Y143_D = CLBLL_L_X4Y143_SLICE_X4Y143_DO6;
  assign CLBLL_L_X4Y143_SLICE_X4Y143_AMUX = CLBLL_L_X4Y143_SLICE_X4Y143_A5Q;
  assign CLBLL_L_X4Y143_SLICE_X4Y143_BMUX = CLBLL_L_X4Y143_SLICE_X4Y143_BO5;
  assign CLBLL_L_X4Y143_SLICE_X4Y143_CMUX = CLBLL_L_X4Y143_SLICE_X4Y143_C5Q;
  assign CLBLL_L_X4Y143_SLICE_X4Y143_DMUX = CLBLL_L_X4Y143_SLICE_X4Y143_D5Q;
  assign CLBLL_L_X4Y143_SLICE_X5Y143_A = CLBLL_L_X4Y143_SLICE_X5Y143_AO6;
  assign CLBLL_L_X4Y143_SLICE_X5Y143_B = CLBLL_L_X4Y143_SLICE_X5Y143_BO6;
  assign CLBLL_L_X4Y143_SLICE_X5Y143_C = CLBLL_L_X4Y143_SLICE_X5Y143_CO6;
  assign CLBLL_L_X4Y143_SLICE_X5Y143_D = CLBLL_L_X4Y143_SLICE_X5Y143_DO6;
  assign CLBLL_L_X4Y143_SLICE_X5Y143_BMUX = CLBLL_L_X4Y143_SLICE_X5Y143_B5Q;
  assign CLBLL_L_X4Y143_SLICE_X5Y143_CMUX = CLBLL_L_X4Y143_SLICE_X5Y143_CO5;
  assign CLBLL_L_X4Y143_SLICE_X5Y143_DMUX = CLBLL_L_X4Y143_SLICE_X5Y143_D5Q;
  assign CLBLL_L_X4Y144_SLICE_X4Y144_A = CLBLL_L_X4Y144_SLICE_X4Y144_AO6;
  assign CLBLL_L_X4Y144_SLICE_X4Y144_B = CLBLL_L_X4Y144_SLICE_X4Y144_BO6;
  assign CLBLL_L_X4Y144_SLICE_X4Y144_C = CLBLL_L_X4Y144_SLICE_X4Y144_CO6;
  assign CLBLL_L_X4Y144_SLICE_X4Y144_D = CLBLL_L_X4Y144_SLICE_X4Y144_DO6;
  assign CLBLL_L_X4Y144_SLICE_X4Y144_BMUX = CLBLL_L_X4Y144_SLICE_X4Y144_B5Q;
  assign CLBLL_L_X4Y144_SLICE_X4Y144_CMUX = CLBLL_L_X4Y144_SLICE_X4Y144_C5Q;
  assign CLBLL_L_X4Y144_SLICE_X4Y144_DMUX = CLBLL_L_X4Y144_SLICE_X4Y144_D5Q;
  assign CLBLL_L_X4Y144_SLICE_X5Y144_A = CLBLL_L_X4Y144_SLICE_X5Y144_AO6;
  assign CLBLL_L_X4Y144_SLICE_X5Y144_B = CLBLL_L_X4Y144_SLICE_X5Y144_BO6;
  assign CLBLL_L_X4Y144_SLICE_X5Y144_C = CLBLL_L_X4Y144_SLICE_X5Y144_CO6;
  assign CLBLL_L_X4Y144_SLICE_X5Y144_D = CLBLL_L_X4Y144_SLICE_X5Y144_DO6;
  assign CLBLL_L_X4Y144_SLICE_X5Y144_DMUX = CLBLL_L_X4Y144_SLICE_X5Y144_D5Q;
  assign CLBLL_L_X4Y145_SLICE_X4Y145_A = CLBLL_L_X4Y145_SLICE_X4Y145_AO6;
  assign CLBLL_L_X4Y145_SLICE_X4Y145_B = CLBLL_L_X4Y145_SLICE_X4Y145_BO6;
  assign CLBLL_L_X4Y145_SLICE_X4Y145_C = CLBLL_L_X4Y145_SLICE_X4Y145_CO6;
  assign CLBLL_L_X4Y145_SLICE_X4Y145_D = CLBLL_L_X4Y145_SLICE_X4Y145_DO6;
  assign CLBLL_L_X4Y145_SLICE_X4Y145_BMUX = CLBLL_L_X4Y145_SLICE_X4Y145_B5Q;
  assign CLBLL_L_X4Y145_SLICE_X4Y145_CMUX = CLBLL_L_X4Y145_SLICE_X4Y145_C5Q;
  assign CLBLL_L_X4Y145_SLICE_X4Y145_DMUX = CLBLL_L_X4Y145_SLICE_X4Y145_DO5;
  assign CLBLL_L_X4Y145_SLICE_X5Y145_A = CLBLL_L_X4Y145_SLICE_X5Y145_AO6;
  assign CLBLL_L_X4Y145_SLICE_X5Y145_B = CLBLL_L_X4Y145_SLICE_X5Y145_BO6;
  assign CLBLL_L_X4Y145_SLICE_X5Y145_C = CLBLL_L_X4Y145_SLICE_X5Y145_CO6;
  assign CLBLL_L_X4Y145_SLICE_X5Y145_D = CLBLL_L_X4Y145_SLICE_X5Y145_DO6;
  assign CLBLL_L_X4Y145_SLICE_X5Y145_CMUX = CLBLL_L_X4Y145_SLICE_X5Y145_C5Q;
  assign CLBLL_L_X4Y146_SLICE_X4Y146_A = CLBLL_L_X4Y146_SLICE_X4Y146_AO6;
  assign CLBLL_L_X4Y146_SLICE_X4Y146_B = CLBLL_L_X4Y146_SLICE_X4Y146_BO6;
  assign CLBLL_L_X4Y146_SLICE_X4Y146_C = CLBLL_L_X4Y146_SLICE_X4Y146_CO6;
  assign CLBLL_L_X4Y146_SLICE_X4Y146_D = CLBLL_L_X4Y146_SLICE_X4Y146_DO6;
  assign CLBLL_L_X4Y146_SLICE_X4Y146_BMUX = CLBLL_L_X4Y146_SLICE_X4Y146_B5Q;
  assign CLBLL_L_X4Y146_SLICE_X4Y146_CMUX = CLBLL_L_X4Y146_SLICE_X4Y146_C5Q;
  assign CLBLL_L_X4Y146_SLICE_X4Y146_DMUX = CLBLL_L_X4Y146_SLICE_X4Y146_DO5;
  assign CLBLL_L_X4Y146_SLICE_X5Y146_A = CLBLL_L_X4Y146_SLICE_X5Y146_AO6;
  assign CLBLL_L_X4Y146_SLICE_X5Y146_B = CLBLL_L_X4Y146_SLICE_X5Y146_BO6;
  assign CLBLL_L_X4Y146_SLICE_X5Y146_C = CLBLL_L_X4Y146_SLICE_X5Y146_CO6;
  assign CLBLL_L_X4Y146_SLICE_X5Y146_D = CLBLL_L_X4Y146_SLICE_X5Y146_DO6;
  assign CLBLL_L_X4Y146_SLICE_X5Y146_AMUX = CLBLL_L_X4Y146_SLICE_X5Y146_AO5;
  assign CLBLL_L_X4Y147_SLICE_X4Y147_A = CLBLL_L_X4Y147_SLICE_X4Y147_AO6;
  assign CLBLL_L_X4Y147_SLICE_X4Y147_B = CLBLL_L_X4Y147_SLICE_X4Y147_BO6;
  assign CLBLL_L_X4Y147_SLICE_X4Y147_C = CLBLL_L_X4Y147_SLICE_X4Y147_CO6;
  assign CLBLL_L_X4Y147_SLICE_X4Y147_D = CLBLL_L_X4Y147_SLICE_X4Y147_DO6;
  assign CLBLL_L_X4Y147_SLICE_X4Y147_BMUX = CLBLL_L_X4Y147_SLICE_X4Y147_B5Q;
  assign CLBLL_L_X4Y147_SLICE_X4Y147_CMUX = CLBLL_L_X4Y147_SLICE_X4Y147_C5Q;
  assign CLBLL_L_X4Y147_SLICE_X4Y147_DMUX = CLBLL_L_X4Y147_SLICE_X4Y147_D5Q;
  assign CLBLL_L_X4Y147_SLICE_X5Y147_A = CLBLL_L_X4Y147_SLICE_X5Y147_AO6;
  assign CLBLL_L_X4Y147_SLICE_X5Y147_B = CLBLL_L_X4Y147_SLICE_X5Y147_BO6;
  assign CLBLL_L_X4Y147_SLICE_X5Y147_C = CLBLL_L_X4Y147_SLICE_X5Y147_CO6;
  assign CLBLL_L_X4Y147_SLICE_X5Y147_D = CLBLL_L_X4Y147_SLICE_X5Y147_DO6;
  assign CLBLL_L_X4Y147_SLICE_X5Y147_BMUX = CLBLL_L_X4Y147_SLICE_X5Y147_B5Q;
  assign CLBLL_L_X4Y147_SLICE_X5Y147_CMUX = CLBLL_L_X4Y147_SLICE_X5Y147_C5Q;
  assign CLBLL_L_X4Y147_SLICE_X5Y147_DMUX = CLBLL_L_X4Y147_SLICE_X5Y147_DO6;
  assign CLBLL_L_X4Y148_SLICE_X4Y148_A = CLBLL_L_X4Y148_SLICE_X4Y148_AO6;
  assign CLBLL_L_X4Y148_SLICE_X4Y148_B = CLBLL_L_X4Y148_SLICE_X4Y148_BO6;
  assign CLBLL_L_X4Y148_SLICE_X4Y148_C = CLBLL_L_X4Y148_SLICE_X4Y148_CO6;
  assign CLBLL_L_X4Y148_SLICE_X4Y148_D = CLBLL_L_X4Y148_SLICE_X4Y148_DO6;
  assign CLBLL_L_X4Y148_SLICE_X4Y148_CMUX = CLBLL_L_X4Y148_SLICE_X4Y148_C5Q;
  assign CLBLL_L_X4Y148_SLICE_X5Y148_A = CLBLL_L_X4Y148_SLICE_X5Y148_AO6;
  assign CLBLL_L_X4Y148_SLICE_X5Y148_B = CLBLL_L_X4Y148_SLICE_X5Y148_BO6;
  assign CLBLL_L_X4Y148_SLICE_X5Y148_C = CLBLL_L_X4Y148_SLICE_X5Y148_CO6;
  assign CLBLL_L_X4Y148_SLICE_X5Y148_D = CLBLL_L_X4Y148_SLICE_X5Y148_DO6;
  assign CLBLL_L_X4Y148_SLICE_X5Y148_AMUX = CLBLL_L_X4Y148_SLICE_X5Y148_A5Q;
  assign CLBLL_L_X4Y148_SLICE_X5Y148_BMUX = CLBLL_L_X4Y148_SLICE_X5Y148_B5Q;
  assign CLBLL_L_X4Y148_SLICE_X5Y148_DMUX = CLBLL_L_X4Y148_SLICE_X5Y148_D5Q;
  assign CLBLL_L_X4Y149_SLICE_X4Y149_A = CLBLL_L_X4Y149_SLICE_X4Y149_AO6;
  assign CLBLL_L_X4Y149_SLICE_X4Y149_B = CLBLL_L_X4Y149_SLICE_X4Y149_BO6;
  assign CLBLL_L_X4Y149_SLICE_X4Y149_C = CLBLL_L_X4Y149_SLICE_X4Y149_CO6;
  assign CLBLL_L_X4Y149_SLICE_X4Y149_D = CLBLL_L_X4Y149_SLICE_X4Y149_DO6;
  assign CLBLL_L_X4Y149_SLICE_X4Y149_BMUX = CLBLL_L_X4Y149_SLICE_X4Y149_B5Q;
  assign CLBLL_L_X4Y149_SLICE_X4Y149_DMUX = CLBLL_L_X4Y149_SLICE_X4Y149_D5Q;
  assign CLBLL_L_X4Y149_SLICE_X5Y149_A = CLBLL_L_X4Y149_SLICE_X5Y149_AO6;
  assign CLBLL_L_X4Y149_SLICE_X5Y149_B = CLBLL_L_X4Y149_SLICE_X5Y149_BO6;
  assign CLBLL_L_X4Y149_SLICE_X5Y149_C = CLBLL_L_X4Y149_SLICE_X5Y149_CO6;
  assign CLBLL_L_X4Y149_SLICE_X5Y149_D = CLBLL_L_X4Y149_SLICE_X5Y149_DO6;
  assign CLBLL_L_X4Y149_SLICE_X5Y149_CMUX = CLBLL_L_X4Y149_SLICE_X5Y149_C5Q;
  assign CLBLL_L_X4Y150_SLICE_X4Y150_A = CLBLL_L_X4Y150_SLICE_X4Y150_AO6;
  assign CLBLL_L_X4Y150_SLICE_X4Y150_B = CLBLL_L_X4Y150_SLICE_X4Y150_BO6;
  assign CLBLL_L_X4Y150_SLICE_X4Y150_C = CLBLL_L_X4Y150_SLICE_X4Y150_CO6;
  assign CLBLL_L_X4Y150_SLICE_X4Y150_D = CLBLL_L_X4Y150_SLICE_X4Y150_DO6;
  assign CLBLL_L_X4Y150_SLICE_X4Y150_AMUX = CLBLL_L_X4Y150_SLICE_X4Y150_A5Q;
  assign CLBLL_L_X4Y150_SLICE_X4Y150_BMUX = CLBLL_L_X4Y150_SLICE_X4Y150_B5Q;
  assign CLBLL_L_X4Y150_SLICE_X4Y150_CMUX = CLBLL_L_X4Y150_SLICE_X4Y150_C5Q;
  assign CLBLL_L_X4Y150_SLICE_X5Y150_A = CLBLL_L_X4Y150_SLICE_X5Y150_AO6;
  assign CLBLL_L_X4Y150_SLICE_X5Y150_B = CLBLL_L_X4Y150_SLICE_X5Y150_BO6;
  assign CLBLL_L_X4Y150_SLICE_X5Y150_C = CLBLL_L_X4Y150_SLICE_X5Y150_CO6;
  assign CLBLL_L_X4Y150_SLICE_X5Y150_D = CLBLL_L_X4Y150_SLICE_X5Y150_DO6;
  assign CLBLL_L_X4Y150_SLICE_X5Y150_AMUX = CLBLL_L_X4Y150_SLICE_X5Y150_A5Q;
  assign CLBLL_L_X4Y150_SLICE_X5Y150_CMUX = CLBLL_L_X4Y150_SLICE_X5Y150_CO5;
  assign CLBLL_L_X4Y151_SLICE_X4Y151_A = CLBLL_L_X4Y151_SLICE_X4Y151_AO6;
  assign CLBLL_L_X4Y151_SLICE_X4Y151_B = CLBLL_L_X4Y151_SLICE_X4Y151_BO6;
  assign CLBLL_L_X4Y151_SLICE_X4Y151_C = CLBLL_L_X4Y151_SLICE_X4Y151_CO6;
  assign CLBLL_L_X4Y151_SLICE_X4Y151_D = CLBLL_L_X4Y151_SLICE_X4Y151_DO6;
  assign CLBLL_L_X4Y151_SLICE_X4Y151_AMUX = CLBLL_L_X4Y151_SLICE_X4Y151_A5Q;
  assign CLBLL_L_X4Y151_SLICE_X4Y151_BMUX = CLBLL_L_X4Y151_SLICE_X4Y151_B5Q;
  assign CLBLL_L_X4Y151_SLICE_X4Y151_CMUX = CLBLL_L_X4Y151_SLICE_X4Y151_C5Q;
  assign CLBLL_L_X4Y151_SLICE_X5Y151_A = CLBLL_L_X4Y151_SLICE_X5Y151_AO6;
  assign CLBLL_L_X4Y151_SLICE_X5Y151_B = CLBLL_L_X4Y151_SLICE_X5Y151_BO6;
  assign CLBLL_L_X4Y151_SLICE_X5Y151_C = CLBLL_L_X4Y151_SLICE_X5Y151_CO6;
  assign CLBLL_L_X4Y151_SLICE_X5Y151_D = CLBLL_L_X4Y151_SLICE_X5Y151_DO6;
  assign CLBLL_L_X4Y151_SLICE_X5Y151_BMUX = CLBLL_L_X4Y151_SLICE_X5Y151_B5Q;
  assign CLBLL_L_X4Y151_SLICE_X5Y151_DMUX = CLBLL_L_X4Y151_SLICE_X5Y151_D5Q;
  assign CLBLL_L_X4Y152_SLICE_X4Y152_A = CLBLL_L_X4Y152_SLICE_X4Y152_AO6;
  assign CLBLL_L_X4Y152_SLICE_X4Y152_B = CLBLL_L_X4Y152_SLICE_X4Y152_BO6;
  assign CLBLL_L_X4Y152_SLICE_X4Y152_C = CLBLL_L_X4Y152_SLICE_X4Y152_CO6;
  assign CLBLL_L_X4Y152_SLICE_X4Y152_D = CLBLL_L_X4Y152_SLICE_X4Y152_DO6;
  assign CLBLL_L_X4Y152_SLICE_X4Y152_BMUX = CLBLL_L_X4Y152_SLICE_X4Y152_B5Q;
  assign CLBLL_L_X4Y152_SLICE_X5Y152_A = CLBLL_L_X4Y152_SLICE_X5Y152_AO6;
  assign CLBLL_L_X4Y152_SLICE_X5Y152_B = CLBLL_L_X4Y152_SLICE_X5Y152_BO6;
  assign CLBLL_L_X4Y152_SLICE_X5Y152_C = CLBLL_L_X4Y152_SLICE_X5Y152_CO6;
  assign CLBLL_L_X4Y152_SLICE_X5Y152_D = CLBLL_L_X4Y152_SLICE_X5Y152_DO6;
  assign CLBLL_L_X4Y152_SLICE_X5Y152_AMUX = CLBLL_L_X4Y152_SLICE_X5Y152_A5Q;
  assign CLBLL_L_X4Y152_SLICE_X5Y152_CMUX = CLBLL_L_X4Y152_SLICE_X5Y152_CO5;
  assign CLBLL_L_X4Y153_SLICE_X4Y153_A = CLBLL_L_X4Y153_SLICE_X4Y153_AO6;
  assign CLBLL_L_X4Y153_SLICE_X4Y153_B = CLBLL_L_X4Y153_SLICE_X4Y153_BO6;
  assign CLBLL_L_X4Y153_SLICE_X4Y153_C = CLBLL_L_X4Y153_SLICE_X4Y153_CO6;
  assign CLBLL_L_X4Y153_SLICE_X4Y153_D = CLBLL_L_X4Y153_SLICE_X4Y153_DO6;
  assign CLBLL_L_X4Y153_SLICE_X4Y153_AMUX = CLBLL_L_X4Y153_SLICE_X4Y153_A5Q;
  assign CLBLL_L_X4Y153_SLICE_X4Y153_BMUX = CLBLL_L_X4Y153_SLICE_X4Y153_B5Q;
  assign CLBLL_L_X4Y153_SLICE_X4Y153_CMUX = CLBLL_L_X4Y153_SLICE_X4Y153_CO5;
  assign CLBLL_L_X4Y153_SLICE_X4Y153_DMUX = CLBLL_L_X4Y153_SLICE_X4Y153_DO5;
  assign CLBLL_L_X4Y153_SLICE_X5Y153_A = CLBLL_L_X4Y153_SLICE_X5Y153_AO6;
  assign CLBLL_L_X4Y153_SLICE_X5Y153_B = CLBLL_L_X4Y153_SLICE_X5Y153_BO6;
  assign CLBLL_L_X4Y153_SLICE_X5Y153_C = CLBLL_L_X4Y153_SLICE_X5Y153_CO6;
  assign CLBLL_L_X4Y153_SLICE_X5Y153_D = CLBLL_L_X4Y153_SLICE_X5Y153_DO6;
  assign CLBLL_L_X4Y153_SLICE_X5Y153_AMUX = CLBLL_L_X4Y153_SLICE_X5Y153_A5Q;
  assign CLBLL_L_X4Y153_SLICE_X5Y153_BMUX = CLBLL_L_X4Y153_SLICE_X5Y153_BO5;
  assign CLBLM_L_X8Y142_SLICE_X10Y142_A = CLBLM_L_X8Y142_SLICE_X10Y142_AO6;
  assign CLBLM_L_X8Y142_SLICE_X10Y142_B = CLBLM_L_X8Y142_SLICE_X10Y142_BO6;
  assign CLBLM_L_X8Y142_SLICE_X10Y142_C = CLBLM_L_X8Y142_SLICE_X10Y142_CO6;
  assign CLBLM_L_X8Y142_SLICE_X10Y142_D = CLBLM_L_X8Y142_SLICE_X10Y142_DO6;
  assign CLBLM_L_X8Y142_SLICE_X10Y142_AMUX = CLBLM_L_X8Y142_SLICE_X10Y142_A5Q;
  assign CLBLM_L_X8Y142_SLICE_X11Y142_A = CLBLM_L_X8Y142_SLICE_X11Y142_AO6;
  assign CLBLM_L_X8Y142_SLICE_X11Y142_B = CLBLM_L_X8Y142_SLICE_X11Y142_BO6;
  assign CLBLM_L_X8Y142_SLICE_X11Y142_C = CLBLM_L_X8Y142_SLICE_X11Y142_CO6;
  assign CLBLM_L_X8Y142_SLICE_X11Y142_D = CLBLM_L_X8Y142_SLICE_X11Y142_DO6;
  assign CLBLM_L_X8Y142_SLICE_X11Y142_CMUX = CLBLM_L_X8Y142_SLICE_X11Y142_CO5;
  assign CLBLM_L_X8Y142_SLICE_X11Y142_DMUX = CLBLM_L_X8Y142_SLICE_X11Y142_DO6;
  assign CLBLM_L_X8Y143_SLICE_X10Y143_A = CLBLM_L_X8Y143_SLICE_X10Y143_AO6;
  assign CLBLM_L_X8Y143_SLICE_X10Y143_B = CLBLM_L_X8Y143_SLICE_X10Y143_BO6;
  assign CLBLM_L_X8Y143_SLICE_X10Y143_C = CLBLM_L_X8Y143_SLICE_X10Y143_CO6;
  assign CLBLM_L_X8Y143_SLICE_X10Y143_D = CLBLM_L_X8Y143_SLICE_X10Y143_DO6;
  assign CLBLM_L_X8Y143_SLICE_X11Y143_A = CLBLM_L_X8Y143_SLICE_X11Y143_AO6;
  assign CLBLM_L_X8Y143_SLICE_X11Y143_B = CLBLM_L_X8Y143_SLICE_X11Y143_BO6;
  assign CLBLM_L_X8Y143_SLICE_X11Y143_C = CLBLM_L_X8Y143_SLICE_X11Y143_CO6;
  assign CLBLM_L_X8Y143_SLICE_X11Y143_D = CLBLM_L_X8Y143_SLICE_X11Y143_DO6;
  assign CLBLM_L_X8Y143_SLICE_X11Y143_DMUX = CLBLM_L_X8Y143_SLICE_X11Y143_D5Q;
  assign CLBLM_L_X8Y144_SLICE_X10Y144_A = CLBLM_L_X8Y144_SLICE_X10Y144_AO6;
  assign CLBLM_L_X8Y144_SLICE_X10Y144_B = CLBLM_L_X8Y144_SLICE_X10Y144_BO6;
  assign CLBLM_L_X8Y144_SLICE_X10Y144_C = CLBLM_L_X8Y144_SLICE_X10Y144_CO6;
  assign CLBLM_L_X8Y144_SLICE_X10Y144_D = CLBLM_L_X8Y144_SLICE_X10Y144_DO6;
  assign CLBLM_L_X8Y144_SLICE_X10Y144_AMUX = CLBLM_L_X8Y144_SLICE_X10Y144_AO5;
  assign CLBLM_L_X8Y144_SLICE_X10Y144_BMUX = CLBLM_L_X8Y144_SLICE_X10Y144_BO5;
  assign CLBLM_L_X8Y144_SLICE_X11Y144_A = CLBLM_L_X8Y144_SLICE_X11Y144_AO6;
  assign CLBLM_L_X8Y144_SLICE_X11Y144_B = CLBLM_L_X8Y144_SLICE_X11Y144_BO6;
  assign CLBLM_L_X8Y144_SLICE_X11Y144_C = CLBLM_L_X8Y144_SLICE_X11Y144_CO6;
  assign CLBLM_L_X8Y144_SLICE_X11Y144_D = CLBLM_L_X8Y144_SLICE_X11Y144_DO6;
  assign CLBLM_L_X8Y144_SLICE_X11Y144_BMUX = CLBLM_L_X8Y144_SLICE_X11Y144_B5Q;
  assign CLBLM_L_X8Y145_SLICE_X10Y145_A = CLBLM_L_X8Y145_SLICE_X10Y145_AO6;
  assign CLBLM_L_X8Y145_SLICE_X10Y145_B = CLBLM_L_X8Y145_SLICE_X10Y145_BO6;
  assign CLBLM_L_X8Y145_SLICE_X10Y145_C = CLBLM_L_X8Y145_SLICE_X10Y145_CO6;
  assign CLBLM_L_X8Y145_SLICE_X10Y145_D = CLBLM_L_X8Y145_SLICE_X10Y145_DO6;
  assign CLBLM_L_X8Y145_SLICE_X10Y145_AMUX = CLBLM_L_X8Y145_SLICE_X10Y145_A5Q;
  assign CLBLM_L_X8Y145_SLICE_X11Y145_A = CLBLM_L_X8Y145_SLICE_X11Y145_AO6;
  assign CLBLM_L_X8Y145_SLICE_X11Y145_B = CLBLM_L_X8Y145_SLICE_X11Y145_BO6;
  assign CLBLM_L_X8Y145_SLICE_X11Y145_C = CLBLM_L_X8Y145_SLICE_X11Y145_CO6;
  assign CLBLM_L_X8Y145_SLICE_X11Y145_D = CLBLM_L_X8Y145_SLICE_X11Y145_DO6;
  assign CLBLM_L_X8Y145_SLICE_X11Y145_CMUX = CLBLM_L_X8Y145_SLICE_X11Y145_C5Q;
  assign CLBLM_L_X8Y146_SLICE_X10Y146_A = CLBLM_L_X8Y146_SLICE_X10Y146_AO6;
  assign CLBLM_L_X8Y146_SLICE_X10Y146_B = CLBLM_L_X8Y146_SLICE_X10Y146_BO6;
  assign CLBLM_L_X8Y146_SLICE_X10Y146_C = CLBLM_L_X8Y146_SLICE_X10Y146_CO6;
  assign CLBLM_L_X8Y146_SLICE_X10Y146_D = CLBLM_L_X8Y146_SLICE_X10Y146_DO6;
  assign CLBLM_L_X8Y146_SLICE_X10Y146_AMUX = CLBLM_L_X8Y146_SLICE_X10Y146_AO5;
  assign CLBLM_L_X8Y146_SLICE_X10Y146_BMUX = CLBLM_L_X8Y146_SLICE_X10Y146_BO5;
  assign CLBLM_L_X8Y146_SLICE_X10Y146_CMUX = CLBLM_L_X8Y146_SLICE_X10Y146_CO6;
  assign CLBLM_L_X8Y146_SLICE_X11Y146_A = CLBLM_L_X8Y146_SLICE_X11Y146_AO6;
  assign CLBLM_L_X8Y146_SLICE_X11Y146_B = CLBLM_L_X8Y146_SLICE_X11Y146_BO6;
  assign CLBLM_L_X8Y146_SLICE_X11Y146_C = CLBLM_L_X8Y146_SLICE_X11Y146_CO6;
  assign CLBLM_L_X8Y146_SLICE_X11Y146_D = CLBLM_L_X8Y146_SLICE_X11Y146_DO6;
  assign CLBLM_L_X8Y146_SLICE_X11Y146_BMUX = CLBLM_L_X8Y146_SLICE_X11Y146_B5Q;
  assign CLBLM_L_X8Y146_SLICE_X11Y146_CMUX = CLBLM_L_X8Y146_SLICE_X11Y146_C5Q;
  assign CLBLM_L_X8Y146_SLICE_X11Y146_DMUX = CLBLM_L_X8Y146_SLICE_X11Y146_D5Q;
  assign CLBLM_L_X8Y147_SLICE_X10Y147_A = CLBLM_L_X8Y147_SLICE_X10Y147_AO6;
  assign CLBLM_L_X8Y147_SLICE_X10Y147_B = CLBLM_L_X8Y147_SLICE_X10Y147_BO6;
  assign CLBLM_L_X8Y147_SLICE_X10Y147_C = CLBLM_L_X8Y147_SLICE_X10Y147_CO6;
  assign CLBLM_L_X8Y147_SLICE_X10Y147_D = CLBLM_L_X8Y147_SLICE_X10Y147_DO6;
  assign CLBLM_L_X8Y147_SLICE_X10Y147_CMUX = CLBLM_L_X8Y147_SLICE_X10Y147_C5Q;
  assign CLBLM_L_X8Y147_SLICE_X11Y147_A = CLBLM_L_X8Y147_SLICE_X11Y147_AO6;
  assign CLBLM_L_X8Y147_SLICE_X11Y147_B = CLBLM_L_X8Y147_SLICE_X11Y147_BO6;
  assign CLBLM_L_X8Y147_SLICE_X11Y147_C = CLBLM_L_X8Y147_SLICE_X11Y147_CO6;
  assign CLBLM_L_X8Y147_SLICE_X11Y147_D = CLBLM_L_X8Y147_SLICE_X11Y147_DO6;
  assign CLBLM_L_X8Y147_SLICE_X11Y147_CMUX = CLBLM_L_X8Y147_SLICE_X11Y147_C5Q;
  assign CLBLM_L_X8Y148_SLICE_X10Y148_A = CLBLM_L_X8Y148_SLICE_X10Y148_AO6;
  assign CLBLM_L_X8Y148_SLICE_X10Y148_B = CLBLM_L_X8Y148_SLICE_X10Y148_BO6;
  assign CLBLM_L_X8Y148_SLICE_X10Y148_C = CLBLM_L_X8Y148_SLICE_X10Y148_CO6;
  assign CLBLM_L_X8Y148_SLICE_X10Y148_D = CLBLM_L_X8Y148_SLICE_X10Y148_DO6;
  assign CLBLM_L_X8Y148_SLICE_X10Y148_BMUX = CLBLM_L_X8Y148_SLICE_X10Y148_B5Q;
  assign CLBLM_L_X8Y148_SLICE_X11Y148_A = CLBLM_L_X8Y148_SLICE_X11Y148_AO6;
  assign CLBLM_L_X8Y148_SLICE_X11Y148_B = CLBLM_L_X8Y148_SLICE_X11Y148_BO6;
  assign CLBLM_L_X8Y148_SLICE_X11Y148_C = CLBLM_L_X8Y148_SLICE_X11Y148_CO6;
  assign CLBLM_L_X8Y148_SLICE_X11Y148_D = CLBLM_L_X8Y148_SLICE_X11Y148_DO6;
  assign CLBLM_L_X8Y148_SLICE_X11Y148_BMUX = CLBLM_L_X8Y148_SLICE_X11Y148_B5Q;
  assign CLBLM_L_X8Y149_SLICE_X10Y149_A = CLBLM_L_X8Y149_SLICE_X10Y149_AO6;
  assign CLBLM_L_X8Y149_SLICE_X10Y149_B = CLBLM_L_X8Y149_SLICE_X10Y149_BO6;
  assign CLBLM_L_X8Y149_SLICE_X10Y149_C = CLBLM_L_X8Y149_SLICE_X10Y149_CO6;
  assign CLBLM_L_X8Y149_SLICE_X10Y149_D = CLBLM_L_X8Y149_SLICE_X10Y149_DO6;
  assign CLBLM_L_X8Y149_SLICE_X11Y149_A = CLBLM_L_X8Y149_SLICE_X11Y149_AO6;
  assign CLBLM_L_X8Y149_SLICE_X11Y149_B = CLBLM_L_X8Y149_SLICE_X11Y149_BO6;
  assign CLBLM_L_X8Y149_SLICE_X11Y149_C = CLBLM_L_X8Y149_SLICE_X11Y149_CO6;
  assign CLBLM_L_X8Y149_SLICE_X11Y149_D = CLBLM_L_X8Y149_SLICE_X11Y149_DO6;
  assign CLBLM_L_X8Y149_SLICE_X11Y149_AMUX = CLBLM_L_X8Y149_SLICE_X11Y149_A5Q;
  assign CLBLM_L_X8Y150_SLICE_X10Y150_A = CLBLM_L_X8Y150_SLICE_X10Y150_AO6;
  assign CLBLM_L_X8Y150_SLICE_X10Y150_B = CLBLM_L_X8Y150_SLICE_X10Y150_BO6;
  assign CLBLM_L_X8Y150_SLICE_X10Y150_C = CLBLM_L_X8Y150_SLICE_X10Y150_CO6;
  assign CLBLM_L_X8Y150_SLICE_X10Y150_D = CLBLM_L_X8Y150_SLICE_X10Y150_DO6;
  assign CLBLM_L_X8Y150_SLICE_X10Y150_BMUX = CLBLM_L_X8Y150_SLICE_X10Y150_BO5;
  assign CLBLM_L_X8Y150_SLICE_X10Y150_CMUX = CLBLM_L_X8Y150_SLICE_X10Y150_CO6;
  assign CLBLM_L_X8Y150_SLICE_X11Y150_A = CLBLM_L_X8Y150_SLICE_X11Y150_AO6;
  assign CLBLM_L_X8Y150_SLICE_X11Y150_B = CLBLM_L_X8Y150_SLICE_X11Y150_BO6;
  assign CLBLM_L_X8Y150_SLICE_X11Y150_C = CLBLM_L_X8Y150_SLICE_X11Y150_CO6;
  assign CLBLM_L_X8Y150_SLICE_X11Y150_D = CLBLM_L_X8Y150_SLICE_X11Y150_DO6;
  assign CLBLM_L_X8Y150_SLICE_X11Y150_BMUX = CLBLM_L_X8Y150_SLICE_X11Y150_BO5;
  assign CLBLM_L_X8Y151_SLICE_X10Y151_A = CLBLM_L_X8Y151_SLICE_X10Y151_AO6;
  assign CLBLM_L_X8Y151_SLICE_X10Y151_B = CLBLM_L_X8Y151_SLICE_X10Y151_BO6;
  assign CLBLM_L_X8Y151_SLICE_X10Y151_C = CLBLM_L_X8Y151_SLICE_X10Y151_CO6;
  assign CLBLM_L_X8Y151_SLICE_X10Y151_D = CLBLM_L_X8Y151_SLICE_X10Y151_DO6;
  assign CLBLM_L_X8Y151_SLICE_X10Y151_AMUX = CLBLM_L_X8Y151_SLICE_X10Y151_A5Q;
  assign CLBLM_L_X8Y151_SLICE_X10Y151_BMUX = CLBLM_L_X8Y151_SLICE_X10Y151_B5Q;
  assign CLBLM_L_X8Y151_SLICE_X10Y151_CMUX = CLBLM_L_X8Y151_SLICE_X10Y151_C5Q;
  assign CLBLM_L_X8Y151_SLICE_X11Y151_A = CLBLM_L_X8Y151_SLICE_X11Y151_AO6;
  assign CLBLM_L_X8Y151_SLICE_X11Y151_B = CLBLM_L_X8Y151_SLICE_X11Y151_BO6;
  assign CLBLM_L_X8Y151_SLICE_X11Y151_C = CLBLM_L_X8Y151_SLICE_X11Y151_CO6;
  assign CLBLM_L_X8Y151_SLICE_X11Y151_D = CLBLM_L_X8Y151_SLICE_X11Y151_DO6;
  assign CLBLM_L_X8Y152_SLICE_X10Y152_A = CLBLM_L_X8Y152_SLICE_X10Y152_AO6;
  assign CLBLM_L_X8Y152_SLICE_X10Y152_B = CLBLM_L_X8Y152_SLICE_X10Y152_BO6;
  assign CLBLM_L_X8Y152_SLICE_X10Y152_C = CLBLM_L_X8Y152_SLICE_X10Y152_CO6;
  assign CLBLM_L_X8Y152_SLICE_X10Y152_D = CLBLM_L_X8Y152_SLICE_X10Y152_DO6;
  assign CLBLM_L_X8Y152_SLICE_X10Y152_AMUX = CLBLM_L_X8Y152_SLICE_X10Y152_A5Q;
  assign CLBLM_L_X8Y152_SLICE_X10Y152_CMUX = CLBLM_L_X8Y152_SLICE_X10Y152_C5Q;
  assign CLBLM_L_X8Y152_SLICE_X11Y152_A = CLBLM_L_X8Y152_SLICE_X11Y152_AO6;
  assign CLBLM_L_X8Y152_SLICE_X11Y152_B = CLBLM_L_X8Y152_SLICE_X11Y152_BO6;
  assign CLBLM_L_X8Y152_SLICE_X11Y152_C = CLBLM_L_X8Y152_SLICE_X11Y152_CO6;
  assign CLBLM_L_X8Y152_SLICE_X11Y152_D = CLBLM_L_X8Y152_SLICE_X11Y152_DO6;
  assign CLBLM_L_X8Y152_SLICE_X11Y152_DMUX = CLBLM_L_X8Y152_SLICE_X11Y152_D5Q;
  assign CLBLM_L_X8Y153_SLICE_X10Y153_A = CLBLM_L_X8Y153_SLICE_X10Y153_AO6;
  assign CLBLM_L_X8Y153_SLICE_X10Y153_B = CLBLM_L_X8Y153_SLICE_X10Y153_BO6;
  assign CLBLM_L_X8Y153_SLICE_X10Y153_C = CLBLM_L_X8Y153_SLICE_X10Y153_CO6;
  assign CLBLM_L_X8Y153_SLICE_X10Y153_D = CLBLM_L_X8Y153_SLICE_X10Y153_DO6;
  assign CLBLM_L_X8Y153_SLICE_X10Y153_AMUX = CLBLM_L_X8Y153_SLICE_X10Y153_A5Q;
  assign CLBLM_L_X8Y153_SLICE_X10Y153_BMUX = CLBLM_L_X8Y153_SLICE_X10Y153_B5Q;
  assign CLBLM_L_X8Y153_SLICE_X10Y153_CMUX = CLBLM_L_X8Y153_SLICE_X10Y153_C5Q;
  assign CLBLM_L_X8Y153_SLICE_X10Y153_DMUX = CLBLM_L_X8Y153_SLICE_X10Y153_D5Q;
  assign CLBLM_L_X8Y153_SLICE_X11Y153_A = CLBLM_L_X8Y153_SLICE_X11Y153_AO6;
  assign CLBLM_L_X8Y153_SLICE_X11Y153_B = CLBLM_L_X8Y153_SLICE_X11Y153_BO6;
  assign CLBLM_L_X8Y153_SLICE_X11Y153_C = CLBLM_L_X8Y153_SLICE_X11Y153_CO6;
  assign CLBLM_L_X8Y153_SLICE_X11Y153_D = CLBLM_L_X8Y153_SLICE_X11Y153_DO6;
  assign CLBLM_L_X8Y154_SLICE_X10Y154_A = CLBLM_L_X8Y154_SLICE_X10Y154_AO6;
  assign CLBLM_L_X8Y154_SLICE_X10Y154_B = CLBLM_L_X8Y154_SLICE_X10Y154_BO6;
  assign CLBLM_L_X8Y154_SLICE_X10Y154_C = CLBLM_L_X8Y154_SLICE_X10Y154_CO6;
  assign CLBLM_L_X8Y154_SLICE_X10Y154_D = CLBLM_L_X8Y154_SLICE_X10Y154_DO6;
  assign CLBLM_L_X8Y154_SLICE_X10Y154_BMUX = CLBLM_L_X8Y154_SLICE_X10Y154_BO5;
  assign CLBLM_L_X8Y154_SLICE_X11Y154_A = CLBLM_L_X8Y154_SLICE_X11Y154_AO6;
  assign CLBLM_L_X8Y154_SLICE_X11Y154_B = CLBLM_L_X8Y154_SLICE_X11Y154_BO6;
  assign CLBLM_L_X8Y154_SLICE_X11Y154_C = CLBLM_L_X8Y154_SLICE_X11Y154_CO6;
  assign CLBLM_L_X8Y154_SLICE_X11Y154_D = CLBLM_L_X8Y154_SLICE_X11Y154_DO6;
  assign CLBLM_L_X10Y142_SLICE_X12Y142_A = CLBLM_L_X10Y142_SLICE_X12Y142_AO6;
  assign CLBLM_L_X10Y142_SLICE_X12Y142_B = CLBLM_L_X10Y142_SLICE_X12Y142_BO6;
  assign CLBLM_L_X10Y142_SLICE_X12Y142_C = CLBLM_L_X10Y142_SLICE_X12Y142_CO6;
  assign CLBLM_L_X10Y142_SLICE_X12Y142_D = CLBLM_L_X10Y142_SLICE_X12Y142_DO6;
  assign CLBLM_L_X10Y142_SLICE_X13Y142_A = CLBLM_L_X10Y142_SLICE_X13Y142_AO6;
  assign CLBLM_L_X10Y142_SLICE_X13Y142_B = CLBLM_L_X10Y142_SLICE_X13Y142_BO6;
  assign CLBLM_L_X10Y142_SLICE_X13Y142_C = CLBLM_L_X10Y142_SLICE_X13Y142_CO6;
  assign CLBLM_L_X10Y142_SLICE_X13Y142_D = CLBLM_L_X10Y142_SLICE_X13Y142_DO6;
  assign CLBLM_L_X10Y143_SLICE_X12Y143_A = CLBLM_L_X10Y143_SLICE_X12Y143_AO6;
  assign CLBLM_L_X10Y143_SLICE_X12Y143_B = CLBLM_L_X10Y143_SLICE_X12Y143_BO6;
  assign CLBLM_L_X10Y143_SLICE_X12Y143_C = CLBLM_L_X10Y143_SLICE_X12Y143_CO6;
  assign CLBLM_L_X10Y143_SLICE_X12Y143_D = CLBLM_L_X10Y143_SLICE_X12Y143_DO6;
  assign CLBLM_L_X10Y143_SLICE_X12Y143_CMUX = CLBLM_L_X10Y143_SLICE_X12Y143_CO5;
  assign CLBLM_L_X10Y143_SLICE_X13Y143_A = CLBLM_L_X10Y143_SLICE_X13Y143_AO6;
  assign CLBLM_L_X10Y143_SLICE_X13Y143_B = CLBLM_L_X10Y143_SLICE_X13Y143_BO6;
  assign CLBLM_L_X10Y143_SLICE_X13Y143_C = CLBLM_L_X10Y143_SLICE_X13Y143_CO6;
  assign CLBLM_L_X10Y143_SLICE_X13Y143_D = CLBLM_L_X10Y143_SLICE_X13Y143_DO6;
  assign CLBLM_L_X10Y143_SLICE_X13Y143_CMUX = CLBLM_L_X10Y143_SLICE_X13Y143_C5Q;
  assign CLBLM_L_X10Y143_SLICE_X13Y143_DMUX = CLBLM_L_X10Y143_SLICE_X13Y143_DO5;
  assign CLBLM_L_X10Y144_SLICE_X12Y144_A = CLBLM_L_X10Y144_SLICE_X12Y144_AO6;
  assign CLBLM_L_X10Y144_SLICE_X12Y144_B = CLBLM_L_X10Y144_SLICE_X12Y144_BO6;
  assign CLBLM_L_X10Y144_SLICE_X12Y144_C = CLBLM_L_X10Y144_SLICE_X12Y144_CO6;
  assign CLBLM_L_X10Y144_SLICE_X12Y144_D = CLBLM_L_X10Y144_SLICE_X12Y144_DO6;
  assign CLBLM_L_X10Y144_SLICE_X12Y144_AMUX = CLBLM_L_X10Y144_SLICE_X12Y144_AO5;
  assign CLBLM_L_X10Y144_SLICE_X12Y144_BMUX = CLBLM_L_X10Y144_SLICE_X12Y144_BO5;
  assign CLBLM_L_X10Y144_SLICE_X13Y144_A = CLBLM_L_X10Y144_SLICE_X13Y144_AO6;
  assign CLBLM_L_X10Y144_SLICE_X13Y144_B = CLBLM_L_X10Y144_SLICE_X13Y144_BO6;
  assign CLBLM_L_X10Y144_SLICE_X13Y144_C = CLBLM_L_X10Y144_SLICE_X13Y144_CO6;
  assign CLBLM_L_X10Y144_SLICE_X13Y144_D = CLBLM_L_X10Y144_SLICE_X13Y144_DO6;
  assign CLBLM_L_X10Y144_SLICE_X13Y144_AMUX = CLBLM_L_X10Y144_SLICE_X13Y144_A5Q;
  assign CLBLM_L_X10Y144_SLICE_X13Y144_CMUX = CLBLM_L_X10Y144_SLICE_X13Y144_C5Q;
  assign CLBLM_L_X10Y145_SLICE_X12Y145_A = CLBLM_L_X10Y145_SLICE_X12Y145_AO6;
  assign CLBLM_L_X10Y145_SLICE_X12Y145_B = CLBLM_L_X10Y145_SLICE_X12Y145_BO6;
  assign CLBLM_L_X10Y145_SLICE_X12Y145_C = CLBLM_L_X10Y145_SLICE_X12Y145_CO6;
  assign CLBLM_L_X10Y145_SLICE_X12Y145_D = CLBLM_L_X10Y145_SLICE_X12Y145_DO6;
  assign CLBLM_L_X10Y145_SLICE_X12Y145_AMUX = CLBLM_L_X10Y145_SLICE_X12Y145_A5Q;
  assign CLBLM_L_X10Y145_SLICE_X13Y145_A = CLBLM_L_X10Y145_SLICE_X13Y145_AO6;
  assign CLBLM_L_X10Y145_SLICE_X13Y145_B = CLBLM_L_X10Y145_SLICE_X13Y145_BO6;
  assign CLBLM_L_X10Y145_SLICE_X13Y145_C = CLBLM_L_X10Y145_SLICE_X13Y145_CO6;
  assign CLBLM_L_X10Y145_SLICE_X13Y145_D = CLBLM_L_X10Y145_SLICE_X13Y145_DO6;
  assign CLBLM_L_X10Y146_SLICE_X12Y146_A = CLBLM_L_X10Y146_SLICE_X12Y146_AO6;
  assign CLBLM_L_X10Y146_SLICE_X12Y146_B = CLBLM_L_X10Y146_SLICE_X12Y146_BO6;
  assign CLBLM_L_X10Y146_SLICE_X12Y146_C = CLBLM_L_X10Y146_SLICE_X12Y146_CO6;
  assign CLBLM_L_X10Y146_SLICE_X12Y146_D = CLBLM_L_X10Y146_SLICE_X12Y146_DO6;
  assign CLBLM_L_X10Y146_SLICE_X12Y146_DMUX = CLBLM_L_X10Y146_SLICE_X12Y146_D5Q;
  assign CLBLM_L_X10Y146_SLICE_X13Y146_A = CLBLM_L_X10Y146_SLICE_X13Y146_AO6;
  assign CLBLM_L_X10Y146_SLICE_X13Y146_B = CLBLM_L_X10Y146_SLICE_X13Y146_BO6;
  assign CLBLM_L_X10Y146_SLICE_X13Y146_C = CLBLM_L_X10Y146_SLICE_X13Y146_CO6;
  assign CLBLM_L_X10Y146_SLICE_X13Y146_D = CLBLM_L_X10Y146_SLICE_X13Y146_DO6;
  assign CLBLM_L_X10Y146_SLICE_X13Y146_DMUX = CLBLM_L_X10Y146_SLICE_X13Y146_DO5;
  assign CLBLM_L_X10Y147_SLICE_X12Y147_A = CLBLM_L_X10Y147_SLICE_X12Y147_AO6;
  assign CLBLM_L_X10Y147_SLICE_X12Y147_B = CLBLM_L_X10Y147_SLICE_X12Y147_BO6;
  assign CLBLM_L_X10Y147_SLICE_X12Y147_C = CLBLM_L_X10Y147_SLICE_X12Y147_CO6;
  assign CLBLM_L_X10Y147_SLICE_X12Y147_D = CLBLM_L_X10Y147_SLICE_X12Y147_DO6;
  assign CLBLM_L_X10Y147_SLICE_X12Y147_AMUX = CLBLM_L_X10Y147_SLICE_X12Y147_AO5;
  assign CLBLM_L_X10Y147_SLICE_X12Y147_BMUX = CLBLM_L_X10Y147_SLICE_X12Y147_BO5;
  assign CLBLM_L_X10Y147_SLICE_X13Y147_A = CLBLM_L_X10Y147_SLICE_X13Y147_AO6;
  assign CLBLM_L_X10Y147_SLICE_X13Y147_B = CLBLM_L_X10Y147_SLICE_X13Y147_BO6;
  assign CLBLM_L_X10Y147_SLICE_X13Y147_C = CLBLM_L_X10Y147_SLICE_X13Y147_CO6;
  assign CLBLM_L_X10Y147_SLICE_X13Y147_D = CLBLM_L_X10Y147_SLICE_X13Y147_DO6;
  assign CLBLM_L_X10Y148_SLICE_X12Y148_A = CLBLM_L_X10Y148_SLICE_X12Y148_AO6;
  assign CLBLM_L_X10Y148_SLICE_X12Y148_B = CLBLM_L_X10Y148_SLICE_X12Y148_BO6;
  assign CLBLM_L_X10Y148_SLICE_X12Y148_C = CLBLM_L_X10Y148_SLICE_X12Y148_CO6;
  assign CLBLM_L_X10Y148_SLICE_X12Y148_D = CLBLM_L_X10Y148_SLICE_X12Y148_DO6;
  assign CLBLM_L_X10Y148_SLICE_X12Y148_AMUX = CLBLM_L_X10Y148_SLICE_X12Y148_AO5;
  assign CLBLM_L_X10Y148_SLICE_X13Y148_A = CLBLM_L_X10Y148_SLICE_X13Y148_AO6;
  assign CLBLM_L_X10Y148_SLICE_X13Y148_B = CLBLM_L_X10Y148_SLICE_X13Y148_BO6;
  assign CLBLM_L_X10Y148_SLICE_X13Y148_C = CLBLM_L_X10Y148_SLICE_X13Y148_CO6;
  assign CLBLM_L_X10Y148_SLICE_X13Y148_D = CLBLM_L_X10Y148_SLICE_X13Y148_DO6;
  assign CLBLM_L_X10Y148_SLICE_X13Y148_CMUX = CLBLM_L_X10Y148_SLICE_X13Y148_C5Q;
  assign CLBLM_L_X10Y149_SLICE_X12Y149_A = CLBLM_L_X10Y149_SLICE_X12Y149_AO6;
  assign CLBLM_L_X10Y149_SLICE_X12Y149_B = CLBLM_L_X10Y149_SLICE_X12Y149_BO6;
  assign CLBLM_L_X10Y149_SLICE_X12Y149_C = CLBLM_L_X10Y149_SLICE_X12Y149_CO6;
  assign CLBLM_L_X10Y149_SLICE_X12Y149_D = CLBLM_L_X10Y149_SLICE_X12Y149_DO6;
  assign CLBLM_L_X10Y149_SLICE_X12Y149_AMUX = CLBLM_L_X10Y149_SLICE_X12Y149_A5Q;
  assign CLBLM_L_X10Y149_SLICE_X12Y149_BMUX = CLBLM_L_X10Y149_SLICE_X12Y149_BO5;
  assign CLBLM_L_X10Y149_SLICE_X12Y149_CMUX = CLBLM_L_X10Y149_SLICE_X12Y149_CO6;
  assign CLBLM_L_X10Y149_SLICE_X13Y149_A = CLBLM_L_X10Y149_SLICE_X13Y149_AO6;
  assign CLBLM_L_X10Y149_SLICE_X13Y149_B = CLBLM_L_X10Y149_SLICE_X13Y149_BO6;
  assign CLBLM_L_X10Y149_SLICE_X13Y149_C = CLBLM_L_X10Y149_SLICE_X13Y149_CO6;
  assign CLBLM_L_X10Y149_SLICE_X13Y149_D = CLBLM_L_X10Y149_SLICE_X13Y149_DO6;
  assign CLBLM_L_X10Y149_SLICE_X13Y149_AMUX = CLBLM_L_X10Y149_SLICE_X13Y149_AO5;
  assign CLBLM_L_X10Y149_SLICE_X13Y149_DMUX = CLBLM_L_X10Y149_SLICE_X13Y149_DO6;
  assign CLBLM_L_X10Y150_SLICE_X12Y150_A = CLBLM_L_X10Y150_SLICE_X12Y150_AO6;
  assign CLBLM_L_X10Y150_SLICE_X12Y150_B = CLBLM_L_X10Y150_SLICE_X12Y150_BO6;
  assign CLBLM_L_X10Y150_SLICE_X12Y150_C = CLBLM_L_X10Y150_SLICE_X12Y150_CO6;
  assign CLBLM_L_X10Y150_SLICE_X12Y150_D = CLBLM_L_X10Y150_SLICE_X12Y150_DO6;
  assign CLBLM_L_X10Y150_SLICE_X12Y150_AMUX = CLBLM_L_X10Y150_SLICE_X12Y150_AO5;
  assign CLBLM_L_X10Y150_SLICE_X12Y150_BMUX = CLBLM_L_X10Y150_SLICE_X12Y150_BO5;
  assign CLBLM_L_X10Y150_SLICE_X13Y150_A = CLBLM_L_X10Y150_SLICE_X13Y150_AO6;
  assign CLBLM_L_X10Y150_SLICE_X13Y150_B = CLBLM_L_X10Y150_SLICE_X13Y150_BO6;
  assign CLBLM_L_X10Y150_SLICE_X13Y150_C = CLBLM_L_X10Y150_SLICE_X13Y150_CO6;
  assign CLBLM_L_X10Y150_SLICE_X13Y150_D = CLBLM_L_X10Y150_SLICE_X13Y150_DO6;
  assign CLBLM_L_X10Y150_SLICE_X13Y150_BMUX = CLBLM_L_X10Y150_SLICE_X13Y150_BO5;
  assign CLBLM_L_X10Y151_SLICE_X12Y151_A = CLBLM_L_X10Y151_SLICE_X12Y151_AO6;
  assign CLBLM_L_X10Y151_SLICE_X12Y151_B = CLBLM_L_X10Y151_SLICE_X12Y151_BO6;
  assign CLBLM_L_X10Y151_SLICE_X12Y151_C = CLBLM_L_X10Y151_SLICE_X12Y151_CO6;
  assign CLBLM_L_X10Y151_SLICE_X12Y151_D = CLBLM_L_X10Y151_SLICE_X12Y151_DO6;
  assign CLBLM_L_X10Y151_SLICE_X13Y151_A = CLBLM_L_X10Y151_SLICE_X13Y151_AO6;
  assign CLBLM_L_X10Y151_SLICE_X13Y151_B = CLBLM_L_X10Y151_SLICE_X13Y151_BO6;
  assign CLBLM_L_X10Y151_SLICE_X13Y151_C = CLBLM_L_X10Y151_SLICE_X13Y151_CO6;
  assign CLBLM_L_X10Y151_SLICE_X13Y151_D = CLBLM_L_X10Y151_SLICE_X13Y151_DO6;
  assign CLBLM_L_X10Y151_SLICE_X13Y151_AMUX = CLBLM_L_X10Y151_SLICE_X13Y151_A5Q;
  assign CLBLM_L_X10Y151_SLICE_X13Y151_BMUX = CLBLM_L_X10Y151_SLICE_X13Y151_BO5;
  assign CLBLM_L_X10Y152_SLICE_X12Y152_A = CLBLM_L_X10Y152_SLICE_X12Y152_AO6;
  assign CLBLM_L_X10Y152_SLICE_X12Y152_B = CLBLM_L_X10Y152_SLICE_X12Y152_BO6;
  assign CLBLM_L_X10Y152_SLICE_X12Y152_C = CLBLM_L_X10Y152_SLICE_X12Y152_CO6;
  assign CLBLM_L_X10Y152_SLICE_X12Y152_D = CLBLM_L_X10Y152_SLICE_X12Y152_DO6;
  assign CLBLM_L_X10Y152_SLICE_X13Y152_A = CLBLM_L_X10Y152_SLICE_X13Y152_AO6;
  assign CLBLM_L_X10Y152_SLICE_X13Y152_B = CLBLM_L_X10Y152_SLICE_X13Y152_BO6;
  assign CLBLM_L_X10Y152_SLICE_X13Y152_C = CLBLM_L_X10Y152_SLICE_X13Y152_CO6;
  assign CLBLM_L_X10Y152_SLICE_X13Y152_D = CLBLM_L_X10Y152_SLICE_X13Y152_DO6;
  assign CLBLM_L_X10Y152_SLICE_X13Y152_DMUX = CLBLM_L_X10Y152_SLICE_X13Y152_DO6;
  assign CLBLM_L_X10Y153_SLICE_X12Y153_A = CLBLM_L_X10Y153_SLICE_X12Y153_AO6;
  assign CLBLM_L_X10Y153_SLICE_X12Y153_B = CLBLM_L_X10Y153_SLICE_X12Y153_BO6;
  assign CLBLM_L_X10Y153_SLICE_X12Y153_C = CLBLM_L_X10Y153_SLICE_X12Y153_CO6;
  assign CLBLM_L_X10Y153_SLICE_X12Y153_D = CLBLM_L_X10Y153_SLICE_X12Y153_DO6;
  assign CLBLM_L_X10Y153_SLICE_X12Y153_AMUX = CLBLM_L_X10Y153_SLICE_X12Y153_A5Q;
  assign CLBLM_L_X10Y153_SLICE_X12Y153_CMUX = CLBLM_L_X10Y153_SLICE_X12Y153_CO5;
  assign CLBLM_L_X10Y153_SLICE_X13Y153_A = CLBLM_L_X10Y153_SLICE_X13Y153_AO6;
  assign CLBLM_L_X10Y153_SLICE_X13Y153_B = CLBLM_L_X10Y153_SLICE_X13Y153_BO6;
  assign CLBLM_L_X10Y153_SLICE_X13Y153_C = CLBLM_L_X10Y153_SLICE_X13Y153_CO6;
  assign CLBLM_L_X10Y153_SLICE_X13Y153_D = CLBLM_L_X10Y153_SLICE_X13Y153_DO6;
  assign CLBLM_L_X10Y153_SLICE_X13Y153_AMUX = CLBLM_L_X10Y153_SLICE_X13Y153_A5Q;
  assign CLBLM_L_X10Y153_SLICE_X13Y153_DMUX = CLBLM_L_X10Y153_SLICE_X13Y153_DO6;
  assign CLBLM_L_X10Y154_SLICE_X12Y154_A = CLBLM_L_X10Y154_SLICE_X12Y154_AO6;
  assign CLBLM_L_X10Y154_SLICE_X12Y154_B = CLBLM_L_X10Y154_SLICE_X12Y154_BO6;
  assign CLBLM_L_X10Y154_SLICE_X12Y154_C = CLBLM_L_X10Y154_SLICE_X12Y154_CO6;
  assign CLBLM_L_X10Y154_SLICE_X12Y154_D = CLBLM_L_X10Y154_SLICE_X12Y154_DO6;
  assign CLBLM_L_X10Y154_SLICE_X12Y154_AMUX = CLBLM_L_X10Y154_SLICE_X12Y154_A5Q;
  assign CLBLM_L_X10Y154_SLICE_X12Y154_BMUX = CLBLM_L_X10Y154_SLICE_X12Y154_B5Q;
  assign CLBLM_L_X10Y154_SLICE_X12Y154_CMUX = CLBLM_L_X10Y154_SLICE_X12Y154_CO5;
  assign CLBLM_L_X10Y154_SLICE_X12Y154_DMUX = CLBLM_L_X10Y154_SLICE_X12Y154_DO5;
  assign CLBLM_L_X10Y154_SLICE_X13Y154_A = CLBLM_L_X10Y154_SLICE_X13Y154_AO6;
  assign CLBLM_L_X10Y154_SLICE_X13Y154_B = CLBLM_L_X10Y154_SLICE_X13Y154_BO6;
  assign CLBLM_L_X10Y154_SLICE_X13Y154_C = CLBLM_L_X10Y154_SLICE_X13Y154_CO6;
  assign CLBLM_L_X10Y154_SLICE_X13Y154_D = CLBLM_L_X10Y154_SLICE_X13Y154_DO6;
  assign CLBLM_L_X10Y154_SLICE_X13Y154_BMUX = CLBLM_L_X10Y154_SLICE_X13Y154_BO5;
  assign CLBLM_L_X10Y154_SLICE_X13Y154_CMUX = CLBLM_L_X10Y154_SLICE_X13Y154_CO5;
  assign CLBLM_L_X10Y155_SLICE_X12Y155_A = CLBLM_L_X10Y155_SLICE_X12Y155_AO6;
  assign CLBLM_L_X10Y155_SLICE_X12Y155_B = CLBLM_L_X10Y155_SLICE_X12Y155_BO6;
  assign CLBLM_L_X10Y155_SLICE_X12Y155_C = CLBLM_L_X10Y155_SLICE_X12Y155_CO6;
  assign CLBLM_L_X10Y155_SLICE_X12Y155_D = CLBLM_L_X10Y155_SLICE_X12Y155_DO6;
  assign CLBLM_L_X10Y155_SLICE_X12Y155_BMUX = CLBLM_L_X10Y155_SLICE_X12Y155_BO5;
  assign CLBLM_L_X10Y155_SLICE_X13Y155_A = CLBLM_L_X10Y155_SLICE_X13Y155_AO6;
  assign CLBLM_L_X10Y155_SLICE_X13Y155_B = CLBLM_L_X10Y155_SLICE_X13Y155_BO6;
  assign CLBLM_L_X10Y155_SLICE_X13Y155_C = CLBLM_L_X10Y155_SLICE_X13Y155_CO6;
  assign CLBLM_L_X10Y155_SLICE_X13Y155_D = CLBLM_L_X10Y155_SLICE_X13Y155_DO6;
  assign CLBLM_L_X10Y155_SLICE_X13Y155_AMUX = CLBLM_L_X10Y155_SLICE_X13Y155_AO5;
  assign CLBLM_L_X12Y145_SLICE_X16Y145_A = CLBLM_L_X12Y145_SLICE_X16Y145_AO6;
  assign CLBLM_L_X12Y145_SLICE_X16Y145_B = CLBLM_L_X12Y145_SLICE_X16Y145_BO6;
  assign CLBLM_L_X12Y145_SLICE_X16Y145_C = CLBLM_L_X12Y145_SLICE_X16Y145_CO6;
  assign CLBLM_L_X12Y145_SLICE_X16Y145_D = CLBLM_L_X12Y145_SLICE_X16Y145_DO6;
  assign CLBLM_L_X12Y145_SLICE_X16Y145_AMUX = CLBLM_L_X12Y145_SLICE_X16Y145_AO5;
  assign CLBLM_L_X12Y145_SLICE_X17Y145_A = CLBLM_L_X12Y145_SLICE_X17Y145_AO6;
  assign CLBLM_L_X12Y145_SLICE_X17Y145_B = CLBLM_L_X12Y145_SLICE_X17Y145_BO6;
  assign CLBLM_L_X12Y145_SLICE_X17Y145_C = CLBLM_L_X12Y145_SLICE_X17Y145_CO6;
  assign CLBLM_L_X12Y145_SLICE_X17Y145_D = CLBLM_L_X12Y145_SLICE_X17Y145_DO6;
  assign CLBLM_L_X12Y145_SLICE_X17Y145_AMUX = CLBLM_L_X12Y145_SLICE_X17Y145_AO5;
  assign CLBLM_L_X12Y145_SLICE_X17Y145_CMUX = CLBLM_L_X12Y145_SLICE_X17Y145_CO6;
  assign CLBLM_L_X12Y146_SLICE_X16Y146_A = CLBLM_L_X12Y146_SLICE_X16Y146_AO6;
  assign CLBLM_L_X12Y146_SLICE_X16Y146_B = CLBLM_L_X12Y146_SLICE_X16Y146_BO6;
  assign CLBLM_L_X12Y146_SLICE_X16Y146_C = CLBLM_L_X12Y146_SLICE_X16Y146_CO6;
  assign CLBLM_L_X12Y146_SLICE_X16Y146_D = CLBLM_L_X12Y146_SLICE_X16Y146_DO6;
  assign CLBLM_L_X12Y146_SLICE_X16Y146_AMUX = CLBLM_L_X12Y146_SLICE_X16Y146_AO5;
  assign CLBLM_L_X12Y146_SLICE_X17Y146_A = CLBLM_L_X12Y146_SLICE_X17Y146_AO6;
  assign CLBLM_L_X12Y146_SLICE_X17Y146_B = CLBLM_L_X12Y146_SLICE_X17Y146_BO6;
  assign CLBLM_L_X12Y146_SLICE_X17Y146_C = CLBLM_L_X12Y146_SLICE_X17Y146_CO6;
  assign CLBLM_L_X12Y146_SLICE_X17Y146_D = CLBLM_L_X12Y146_SLICE_X17Y146_DO6;
  assign CLBLM_L_X12Y146_SLICE_X17Y146_CMUX = CLBLM_L_X12Y146_SLICE_X17Y146_CO6;
  assign CLBLM_L_X12Y147_SLICE_X16Y147_A = CLBLM_L_X12Y147_SLICE_X16Y147_AO6;
  assign CLBLM_L_X12Y147_SLICE_X16Y147_B = CLBLM_L_X12Y147_SLICE_X16Y147_BO6;
  assign CLBLM_L_X12Y147_SLICE_X16Y147_C = CLBLM_L_X12Y147_SLICE_X16Y147_CO6;
  assign CLBLM_L_X12Y147_SLICE_X16Y147_D = CLBLM_L_X12Y147_SLICE_X16Y147_DO6;
  assign CLBLM_L_X12Y147_SLICE_X16Y147_AMUX = CLBLM_L_X12Y147_SLICE_X16Y147_AO5;
  assign CLBLM_L_X12Y147_SLICE_X16Y147_CMUX = CLBLM_L_X12Y147_SLICE_X16Y147_CO6;
  assign CLBLM_L_X12Y147_SLICE_X16Y147_DMUX = CLBLM_L_X12Y147_SLICE_X16Y147_DO6;
  assign CLBLM_L_X12Y147_SLICE_X17Y147_A = CLBLM_L_X12Y147_SLICE_X17Y147_AO6;
  assign CLBLM_L_X12Y147_SLICE_X17Y147_B = CLBLM_L_X12Y147_SLICE_X17Y147_BO6;
  assign CLBLM_L_X12Y147_SLICE_X17Y147_C = CLBLM_L_X12Y147_SLICE_X17Y147_CO6;
  assign CLBLM_L_X12Y147_SLICE_X17Y147_D = CLBLM_L_X12Y147_SLICE_X17Y147_DO6;
  assign CLBLM_L_X12Y147_SLICE_X17Y147_AMUX = CLBLM_L_X12Y147_SLICE_X17Y147_AO5;
  assign CLBLM_L_X12Y148_SLICE_X16Y148_A = CLBLM_L_X12Y148_SLICE_X16Y148_AO6;
  assign CLBLM_L_X12Y148_SLICE_X16Y148_B = CLBLM_L_X12Y148_SLICE_X16Y148_BO6;
  assign CLBLM_L_X12Y148_SLICE_X16Y148_C = CLBLM_L_X12Y148_SLICE_X16Y148_CO6;
  assign CLBLM_L_X12Y148_SLICE_X16Y148_D = CLBLM_L_X12Y148_SLICE_X16Y148_DO6;
  assign CLBLM_L_X12Y148_SLICE_X16Y148_AMUX = CLBLM_L_X12Y148_SLICE_X16Y148_AO5;
  assign CLBLM_L_X12Y148_SLICE_X17Y148_A = CLBLM_L_X12Y148_SLICE_X17Y148_AO6;
  assign CLBLM_L_X12Y148_SLICE_X17Y148_B = CLBLM_L_X12Y148_SLICE_X17Y148_BO6;
  assign CLBLM_L_X12Y148_SLICE_X17Y148_C = CLBLM_L_X12Y148_SLICE_X17Y148_CO6;
  assign CLBLM_L_X12Y148_SLICE_X17Y148_D = CLBLM_L_X12Y148_SLICE_X17Y148_DO6;
  assign CLBLM_L_X12Y149_SLICE_X16Y149_A = CLBLM_L_X12Y149_SLICE_X16Y149_AO6;
  assign CLBLM_L_X12Y149_SLICE_X16Y149_B = CLBLM_L_X12Y149_SLICE_X16Y149_BO6;
  assign CLBLM_L_X12Y149_SLICE_X16Y149_C = CLBLM_L_X12Y149_SLICE_X16Y149_CO6;
  assign CLBLM_L_X12Y149_SLICE_X16Y149_D = CLBLM_L_X12Y149_SLICE_X16Y149_DO6;
  assign CLBLM_L_X12Y149_SLICE_X17Y149_A = CLBLM_L_X12Y149_SLICE_X17Y149_AO6;
  assign CLBLM_L_X12Y149_SLICE_X17Y149_B = CLBLM_L_X12Y149_SLICE_X17Y149_BO6;
  assign CLBLM_L_X12Y149_SLICE_X17Y149_C = CLBLM_L_X12Y149_SLICE_X17Y149_CO6;
  assign CLBLM_L_X12Y149_SLICE_X17Y149_D = CLBLM_L_X12Y149_SLICE_X17Y149_DO6;
  assign CLBLM_L_X12Y149_SLICE_X17Y149_AMUX = CLBLM_L_X12Y149_SLICE_X17Y149_AO5;
  assign CLBLM_L_X12Y149_SLICE_X17Y149_BMUX = CLBLM_L_X12Y149_SLICE_X17Y149_BO5;
  assign CLBLM_L_X12Y149_SLICE_X17Y149_DMUX = CLBLM_L_X12Y149_SLICE_X17Y149_DO6;
  assign CLBLM_L_X12Y150_SLICE_X16Y150_A = CLBLM_L_X12Y150_SLICE_X16Y150_AO6;
  assign CLBLM_L_X12Y150_SLICE_X16Y150_B = CLBLM_L_X12Y150_SLICE_X16Y150_BO6;
  assign CLBLM_L_X12Y150_SLICE_X16Y150_C = CLBLM_L_X12Y150_SLICE_X16Y150_CO6;
  assign CLBLM_L_X12Y150_SLICE_X16Y150_D = CLBLM_L_X12Y150_SLICE_X16Y150_DO6;
  assign CLBLM_L_X12Y150_SLICE_X16Y150_AMUX = CLBLM_L_X12Y150_SLICE_X16Y150_AO5;
  assign CLBLM_L_X12Y150_SLICE_X17Y150_A = CLBLM_L_X12Y150_SLICE_X17Y150_AO6;
  assign CLBLM_L_X12Y150_SLICE_X17Y150_B = CLBLM_L_X12Y150_SLICE_X17Y150_BO6;
  assign CLBLM_L_X12Y150_SLICE_X17Y150_C = CLBLM_L_X12Y150_SLICE_X17Y150_CO6;
  assign CLBLM_L_X12Y150_SLICE_X17Y150_D = CLBLM_L_X12Y150_SLICE_X17Y150_DO6;
  assign CLBLM_L_X12Y151_SLICE_X16Y151_A = CLBLM_L_X12Y151_SLICE_X16Y151_AO6;
  assign CLBLM_L_X12Y151_SLICE_X16Y151_B = CLBLM_L_X12Y151_SLICE_X16Y151_BO6;
  assign CLBLM_L_X12Y151_SLICE_X16Y151_C = CLBLM_L_X12Y151_SLICE_X16Y151_CO6;
  assign CLBLM_L_X12Y151_SLICE_X16Y151_D = CLBLM_L_X12Y151_SLICE_X16Y151_DO6;
  assign CLBLM_L_X12Y151_SLICE_X16Y151_AMUX = CLBLM_L_X12Y151_SLICE_X16Y151_AO5;
  assign CLBLM_L_X12Y151_SLICE_X16Y151_BMUX = CLBLM_L_X12Y151_SLICE_X16Y151_BO5;
  assign CLBLM_L_X12Y151_SLICE_X17Y151_A = CLBLM_L_X12Y151_SLICE_X17Y151_AO6;
  assign CLBLM_L_X12Y151_SLICE_X17Y151_B = CLBLM_L_X12Y151_SLICE_X17Y151_BO6;
  assign CLBLM_L_X12Y151_SLICE_X17Y151_C = CLBLM_L_X12Y151_SLICE_X17Y151_CO6;
  assign CLBLM_L_X12Y151_SLICE_X17Y151_D = CLBLM_L_X12Y151_SLICE_X17Y151_DO6;
  assign CLBLM_L_X12Y152_SLICE_X16Y152_A = CLBLM_L_X12Y152_SLICE_X16Y152_AO6;
  assign CLBLM_L_X12Y152_SLICE_X16Y152_B = CLBLM_L_X12Y152_SLICE_X16Y152_BO6;
  assign CLBLM_L_X12Y152_SLICE_X16Y152_C = CLBLM_L_X12Y152_SLICE_X16Y152_CO6;
  assign CLBLM_L_X12Y152_SLICE_X16Y152_D = CLBLM_L_X12Y152_SLICE_X16Y152_DO6;
  assign CLBLM_L_X12Y152_SLICE_X16Y152_AMUX = CLBLM_L_X12Y152_SLICE_X16Y152_AO5;
  assign CLBLM_L_X12Y152_SLICE_X17Y152_A = CLBLM_L_X12Y152_SLICE_X17Y152_AO6;
  assign CLBLM_L_X12Y152_SLICE_X17Y152_B = CLBLM_L_X12Y152_SLICE_X17Y152_BO6;
  assign CLBLM_L_X12Y152_SLICE_X17Y152_C = CLBLM_L_X12Y152_SLICE_X17Y152_CO6;
  assign CLBLM_L_X12Y152_SLICE_X17Y152_D = CLBLM_L_X12Y152_SLICE_X17Y152_DO6;
  assign CLBLM_L_X12Y153_SLICE_X16Y153_A = CLBLM_L_X12Y153_SLICE_X16Y153_AO6;
  assign CLBLM_L_X12Y153_SLICE_X16Y153_B = CLBLM_L_X12Y153_SLICE_X16Y153_BO6;
  assign CLBLM_L_X12Y153_SLICE_X16Y153_C = CLBLM_L_X12Y153_SLICE_X16Y153_CO6;
  assign CLBLM_L_X12Y153_SLICE_X16Y153_D = CLBLM_L_X12Y153_SLICE_X16Y153_DO6;
  assign CLBLM_L_X12Y153_SLICE_X16Y153_AMUX = CLBLM_L_X12Y153_SLICE_X16Y153_AO5;
  assign CLBLM_L_X12Y153_SLICE_X17Y153_A = CLBLM_L_X12Y153_SLICE_X17Y153_AO6;
  assign CLBLM_L_X12Y153_SLICE_X17Y153_B = CLBLM_L_X12Y153_SLICE_X17Y153_BO6;
  assign CLBLM_L_X12Y153_SLICE_X17Y153_C = CLBLM_L_X12Y153_SLICE_X17Y153_CO6;
  assign CLBLM_L_X12Y153_SLICE_X17Y153_D = CLBLM_L_X12Y153_SLICE_X17Y153_DO6;
  assign CLBLM_R_X3Y142_SLICE_X2Y142_A = CLBLM_R_X3Y142_SLICE_X2Y142_AO6;
  assign CLBLM_R_X3Y142_SLICE_X2Y142_B = CLBLM_R_X3Y142_SLICE_X2Y142_BO6;
  assign CLBLM_R_X3Y142_SLICE_X2Y142_C = CLBLM_R_X3Y142_SLICE_X2Y142_CO6;
  assign CLBLM_R_X3Y142_SLICE_X2Y142_D = CLBLM_R_X3Y142_SLICE_X2Y142_DO6;
  assign CLBLM_R_X3Y142_SLICE_X2Y142_BMUX = CLBLM_R_X3Y142_SLICE_X2Y142_BO5;
  assign CLBLM_R_X3Y142_SLICE_X3Y142_A = CLBLM_R_X3Y142_SLICE_X3Y142_AO6;
  assign CLBLM_R_X3Y142_SLICE_X3Y142_B = CLBLM_R_X3Y142_SLICE_X3Y142_BO6;
  assign CLBLM_R_X3Y142_SLICE_X3Y142_C = CLBLM_R_X3Y142_SLICE_X3Y142_CO6;
  assign CLBLM_R_X3Y142_SLICE_X3Y142_D = CLBLM_R_X3Y142_SLICE_X3Y142_DO6;
  assign CLBLM_R_X3Y143_SLICE_X2Y143_A = CLBLM_R_X3Y143_SLICE_X2Y143_AO6;
  assign CLBLM_R_X3Y143_SLICE_X2Y143_B = CLBLM_R_X3Y143_SLICE_X2Y143_BO6;
  assign CLBLM_R_X3Y143_SLICE_X2Y143_C = CLBLM_R_X3Y143_SLICE_X2Y143_CO6;
  assign CLBLM_R_X3Y143_SLICE_X2Y143_D = CLBLM_R_X3Y143_SLICE_X2Y143_DO6;
  assign CLBLM_R_X3Y143_SLICE_X2Y143_AMUX = CLBLM_R_X3Y143_SLICE_X2Y143_A5Q;
  assign CLBLM_R_X3Y143_SLICE_X2Y143_BMUX = CLBLM_R_X3Y143_SLICE_X2Y143_BO5;
  assign CLBLM_R_X3Y143_SLICE_X2Y143_CMUX = CLBLM_R_X3Y143_SLICE_X2Y143_CO5;
  assign CLBLM_R_X3Y143_SLICE_X3Y143_A = CLBLM_R_X3Y143_SLICE_X3Y143_AO6;
  assign CLBLM_R_X3Y143_SLICE_X3Y143_B = CLBLM_R_X3Y143_SLICE_X3Y143_BO6;
  assign CLBLM_R_X3Y143_SLICE_X3Y143_C = CLBLM_R_X3Y143_SLICE_X3Y143_CO6;
  assign CLBLM_R_X3Y143_SLICE_X3Y143_D = CLBLM_R_X3Y143_SLICE_X3Y143_DO6;
  assign CLBLM_R_X3Y143_SLICE_X3Y143_CMUX = CLBLM_R_X3Y143_SLICE_X3Y143_C5Q;
  assign CLBLM_R_X3Y144_SLICE_X2Y144_A = CLBLM_R_X3Y144_SLICE_X2Y144_AO6;
  assign CLBLM_R_X3Y144_SLICE_X2Y144_B = CLBLM_R_X3Y144_SLICE_X2Y144_BO6;
  assign CLBLM_R_X3Y144_SLICE_X2Y144_C = CLBLM_R_X3Y144_SLICE_X2Y144_CO6;
  assign CLBLM_R_X3Y144_SLICE_X2Y144_D = CLBLM_R_X3Y144_SLICE_X2Y144_DO6;
  assign CLBLM_R_X3Y144_SLICE_X2Y144_AMUX = CLBLM_R_X3Y144_SLICE_X2Y144_AO5;
  assign CLBLM_R_X3Y144_SLICE_X2Y144_BMUX = CLBLM_R_X3Y144_SLICE_X2Y144_BO5;
  assign CLBLM_R_X3Y144_SLICE_X3Y144_A = CLBLM_R_X3Y144_SLICE_X3Y144_AO6;
  assign CLBLM_R_X3Y144_SLICE_X3Y144_B = CLBLM_R_X3Y144_SLICE_X3Y144_BO6;
  assign CLBLM_R_X3Y144_SLICE_X3Y144_C = CLBLM_R_X3Y144_SLICE_X3Y144_CO6;
  assign CLBLM_R_X3Y144_SLICE_X3Y144_D = CLBLM_R_X3Y144_SLICE_X3Y144_DO6;
  assign CLBLM_R_X3Y145_SLICE_X2Y145_A = CLBLM_R_X3Y145_SLICE_X2Y145_AO6;
  assign CLBLM_R_X3Y145_SLICE_X2Y145_B = CLBLM_R_X3Y145_SLICE_X2Y145_BO6;
  assign CLBLM_R_X3Y145_SLICE_X2Y145_C = CLBLM_R_X3Y145_SLICE_X2Y145_CO6;
  assign CLBLM_R_X3Y145_SLICE_X2Y145_D = CLBLM_R_X3Y145_SLICE_X2Y145_DO6;
  assign CLBLM_R_X3Y145_SLICE_X2Y145_BMUX = CLBLM_R_X3Y145_SLICE_X2Y145_B5Q;
  assign CLBLM_R_X3Y145_SLICE_X2Y145_CMUX = CLBLM_R_X3Y145_SLICE_X2Y145_C5Q;
  assign CLBLM_R_X3Y145_SLICE_X3Y145_A = CLBLM_R_X3Y145_SLICE_X3Y145_AO6;
  assign CLBLM_R_X3Y145_SLICE_X3Y145_B = CLBLM_R_X3Y145_SLICE_X3Y145_BO6;
  assign CLBLM_R_X3Y145_SLICE_X3Y145_C = CLBLM_R_X3Y145_SLICE_X3Y145_CO6;
  assign CLBLM_R_X3Y145_SLICE_X3Y145_D = CLBLM_R_X3Y145_SLICE_X3Y145_DO6;
  assign CLBLM_R_X3Y145_SLICE_X3Y145_CMUX = CLBLM_R_X3Y145_SLICE_X3Y145_C5Q;
  assign CLBLM_R_X3Y145_SLICE_X3Y145_DMUX = CLBLM_R_X3Y145_SLICE_X3Y145_D5Q;
  assign CLBLM_R_X3Y146_SLICE_X2Y146_A = CLBLM_R_X3Y146_SLICE_X2Y146_AO6;
  assign CLBLM_R_X3Y146_SLICE_X2Y146_B = CLBLM_R_X3Y146_SLICE_X2Y146_BO6;
  assign CLBLM_R_X3Y146_SLICE_X2Y146_C = CLBLM_R_X3Y146_SLICE_X2Y146_CO6;
  assign CLBLM_R_X3Y146_SLICE_X2Y146_D = CLBLM_R_X3Y146_SLICE_X2Y146_DO6;
  assign CLBLM_R_X3Y146_SLICE_X2Y146_CMUX = CLBLM_R_X3Y146_SLICE_X2Y146_C5Q;
  assign CLBLM_R_X3Y146_SLICE_X2Y146_DMUX = CLBLM_R_X3Y146_SLICE_X2Y146_D5Q;
  assign CLBLM_R_X3Y146_SLICE_X3Y146_A = CLBLM_R_X3Y146_SLICE_X3Y146_AO6;
  assign CLBLM_R_X3Y146_SLICE_X3Y146_B = CLBLM_R_X3Y146_SLICE_X3Y146_BO6;
  assign CLBLM_R_X3Y146_SLICE_X3Y146_C = CLBLM_R_X3Y146_SLICE_X3Y146_CO6;
  assign CLBLM_R_X3Y146_SLICE_X3Y146_D = CLBLM_R_X3Y146_SLICE_X3Y146_DO6;
  assign CLBLM_R_X3Y147_SLICE_X2Y147_A = CLBLM_R_X3Y147_SLICE_X2Y147_AO6;
  assign CLBLM_R_X3Y147_SLICE_X2Y147_B = CLBLM_R_X3Y147_SLICE_X2Y147_BO6;
  assign CLBLM_R_X3Y147_SLICE_X2Y147_C = CLBLM_R_X3Y147_SLICE_X2Y147_CO6;
  assign CLBLM_R_X3Y147_SLICE_X2Y147_D = CLBLM_R_X3Y147_SLICE_X2Y147_DO6;
  assign CLBLM_R_X3Y147_SLICE_X2Y147_DMUX = CLBLM_R_X3Y147_SLICE_X2Y147_D5Q;
  assign CLBLM_R_X3Y147_SLICE_X3Y147_A = CLBLM_R_X3Y147_SLICE_X3Y147_AO6;
  assign CLBLM_R_X3Y147_SLICE_X3Y147_B = CLBLM_R_X3Y147_SLICE_X3Y147_BO6;
  assign CLBLM_R_X3Y147_SLICE_X3Y147_C = CLBLM_R_X3Y147_SLICE_X3Y147_CO6;
  assign CLBLM_R_X3Y147_SLICE_X3Y147_D = CLBLM_R_X3Y147_SLICE_X3Y147_DO6;
  assign CLBLM_R_X3Y147_SLICE_X3Y147_BMUX = CLBLM_R_X3Y147_SLICE_X3Y147_B5Q;
  assign CLBLM_R_X3Y147_SLICE_X3Y147_CMUX = CLBLM_R_X3Y147_SLICE_X3Y147_C5Q;
  assign CLBLM_R_X3Y148_SLICE_X2Y148_A = CLBLM_R_X3Y148_SLICE_X2Y148_AO6;
  assign CLBLM_R_X3Y148_SLICE_X2Y148_B = CLBLM_R_X3Y148_SLICE_X2Y148_BO6;
  assign CLBLM_R_X3Y148_SLICE_X2Y148_C = CLBLM_R_X3Y148_SLICE_X2Y148_CO6;
  assign CLBLM_R_X3Y148_SLICE_X2Y148_D = CLBLM_R_X3Y148_SLICE_X2Y148_DO6;
  assign CLBLM_R_X3Y148_SLICE_X2Y148_AMUX = CLBLM_R_X3Y148_SLICE_X2Y148_A5Q;
  assign CLBLM_R_X3Y148_SLICE_X2Y148_BMUX = CLBLM_R_X3Y148_SLICE_X2Y148_B5Q;
  assign CLBLM_R_X3Y148_SLICE_X2Y148_CMUX = CLBLM_R_X3Y148_SLICE_X2Y148_CO5;
  assign CLBLM_R_X3Y148_SLICE_X3Y148_A = CLBLM_R_X3Y148_SLICE_X3Y148_AO6;
  assign CLBLM_R_X3Y148_SLICE_X3Y148_B = CLBLM_R_X3Y148_SLICE_X3Y148_BO6;
  assign CLBLM_R_X3Y148_SLICE_X3Y148_C = CLBLM_R_X3Y148_SLICE_X3Y148_CO6;
  assign CLBLM_R_X3Y148_SLICE_X3Y148_D = CLBLM_R_X3Y148_SLICE_X3Y148_DO6;
  assign CLBLM_R_X3Y148_SLICE_X3Y148_BMUX = CLBLM_R_X3Y148_SLICE_X3Y148_B5Q;
  assign CLBLM_R_X3Y148_SLICE_X3Y148_CMUX = CLBLM_R_X3Y148_SLICE_X3Y148_C5Q;
  assign CLBLM_R_X3Y148_SLICE_X3Y148_DMUX = CLBLM_R_X3Y148_SLICE_X3Y148_DO5;
  assign CLBLM_R_X3Y149_SLICE_X2Y149_A = CLBLM_R_X3Y149_SLICE_X2Y149_AO6;
  assign CLBLM_R_X3Y149_SLICE_X2Y149_B = CLBLM_R_X3Y149_SLICE_X2Y149_BO6;
  assign CLBLM_R_X3Y149_SLICE_X2Y149_C = CLBLM_R_X3Y149_SLICE_X2Y149_CO6;
  assign CLBLM_R_X3Y149_SLICE_X2Y149_D = CLBLM_R_X3Y149_SLICE_X2Y149_DO6;
  assign CLBLM_R_X3Y149_SLICE_X2Y149_CMUX = CLBLM_R_X3Y149_SLICE_X2Y149_C5Q;
  assign CLBLM_R_X3Y149_SLICE_X3Y149_A = CLBLM_R_X3Y149_SLICE_X3Y149_AO6;
  assign CLBLM_R_X3Y149_SLICE_X3Y149_B = CLBLM_R_X3Y149_SLICE_X3Y149_BO6;
  assign CLBLM_R_X3Y149_SLICE_X3Y149_C = CLBLM_R_X3Y149_SLICE_X3Y149_CO6;
  assign CLBLM_R_X3Y149_SLICE_X3Y149_D = CLBLM_R_X3Y149_SLICE_X3Y149_DO6;
  assign CLBLM_R_X3Y149_SLICE_X3Y149_DMUX = CLBLM_R_X3Y149_SLICE_X3Y149_D5Q;
  assign CLBLM_R_X3Y150_SLICE_X2Y150_A = CLBLM_R_X3Y150_SLICE_X2Y150_AO6;
  assign CLBLM_R_X3Y150_SLICE_X2Y150_B = CLBLM_R_X3Y150_SLICE_X2Y150_BO6;
  assign CLBLM_R_X3Y150_SLICE_X2Y150_C = CLBLM_R_X3Y150_SLICE_X2Y150_CO6;
  assign CLBLM_R_X3Y150_SLICE_X2Y150_D = CLBLM_R_X3Y150_SLICE_X2Y150_DO6;
  assign CLBLM_R_X3Y150_SLICE_X2Y150_DMUX = CLBLM_R_X3Y150_SLICE_X2Y150_D5Q;
  assign CLBLM_R_X3Y150_SLICE_X3Y150_A = CLBLM_R_X3Y150_SLICE_X3Y150_AO6;
  assign CLBLM_R_X3Y150_SLICE_X3Y150_B = CLBLM_R_X3Y150_SLICE_X3Y150_BO6;
  assign CLBLM_R_X3Y150_SLICE_X3Y150_C = CLBLM_R_X3Y150_SLICE_X3Y150_CO6;
  assign CLBLM_R_X3Y150_SLICE_X3Y150_D = CLBLM_R_X3Y150_SLICE_X3Y150_DO6;
  assign CLBLM_R_X3Y150_SLICE_X3Y150_AMUX = CLBLM_R_X3Y150_SLICE_X3Y150_A5Q;
  assign CLBLM_R_X3Y150_SLICE_X3Y150_BMUX = CLBLM_R_X3Y150_SLICE_X3Y150_B5Q;
  assign CLBLM_R_X3Y150_SLICE_X3Y150_DMUX = CLBLM_R_X3Y150_SLICE_X3Y150_D5Q;
  assign CLBLM_R_X3Y151_SLICE_X2Y151_A = CLBLM_R_X3Y151_SLICE_X2Y151_AO6;
  assign CLBLM_R_X3Y151_SLICE_X2Y151_B = CLBLM_R_X3Y151_SLICE_X2Y151_BO6;
  assign CLBLM_R_X3Y151_SLICE_X2Y151_C = CLBLM_R_X3Y151_SLICE_X2Y151_CO6;
  assign CLBLM_R_X3Y151_SLICE_X2Y151_D = CLBLM_R_X3Y151_SLICE_X2Y151_DO6;
  assign CLBLM_R_X3Y151_SLICE_X2Y151_AMUX = CLBLM_R_X3Y151_SLICE_X2Y151_AO5;
  assign CLBLM_R_X3Y151_SLICE_X2Y151_BMUX = CLBLM_R_X3Y151_SLICE_X2Y151_BO5;
  assign CLBLM_R_X3Y151_SLICE_X3Y151_A = CLBLM_R_X3Y151_SLICE_X3Y151_AO6;
  assign CLBLM_R_X3Y151_SLICE_X3Y151_B = CLBLM_R_X3Y151_SLICE_X3Y151_BO6;
  assign CLBLM_R_X3Y151_SLICE_X3Y151_C = CLBLM_R_X3Y151_SLICE_X3Y151_CO6;
  assign CLBLM_R_X3Y151_SLICE_X3Y151_D = CLBLM_R_X3Y151_SLICE_X3Y151_DO6;
  assign CLBLM_R_X3Y151_SLICE_X3Y151_AMUX = CLBLM_R_X3Y151_SLICE_X3Y151_A5Q;
  assign CLBLM_R_X3Y151_SLICE_X3Y151_DMUX = CLBLM_R_X3Y151_SLICE_X3Y151_DO5;
  assign CLBLM_R_X3Y152_SLICE_X2Y152_A = CLBLM_R_X3Y152_SLICE_X2Y152_AO6;
  assign CLBLM_R_X3Y152_SLICE_X2Y152_B = CLBLM_R_X3Y152_SLICE_X2Y152_BO6;
  assign CLBLM_R_X3Y152_SLICE_X2Y152_C = CLBLM_R_X3Y152_SLICE_X2Y152_CO6;
  assign CLBLM_R_X3Y152_SLICE_X2Y152_D = CLBLM_R_X3Y152_SLICE_X2Y152_DO6;
  assign CLBLM_R_X3Y152_SLICE_X3Y152_A = CLBLM_R_X3Y152_SLICE_X3Y152_AO6;
  assign CLBLM_R_X3Y152_SLICE_X3Y152_B = CLBLM_R_X3Y152_SLICE_X3Y152_BO6;
  assign CLBLM_R_X3Y152_SLICE_X3Y152_C = CLBLM_R_X3Y152_SLICE_X3Y152_CO6;
  assign CLBLM_R_X3Y152_SLICE_X3Y152_D = CLBLM_R_X3Y152_SLICE_X3Y152_DO6;
  assign CLBLM_R_X3Y153_SLICE_X2Y153_A = CLBLM_R_X3Y153_SLICE_X2Y153_AO6;
  assign CLBLM_R_X3Y153_SLICE_X2Y153_B = CLBLM_R_X3Y153_SLICE_X2Y153_BO6;
  assign CLBLM_R_X3Y153_SLICE_X2Y153_C = CLBLM_R_X3Y153_SLICE_X2Y153_CO6;
  assign CLBLM_R_X3Y153_SLICE_X2Y153_D = CLBLM_R_X3Y153_SLICE_X2Y153_DO6;
  assign CLBLM_R_X3Y153_SLICE_X3Y153_A = CLBLM_R_X3Y153_SLICE_X3Y153_AO6;
  assign CLBLM_R_X3Y153_SLICE_X3Y153_B = CLBLM_R_X3Y153_SLICE_X3Y153_BO6;
  assign CLBLM_R_X3Y153_SLICE_X3Y153_C = CLBLM_R_X3Y153_SLICE_X3Y153_CO6;
  assign CLBLM_R_X3Y153_SLICE_X3Y153_D = CLBLM_R_X3Y153_SLICE_X3Y153_DO6;
  assign CLBLM_R_X5Y140_SLICE_X6Y140_A = CLBLM_R_X5Y140_SLICE_X6Y140_AO6;
  assign CLBLM_R_X5Y140_SLICE_X6Y140_B = CLBLM_R_X5Y140_SLICE_X6Y140_BO6;
  assign CLBLM_R_X5Y140_SLICE_X6Y140_C = CLBLM_R_X5Y140_SLICE_X6Y140_CO6;
  assign CLBLM_R_X5Y140_SLICE_X6Y140_D = CLBLM_R_X5Y140_SLICE_X6Y140_DO6;
  assign CLBLM_R_X5Y140_SLICE_X6Y140_AMUX = CLBLM_R_X5Y140_SLICE_X6Y140_A5Q;
  assign CLBLM_R_X5Y140_SLICE_X6Y140_DMUX = CLBLM_R_X5Y140_SLICE_X6Y140_DO5;
  assign CLBLM_R_X5Y140_SLICE_X7Y140_A = CLBLM_R_X5Y140_SLICE_X7Y140_AO6;
  assign CLBLM_R_X5Y140_SLICE_X7Y140_B = CLBLM_R_X5Y140_SLICE_X7Y140_BO6;
  assign CLBLM_R_X5Y140_SLICE_X7Y140_C = CLBLM_R_X5Y140_SLICE_X7Y140_CO6;
  assign CLBLM_R_X5Y140_SLICE_X7Y140_D = CLBLM_R_X5Y140_SLICE_X7Y140_DO6;
  assign CLBLM_R_X5Y141_SLICE_X6Y141_A = CLBLM_R_X5Y141_SLICE_X6Y141_AO6;
  assign CLBLM_R_X5Y141_SLICE_X6Y141_B = CLBLM_R_X5Y141_SLICE_X6Y141_BO6;
  assign CLBLM_R_X5Y141_SLICE_X6Y141_C = CLBLM_R_X5Y141_SLICE_X6Y141_CO6;
  assign CLBLM_R_X5Y141_SLICE_X6Y141_D = CLBLM_R_X5Y141_SLICE_X6Y141_DO6;
  assign CLBLM_R_X5Y141_SLICE_X6Y141_BMUX = CLBLM_R_X5Y141_SLICE_X6Y141_B5Q;
  assign CLBLM_R_X5Y141_SLICE_X6Y141_CMUX = CLBLM_R_X5Y141_SLICE_X6Y141_CO5;
  assign CLBLM_R_X5Y141_SLICE_X6Y141_DMUX = CLBLM_R_X5Y141_SLICE_X6Y141_D5Q;
  assign CLBLM_R_X5Y141_SLICE_X7Y141_A = CLBLM_R_X5Y141_SLICE_X7Y141_AO6;
  assign CLBLM_R_X5Y141_SLICE_X7Y141_B = CLBLM_R_X5Y141_SLICE_X7Y141_BO6;
  assign CLBLM_R_X5Y141_SLICE_X7Y141_C = CLBLM_R_X5Y141_SLICE_X7Y141_CO6;
  assign CLBLM_R_X5Y141_SLICE_X7Y141_D = CLBLM_R_X5Y141_SLICE_X7Y141_DO6;
  assign CLBLM_R_X5Y142_SLICE_X6Y142_A = CLBLM_R_X5Y142_SLICE_X6Y142_AO6;
  assign CLBLM_R_X5Y142_SLICE_X6Y142_B = CLBLM_R_X5Y142_SLICE_X6Y142_BO6;
  assign CLBLM_R_X5Y142_SLICE_X6Y142_C = CLBLM_R_X5Y142_SLICE_X6Y142_CO6;
  assign CLBLM_R_X5Y142_SLICE_X6Y142_D = CLBLM_R_X5Y142_SLICE_X6Y142_DO6;
  assign CLBLM_R_X5Y142_SLICE_X6Y142_DMUX = CLBLM_R_X5Y142_SLICE_X6Y142_D5Q;
  assign CLBLM_R_X5Y142_SLICE_X7Y142_A = CLBLM_R_X5Y142_SLICE_X7Y142_AO6;
  assign CLBLM_R_X5Y142_SLICE_X7Y142_B = CLBLM_R_X5Y142_SLICE_X7Y142_BO6;
  assign CLBLM_R_X5Y142_SLICE_X7Y142_C = CLBLM_R_X5Y142_SLICE_X7Y142_CO6;
  assign CLBLM_R_X5Y142_SLICE_X7Y142_D = CLBLM_R_X5Y142_SLICE_X7Y142_DO6;
  assign CLBLM_R_X5Y142_SLICE_X7Y142_AMUX = CLBLM_R_X5Y142_SLICE_X7Y142_A5Q;
  assign CLBLM_R_X5Y143_SLICE_X6Y143_A = CLBLM_R_X5Y143_SLICE_X6Y143_AO6;
  assign CLBLM_R_X5Y143_SLICE_X6Y143_B = CLBLM_R_X5Y143_SLICE_X6Y143_BO6;
  assign CLBLM_R_X5Y143_SLICE_X6Y143_C = CLBLM_R_X5Y143_SLICE_X6Y143_CO6;
  assign CLBLM_R_X5Y143_SLICE_X6Y143_D = CLBLM_R_X5Y143_SLICE_X6Y143_DO6;
  assign CLBLM_R_X5Y143_SLICE_X6Y143_CMUX = CLBLM_R_X5Y143_SLICE_X6Y143_C5Q;
  assign CLBLM_R_X5Y143_SLICE_X6Y143_DMUX = CLBLM_R_X5Y143_SLICE_X6Y143_D5Q;
  assign CLBLM_R_X5Y143_SLICE_X7Y143_A = CLBLM_R_X5Y143_SLICE_X7Y143_AO6;
  assign CLBLM_R_X5Y143_SLICE_X7Y143_B = CLBLM_R_X5Y143_SLICE_X7Y143_BO6;
  assign CLBLM_R_X5Y143_SLICE_X7Y143_C = CLBLM_R_X5Y143_SLICE_X7Y143_CO6;
  assign CLBLM_R_X5Y143_SLICE_X7Y143_D = CLBLM_R_X5Y143_SLICE_X7Y143_DO6;
  assign CLBLM_R_X5Y143_SLICE_X7Y143_CMUX = CLBLM_R_X5Y143_SLICE_X7Y143_C5Q;
  assign CLBLM_R_X5Y143_SLICE_X7Y143_DMUX = CLBLM_R_X5Y143_SLICE_X7Y143_DO6;
  assign CLBLM_R_X5Y144_SLICE_X6Y144_A = CLBLM_R_X5Y144_SLICE_X6Y144_AO6;
  assign CLBLM_R_X5Y144_SLICE_X6Y144_B = CLBLM_R_X5Y144_SLICE_X6Y144_BO6;
  assign CLBLM_R_X5Y144_SLICE_X6Y144_C = CLBLM_R_X5Y144_SLICE_X6Y144_CO6;
  assign CLBLM_R_X5Y144_SLICE_X6Y144_D = CLBLM_R_X5Y144_SLICE_X6Y144_DO6;
  assign CLBLM_R_X5Y144_SLICE_X6Y144_DMUX = CLBLM_R_X5Y144_SLICE_X6Y144_D5Q;
  assign CLBLM_R_X5Y144_SLICE_X7Y144_A = CLBLM_R_X5Y144_SLICE_X7Y144_AO6;
  assign CLBLM_R_X5Y144_SLICE_X7Y144_B = CLBLM_R_X5Y144_SLICE_X7Y144_BO6;
  assign CLBLM_R_X5Y144_SLICE_X7Y144_C = CLBLM_R_X5Y144_SLICE_X7Y144_CO6;
  assign CLBLM_R_X5Y144_SLICE_X7Y144_D = CLBLM_R_X5Y144_SLICE_X7Y144_DO6;
  assign CLBLM_R_X5Y144_SLICE_X7Y144_BMUX = CLBLM_R_X5Y144_SLICE_X7Y144_B5Q;
  assign CLBLM_R_X5Y144_SLICE_X7Y144_CMUX = CLBLM_R_X5Y144_SLICE_X7Y144_C5Q;
  assign CLBLM_R_X5Y144_SLICE_X7Y144_DMUX = CLBLM_R_X5Y144_SLICE_X7Y144_DO6;
  assign CLBLM_R_X5Y145_SLICE_X6Y145_A = CLBLM_R_X5Y145_SLICE_X6Y145_AO6;
  assign CLBLM_R_X5Y145_SLICE_X6Y145_B = CLBLM_R_X5Y145_SLICE_X6Y145_BO6;
  assign CLBLM_R_X5Y145_SLICE_X6Y145_C = CLBLM_R_X5Y145_SLICE_X6Y145_CO6;
  assign CLBLM_R_X5Y145_SLICE_X6Y145_D = CLBLM_R_X5Y145_SLICE_X6Y145_DO6;
  assign CLBLM_R_X5Y145_SLICE_X6Y145_BMUX = CLBLM_R_X5Y145_SLICE_X6Y145_B5Q;
  assign CLBLM_R_X5Y145_SLICE_X6Y145_CMUX = CLBLM_R_X5Y145_SLICE_X6Y145_C5Q;
  assign CLBLM_R_X5Y145_SLICE_X6Y145_DMUX = CLBLM_R_X5Y145_SLICE_X6Y145_D5Q;
  assign CLBLM_R_X5Y145_SLICE_X7Y145_A = CLBLM_R_X5Y145_SLICE_X7Y145_AO6;
  assign CLBLM_R_X5Y145_SLICE_X7Y145_B = CLBLM_R_X5Y145_SLICE_X7Y145_BO6;
  assign CLBLM_R_X5Y145_SLICE_X7Y145_C = CLBLM_R_X5Y145_SLICE_X7Y145_CO6;
  assign CLBLM_R_X5Y145_SLICE_X7Y145_D = CLBLM_R_X5Y145_SLICE_X7Y145_DO6;
  assign CLBLM_R_X5Y145_SLICE_X7Y145_AMUX = CLBLM_R_X5Y145_SLICE_X7Y145_A5Q;
  assign CLBLM_R_X5Y145_SLICE_X7Y145_BMUX = CLBLM_R_X5Y145_SLICE_X7Y145_B5Q;
  assign CLBLM_R_X5Y146_SLICE_X6Y146_A = CLBLM_R_X5Y146_SLICE_X6Y146_AO6;
  assign CLBLM_R_X5Y146_SLICE_X6Y146_B = CLBLM_R_X5Y146_SLICE_X6Y146_BO6;
  assign CLBLM_R_X5Y146_SLICE_X6Y146_C = CLBLM_R_X5Y146_SLICE_X6Y146_CO6;
  assign CLBLM_R_X5Y146_SLICE_X6Y146_D = CLBLM_R_X5Y146_SLICE_X6Y146_DO6;
  assign CLBLM_R_X5Y146_SLICE_X6Y146_BMUX = CLBLM_R_X5Y146_SLICE_X6Y146_B5Q;
  assign CLBLM_R_X5Y146_SLICE_X7Y146_A = CLBLM_R_X5Y146_SLICE_X7Y146_AO6;
  assign CLBLM_R_X5Y146_SLICE_X7Y146_B = CLBLM_R_X5Y146_SLICE_X7Y146_BO6;
  assign CLBLM_R_X5Y146_SLICE_X7Y146_C = CLBLM_R_X5Y146_SLICE_X7Y146_CO6;
  assign CLBLM_R_X5Y146_SLICE_X7Y146_D = CLBLM_R_X5Y146_SLICE_X7Y146_DO6;
  assign CLBLM_R_X5Y146_SLICE_X7Y146_CMUX = CLBLM_R_X5Y146_SLICE_X7Y146_C5Q;
  assign CLBLM_R_X5Y146_SLICE_X7Y146_DMUX = CLBLM_R_X5Y146_SLICE_X7Y146_D5Q;
  assign CLBLM_R_X5Y147_SLICE_X6Y147_A = CLBLM_R_X5Y147_SLICE_X6Y147_AO6;
  assign CLBLM_R_X5Y147_SLICE_X6Y147_B = CLBLM_R_X5Y147_SLICE_X6Y147_BO6;
  assign CLBLM_R_X5Y147_SLICE_X6Y147_C = CLBLM_R_X5Y147_SLICE_X6Y147_CO6;
  assign CLBLM_R_X5Y147_SLICE_X6Y147_D = CLBLM_R_X5Y147_SLICE_X6Y147_DO6;
  assign CLBLM_R_X5Y147_SLICE_X6Y147_BMUX = CLBLM_R_X5Y147_SLICE_X6Y147_B5Q;
  assign CLBLM_R_X5Y147_SLICE_X6Y147_CMUX = CLBLM_R_X5Y147_SLICE_X6Y147_C5Q;
  assign CLBLM_R_X5Y147_SLICE_X7Y147_A = CLBLM_R_X5Y147_SLICE_X7Y147_AO6;
  assign CLBLM_R_X5Y147_SLICE_X7Y147_B = CLBLM_R_X5Y147_SLICE_X7Y147_BO6;
  assign CLBLM_R_X5Y147_SLICE_X7Y147_C = CLBLM_R_X5Y147_SLICE_X7Y147_CO6;
  assign CLBLM_R_X5Y147_SLICE_X7Y147_D = CLBLM_R_X5Y147_SLICE_X7Y147_DO6;
  assign CLBLM_R_X5Y147_SLICE_X7Y147_BMUX = CLBLM_R_X5Y147_SLICE_X7Y147_B5Q;
  assign CLBLM_R_X5Y147_SLICE_X7Y147_CMUX = CLBLM_R_X5Y147_SLICE_X7Y147_C5Q;
  assign CLBLM_R_X5Y148_SLICE_X6Y148_A = CLBLM_R_X5Y148_SLICE_X6Y148_AO6;
  assign CLBLM_R_X5Y148_SLICE_X6Y148_B = CLBLM_R_X5Y148_SLICE_X6Y148_BO6;
  assign CLBLM_R_X5Y148_SLICE_X6Y148_C = CLBLM_R_X5Y148_SLICE_X6Y148_CO6;
  assign CLBLM_R_X5Y148_SLICE_X6Y148_D = CLBLM_R_X5Y148_SLICE_X6Y148_DO6;
  assign CLBLM_R_X5Y148_SLICE_X6Y148_AMUX = CLBLM_R_X5Y148_SLICE_X6Y148_AO5;
  assign CLBLM_R_X5Y148_SLICE_X7Y148_A = CLBLM_R_X5Y148_SLICE_X7Y148_AO6;
  assign CLBLM_R_X5Y148_SLICE_X7Y148_B = CLBLM_R_X5Y148_SLICE_X7Y148_BO6;
  assign CLBLM_R_X5Y148_SLICE_X7Y148_C = CLBLM_R_X5Y148_SLICE_X7Y148_CO6;
  assign CLBLM_R_X5Y148_SLICE_X7Y148_D = CLBLM_R_X5Y148_SLICE_X7Y148_DO6;
  assign CLBLM_R_X5Y148_SLICE_X7Y148_CMUX = CLBLM_R_X5Y148_SLICE_X7Y148_C5Q;
  assign CLBLM_R_X5Y148_SLICE_X7Y148_DMUX = CLBLM_R_X5Y148_SLICE_X7Y148_DO6;
  assign CLBLM_R_X5Y149_SLICE_X6Y149_A = CLBLM_R_X5Y149_SLICE_X6Y149_AO6;
  assign CLBLM_R_X5Y149_SLICE_X6Y149_B = CLBLM_R_X5Y149_SLICE_X6Y149_BO6;
  assign CLBLM_R_X5Y149_SLICE_X6Y149_C = CLBLM_R_X5Y149_SLICE_X6Y149_CO6;
  assign CLBLM_R_X5Y149_SLICE_X6Y149_D = CLBLM_R_X5Y149_SLICE_X6Y149_DO6;
  assign CLBLM_R_X5Y149_SLICE_X6Y149_BMUX = CLBLM_R_X5Y149_SLICE_X6Y149_B5Q;
  assign CLBLM_R_X5Y149_SLICE_X6Y149_CMUX = CLBLM_R_X5Y149_SLICE_X6Y149_C5Q;
  assign CLBLM_R_X5Y149_SLICE_X7Y149_A = CLBLM_R_X5Y149_SLICE_X7Y149_AO6;
  assign CLBLM_R_X5Y149_SLICE_X7Y149_B = CLBLM_R_X5Y149_SLICE_X7Y149_BO6;
  assign CLBLM_R_X5Y149_SLICE_X7Y149_C = CLBLM_R_X5Y149_SLICE_X7Y149_CO6;
  assign CLBLM_R_X5Y149_SLICE_X7Y149_D = CLBLM_R_X5Y149_SLICE_X7Y149_DO6;
  assign CLBLM_R_X5Y149_SLICE_X7Y149_CMUX = CLBLM_R_X5Y149_SLICE_X7Y149_C5Q;
  assign CLBLM_R_X5Y149_SLICE_X7Y149_DMUX = CLBLM_R_X5Y149_SLICE_X7Y149_D5Q;
  assign CLBLM_R_X5Y150_SLICE_X6Y150_A = CLBLM_R_X5Y150_SLICE_X6Y150_AO6;
  assign CLBLM_R_X5Y150_SLICE_X6Y150_B = CLBLM_R_X5Y150_SLICE_X6Y150_BO6;
  assign CLBLM_R_X5Y150_SLICE_X6Y150_C = CLBLM_R_X5Y150_SLICE_X6Y150_CO6;
  assign CLBLM_R_X5Y150_SLICE_X6Y150_D = CLBLM_R_X5Y150_SLICE_X6Y150_DO6;
  assign CLBLM_R_X5Y150_SLICE_X6Y150_AMUX = CLBLM_R_X5Y150_SLICE_X6Y150_A5Q;
  assign CLBLM_R_X5Y150_SLICE_X6Y150_BMUX = CLBLM_R_X5Y150_SLICE_X6Y150_B5Q;
  assign CLBLM_R_X5Y150_SLICE_X6Y150_CMUX = CLBLM_R_X5Y150_SLICE_X6Y150_C5Q;
  assign CLBLM_R_X5Y150_SLICE_X7Y150_A = CLBLM_R_X5Y150_SLICE_X7Y150_AO6;
  assign CLBLM_R_X5Y150_SLICE_X7Y150_B = CLBLM_R_X5Y150_SLICE_X7Y150_BO6;
  assign CLBLM_R_X5Y150_SLICE_X7Y150_C = CLBLM_R_X5Y150_SLICE_X7Y150_CO6;
  assign CLBLM_R_X5Y150_SLICE_X7Y150_D = CLBLM_R_X5Y150_SLICE_X7Y150_DO6;
  assign CLBLM_R_X5Y150_SLICE_X7Y150_AMUX = CLBLM_R_X5Y150_SLICE_X7Y150_A5Q;
  assign CLBLM_R_X5Y150_SLICE_X7Y150_DMUX = CLBLM_R_X5Y150_SLICE_X7Y150_DO6;
  assign CLBLM_R_X5Y151_SLICE_X6Y151_A = CLBLM_R_X5Y151_SLICE_X6Y151_AO6;
  assign CLBLM_R_X5Y151_SLICE_X6Y151_B = CLBLM_R_X5Y151_SLICE_X6Y151_BO6;
  assign CLBLM_R_X5Y151_SLICE_X6Y151_C = CLBLM_R_X5Y151_SLICE_X6Y151_CO6;
  assign CLBLM_R_X5Y151_SLICE_X6Y151_D = CLBLM_R_X5Y151_SLICE_X6Y151_DO6;
  assign CLBLM_R_X5Y151_SLICE_X6Y151_CMUX = CLBLM_R_X5Y151_SLICE_X6Y151_C5Q;
  assign CLBLM_R_X5Y151_SLICE_X7Y151_A = CLBLM_R_X5Y151_SLICE_X7Y151_AO6;
  assign CLBLM_R_X5Y151_SLICE_X7Y151_B = CLBLM_R_X5Y151_SLICE_X7Y151_BO6;
  assign CLBLM_R_X5Y151_SLICE_X7Y151_C = CLBLM_R_X5Y151_SLICE_X7Y151_CO6;
  assign CLBLM_R_X5Y151_SLICE_X7Y151_D = CLBLM_R_X5Y151_SLICE_X7Y151_DO6;
  assign CLBLM_R_X5Y151_SLICE_X7Y151_BMUX = CLBLM_R_X5Y151_SLICE_X7Y151_B5Q;
  assign CLBLM_R_X5Y151_SLICE_X7Y151_DMUX = CLBLM_R_X5Y151_SLICE_X7Y151_DO6;
  assign CLBLM_R_X5Y152_SLICE_X6Y152_A = CLBLM_R_X5Y152_SLICE_X6Y152_AO6;
  assign CLBLM_R_X5Y152_SLICE_X6Y152_B = CLBLM_R_X5Y152_SLICE_X6Y152_BO6;
  assign CLBLM_R_X5Y152_SLICE_X6Y152_C = CLBLM_R_X5Y152_SLICE_X6Y152_CO6;
  assign CLBLM_R_X5Y152_SLICE_X6Y152_D = CLBLM_R_X5Y152_SLICE_X6Y152_DO6;
  assign CLBLM_R_X5Y152_SLICE_X6Y152_BMUX = CLBLM_R_X5Y152_SLICE_X6Y152_B5Q;
  assign CLBLM_R_X5Y152_SLICE_X7Y152_A = CLBLM_R_X5Y152_SLICE_X7Y152_AO6;
  assign CLBLM_R_X5Y152_SLICE_X7Y152_B = CLBLM_R_X5Y152_SLICE_X7Y152_BO6;
  assign CLBLM_R_X5Y152_SLICE_X7Y152_C = CLBLM_R_X5Y152_SLICE_X7Y152_CO6;
  assign CLBLM_R_X5Y152_SLICE_X7Y152_D = CLBLM_R_X5Y152_SLICE_X7Y152_DO6;
  assign CLBLM_R_X5Y152_SLICE_X7Y152_AMUX = CLBLM_R_X5Y152_SLICE_X7Y152_A5Q;
  assign CLBLM_R_X5Y152_SLICE_X7Y152_BMUX = CLBLM_R_X5Y152_SLICE_X7Y152_B5Q;
  assign CLBLM_R_X5Y152_SLICE_X7Y152_CMUX = CLBLM_R_X5Y152_SLICE_X7Y152_C5Q;
  assign CLBLM_R_X5Y153_SLICE_X6Y153_A = CLBLM_R_X5Y153_SLICE_X6Y153_AO6;
  assign CLBLM_R_X5Y153_SLICE_X6Y153_B = CLBLM_R_X5Y153_SLICE_X6Y153_BO6;
  assign CLBLM_R_X5Y153_SLICE_X6Y153_C = CLBLM_R_X5Y153_SLICE_X6Y153_CO6;
  assign CLBLM_R_X5Y153_SLICE_X6Y153_D = CLBLM_R_X5Y153_SLICE_X6Y153_DO6;
  assign CLBLM_R_X5Y153_SLICE_X6Y153_AMUX = CLBLM_R_X5Y153_SLICE_X6Y153_A5Q;
  assign CLBLM_R_X5Y153_SLICE_X6Y153_BMUX = CLBLM_R_X5Y153_SLICE_X6Y153_B5Q;
  assign CLBLM_R_X5Y153_SLICE_X6Y153_DMUX = CLBLM_R_X5Y153_SLICE_X6Y153_D5Q;
  assign CLBLM_R_X5Y153_SLICE_X7Y153_A = CLBLM_R_X5Y153_SLICE_X7Y153_AO6;
  assign CLBLM_R_X5Y153_SLICE_X7Y153_B = CLBLM_R_X5Y153_SLICE_X7Y153_BO6;
  assign CLBLM_R_X5Y153_SLICE_X7Y153_C = CLBLM_R_X5Y153_SLICE_X7Y153_CO6;
  assign CLBLM_R_X5Y153_SLICE_X7Y153_D = CLBLM_R_X5Y153_SLICE_X7Y153_DO6;
  assign CLBLM_R_X5Y153_SLICE_X7Y153_DMUX = CLBLM_R_X5Y153_SLICE_X7Y153_DO5;
  assign CLBLM_R_X5Y154_SLICE_X6Y154_A = CLBLM_R_X5Y154_SLICE_X6Y154_AO6;
  assign CLBLM_R_X5Y154_SLICE_X6Y154_B = CLBLM_R_X5Y154_SLICE_X6Y154_BO6;
  assign CLBLM_R_X5Y154_SLICE_X6Y154_C = CLBLM_R_X5Y154_SLICE_X6Y154_CO6;
  assign CLBLM_R_X5Y154_SLICE_X6Y154_D = CLBLM_R_X5Y154_SLICE_X6Y154_DO6;
  assign CLBLM_R_X5Y154_SLICE_X7Y154_A = CLBLM_R_X5Y154_SLICE_X7Y154_AO6;
  assign CLBLM_R_X5Y154_SLICE_X7Y154_B = CLBLM_R_X5Y154_SLICE_X7Y154_BO6;
  assign CLBLM_R_X5Y154_SLICE_X7Y154_C = CLBLM_R_X5Y154_SLICE_X7Y154_CO6;
  assign CLBLM_R_X5Y154_SLICE_X7Y154_D = CLBLM_R_X5Y154_SLICE_X7Y154_DO6;
  assign CLBLM_R_X7Y141_SLICE_X8Y141_A = CLBLM_R_X7Y141_SLICE_X8Y141_AO6;
  assign CLBLM_R_X7Y141_SLICE_X8Y141_B = CLBLM_R_X7Y141_SLICE_X8Y141_BO6;
  assign CLBLM_R_X7Y141_SLICE_X8Y141_C = CLBLM_R_X7Y141_SLICE_X8Y141_CO6;
  assign CLBLM_R_X7Y141_SLICE_X8Y141_D = CLBLM_R_X7Y141_SLICE_X8Y141_DO6;
  assign CLBLM_R_X7Y141_SLICE_X8Y141_AMUX = CLBLM_R_X7Y141_SLICE_X8Y141_AO5;
  assign CLBLM_R_X7Y141_SLICE_X9Y141_A = CLBLM_R_X7Y141_SLICE_X9Y141_AO6;
  assign CLBLM_R_X7Y141_SLICE_X9Y141_B = CLBLM_R_X7Y141_SLICE_X9Y141_BO6;
  assign CLBLM_R_X7Y141_SLICE_X9Y141_C = CLBLM_R_X7Y141_SLICE_X9Y141_CO6;
  assign CLBLM_R_X7Y141_SLICE_X9Y141_D = CLBLM_R_X7Y141_SLICE_X9Y141_DO6;
  assign CLBLM_R_X7Y142_SLICE_X8Y142_A = CLBLM_R_X7Y142_SLICE_X8Y142_AO6;
  assign CLBLM_R_X7Y142_SLICE_X8Y142_B = CLBLM_R_X7Y142_SLICE_X8Y142_BO6;
  assign CLBLM_R_X7Y142_SLICE_X8Y142_C = CLBLM_R_X7Y142_SLICE_X8Y142_CO6;
  assign CLBLM_R_X7Y142_SLICE_X8Y142_D = CLBLM_R_X7Y142_SLICE_X8Y142_DO6;
  assign CLBLM_R_X7Y142_SLICE_X8Y142_CMUX = CLBLM_R_X7Y142_SLICE_X8Y142_C5Q;
  assign CLBLM_R_X7Y142_SLICE_X8Y142_DMUX = CLBLM_R_X7Y142_SLICE_X8Y142_D5Q;
  assign CLBLM_R_X7Y142_SLICE_X9Y142_A = CLBLM_R_X7Y142_SLICE_X9Y142_AO6;
  assign CLBLM_R_X7Y142_SLICE_X9Y142_B = CLBLM_R_X7Y142_SLICE_X9Y142_BO6;
  assign CLBLM_R_X7Y142_SLICE_X9Y142_C = CLBLM_R_X7Y142_SLICE_X9Y142_CO6;
  assign CLBLM_R_X7Y142_SLICE_X9Y142_D = CLBLM_R_X7Y142_SLICE_X9Y142_DO6;
  assign CLBLM_R_X7Y143_SLICE_X8Y143_A = CLBLM_R_X7Y143_SLICE_X8Y143_AO6;
  assign CLBLM_R_X7Y143_SLICE_X8Y143_B = CLBLM_R_X7Y143_SLICE_X8Y143_BO6;
  assign CLBLM_R_X7Y143_SLICE_X8Y143_C = CLBLM_R_X7Y143_SLICE_X8Y143_CO6;
  assign CLBLM_R_X7Y143_SLICE_X8Y143_D = CLBLM_R_X7Y143_SLICE_X8Y143_DO6;
  assign CLBLM_R_X7Y143_SLICE_X8Y143_CMUX = CLBLM_R_X7Y143_SLICE_X8Y143_CO5;
  assign CLBLM_R_X7Y143_SLICE_X9Y143_A = CLBLM_R_X7Y143_SLICE_X9Y143_AO6;
  assign CLBLM_R_X7Y143_SLICE_X9Y143_B = CLBLM_R_X7Y143_SLICE_X9Y143_BO6;
  assign CLBLM_R_X7Y143_SLICE_X9Y143_C = CLBLM_R_X7Y143_SLICE_X9Y143_CO6;
  assign CLBLM_R_X7Y143_SLICE_X9Y143_D = CLBLM_R_X7Y143_SLICE_X9Y143_DO6;
  assign CLBLM_R_X7Y143_SLICE_X9Y143_BMUX = CLBLM_R_X7Y143_SLICE_X9Y143_B5Q;
  assign CLBLM_R_X7Y144_SLICE_X8Y144_A = CLBLM_R_X7Y144_SLICE_X8Y144_AO6;
  assign CLBLM_R_X7Y144_SLICE_X8Y144_B = CLBLM_R_X7Y144_SLICE_X8Y144_BO6;
  assign CLBLM_R_X7Y144_SLICE_X8Y144_C = CLBLM_R_X7Y144_SLICE_X8Y144_CO6;
  assign CLBLM_R_X7Y144_SLICE_X8Y144_D = CLBLM_R_X7Y144_SLICE_X8Y144_DO6;
  assign CLBLM_R_X7Y144_SLICE_X8Y144_BMUX = CLBLM_R_X7Y144_SLICE_X8Y144_B5Q;
  assign CLBLM_R_X7Y144_SLICE_X8Y144_CMUX = CLBLM_R_X7Y144_SLICE_X8Y144_C5Q;
  assign CLBLM_R_X7Y144_SLICE_X8Y144_DMUX = CLBLM_R_X7Y144_SLICE_X8Y144_D5Q;
  assign CLBLM_R_X7Y144_SLICE_X9Y144_A = CLBLM_R_X7Y144_SLICE_X9Y144_AO6;
  assign CLBLM_R_X7Y144_SLICE_X9Y144_B = CLBLM_R_X7Y144_SLICE_X9Y144_BO6;
  assign CLBLM_R_X7Y144_SLICE_X9Y144_C = CLBLM_R_X7Y144_SLICE_X9Y144_CO6;
  assign CLBLM_R_X7Y144_SLICE_X9Y144_D = CLBLM_R_X7Y144_SLICE_X9Y144_DO6;
  assign CLBLM_R_X7Y144_SLICE_X9Y144_AMUX = CLBLM_R_X7Y144_SLICE_X9Y144_A5Q;
  assign CLBLM_R_X7Y144_SLICE_X9Y144_BMUX = CLBLM_R_X7Y144_SLICE_X9Y144_B5Q;
  assign CLBLM_R_X7Y145_SLICE_X8Y145_A = CLBLM_R_X7Y145_SLICE_X8Y145_AO6;
  assign CLBLM_R_X7Y145_SLICE_X8Y145_B = CLBLM_R_X7Y145_SLICE_X8Y145_BO6;
  assign CLBLM_R_X7Y145_SLICE_X8Y145_C = CLBLM_R_X7Y145_SLICE_X8Y145_CO6;
  assign CLBLM_R_X7Y145_SLICE_X8Y145_D = CLBLM_R_X7Y145_SLICE_X8Y145_DO6;
  assign CLBLM_R_X7Y145_SLICE_X8Y145_AMUX = CLBLM_R_X7Y145_SLICE_X8Y145_A5Q;
  assign CLBLM_R_X7Y145_SLICE_X8Y145_BMUX = CLBLM_R_X7Y145_SLICE_X8Y145_B5Q;
  assign CLBLM_R_X7Y145_SLICE_X8Y145_CMUX = CLBLM_R_X7Y145_SLICE_X8Y145_C5Q;
  assign CLBLM_R_X7Y145_SLICE_X8Y145_DMUX = CLBLM_R_X7Y145_SLICE_X8Y145_D5Q;
  assign CLBLM_R_X7Y145_SLICE_X9Y145_A = CLBLM_R_X7Y145_SLICE_X9Y145_AO6;
  assign CLBLM_R_X7Y145_SLICE_X9Y145_B = CLBLM_R_X7Y145_SLICE_X9Y145_BO6;
  assign CLBLM_R_X7Y145_SLICE_X9Y145_C = CLBLM_R_X7Y145_SLICE_X9Y145_CO6;
  assign CLBLM_R_X7Y145_SLICE_X9Y145_D = CLBLM_R_X7Y145_SLICE_X9Y145_DO6;
  assign CLBLM_R_X7Y145_SLICE_X9Y145_DMUX = CLBLM_R_X7Y145_SLICE_X9Y145_DO6;
  assign CLBLM_R_X7Y146_SLICE_X8Y146_A = CLBLM_R_X7Y146_SLICE_X8Y146_AO6;
  assign CLBLM_R_X7Y146_SLICE_X8Y146_B = CLBLM_R_X7Y146_SLICE_X8Y146_BO6;
  assign CLBLM_R_X7Y146_SLICE_X8Y146_C = CLBLM_R_X7Y146_SLICE_X8Y146_CO6;
  assign CLBLM_R_X7Y146_SLICE_X8Y146_D = CLBLM_R_X7Y146_SLICE_X8Y146_DO6;
  assign CLBLM_R_X7Y146_SLICE_X8Y146_AMUX = CLBLM_R_X7Y146_SLICE_X8Y146_A5Q;
  assign CLBLM_R_X7Y146_SLICE_X8Y146_BMUX = CLBLM_R_X7Y146_SLICE_X8Y146_B5Q;
  assign CLBLM_R_X7Y146_SLICE_X8Y146_CMUX = CLBLM_R_X7Y146_SLICE_X8Y146_C5Q;
  assign CLBLM_R_X7Y146_SLICE_X8Y146_DMUX = CLBLM_R_X7Y146_SLICE_X8Y146_D5Q;
  assign CLBLM_R_X7Y146_SLICE_X9Y146_A = CLBLM_R_X7Y146_SLICE_X9Y146_AO6;
  assign CLBLM_R_X7Y146_SLICE_X9Y146_B = CLBLM_R_X7Y146_SLICE_X9Y146_BO6;
  assign CLBLM_R_X7Y146_SLICE_X9Y146_C = CLBLM_R_X7Y146_SLICE_X9Y146_CO6;
  assign CLBLM_R_X7Y146_SLICE_X9Y146_D = CLBLM_R_X7Y146_SLICE_X9Y146_DO6;
  assign CLBLM_R_X7Y146_SLICE_X9Y146_CMUX = CLBLM_R_X7Y146_SLICE_X9Y146_CO5;
  assign CLBLM_R_X7Y147_SLICE_X8Y147_A = CLBLM_R_X7Y147_SLICE_X8Y147_AO6;
  assign CLBLM_R_X7Y147_SLICE_X8Y147_B = CLBLM_R_X7Y147_SLICE_X8Y147_BO6;
  assign CLBLM_R_X7Y147_SLICE_X8Y147_C = CLBLM_R_X7Y147_SLICE_X8Y147_CO6;
  assign CLBLM_R_X7Y147_SLICE_X8Y147_D = CLBLM_R_X7Y147_SLICE_X8Y147_DO6;
  assign CLBLM_R_X7Y147_SLICE_X8Y147_BMUX = CLBLM_R_X7Y147_SLICE_X8Y147_BO6;
  assign CLBLM_R_X7Y147_SLICE_X8Y147_CMUX = CLBLM_R_X7Y147_SLICE_X8Y147_CO6;
  assign CLBLM_R_X7Y147_SLICE_X9Y147_A = CLBLM_R_X7Y147_SLICE_X9Y147_AO6;
  assign CLBLM_R_X7Y147_SLICE_X9Y147_B = CLBLM_R_X7Y147_SLICE_X9Y147_BO6;
  assign CLBLM_R_X7Y147_SLICE_X9Y147_C = CLBLM_R_X7Y147_SLICE_X9Y147_CO6;
  assign CLBLM_R_X7Y147_SLICE_X9Y147_D = CLBLM_R_X7Y147_SLICE_X9Y147_DO6;
  assign CLBLM_R_X7Y147_SLICE_X9Y147_AMUX = CLBLM_R_X7Y147_SLICE_X9Y147_A5Q;
  assign CLBLM_R_X7Y147_SLICE_X9Y147_CMUX = CLBLM_R_X7Y147_SLICE_X9Y147_C5Q;
  assign CLBLM_R_X7Y147_SLICE_X9Y147_DMUX = CLBLM_R_X7Y147_SLICE_X9Y147_D5Q;
  assign CLBLM_R_X7Y148_SLICE_X8Y148_A = CLBLM_R_X7Y148_SLICE_X8Y148_AO6;
  assign CLBLM_R_X7Y148_SLICE_X8Y148_B = CLBLM_R_X7Y148_SLICE_X8Y148_BO6;
  assign CLBLM_R_X7Y148_SLICE_X8Y148_C = CLBLM_R_X7Y148_SLICE_X8Y148_CO6;
  assign CLBLM_R_X7Y148_SLICE_X8Y148_D = CLBLM_R_X7Y148_SLICE_X8Y148_DO6;
  assign CLBLM_R_X7Y148_SLICE_X8Y148_AMUX = CLBLM_R_X7Y148_SLICE_X8Y148_AO5;
  assign CLBLM_R_X7Y148_SLICE_X9Y148_A = CLBLM_R_X7Y148_SLICE_X9Y148_AO6;
  assign CLBLM_R_X7Y148_SLICE_X9Y148_B = CLBLM_R_X7Y148_SLICE_X9Y148_BO6;
  assign CLBLM_R_X7Y148_SLICE_X9Y148_C = CLBLM_R_X7Y148_SLICE_X9Y148_CO6;
  assign CLBLM_R_X7Y148_SLICE_X9Y148_D = CLBLM_R_X7Y148_SLICE_X9Y148_DO6;
  assign CLBLM_R_X7Y148_SLICE_X9Y148_AMUX = CLBLM_R_X7Y148_SLICE_X9Y148_A5Q;
  assign CLBLM_R_X7Y148_SLICE_X9Y148_CMUX = CLBLM_R_X7Y148_SLICE_X9Y148_C5Q;
  assign CLBLM_R_X7Y148_SLICE_X9Y148_DMUX = CLBLM_R_X7Y148_SLICE_X9Y148_DO6;
  assign CLBLM_R_X7Y149_SLICE_X8Y149_A = CLBLM_R_X7Y149_SLICE_X8Y149_AO6;
  assign CLBLM_R_X7Y149_SLICE_X8Y149_B = CLBLM_R_X7Y149_SLICE_X8Y149_BO6;
  assign CLBLM_R_X7Y149_SLICE_X8Y149_C = CLBLM_R_X7Y149_SLICE_X8Y149_CO6;
  assign CLBLM_R_X7Y149_SLICE_X8Y149_D = CLBLM_R_X7Y149_SLICE_X8Y149_DO6;
  assign CLBLM_R_X7Y149_SLICE_X8Y149_AMUX = CLBLM_R_X7Y149_SLICE_X8Y149_A5Q;
  assign CLBLM_R_X7Y149_SLICE_X9Y149_A = CLBLM_R_X7Y149_SLICE_X9Y149_AO6;
  assign CLBLM_R_X7Y149_SLICE_X9Y149_B = CLBLM_R_X7Y149_SLICE_X9Y149_BO6;
  assign CLBLM_R_X7Y149_SLICE_X9Y149_C = CLBLM_R_X7Y149_SLICE_X9Y149_CO6;
  assign CLBLM_R_X7Y149_SLICE_X9Y149_D = CLBLM_R_X7Y149_SLICE_X9Y149_DO6;
  assign CLBLM_R_X7Y149_SLICE_X9Y149_AMUX = CLBLM_R_X7Y149_SLICE_X9Y149_A5Q;
  assign CLBLM_R_X7Y149_SLICE_X9Y149_BMUX = CLBLM_R_X7Y149_SLICE_X9Y149_B5Q;
  assign CLBLM_R_X7Y149_SLICE_X9Y149_CMUX = CLBLM_R_X7Y149_SLICE_X9Y149_C5Q;
  assign CLBLM_R_X7Y150_SLICE_X8Y150_A = CLBLM_R_X7Y150_SLICE_X8Y150_AO6;
  assign CLBLM_R_X7Y150_SLICE_X8Y150_B = CLBLM_R_X7Y150_SLICE_X8Y150_BO6;
  assign CLBLM_R_X7Y150_SLICE_X8Y150_C = CLBLM_R_X7Y150_SLICE_X8Y150_CO6;
  assign CLBLM_R_X7Y150_SLICE_X8Y150_D = CLBLM_R_X7Y150_SLICE_X8Y150_DO6;
  assign CLBLM_R_X7Y150_SLICE_X8Y150_BMUX = CLBLM_R_X7Y150_SLICE_X8Y150_BO5;
  assign CLBLM_R_X7Y150_SLICE_X9Y150_A = CLBLM_R_X7Y150_SLICE_X9Y150_AO6;
  assign CLBLM_R_X7Y150_SLICE_X9Y150_B = CLBLM_R_X7Y150_SLICE_X9Y150_BO6;
  assign CLBLM_R_X7Y150_SLICE_X9Y150_C = CLBLM_R_X7Y150_SLICE_X9Y150_CO6;
  assign CLBLM_R_X7Y150_SLICE_X9Y150_D = CLBLM_R_X7Y150_SLICE_X9Y150_DO6;
  assign CLBLM_R_X7Y151_SLICE_X8Y151_A = CLBLM_R_X7Y151_SLICE_X8Y151_AO6;
  assign CLBLM_R_X7Y151_SLICE_X8Y151_B = CLBLM_R_X7Y151_SLICE_X8Y151_BO6;
  assign CLBLM_R_X7Y151_SLICE_X8Y151_C = CLBLM_R_X7Y151_SLICE_X8Y151_CO6;
  assign CLBLM_R_X7Y151_SLICE_X8Y151_D = CLBLM_R_X7Y151_SLICE_X8Y151_DO6;
  assign CLBLM_R_X7Y151_SLICE_X8Y151_CMUX = CLBLM_R_X7Y151_SLICE_X8Y151_C5Q;
  assign CLBLM_R_X7Y151_SLICE_X8Y151_DMUX = CLBLM_R_X7Y151_SLICE_X8Y151_D5Q;
  assign CLBLM_R_X7Y151_SLICE_X9Y151_A = CLBLM_R_X7Y151_SLICE_X9Y151_AO6;
  assign CLBLM_R_X7Y151_SLICE_X9Y151_B = CLBLM_R_X7Y151_SLICE_X9Y151_BO6;
  assign CLBLM_R_X7Y151_SLICE_X9Y151_C = CLBLM_R_X7Y151_SLICE_X9Y151_CO6;
  assign CLBLM_R_X7Y151_SLICE_X9Y151_D = CLBLM_R_X7Y151_SLICE_X9Y151_DO6;
  assign CLBLM_R_X7Y151_SLICE_X9Y151_AMUX = CLBLM_R_X7Y151_SLICE_X9Y151_A5Q;
  assign CLBLM_R_X7Y151_SLICE_X9Y151_CMUX = CLBLM_R_X7Y151_SLICE_X9Y151_C5Q;
  assign CLBLM_R_X7Y151_SLICE_X9Y151_DMUX = CLBLM_R_X7Y151_SLICE_X9Y151_D5Q;
  assign CLBLM_R_X7Y152_SLICE_X8Y152_A = CLBLM_R_X7Y152_SLICE_X8Y152_AO6;
  assign CLBLM_R_X7Y152_SLICE_X8Y152_B = CLBLM_R_X7Y152_SLICE_X8Y152_BO6;
  assign CLBLM_R_X7Y152_SLICE_X8Y152_C = CLBLM_R_X7Y152_SLICE_X8Y152_CO6;
  assign CLBLM_R_X7Y152_SLICE_X8Y152_D = CLBLM_R_X7Y152_SLICE_X8Y152_DO6;
  assign CLBLM_R_X7Y152_SLICE_X8Y152_BMUX = CLBLM_R_X7Y152_SLICE_X8Y152_B5Q;
  assign CLBLM_R_X7Y152_SLICE_X8Y152_DMUX = CLBLM_R_X7Y152_SLICE_X8Y152_D5Q;
  assign CLBLM_R_X7Y152_SLICE_X9Y152_A = CLBLM_R_X7Y152_SLICE_X9Y152_AO6;
  assign CLBLM_R_X7Y152_SLICE_X9Y152_B = CLBLM_R_X7Y152_SLICE_X9Y152_BO6;
  assign CLBLM_R_X7Y152_SLICE_X9Y152_C = CLBLM_R_X7Y152_SLICE_X9Y152_CO6;
  assign CLBLM_R_X7Y152_SLICE_X9Y152_D = CLBLM_R_X7Y152_SLICE_X9Y152_DO6;
  assign CLBLM_R_X7Y152_SLICE_X9Y152_BMUX = CLBLM_R_X7Y152_SLICE_X9Y152_B5Q;
  assign CLBLM_R_X7Y152_SLICE_X9Y152_CMUX = CLBLM_R_X7Y152_SLICE_X9Y152_C5Q;
  assign CLBLM_R_X7Y152_SLICE_X9Y152_DMUX = CLBLM_R_X7Y152_SLICE_X9Y152_DO5;
  assign CLBLM_R_X7Y153_SLICE_X8Y153_A = CLBLM_R_X7Y153_SLICE_X8Y153_AO6;
  assign CLBLM_R_X7Y153_SLICE_X8Y153_B = CLBLM_R_X7Y153_SLICE_X8Y153_BO6;
  assign CLBLM_R_X7Y153_SLICE_X8Y153_C = CLBLM_R_X7Y153_SLICE_X8Y153_CO6;
  assign CLBLM_R_X7Y153_SLICE_X8Y153_D = CLBLM_R_X7Y153_SLICE_X8Y153_DO6;
  assign CLBLM_R_X7Y153_SLICE_X8Y153_AMUX = CLBLM_R_X7Y153_SLICE_X8Y153_A5Q;
  assign CLBLM_R_X7Y153_SLICE_X9Y153_A = CLBLM_R_X7Y153_SLICE_X9Y153_AO6;
  assign CLBLM_R_X7Y153_SLICE_X9Y153_B = CLBLM_R_X7Y153_SLICE_X9Y153_BO6;
  assign CLBLM_R_X7Y153_SLICE_X9Y153_C = CLBLM_R_X7Y153_SLICE_X9Y153_CO6;
  assign CLBLM_R_X7Y153_SLICE_X9Y153_D = CLBLM_R_X7Y153_SLICE_X9Y153_DO6;
  assign CLBLM_R_X7Y153_SLICE_X9Y153_AMUX = CLBLM_R_X7Y153_SLICE_X9Y153_A5Q;
  assign CLBLM_R_X7Y153_SLICE_X9Y153_CMUX = CLBLM_R_X7Y153_SLICE_X9Y153_C5Q;
  assign CLBLM_R_X7Y153_SLICE_X9Y153_DMUX = CLBLM_R_X7Y153_SLICE_X9Y153_D5Q;
  assign CLBLM_R_X7Y154_SLICE_X8Y154_A = CLBLM_R_X7Y154_SLICE_X8Y154_AO6;
  assign CLBLM_R_X7Y154_SLICE_X8Y154_B = CLBLM_R_X7Y154_SLICE_X8Y154_BO6;
  assign CLBLM_R_X7Y154_SLICE_X8Y154_C = CLBLM_R_X7Y154_SLICE_X8Y154_CO6;
  assign CLBLM_R_X7Y154_SLICE_X8Y154_D = CLBLM_R_X7Y154_SLICE_X8Y154_DO6;
  assign CLBLM_R_X7Y154_SLICE_X8Y154_CMUX = CLBLM_R_X7Y154_SLICE_X8Y154_CO5;
  assign CLBLM_R_X7Y154_SLICE_X9Y154_A = CLBLM_R_X7Y154_SLICE_X9Y154_AO6;
  assign CLBLM_R_X7Y154_SLICE_X9Y154_B = CLBLM_R_X7Y154_SLICE_X9Y154_BO6;
  assign CLBLM_R_X7Y154_SLICE_X9Y154_C = CLBLM_R_X7Y154_SLICE_X9Y154_CO6;
  assign CLBLM_R_X7Y154_SLICE_X9Y154_D = CLBLM_R_X7Y154_SLICE_X9Y154_DO6;
  assign CLBLM_R_X7Y154_SLICE_X9Y154_CMUX = CLBLM_R_X7Y154_SLICE_X9Y154_CO5;
  assign CLBLM_R_X7Y155_SLICE_X8Y155_A = CLBLM_R_X7Y155_SLICE_X8Y155_AO6;
  assign CLBLM_R_X7Y155_SLICE_X8Y155_B = CLBLM_R_X7Y155_SLICE_X8Y155_BO6;
  assign CLBLM_R_X7Y155_SLICE_X8Y155_C = CLBLM_R_X7Y155_SLICE_X8Y155_CO6;
  assign CLBLM_R_X7Y155_SLICE_X8Y155_D = CLBLM_R_X7Y155_SLICE_X8Y155_DO6;
  assign CLBLM_R_X7Y155_SLICE_X8Y155_AMUX = CLBLM_R_X7Y155_SLICE_X8Y155_A5Q;
  assign CLBLM_R_X7Y155_SLICE_X8Y155_BMUX = CLBLM_R_X7Y155_SLICE_X8Y155_BO5;
  assign CLBLM_R_X7Y155_SLICE_X9Y155_A = CLBLM_R_X7Y155_SLICE_X9Y155_AO6;
  assign CLBLM_R_X7Y155_SLICE_X9Y155_B = CLBLM_R_X7Y155_SLICE_X9Y155_BO6;
  assign CLBLM_R_X7Y155_SLICE_X9Y155_C = CLBLM_R_X7Y155_SLICE_X9Y155_CO6;
  assign CLBLM_R_X7Y155_SLICE_X9Y155_D = CLBLM_R_X7Y155_SLICE_X9Y155_DO6;
  assign CLBLM_R_X11Y144_SLICE_X14Y144_A = CLBLM_R_X11Y144_SLICE_X14Y144_AO6;
  assign CLBLM_R_X11Y144_SLICE_X14Y144_B = CLBLM_R_X11Y144_SLICE_X14Y144_BO6;
  assign CLBLM_R_X11Y144_SLICE_X14Y144_C = CLBLM_R_X11Y144_SLICE_X14Y144_CO6;
  assign CLBLM_R_X11Y144_SLICE_X14Y144_D = CLBLM_R_X11Y144_SLICE_X14Y144_DO6;
  assign CLBLM_R_X11Y144_SLICE_X15Y144_A = CLBLM_R_X11Y144_SLICE_X15Y144_AO6;
  assign CLBLM_R_X11Y144_SLICE_X15Y144_B = CLBLM_R_X11Y144_SLICE_X15Y144_BO6;
  assign CLBLM_R_X11Y144_SLICE_X15Y144_C = CLBLM_R_X11Y144_SLICE_X15Y144_CO6;
  assign CLBLM_R_X11Y144_SLICE_X15Y144_D = CLBLM_R_X11Y144_SLICE_X15Y144_DO6;
  assign CLBLM_R_X11Y145_SLICE_X14Y145_A = CLBLM_R_X11Y145_SLICE_X14Y145_AO6;
  assign CLBLM_R_X11Y145_SLICE_X14Y145_B = CLBLM_R_X11Y145_SLICE_X14Y145_BO6;
  assign CLBLM_R_X11Y145_SLICE_X14Y145_C = CLBLM_R_X11Y145_SLICE_X14Y145_CO6;
  assign CLBLM_R_X11Y145_SLICE_X14Y145_D = CLBLM_R_X11Y145_SLICE_X14Y145_DO6;
  assign CLBLM_R_X11Y145_SLICE_X15Y145_A = CLBLM_R_X11Y145_SLICE_X15Y145_AO6;
  assign CLBLM_R_X11Y145_SLICE_X15Y145_B = CLBLM_R_X11Y145_SLICE_X15Y145_BO6;
  assign CLBLM_R_X11Y145_SLICE_X15Y145_C = CLBLM_R_X11Y145_SLICE_X15Y145_CO6;
  assign CLBLM_R_X11Y145_SLICE_X15Y145_D = CLBLM_R_X11Y145_SLICE_X15Y145_DO6;
  assign CLBLM_R_X11Y145_SLICE_X15Y145_BMUX = CLBLM_R_X11Y145_SLICE_X15Y145_BO6;
  assign CLBLM_R_X11Y146_SLICE_X14Y146_A = CLBLM_R_X11Y146_SLICE_X14Y146_AO6;
  assign CLBLM_R_X11Y146_SLICE_X14Y146_B = CLBLM_R_X11Y146_SLICE_X14Y146_BO6;
  assign CLBLM_R_X11Y146_SLICE_X14Y146_C = CLBLM_R_X11Y146_SLICE_X14Y146_CO6;
  assign CLBLM_R_X11Y146_SLICE_X14Y146_D = CLBLM_R_X11Y146_SLICE_X14Y146_DO6;
  assign CLBLM_R_X11Y146_SLICE_X14Y146_BMUX = CLBLM_R_X11Y146_SLICE_X14Y146_BO5;
  assign CLBLM_R_X11Y146_SLICE_X14Y146_CMUX = CLBLM_R_X11Y146_SLICE_X14Y146_CO5;
  assign CLBLM_R_X11Y146_SLICE_X15Y146_A = CLBLM_R_X11Y146_SLICE_X15Y146_AO6;
  assign CLBLM_R_X11Y146_SLICE_X15Y146_B = CLBLM_R_X11Y146_SLICE_X15Y146_BO6;
  assign CLBLM_R_X11Y146_SLICE_X15Y146_C = CLBLM_R_X11Y146_SLICE_X15Y146_CO6;
  assign CLBLM_R_X11Y146_SLICE_X15Y146_D = CLBLM_R_X11Y146_SLICE_X15Y146_DO6;
  assign CLBLM_R_X11Y146_SLICE_X15Y146_AMUX = CLBLM_R_X11Y146_SLICE_X15Y146_AO5;
  assign CLBLM_R_X11Y146_SLICE_X15Y146_BMUX = CLBLM_R_X11Y146_SLICE_X15Y146_BO5;
  assign CLBLM_R_X11Y147_SLICE_X14Y147_A = CLBLM_R_X11Y147_SLICE_X14Y147_AO6;
  assign CLBLM_R_X11Y147_SLICE_X14Y147_B = CLBLM_R_X11Y147_SLICE_X14Y147_BO6;
  assign CLBLM_R_X11Y147_SLICE_X14Y147_C = CLBLM_R_X11Y147_SLICE_X14Y147_CO6;
  assign CLBLM_R_X11Y147_SLICE_X14Y147_D = CLBLM_R_X11Y147_SLICE_X14Y147_DO6;
  assign CLBLM_R_X11Y147_SLICE_X14Y147_AMUX = CLBLM_R_X11Y147_SLICE_X14Y147_AO5;
  assign CLBLM_R_X11Y147_SLICE_X14Y147_BMUX = CLBLM_R_X11Y147_SLICE_X14Y147_BO5;
  assign CLBLM_R_X11Y147_SLICE_X15Y147_A = CLBLM_R_X11Y147_SLICE_X15Y147_AO6;
  assign CLBLM_R_X11Y147_SLICE_X15Y147_B = CLBLM_R_X11Y147_SLICE_X15Y147_BO6;
  assign CLBLM_R_X11Y147_SLICE_X15Y147_C = CLBLM_R_X11Y147_SLICE_X15Y147_CO6;
  assign CLBLM_R_X11Y147_SLICE_X15Y147_D = CLBLM_R_X11Y147_SLICE_X15Y147_DO6;
  assign CLBLM_R_X11Y148_SLICE_X14Y148_A = CLBLM_R_X11Y148_SLICE_X14Y148_AO6;
  assign CLBLM_R_X11Y148_SLICE_X14Y148_B = CLBLM_R_X11Y148_SLICE_X14Y148_BO6;
  assign CLBLM_R_X11Y148_SLICE_X14Y148_C = CLBLM_R_X11Y148_SLICE_X14Y148_CO6;
  assign CLBLM_R_X11Y148_SLICE_X14Y148_D = CLBLM_R_X11Y148_SLICE_X14Y148_DO6;
  assign CLBLM_R_X11Y148_SLICE_X15Y148_A = CLBLM_R_X11Y148_SLICE_X15Y148_AO6;
  assign CLBLM_R_X11Y148_SLICE_X15Y148_B = CLBLM_R_X11Y148_SLICE_X15Y148_BO6;
  assign CLBLM_R_X11Y148_SLICE_X15Y148_C = CLBLM_R_X11Y148_SLICE_X15Y148_CO6;
  assign CLBLM_R_X11Y148_SLICE_X15Y148_D = CLBLM_R_X11Y148_SLICE_X15Y148_DO6;
  assign CLBLM_R_X11Y148_SLICE_X15Y148_BMUX = CLBLM_R_X11Y148_SLICE_X15Y148_BO6;
  assign CLBLM_R_X11Y148_SLICE_X15Y148_CMUX = CLBLM_R_X11Y148_SLICE_X15Y148_CO6;
  assign CLBLM_R_X11Y149_SLICE_X14Y149_A = CLBLM_R_X11Y149_SLICE_X14Y149_AO6;
  assign CLBLM_R_X11Y149_SLICE_X14Y149_B = CLBLM_R_X11Y149_SLICE_X14Y149_BO6;
  assign CLBLM_R_X11Y149_SLICE_X14Y149_C = CLBLM_R_X11Y149_SLICE_X14Y149_CO6;
  assign CLBLM_R_X11Y149_SLICE_X14Y149_D = CLBLM_R_X11Y149_SLICE_X14Y149_DO6;
  assign CLBLM_R_X11Y149_SLICE_X14Y149_DMUX = CLBLM_R_X11Y149_SLICE_X14Y149_DO6;
  assign CLBLM_R_X11Y149_SLICE_X15Y149_A = CLBLM_R_X11Y149_SLICE_X15Y149_AO6;
  assign CLBLM_R_X11Y149_SLICE_X15Y149_B = CLBLM_R_X11Y149_SLICE_X15Y149_BO6;
  assign CLBLM_R_X11Y149_SLICE_X15Y149_C = CLBLM_R_X11Y149_SLICE_X15Y149_CO6;
  assign CLBLM_R_X11Y149_SLICE_X15Y149_D = CLBLM_R_X11Y149_SLICE_X15Y149_DO6;
  assign CLBLM_R_X11Y150_SLICE_X14Y150_A = CLBLM_R_X11Y150_SLICE_X14Y150_AO6;
  assign CLBLM_R_X11Y150_SLICE_X14Y150_B = CLBLM_R_X11Y150_SLICE_X14Y150_BO6;
  assign CLBLM_R_X11Y150_SLICE_X14Y150_C = CLBLM_R_X11Y150_SLICE_X14Y150_CO6;
  assign CLBLM_R_X11Y150_SLICE_X14Y150_D = CLBLM_R_X11Y150_SLICE_X14Y150_DO6;
  assign CLBLM_R_X11Y150_SLICE_X15Y150_A = CLBLM_R_X11Y150_SLICE_X15Y150_AO6;
  assign CLBLM_R_X11Y150_SLICE_X15Y150_B = CLBLM_R_X11Y150_SLICE_X15Y150_BO6;
  assign CLBLM_R_X11Y150_SLICE_X15Y150_C = CLBLM_R_X11Y150_SLICE_X15Y150_CO6;
  assign CLBLM_R_X11Y150_SLICE_X15Y150_D = CLBLM_R_X11Y150_SLICE_X15Y150_DO6;
  assign CLBLM_R_X11Y151_SLICE_X14Y151_A = CLBLM_R_X11Y151_SLICE_X14Y151_AO6;
  assign CLBLM_R_X11Y151_SLICE_X14Y151_B = CLBLM_R_X11Y151_SLICE_X14Y151_BO6;
  assign CLBLM_R_X11Y151_SLICE_X14Y151_C = CLBLM_R_X11Y151_SLICE_X14Y151_CO6;
  assign CLBLM_R_X11Y151_SLICE_X14Y151_D = CLBLM_R_X11Y151_SLICE_X14Y151_DO6;
  assign CLBLM_R_X11Y151_SLICE_X15Y151_A = CLBLM_R_X11Y151_SLICE_X15Y151_AO6;
  assign CLBLM_R_X11Y151_SLICE_X15Y151_B = CLBLM_R_X11Y151_SLICE_X15Y151_BO6;
  assign CLBLM_R_X11Y151_SLICE_X15Y151_C = CLBLM_R_X11Y151_SLICE_X15Y151_CO6;
  assign CLBLM_R_X11Y151_SLICE_X15Y151_D = CLBLM_R_X11Y151_SLICE_X15Y151_DO6;
  assign CLBLM_R_X11Y151_SLICE_X15Y151_AMUX = CLBLM_R_X11Y151_SLICE_X15Y151_A5Q;
  assign CLBLM_R_X11Y152_SLICE_X14Y152_A = CLBLM_R_X11Y152_SLICE_X14Y152_AO6;
  assign CLBLM_R_X11Y152_SLICE_X14Y152_B = CLBLM_R_X11Y152_SLICE_X14Y152_BO6;
  assign CLBLM_R_X11Y152_SLICE_X14Y152_C = CLBLM_R_X11Y152_SLICE_X14Y152_CO6;
  assign CLBLM_R_X11Y152_SLICE_X14Y152_D = CLBLM_R_X11Y152_SLICE_X14Y152_DO6;
  assign CLBLM_R_X11Y152_SLICE_X15Y152_A = CLBLM_R_X11Y152_SLICE_X15Y152_AO6;
  assign CLBLM_R_X11Y152_SLICE_X15Y152_B = CLBLM_R_X11Y152_SLICE_X15Y152_BO6;
  assign CLBLM_R_X11Y152_SLICE_X15Y152_C = CLBLM_R_X11Y152_SLICE_X15Y152_CO6;
  assign CLBLM_R_X11Y152_SLICE_X15Y152_D = CLBLM_R_X11Y152_SLICE_X15Y152_DO6;
  assign CLBLM_R_X11Y152_SLICE_X15Y152_AMUX = CLBLM_R_X11Y152_SLICE_X15Y152_A5Q;
  assign CLBLM_R_X11Y152_SLICE_X15Y152_BMUX = CLBLM_R_X11Y152_SLICE_X15Y152_B5Q;
  assign CLBLM_R_X11Y153_SLICE_X14Y153_A = CLBLM_R_X11Y153_SLICE_X14Y153_AO6;
  assign CLBLM_R_X11Y153_SLICE_X14Y153_B = CLBLM_R_X11Y153_SLICE_X14Y153_BO6;
  assign CLBLM_R_X11Y153_SLICE_X14Y153_C = CLBLM_R_X11Y153_SLICE_X14Y153_CO6;
  assign CLBLM_R_X11Y153_SLICE_X14Y153_D = CLBLM_R_X11Y153_SLICE_X14Y153_DO6;
  assign CLBLM_R_X11Y153_SLICE_X14Y153_AMUX = CLBLM_R_X11Y153_SLICE_X14Y153_A5Q;
  assign CLBLM_R_X11Y153_SLICE_X14Y153_CMUX = CLBLM_R_X11Y153_SLICE_X14Y153_CO6;
  assign CLBLM_R_X11Y153_SLICE_X14Y153_DMUX = CLBLM_R_X11Y153_SLICE_X14Y153_DO6;
  assign CLBLM_R_X11Y153_SLICE_X15Y153_A = CLBLM_R_X11Y153_SLICE_X15Y153_AO6;
  assign CLBLM_R_X11Y153_SLICE_X15Y153_B = CLBLM_R_X11Y153_SLICE_X15Y153_BO6;
  assign CLBLM_R_X11Y153_SLICE_X15Y153_C = CLBLM_R_X11Y153_SLICE_X15Y153_CO6;
  assign CLBLM_R_X11Y153_SLICE_X15Y153_D = CLBLM_R_X11Y153_SLICE_X15Y153_DO6;
  assign CLBLM_R_X11Y153_SLICE_X15Y153_BMUX = CLBLM_R_X11Y153_SLICE_X15Y153_BO5;
  assign CLBLM_R_X13Y146_SLICE_X18Y146_A = CLBLM_R_X13Y146_SLICE_X18Y146_AO6;
  assign CLBLM_R_X13Y146_SLICE_X18Y146_B = CLBLM_R_X13Y146_SLICE_X18Y146_BO6;
  assign CLBLM_R_X13Y146_SLICE_X18Y146_C = CLBLM_R_X13Y146_SLICE_X18Y146_CO6;
  assign CLBLM_R_X13Y146_SLICE_X18Y146_D = CLBLM_R_X13Y146_SLICE_X18Y146_DO6;
  assign CLBLM_R_X13Y146_SLICE_X18Y146_AMUX = CLBLM_R_X13Y146_SLICE_X18Y146_AO5;
  assign CLBLM_R_X13Y146_SLICE_X19Y146_A = CLBLM_R_X13Y146_SLICE_X19Y146_AO6;
  assign CLBLM_R_X13Y146_SLICE_X19Y146_B = CLBLM_R_X13Y146_SLICE_X19Y146_BO6;
  assign CLBLM_R_X13Y146_SLICE_X19Y146_C = CLBLM_R_X13Y146_SLICE_X19Y146_CO6;
  assign CLBLM_R_X13Y146_SLICE_X19Y146_D = CLBLM_R_X13Y146_SLICE_X19Y146_DO6;
  assign CLBLM_R_X13Y149_SLICE_X18Y149_A = CLBLM_R_X13Y149_SLICE_X18Y149_AO6;
  assign CLBLM_R_X13Y149_SLICE_X18Y149_B = CLBLM_R_X13Y149_SLICE_X18Y149_BO6;
  assign CLBLM_R_X13Y149_SLICE_X18Y149_C = CLBLM_R_X13Y149_SLICE_X18Y149_CO6;
  assign CLBLM_R_X13Y149_SLICE_X18Y149_D = CLBLM_R_X13Y149_SLICE_X18Y149_DO6;
  assign CLBLM_R_X13Y149_SLICE_X19Y149_A = CLBLM_R_X13Y149_SLICE_X19Y149_AO6;
  assign CLBLM_R_X13Y149_SLICE_X19Y149_B = CLBLM_R_X13Y149_SLICE_X19Y149_BO6;
  assign CLBLM_R_X13Y149_SLICE_X19Y149_C = CLBLM_R_X13Y149_SLICE_X19Y149_CO6;
  assign CLBLM_R_X13Y149_SLICE_X19Y149_D = CLBLM_R_X13Y149_SLICE_X19Y149_DO6;
  assign CLBLM_R_X103Y178_SLICE_X162Y178_A = CLBLM_R_X103Y178_SLICE_X162Y178_AO6;
  assign CLBLM_R_X103Y178_SLICE_X162Y178_B = CLBLM_R_X103Y178_SLICE_X162Y178_BO6;
  assign CLBLM_R_X103Y178_SLICE_X162Y178_C = CLBLM_R_X103Y178_SLICE_X162Y178_CO6;
  assign CLBLM_R_X103Y178_SLICE_X162Y178_D = CLBLM_R_X103Y178_SLICE_X162Y178_DO6;
  assign CLBLM_R_X103Y178_SLICE_X163Y178_A = CLBLM_R_X103Y178_SLICE_X163Y178_AO6;
  assign CLBLM_R_X103Y178_SLICE_X163Y178_B = CLBLM_R_X103Y178_SLICE_X163Y178_BO6;
  assign CLBLM_R_X103Y178_SLICE_X163Y178_C = CLBLM_R_X103Y178_SLICE_X163Y178_CO6;
  assign CLBLM_R_X103Y178_SLICE_X163Y178_D = CLBLM_R_X103Y178_SLICE_X163Y178_DO6;
  assign LIOI3_X0Y51_ILOGIC_X0Y52_O = LIOB33_X0Y51_IOB_X0Y52_I;
  assign LIOI3_X0Y51_ILOGIC_X0Y51_O = LIOB33_X0Y51_IOB_X0Y51_I;
  assign LIOI3_X0Y53_ILOGIC_X0Y54_O = LIOB33_X0Y53_IOB_X0Y54_I;
  assign LIOI3_X0Y53_ILOGIC_X0Y53_O = LIOB33_X0Y53_IOB_X0Y53_I;
  assign LIOI3_X0Y55_ILOGIC_X0Y56_O = LIOB33_X0Y55_IOB_X0Y56_I;
  assign LIOI3_X0Y55_ILOGIC_X0Y55_O = LIOB33_X0Y55_IOB_X0Y55_I;
  assign LIOI3_X0Y59_ILOGIC_X0Y60_O = LIOB33_X0Y59_IOB_X0Y60_I;
  assign LIOI3_X0Y59_ILOGIC_X0Y59_O = LIOB33_X0Y59_IOB_X0Y59_I;
  assign LIOI3_X0Y61_ILOGIC_X0Y62_O = LIOB33_X0Y61_IOB_X0Y62_I;
  assign LIOI3_X0Y61_ILOGIC_X0Y61_O = LIOB33_X0Y61_IOB_X0Y61_I;
  assign LIOI3_X0Y65_OLOGIC_X0Y66_OQ = CLBLL_L_X4Y151_SLICE_X4Y151_CQ;
  assign LIOI3_X0Y65_OLOGIC_X0Y66_TQ = 1'b1;
  assign LIOI3_X0Y65_OLOGIC_X0Y65_OQ = CLBLM_R_X7Y141_SLICE_X8Y141_BO6;
  assign LIOI3_X0Y65_OLOGIC_X0Y65_TQ = 1'b1;
  assign LIOI3_X0Y77_ILOGIC_X0Y78_O = LIOB33_X0Y77_IOB_X0Y78_I;
  assign LIOI3_X0Y101_OLOGIC_X0Y102_OQ = CLBLM_R_X5Y141_SLICE_X6Y141_DQ;
  assign LIOI3_X0Y101_OLOGIC_X0Y102_TQ = 1'b1;
  assign LIOI3_X0Y101_OLOGIC_X0Y101_OQ = CLBLM_L_X8Y145_SLICE_X11Y145_C5Q;
  assign LIOI3_X0Y101_OLOGIC_X0Y101_TQ = 1'b1;
  assign LIOI3_X0Y103_OLOGIC_X0Y104_OQ = CLBLM_R_X3Y145_SLICE_X2Y145_C5Q;
  assign LIOI3_X0Y103_OLOGIC_X0Y104_TQ = 1'b1;
  assign LIOI3_X0Y103_OLOGIC_X0Y103_OQ = CLBLM_R_X5Y145_SLICE_X7Y145_BQ;
  assign LIOI3_X0Y103_OLOGIC_X0Y103_TQ = 1'b1;
  assign LIOI3_X0Y105_OLOGIC_X0Y106_OQ = CLBLM_R_X3Y146_SLICE_X3Y146_BQ;
  assign LIOI3_X0Y105_OLOGIC_X0Y106_TQ = 1'b1;
  assign LIOI3_X0Y105_OLOGIC_X0Y105_OQ = CLBLL_L_X4Y150_SLICE_X4Y150_C5Q;
  assign LIOI3_X0Y105_OLOGIC_X0Y105_TQ = 1'b1;
  assign LIOI3_X0Y109_OLOGIC_X0Y110_OQ = CLBLM_R_X5Y145_SLICE_X7Y145_AQ;
  assign LIOI3_X0Y109_OLOGIC_X0Y110_TQ = 1'b1;
  assign LIOI3_X0Y109_OLOGIC_X0Y109_OQ = CLBLM_R_X5Y141_SLICE_X6Y141_BQ;
  assign LIOI3_X0Y109_OLOGIC_X0Y109_TQ = 1'b1;
  assign LIOI3_X0Y111_OLOGIC_X0Y112_OQ = CLBLL_L_X4Y146_SLICE_X4Y146_C5Q;
  assign LIOI3_X0Y111_OLOGIC_X0Y112_TQ = 1'b1;
  assign LIOI3_X0Y111_OLOGIC_X0Y111_OQ = CLBLM_R_X3Y145_SLICE_X2Y145_B5Q;
  assign LIOI3_X0Y111_OLOGIC_X0Y111_TQ = 1'b1;
  assign LIOI3_X0Y115_OLOGIC_X0Y116_OQ = CLBLM_R_X7Y143_SLICE_X9Y143_B5Q;
  assign LIOI3_X0Y115_OLOGIC_X0Y116_TQ = 1'b1;
  assign LIOI3_X0Y115_OLOGIC_X0Y115_OQ = CLBLM_R_X5Y147_SLICE_X6Y147_C5Q;
  assign LIOI3_X0Y115_OLOGIC_X0Y115_TQ = 1'b1;
  assign LIOI3_X0Y117_OLOGIC_X0Y118_OQ = CLBLM_R_X7Y142_SLICE_X9Y142_BQ;
  assign LIOI3_X0Y117_OLOGIC_X0Y118_TQ = 1'b1;
  assign LIOI3_X0Y117_OLOGIC_X0Y117_OQ = CLBLM_L_X10Y143_SLICE_X13Y143_C5Q;
  assign LIOI3_X0Y117_OLOGIC_X0Y117_TQ = 1'b1;
  assign LIOI3_X0Y121_OLOGIC_X0Y122_OQ = CLBLL_L_X4Y144_SLICE_X5Y144_CQ;
  assign LIOI3_X0Y121_OLOGIC_X0Y122_TQ = 1'b1;
  assign LIOI3_X0Y121_OLOGIC_X0Y121_OQ = CLBLM_L_X8Y147_SLICE_X10Y147_C5Q;
  assign LIOI3_X0Y121_OLOGIC_X0Y121_TQ = 1'b1;
  assign LIOI3_X0Y123_OLOGIC_X0Y124_OQ = CLBLL_L_X4Y151_SLICE_X4Y151_CQ;
  assign LIOI3_X0Y123_OLOGIC_X0Y124_TQ = 1'b1;
  assign LIOI3_X0Y123_OLOGIC_X0Y123_OQ = CLBLL_L_X2Y146_SLICE_X0Y146_CQ;
  assign LIOI3_X0Y123_OLOGIC_X0Y123_TQ = 1'b1;
  assign LIOI3_X0Y125_OLOGIC_X0Y126_OQ = CLBLL_L_X4Y147_SLICE_X5Y147_CQ;
  assign LIOI3_X0Y125_OLOGIC_X0Y126_TQ = 1'b1;
  assign LIOI3_X0Y125_OLOGIC_X0Y125_OQ = CLBLL_L_X4Y151_SLICE_X4Y151_BQ;
  assign LIOI3_X0Y125_OLOGIC_X0Y125_TQ = 1'b1;
  assign LIOI3_X0Y127_OLOGIC_X0Y128_OQ = CLBLM_L_X10Y145_SLICE_X12Y145_AQ;
  assign LIOI3_X0Y127_OLOGIC_X0Y128_TQ = 1'b1;
  assign LIOI3_X0Y127_OLOGIC_X0Y127_OQ = CLBLM_R_X7Y152_SLICE_X8Y152_D5Q;
  assign LIOI3_X0Y127_OLOGIC_X0Y127_TQ = 1'b1;
  assign LIOI3_X0Y129_OLOGIC_X0Y130_OQ = CLBLL_L_X2Y145_SLICE_X0Y145_BQ;
  assign LIOI3_X0Y129_OLOGIC_X0Y130_TQ = 1'b1;
  assign LIOI3_X0Y129_OLOGIC_X0Y129_OQ = CLBLL_L_X2Y146_SLICE_X0Y146_CQ;
  assign LIOI3_X0Y129_OLOGIC_X0Y129_TQ = 1'b1;
  assign LIOI3_X0Y133_OLOGIC_X0Y134_OQ = CLBLL_L_X2Y145_SLICE_X0Y145_BQ;
  assign LIOI3_X0Y133_OLOGIC_X0Y134_TQ = 1'b1;
  assign LIOI3_X0Y133_OLOGIC_X0Y133_OQ = CLBLL_L_X4Y140_SLICE_X4Y140_BO5;
  assign LIOI3_X0Y133_OLOGIC_X0Y133_TQ = 1'b1;
  assign LIOI3_X0Y135_OLOGIC_X0Y136_OQ = CLBLM_L_X10Y153_SLICE_X13Y153_CQ;
  assign LIOI3_X0Y135_OLOGIC_X0Y136_TQ = 1'b1;
  assign LIOI3_X0Y135_OLOGIC_X0Y135_OQ = CLBLL_L_X2Y145_SLICE_X0Y145_BQ;
  assign LIOI3_X0Y135_OLOGIC_X0Y135_TQ = 1'b1;
  assign LIOI3_X0Y139_OLOGIC_X0Y140_OQ = CLBLL_L_X4Y145_SLICE_X4Y145_C5Q;
  assign LIOI3_X0Y139_OLOGIC_X0Y140_TQ = 1'b1;
  assign LIOI3_X0Y139_OLOGIC_X0Y139_OQ = CLBLM_R_X3Y147_SLICE_X2Y147_DQ;
  assign LIOI3_X0Y139_OLOGIC_X0Y139_TQ = 1'b1;
  assign LIOI3_X0Y141_OLOGIC_X0Y142_OQ = CLBLL_L_X2Y146_SLICE_X0Y146_CQ;
  assign LIOI3_X0Y141_OLOGIC_X0Y142_TQ = 1'b1;
  assign LIOI3_X0Y141_OLOGIC_X0Y141_OQ = CLBLL_L_X4Y145_SLICE_X5Y145_CQ;
  assign LIOI3_X0Y141_OLOGIC_X0Y141_TQ = 1'b1;
  assign LIOI3_X0Y145_OLOGIC_X0Y146_OQ = CLBLM_R_X3Y143_SLICE_X3Y143_DO6;
  assign LIOI3_X0Y145_OLOGIC_X0Y146_TQ = 1'b1;
  assign LIOI3_X0Y145_OLOGIC_X0Y145_OQ = CLBLM_R_X3Y148_SLICE_X3Y148_DO6;
  assign LIOI3_X0Y145_OLOGIC_X0Y145_TQ = 1'b1;
  assign LIOI3_X0Y147_OLOGIC_X0Y148_OQ = CLBLL_L_X2Y147_SLICE_X1Y147_AO6;
  assign LIOI3_X0Y147_OLOGIC_X0Y148_TQ = 1'b1;
  assign LIOI3_X0Y147_OLOGIC_X0Y147_OQ = CLBLM_R_X5Y141_SLICE_X6Y141_CO5;
  assign LIOI3_X0Y147_OLOGIC_X0Y147_TQ = 1'b1;
  assign LIOI3_X0Y151_OLOGIC_X0Y152_OQ = CLBLL_L_X4Y147_SLICE_X5Y147_C5Q;
  assign LIOI3_X0Y151_OLOGIC_X0Y152_TQ = 1'b1;
  assign LIOI3_X0Y151_OLOGIC_X0Y151_OQ = CLBLL_L_X2Y146_SLICE_X0Y146_CQ;
  assign LIOI3_X0Y151_OLOGIC_X0Y151_TQ = 1'b1;
  assign LIOI3_X0Y153_OLOGIC_X0Y154_OQ = CLBLM_R_X7Y153_SLICE_X9Y153_DQ;
  assign LIOI3_X0Y153_OLOGIC_X0Y154_TQ = 1'b1;
  assign LIOI3_X0Y153_OLOGIC_X0Y153_OQ = CLBLM_L_X8Y153_SLICE_X10Y153_A5Q;
  assign LIOI3_X0Y153_OLOGIC_X0Y153_TQ = 1'b1;
  assign LIOI3_X0Y155_OLOGIC_X0Y156_OQ = CLBLM_R_X3Y152_SLICE_X3Y152_CQ;
  assign LIOI3_X0Y155_OLOGIC_X0Y156_TQ = 1'b1;
  assign LIOI3_X0Y155_OLOGIC_X0Y155_OQ = CLBLM_R_X5Y154_SLICE_X7Y154_AQ;
  assign LIOI3_X0Y155_OLOGIC_X0Y155_TQ = 1'b1;
  assign LIOI3_X0Y159_OLOGIC_X0Y160_OQ = CLBLL_L_X2Y148_SLICE_X0Y148_AQ;
  assign LIOI3_X0Y159_OLOGIC_X0Y160_TQ = 1'b1;
  assign LIOI3_X0Y159_OLOGIC_X0Y159_OQ = CLBLL_L_X2Y146_SLICE_X0Y146_CQ;
  assign LIOI3_X0Y159_OLOGIC_X0Y159_TQ = 1'b1;
  assign LIOI3_X0Y161_OLOGIC_X0Y162_OQ = CLBLM_L_X10Y144_SLICE_X12Y144_BO6;
  assign LIOI3_X0Y161_OLOGIC_X0Y162_TQ = 1'b1;
  assign LIOI3_X0Y161_OLOGIC_X0Y161_OQ = CLBLM_R_X5Y152_SLICE_X7Y152_DQ;
  assign LIOI3_X0Y161_OLOGIC_X0Y161_TQ = 1'b1;
  assign LIOI3_X0Y165_OLOGIC_X0Y166_OQ = RIOB33_SING_X105Y100_IOB_X1Y100_I;
  assign LIOI3_X0Y165_OLOGIC_X0Y166_TQ = 1'b1;
  assign LIOI3_X0Y165_OLOGIC_X0Y165_OQ = LIOB33_X0Y57_IOB_X0Y57_I;
  assign LIOI3_X0Y165_OLOGIC_X0Y165_TQ = 1'b1;
  assign LIOI3_X0Y167_OLOGIC_X0Y168_OQ = RIOB33_X105Y101_IOB_X1Y101_I;
  assign LIOI3_X0Y167_OLOGIC_X0Y168_TQ = 1'b1;
  assign LIOI3_X0Y167_OLOGIC_X0Y167_OQ = RIOB33_X105Y105_IOB_X1Y106_I;
  assign LIOI3_X0Y167_OLOGIC_X0Y167_TQ = 1'b1;
  assign LIOI3_X0Y171_OLOGIC_X0Y172_OQ = RIOB33_X105Y119_IOB_X1Y120_I;
  assign LIOI3_X0Y171_OLOGIC_X0Y172_TQ = 1'b1;
  assign LIOI3_X0Y171_OLOGIC_X0Y171_OQ = RIOB33_X105Y119_IOB_X1Y119_I;
  assign LIOI3_X0Y171_OLOGIC_X0Y171_TQ = 1'b1;
  assign LIOI3_X0Y173_OLOGIC_X0Y174_OQ = RIOB33_X105Y121_IOB_X1Y122_I;
  assign LIOI3_X0Y173_OLOGIC_X0Y174_TQ = 1'b1;
  assign LIOI3_X0Y173_OLOGIC_X0Y173_OQ = RIOB33_X105Y121_IOB_X1Y121_I;
  assign LIOI3_X0Y173_OLOGIC_X0Y173_TQ = 1'b1;
  assign LIOI3_X0Y175_OLOGIC_X0Y176_OQ = RIOB33_X105Y115_IOB_X1Y116_I;
  assign LIOI3_X0Y175_OLOGIC_X0Y176_TQ = 1'b1;
  assign LIOI3_X0Y175_OLOGIC_X0Y175_OQ = RIOB33_X105Y123_IOB_X1Y123_I;
  assign LIOI3_X0Y175_OLOGIC_X0Y175_TQ = 1'b1;
  assign LIOI3_X0Y177_OLOGIC_X0Y178_OQ = RIOB33_X105Y125_IOB_X1Y125_I;
  assign LIOI3_X0Y177_OLOGIC_X0Y178_TQ = 1'b1;
  assign LIOI3_X0Y177_OLOGIC_X0Y177_OQ = RIOB33_X105Y123_IOB_X1Y124_I;
  assign LIOI3_X0Y177_OLOGIC_X0Y177_TQ = 1'b1;
  assign LIOI3_X0Y179_OLOGIC_X0Y180_OQ = RIOB33_X105Y127_IOB_X1Y127_I;
  assign LIOI3_X0Y179_OLOGIC_X0Y180_TQ = 1'b1;
  assign LIOI3_X0Y179_OLOGIC_X0Y179_OQ = RIOB33_X105Y125_IOB_X1Y126_I;
  assign LIOI3_X0Y179_OLOGIC_X0Y179_TQ = 1'b1;
  assign LIOI3_X0Y183_OLOGIC_X0Y184_OQ = RIOB33_X105Y131_IOB_X1Y132_I;
  assign LIOI3_X0Y183_OLOGIC_X0Y184_TQ = 1'b1;
  assign LIOI3_X0Y183_OLOGIC_X0Y183_OQ = RIOB33_X105Y129_IOB_X1Y130_I;
  assign LIOI3_X0Y183_OLOGIC_X0Y183_TQ = 1'b1;
  assign LIOI3_X0Y185_OLOGIC_X0Y186_OQ = RIOB33_X105Y119_IOB_X1Y120_I;
  assign LIOI3_X0Y185_OLOGIC_X0Y186_TQ = 1'b1;
  assign LIOI3_X0Y185_OLOGIC_X0Y185_OQ = RIOB33_X105Y133_IOB_X1Y133_I;
  assign LIOI3_X0Y185_OLOGIC_X0Y185_TQ = 1'b1;
  assign LIOI3_X0Y189_OLOGIC_X0Y190_OQ = CLBLM_L_X10Y154_SLICE_X12Y154_CO5;
  assign LIOI3_X0Y189_OLOGIC_X0Y190_TQ = 1'b1;
  assign LIOI3_X0Y189_OLOGIC_X0Y189_OQ = CLBLM_L_X8Y147_SLICE_X10Y147_BQ;
  assign LIOI3_X0Y189_OLOGIC_X0Y189_TQ = 1'b1;
  assign LIOI3_X0Y191_OLOGIC_X0Y192_OQ = CLBLL_L_X4Y153_SLICE_X4Y153_DO5;
  assign LIOI3_X0Y191_OLOGIC_X0Y192_TQ = 1'b1;
  assign LIOI3_X0Y191_OLOGIC_X0Y191_OQ = CLBLL_L_X2Y148_SLICE_X1Y148_CO6;
  assign LIOI3_X0Y191_OLOGIC_X0Y191_TQ = 1'b1;
  assign LIOI3_X0Y195_OLOGIC_X0Y196_OQ = CLBLM_R_X3Y148_SLICE_X3Y148_DO5;
  assign LIOI3_X0Y195_OLOGIC_X0Y196_TQ = 1'b1;
  assign LIOI3_X0Y195_OLOGIC_X0Y195_OQ = CLBLM_R_X3Y151_SLICE_X2Y151_AO5;
  assign LIOI3_X0Y195_OLOGIC_X0Y195_TQ = 1'b1;
  assign LIOI3_X0Y197_OLOGIC_X0Y198_OQ = 1'b1;
  assign LIOI3_X0Y197_OLOGIC_X0Y198_TQ = 1'b1;
  assign LIOI3_X0Y197_OLOGIC_X0Y197_OQ = CLBLL_L_X4Y153_SLICE_X4Y153_CO5;
  assign LIOI3_X0Y197_OLOGIC_X0Y197_TQ = 1'b1;
  assign LIOI3_SING_X0Y50_ILOGIC_X0Y50_O = LIOB33_SING_X0Y50_IOB_X0Y50_I;
  assign LIOI3_SING_X0Y100_OLOGIC_X0Y100_OQ = CLBLM_R_X3Y148_SLICE_X2Y148_B5Q;
  assign LIOI3_SING_X0Y100_OLOGIC_X0Y100_TQ = 1'b1;
  assign LIOI3_SING_X0Y149_OLOGIC_X0Y149_OQ = RIOB33_X105Y115_IOB_X1Y115_I;
  assign LIOI3_SING_X0Y149_OLOGIC_X0Y149_TQ = 1'b1;
  assign LIOI3_SING_X0Y150_OLOGIC_X0Y150_OQ = CLBLM_R_X3Y144_SLICE_X2Y144_AO5;
  assign LIOI3_SING_X0Y150_OLOGIC_X0Y150_TQ = 1'b1;
  assign LIOI3_SING_X0Y199_OLOGIC_X0Y199_OQ = 1'b1;
  assign LIOI3_SING_X0Y199_OLOGIC_X0Y199_TQ = 1'b1;
  assign LIOI3_TBYTESRC_X0Y57_ILOGIC_X0Y58_O = LIOB33_X0Y57_IOB_X0Y58_I;
  assign LIOI3_TBYTESRC_X0Y57_ILOGIC_X0Y57_O = LIOB33_X0Y57_IOB_X0Y57_I;
  assign LIOI3_TBYTESRC_X0Y107_OLOGIC_X0Y108_OQ = CLBLL_L_X4Y143_SLICE_X4Y143_DQ;
  assign LIOI3_TBYTESRC_X0Y107_OLOGIC_X0Y108_TQ = 1'b1;
  assign LIOI3_TBYTESRC_X0Y107_OLOGIC_X0Y107_OQ = CLBLM_R_X7Y146_SLICE_X8Y146_DQ;
  assign LIOI3_TBYTESRC_X0Y107_OLOGIC_X0Y107_TQ = 1'b1;
  assign LIOI3_TBYTESRC_X0Y119_OLOGIC_X0Y120_OQ = CLBLL_L_X4Y147_SLICE_X4Y147_AQ;
  assign LIOI3_TBYTESRC_X0Y119_OLOGIC_X0Y120_TQ = 1'b1;
  assign LIOI3_TBYTESRC_X0Y119_OLOGIC_X0Y119_OQ = CLBLL_L_X2Y146_SLICE_X0Y146_CQ;
  assign LIOI3_TBYTESRC_X0Y119_OLOGIC_X0Y119_TQ = 1'b1;
  assign LIOI3_TBYTESRC_X0Y131_OLOGIC_X0Y132_OQ = CLBLM_R_X3Y143_SLICE_X2Y143_BO5;
  assign LIOI3_TBYTESRC_X0Y131_OLOGIC_X0Y132_TQ = 1'b1;
  assign LIOI3_TBYTESRC_X0Y131_OLOGIC_X0Y131_OQ = CLBLL_L_X2Y75_SLICE_X0Y75_AO6;
  assign LIOI3_TBYTESRC_X0Y131_OLOGIC_X0Y131_TQ = 1'b1;
  assign LIOI3_TBYTESRC_X0Y143_OLOGIC_X0Y144_OQ = CLBLM_R_X5Y147_SLICE_X7Y147_DO6;
  assign LIOI3_TBYTESRC_X0Y143_OLOGIC_X0Y144_TQ = 1'b1;
  assign LIOI3_TBYTESRC_X0Y143_OLOGIC_X0Y143_OQ = CLBLM_R_X3Y151_SLICE_X2Y151_BO5;
  assign LIOI3_TBYTESRC_X0Y143_OLOGIC_X0Y143_TQ = 1'b1;
  assign LIOI3_TBYTESRC_X0Y157_OLOGIC_X0Y158_OQ = RIOB33_X105Y133_IOB_X1Y134_I;
  assign LIOI3_TBYTESRC_X0Y157_OLOGIC_X0Y158_TQ = 1'b1;
  assign LIOI3_TBYTESRC_X0Y157_OLOGIC_X0Y157_OQ = CLBLM_R_X3Y152_SLICE_X3Y152_BQ;
  assign LIOI3_TBYTESRC_X0Y157_OLOGIC_X0Y157_TQ = 1'b1;
  assign LIOI3_TBYTESRC_X0Y169_OLOGIC_X0Y170_OQ = RIOB33_X105Y117_IOB_X1Y118_I;
  assign LIOI3_TBYTESRC_X0Y169_OLOGIC_X0Y170_TQ = 1'b1;
  assign LIOI3_TBYTESRC_X0Y169_OLOGIC_X0Y169_OQ = RIOB33_X105Y117_IOB_X1Y117_I;
  assign LIOI3_TBYTESRC_X0Y169_OLOGIC_X0Y169_TQ = 1'b1;
  assign LIOI3_TBYTESRC_X0Y181_OLOGIC_X0Y182_OQ = RIOB33_X105Y129_IOB_X1Y129_I;
  assign LIOI3_TBYTESRC_X0Y181_OLOGIC_X0Y182_TQ = 1'b1;
  assign LIOI3_TBYTESRC_X0Y181_OLOGIC_X0Y181_OQ = RIOB33_X105Y127_IOB_X1Y128_I;
  assign LIOI3_TBYTESRC_X0Y181_OLOGIC_X0Y181_TQ = 1'b1;
  assign LIOI3_TBYTESRC_X0Y193_OLOGIC_X0Y194_OQ = RIOB33_X105Y103_IOB_X1Y103_I;
  assign LIOI3_TBYTESRC_X0Y193_OLOGIC_X0Y194_TQ = 1'b1;
  assign LIOI3_TBYTESRC_X0Y193_OLOGIC_X0Y193_OQ = CLBLL_L_X2Y166_SLICE_X0Y166_AO6;
  assign LIOI3_TBYTESRC_X0Y193_OLOGIC_X0Y193_TQ = 1'b1;
  assign LIOI3_TBYTETERM_X0Y63_ILOGIC_X0Y63_O = LIOB33_X0Y63_IOB_X0Y63_I;
  assign LIOI3_TBYTETERM_X0Y63_OLOGIC_X0Y64_OQ = CLBLM_R_X7Y141_SLICE_X8Y141_AO5;
  assign LIOI3_TBYTETERM_X0Y63_OLOGIC_X0Y64_TQ = 1'b1;
  assign LIOI3_TBYTETERM_X0Y113_OLOGIC_X0Y114_OQ = CLBLM_L_X8Y142_SLICE_X10Y142_A5Q;
  assign LIOI3_TBYTETERM_X0Y113_OLOGIC_X0Y114_TQ = 1'b1;
  assign LIOI3_TBYTETERM_X0Y113_OLOGIC_X0Y113_OQ = CLBLM_R_X3Y147_SLICE_X3Y147_C5Q;
  assign LIOI3_TBYTETERM_X0Y113_OLOGIC_X0Y113_TQ = 1'b1;
  assign LIOI3_TBYTETERM_X0Y137_OLOGIC_X0Y138_OQ = CLBLM_R_X3Y148_SLICE_X2Y148_A5Q;
  assign LIOI3_TBYTETERM_X0Y137_OLOGIC_X0Y138_TQ = 1'b1;
  assign LIOI3_TBYTETERM_X0Y137_OLOGIC_X0Y137_OQ = CLBLM_R_X5Y153_SLICE_X6Y153_B5Q;
  assign LIOI3_TBYTETERM_X0Y137_OLOGIC_X0Y137_TQ = 1'b1;
  assign LIOI3_TBYTETERM_X0Y163_OLOGIC_X0Y164_OQ = RIOB33_X105Y101_IOB_X1Y102_I;
  assign LIOI3_TBYTETERM_X0Y163_OLOGIC_X0Y164_TQ = 1'b1;
  assign LIOI3_TBYTETERM_X0Y163_OLOGIC_X0Y163_OQ = CLBLM_R_X5Y152_SLICE_X7Y152_DO6;
  assign LIOI3_TBYTETERM_X0Y163_OLOGIC_X0Y163_TQ = 1'b1;
  assign LIOI3_TBYTETERM_X0Y187_OLOGIC_X0Y188_OQ = CLBLM_R_X5Y147_SLICE_X6Y147_AQ;
  assign LIOI3_TBYTETERM_X0Y187_OLOGIC_X0Y188_TQ = 1'b1;
  assign LIOI3_TBYTETERM_X0Y187_OLOGIC_X0Y187_OQ = CLBLM_L_X8Y145_SLICE_X11Y145_DQ;
  assign LIOI3_TBYTETERM_X0Y187_OLOGIC_X0Y187_TQ = 1'b1;
  assign RIOI3_X105Y101_ILOGIC_X1Y102_O = RIOB33_X105Y101_IOB_X1Y102_I;
  assign RIOI3_X105Y101_ILOGIC_X1Y101_O = RIOB33_X105Y101_IOB_X1Y101_I;
  assign RIOI3_X105Y103_ILOGIC_X1Y104_O = RIOB33_X105Y103_IOB_X1Y104_I;
  assign RIOI3_X105Y103_ILOGIC_X1Y103_O = RIOB33_X105Y103_IOB_X1Y103_I;
  assign RIOI3_X105Y105_ILOGIC_X1Y106_O = RIOB33_X105Y105_IOB_X1Y106_I;
  assign RIOI3_X105Y105_ILOGIC_X1Y105_O = RIOB33_X105Y105_IOB_X1Y105_I;
  assign RIOI3_X105Y109_ILOGIC_X1Y110_O = RIOB33_X105Y109_IOB_X1Y110_I;
  assign RIOI3_X105Y109_ILOGIC_X1Y109_O = RIOB33_X105Y109_IOB_X1Y109_I;
  assign RIOI3_X105Y111_ILOGIC_X1Y112_O = RIOB33_X105Y111_IOB_X1Y112_I;
  assign RIOI3_X105Y111_ILOGIC_X1Y111_O = RIOB33_X105Y111_IOB_X1Y111_I;
  assign RIOI3_X105Y115_ILOGIC_X1Y116_O = RIOB33_X105Y115_IOB_X1Y116_I;
  assign RIOI3_X105Y115_ILOGIC_X1Y115_O = RIOB33_X105Y115_IOB_X1Y115_I;
  assign RIOI3_X105Y117_ILOGIC_X1Y118_O = RIOB33_X105Y117_IOB_X1Y118_I;
  assign RIOI3_X105Y117_ILOGIC_X1Y117_O = RIOB33_X105Y117_IOB_X1Y117_I;
  assign RIOI3_X105Y121_ILOGIC_X1Y122_O = RIOB33_X105Y121_IOB_X1Y122_I;
  assign RIOI3_X105Y121_ILOGIC_X1Y121_O = RIOB33_X105Y121_IOB_X1Y121_I;
  assign RIOI3_X105Y123_ILOGIC_X1Y124_O = RIOB33_X105Y123_IOB_X1Y124_I;
  assign RIOI3_X105Y123_ILOGIC_X1Y123_O = RIOB33_X105Y123_IOB_X1Y123_I;
  assign RIOI3_X105Y125_ILOGIC_X1Y126_O = RIOB33_X105Y125_IOB_X1Y126_I;
  assign RIOI3_X105Y125_ILOGIC_X1Y125_O = RIOB33_X105Y125_IOB_X1Y125_I;
  assign RIOI3_X105Y127_ILOGIC_X1Y128_O = RIOB33_X105Y127_IOB_X1Y128_I;
  assign RIOI3_X105Y127_ILOGIC_X1Y127_O = RIOB33_X105Y127_IOB_X1Y127_I;
  assign RIOI3_X105Y129_ILOGIC_X1Y130_O = RIOB33_X105Y129_IOB_X1Y130_I;
  assign RIOI3_X105Y129_ILOGIC_X1Y129_O = RIOB33_X105Y129_IOB_X1Y129_I;
  assign RIOI3_X105Y133_ILOGIC_X1Y134_O = RIOB33_X105Y133_IOB_X1Y134_I;
  assign RIOI3_X105Y133_ILOGIC_X1Y133_O = RIOB33_X105Y133_IOB_X1Y133_I;
  assign RIOI3_X105Y135_ILOGIC_X1Y136_O = RIOB33_X105Y135_IOB_X1Y136_I;
  assign RIOI3_X105Y135_ILOGIC_X1Y135_O = RIOB33_X105Y135_IOB_X1Y135_I;
  assign RIOI3_X105Y139_ILOGIC_X1Y140_O = RIOB33_X105Y139_IOB_X1Y140_I;
  assign RIOI3_X105Y139_ILOGIC_X1Y139_O = RIOB33_X105Y139_IOB_X1Y139_I;
  assign RIOI3_X105Y141_ILOGIC_X1Y142_O = RIOB33_X105Y141_IOB_X1Y142_I;
  assign RIOI3_X105Y141_ILOGIC_X1Y141_O = RIOB33_X105Y141_IOB_X1Y141_I;
  assign RIOI3_X105Y145_ILOGIC_X1Y146_O = RIOB33_X105Y145_IOB_X1Y146_I;
  assign RIOI3_X105Y145_ILOGIC_X1Y145_O = RIOB33_X105Y145_IOB_X1Y145_I;
  assign RIOI3_X105Y147_ILOGIC_X1Y148_O = RIOB33_X105Y147_IOB_X1Y148_I;
  assign RIOI3_X105Y147_ILOGIC_X1Y147_O = RIOB33_X105Y147_IOB_X1Y147_I;
  assign RIOI3_X105Y151_OLOGIC_X1Y152_OQ = 1'b1;
  assign RIOI3_X105Y151_OLOGIC_X1Y152_TQ = 1'b1;
  assign RIOI3_X105Y151_OLOGIC_X1Y151_OQ = 1'b1;
  assign RIOI3_X105Y151_OLOGIC_X1Y151_TQ = 1'b1;
  assign RIOI3_X105Y153_OLOGIC_X1Y154_OQ = 1'b1;
  assign RIOI3_X105Y153_OLOGIC_X1Y154_TQ = 1'b1;
  assign RIOI3_X105Y153_OLOGIC_X1Y153_OQ = 1'b1;
  assign RIOI3_X105Y153_OLOGIC_X1Y153_TQ = 1'b1;
  assign RIOI3_X105Y155_OLOGIC_X1Y156_OQ = 1'b1;
  assign RIOI3_X105Y155_OLOGIC_X1Y156_TQ = 1'b1;
  assign RIOI3_X105Y155_OLOGIC_X1Y155_OQ = 1'b1;
  assign RIOI3_X105Y155_OLOGIC_X1Y155_TQ = 1'b1;
  assign RIOI3_X105Y159_OLOGIC_X1Y160_OQ = 1'b1;
  assign RIOI3_X105Y159_OLOGIC_X1Y160_TQ = 1'b1;
  assign RIOI3_X105Y159_OLOGIC_X1Y159_OQ = 1'b1;
  assign RIOI3_X105Y159_OLOGIC_X1Y159_TQ = 1'b1;
  assign RIOI3_X105Y161_OLOGIC_X1Y162_OQ = CLBLM_R_X7Y153_SLICE_X9Y153_C5Q;
  assign RIOI3_X105Y161_OLOGIC_X1Y162_TQ = 1'b1;
  assign RIOI3_X105Y161_OLOGIC_X1Y161_OQ = CLBLM_L_X10Y154_SLICE_X12Y154_DO5;
  assign RIOI3_X105Y161_OLOGIC_X1Y161_TQ = 1'b1;
  assign RIOI3_X105Y165_OLOGIC_X1Y166_OQ = CLBLM_L_X8Y153_SLICE_X10Y153_A5Q;
  assign RIOI3_X105Y165_OLOGIC_X1Y166_TQ = 1'b1;
  assign RIOI3_X105Y165_OLOGIC_X1Y165_OQ = CLBLM_L_X12Y152_SLICE_X16Y152_AO6;
  assign RIOI3_X105Y165_OLOGIC_X1Y165_TQ = 1'b1;
  assign RIOI3_X105Y167_OLOGIC_X1Y168_OQ = CLBLM_R_X5Y154_SLICE_X7Y154_AQ;
  assign RIOI3_X105Y167_OLOGIC_X1Y168_TQ = 1'b1;
  assign RIOI3_X105Y167_OLOGIC_X1Y167_OQ = CLBLM_R_X7Y153_SLICE_X9Y153_DQ;
  assign RIOI3_X105Y167_OLOGIC_X1Y167_TQ = 1'b1;
  assign RIOI3_X105Y171_OLOGIC_X1Y172_OQ = CLBLL_L_X2Y148_SLICE_X0Y148_AQ;
  assign RIOI3_X105Y171_OLOGIC_X1Y172_TQ = 1'b1;
  assign RIOI3_X105Y171_OLOGIC_X1Y171_OQ = CLBLM_L_X8Y153_SLICE_X11Y153_DO6;
  assign RIOI3_X105Y171_OLOGIC_X1Y171_TQ = 1'b1;
  assign RIOI3_X105Y173_OLOGIC_X1Y174_OQ = CLBLM_R_X5Y152_SLICE_X7Y152_DO6;
  assign RIOI3_X105Y173_OLOGIC_X1Y174_TQ = 1'b1;
  assign RIOI3_X105Y173_OLOGIC_X1Y173_OQ = CLBLM_R_X5Y152_SLICE_X7Y152_DQ;
  assign RIOI3_X105Y173_OLOGIC_X1Y173_TQ = 1'b1;
  assign RIOI3_X105Y175_OLOGIC_X1Y176_OQ = CLBLL_L_X2Y148_SLICE_X1Y148_BO6;
  assign RIOI3_X105Y175_OLOGIC_X1Y176_TQ = 1'b1;
  assign RIOI3_X105Y175_OLOGIC_X1Y175_OQ = CLBLM_L_X10Y144_SLICE_X12Y144_BO6;
  assign RIOI3_X105Y175_OLOGIC_X1Y175_TQ = 1'b1;
  assign RIOI3_X105Y177_OLOGIC_X1Y178_OQ = CLBLM_R_X5Y147_SLICE_X6Y147_AQ;
  assign RIOI3_X105Y177_OLOGIC_X1Y178_TQ = 1'b1;
  assign RIOI3_X105Y177_OLOGIC_X1Y177_OQ = CLBLL_L_X2Y146_SLICE_X1Y146_B5Q;
  assign RIOI3_X105Y177_OLOGIC_X1Y177_TQ = 1'b1;
  assign RIOI3_X105Y179_OLOGIC_X1Y180_OQ = CLBLM_L_X8Y145_SLICE_X11Y145_DQ;
  assign RIOI3_X105Y179_OLOGIC_X1Y180_TQ = 1'b1;
  assign RIOI3_X105Y179_OLOGIC_X1Y179_OQ = CLBLM_L_X8Y147_SLICE_X10Y147_BQ;
  assign RIOI3_X105Y179_OLOGIC_X1Y179_TQ = 1'b1;
  assign RIOI3_X105Y183_OLOGIC_X1Y184_OQ = CLBLM_R_X3Y148_SLICE_X3Y148_DO5;
  assign RIOI3_X105Y183_OLOGIC_X1Y184_TQ = 1'b1;
  assign RIOI3_X105Y183_OLOGIC_X1Y183_OQ = 1'b0;
  assign RIOI3_X105Y183_OLOGIC_X1Y183_TQ = 1'b1;
  assign RIOI3_X105Y185_OLOGIC_X1Y186_OQ = CLBLM_L_X10Y149_SLICE_X13Y149_BO6;
  assign RIOI3_X105Y185_OLOGIC_X1Y186_TQ = 1'b1;
  assign RIOI3_X105Y185_OLOGIC_X1Y185_OQ = CLBLM_L_X10Y153_SLICE_X12Y153_DO6;
  assign RIOI3_X105Y185_OLOGIC_X1Y185_TQ = 1'b1;
  assign RIOI3_X105Y189_OLOGIC_X1Y190_OQ = CLBLM_L_X12Y151_SLICE_X16Y151_AO5;
  assign RIOI3_X105Y189_OLOGIC_X1Y190_TQ = 1'b1;
  assign RIOI3_X105Y189_OLOGIC_X1Y189_OQ = CLBLM_R_X103Y178_SLICE_X163Y178_AO6;
  assign RIOI3_X105Y189_OLOGIC_X1Y189_TQ = 1'b1;
  assign RIOI3_X105Y191_OLOGIC_X1Y192_OQ = CLBLM_L_X12Y153_SLICE_X16Y153_AO6;
  assign RIOI3_X105Y191_OLOGIC_X1Y192_TQ = 1'b1;
  assign RIOI3_X105Y191_OLOGIC_X1Y191_OQ = CLBLM_L_X12Y149_SLICE_X17Y149_AO5;
  assign RIOI3_X105Y191_OLOGIC_X1Y191_TQ = 1'b1;
  assign RIOI3_X105Y195_OLOGIC_X1Y196_OQ = CLBLM_L_X12Y150_SLICE_X16Y150_AO6;
  assign RIOI3_X105Y195_OLOGIC_X1Y196_TQ = 1'b1;
  assign RIOI3_X105Y195_OLOGIC_X1Y195_OQ = CLBLM_L_X10Y149_SLICE_X13Y149_AO5;
  assign RIOI3_X105Y195_OLOGIC_X1Y195_TQ = 1'b1;
  assign RIOI3_X105Y197_OLOGIC_X1Y198_OQ = CLBLM_L_X12Y150_SLICE_X16Y150_AO5;
  assign RIOI3_X105Y197_OLOGIC_X1Y198_TQ = 1'b1;
  assign RIOI3_X105Y197_OLOGIC_X1Y197_OQ = CLBLM_L_X12Y152_SLICE_X16Y152_AO5;
  assign RIOI3_X105Y197_OLOGIC_X1Y197_TQ = 1'b1;
  assign RIOI3_SING_X105Y100_ILOGIC_X1Y100_O = RIOB33_SING_X105Y100_IOB_X1Y100_I;
  assign RIOI3_SING_X105Y149_ILOGIC_X1Y149_O = RIOB33_SING_X105Y149_IOB_X1Y149_I;
  assign RIOI3_SING_X105Y150_OLOGIC_X1Y150_OQ = 1'b1;
  assign RIOI3_SING_X105Y150_OLOGIC_X1Y150_TQ = 1'b1;
  assign RIOI3_SING_X105Y199_OLOGIC_X1Y199_OQ = CLBLM_R_X7Y153_SLICE_X8Y153_A5Q;
  assign RIOI3_SING_X105Y199_OLOGIC_X1Y199_TQ = 1'b1;
  assign RIOI3_TBYTESRC_X105Y107_ILOGIC_X1Y108_O = RIOB33_X105Y107_IOB_X1Y108_I;
  assign RIOI3_TBYTESRC_X105Y107_ILOGIC_X1Y107_O = RIOB33_X105Y107_IOB_X1Y107_I;
  assign RIOI3_TBYTESRC_X105Y119_ILOGIC_X1Y120_O = RIOB33_X105Y119_IOB_X1Y120_I;
  assign RIOI3_TBYTESRC_X105Y119_ILOGIC_X1Y119_O = RIOB33_X105Y119_IOB_X1Y119_I;
  assign RIOI3_TBYTESRC_X105Y131_ILOGIC_X1Y132_O = RIOB33_X105Y131_IOB_X1Y132_I;
  assign RIOI3_TBYTESRC_X105Y131_ILOGIC_X1Y131_O = RIOB33_X105Y131_IOB_X1Y131_I;
  assign RIOI3_TBYTESRC_X105Y143_ILOGIC_X1Y144_O = RIOB33_X105Y143_IOB_X1Y144_I;
  assign RIOI3_TBYTESRC_X105Y143_ILOGIC_X1Y143_O = RIOB33_X105Y143_IOB_X1Y143_I;
  assign RIOI3_TBYTESRC_X105Y157_OLOGIC_X1Y158_OQ = 1'b1;
  assign RIOI3_TBYTESRC_X105Y157_OLOGIC_X1Y158_TQ = 1'b1;
  assign RIOI3_TBYTESRC_X105Y157_OLOGIC_X1Y157_OQ = 1'b1;
  assign RIOI3_TBYTESRC_X105Y157_OLOGIC_X1Y157_TQ = 1'b1;
  assign RIOI3_TBYTESRC_X105Y169_OLOGIC_X1Y170_OQ = CLBLM_R_X3Y152_SLICE_X3Y152_BQ;
  assign RIOI3_TBYTESRC_X105Y169_OLOGIC_X1Y170_TQ = 1'b1;
  assign RIOI3_TBYTESRC_X105Y169_OLOGIC_X1Y169_OQ = CLBLM_R_X3Y152_SLICE_X3Y152_CQ;
  assign RIOI3_TBYTESRC_X105Y169_OLOGIC_X1Y169_TQ = 1'b1;
  assign RIOI3_TBYTESRC_X105Y181_OLOGIC_X1Y182_OQ = CLBLM_R_X11Y146_SLICE_X14Y146_BO5;
  assign RIOI3_TBYTESRC_X105Y181_OLOGIC_X1Y182_TQ = 1'b1;
  assign RIOI3_TBYTESRC_X105Y181_OLOGIC_X1Y181_OQ = CLBLM_L_X10Y154_SLICE_X12Y154_CO5;
  assign RIOI3_TBYTESRC_X105Y181_OLOGIC_X1Y181_TQ = 1'b1;
  assign RIOI3_TBYTESRC_X105Y193_OLOGIC_X1Y194_OQ = CLBLM_L_X12Y151_SLICE_X16Y151_BO6;
  assign RIOI3_TBYTESRC_X105Y193_OLOGIC_X1Y194_TQ = 1'b1;
  assign RIOI3_TBYTESRC_X105Y193_OLOGIC_X1Y193_OQ = CLBLM_L_X12Y151_SLICE_X16Y151_BO5;
  assign RIOI3_TBYTESRC_X105Y193_OLOGIC_X1Y193_TQ = 1'b1;
  assign RIOI3_TBYTETERM_X105Y113_ILOGIC_X1Y113_O = RIOB33_X105Y113_IOB_X1Y113_I;
  assign RIOI3_TBYTETERM_X105Y137_ILOGIC_X1Y138_O = RIOB33_X105Y137_IOB_X1Y138_I;
  assign RIOI3_TBYTETERM_X105Y137_ILOGIC_X1Y137_O = RIOB33_X105Y137_IOB_X1Y137_I;
  assign RIOI3_TBYTETERM_X105Y163_OLOGIC_X1Y164_OQ = CLBLM_L_X10Y153_SLICE_X12Y153_AQ;
  assign RIOI3_TBYTETERM_X105Y163_OLOGIC_X1Y164_TQ = 1'b1;
  assign RIOI3_TBYTETERM_X105Y163_OLOGIC_X1Y163_OQ = CLBLM_R_X7Y151_SLICE_X9Y151_D5Q;
  assign RIOI3_TBYTETERM_X105Y163_OLOGIC_X1Y163_TQ = 1'b1;
  assign RIOI3_TBYTETERM_X105Y187_OLOGIC_X1Y188_OQ = CLBLM_R_X11Y146_SLICE_X14Y146_BO5;
  assign RIOI3_TBYTETERM_X105Y187_OLOGIC_X1Y188_TQ = 1'b1;
  assign RIOI3_TBYTETERM_X105Y187_OLOGIC_X1Y187_OQ = CLBLM_R_X103Y178_SLICE_X163Y178_AO6;
  assign RIOI3_TBYTETERM_X105Y187_OLOGIC_X1Y187_TQ = 1'b1;
  assign CLBLM_L_X8Y145_SLICE_X10Y145_B1 = CLBLM_R_X7Y144_SLICE_X9Y144_DO6;
  assign CLBLM_L_X8Y145_SLICE_X10Y145_B2 = CLBLM_R_X7Y144_SLICE_X9Y144_BQ;
  assign CLBLM_L_X8Y145_SLICE_X10Y145_B3 = CLBLM_L_X8Y146_SLICE_X10Y146_AO6;
  assign CLBLM_L_X8Y145_SLICE_X10Y145_B4 = CLBLM_L_X10Y148_SLICE_X12Y148_AO5;
  assign CLBLM_L_X8Y145_SLICE_X10Y145_B5 = CLBLM_L_X12Y151_SLICE_X16Y151_AQ;
  assign CLBLM_L_X8Y145_SLICE_X10Y145_B6 = CLBLM_L_X8Y144_SLICE_X10Y144_CO6;
  assign CLBLM_L_X10Y155_SLICE_X12Y155_CLK = CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O;
  assign CLBLM_L_X10Y155_SLICE_X12Y155_D1 = 1'b1;
  assign CLBLM_L_X10Y155_SLICE_X12Y155_D2 = 1'b1;
  assign CLBLM_L_X8Y145_SLICE_X10Y145_C1 = CLBLM_L_X8Y144_SLICE_X11Y144_BQ;
  assign CLBLM_L_X8Y145_SLICE_X10Y145_C2 = CLBLM_R_X7Y145_SLICE_X9Y145_BO6;
  assign CLBLM_L_X8Y145_SLICE_X10Y145_C3 = CLBLM_L_X10Y148_SLICE_X12Y148_AO5;
  assign CLBLM_L_X8Y145_SLICE_X10Y145_C4 = CLBLM_L_X10Y149_SLICE_X13Y149_AQ;
  assign CLBLM_L_X8Y145_SLICE_X10Y145_C5 = CLBLM_L_X12Y146_SLICE_X16Y146_CO6;
  assign CLBLM_L_X8Y145_SLICE_X10Y145_C6 = CLBLL_L_X4Y148_SLICE_X4Y148_CQ;
  assign CLBLM_L_X10Y155_SLICE_X12Y155_D3 = 1'b1;
  assign CLBLM_L_X10Y155_SLICE_X12Y155_D4 = 1'b1;
  assign CLBLM_L_X10Y155_SLICE_X12Y155_D5 = 1'b1;
  assign CLBLM_L_X8Y145_SLICE_X10Y145_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X10Y155_SLICE_X12Y155_D6 = 1'b1;
  assign CLBLM_L_X8Y145_SLICE_X10Y145_D1 = CLBLL_L_X4Y148_SLICE_X4Y148_CQ;
  assign CLBLM_L_X8Y145_SLICE_X10Y145_D2 = CLBLM_L_X10Y148_SLICE_X12Y148_AO5;
  assign CLBLM_L_X8Y145_SLICE_X10Y145_D3 = CLBLM_R_X7Y145_SLICE_X9Y145_CO6;
  assign CLBLM_L_X8Y145_SLICE_X10Y145_D4 = CLBLM_R_X7Y142_SLICE_X8Y142_DQ;
  assign CLBLM_L_X8Y145_SLICE_X10Y145_D5 = CLBLM_L_X12Y146_SLICE_X16Y146_CO6;
  assign CLBLM_L_X8Y145_SLICE_X10Y145_D6 = CLBLL_L_X4Y149_SLICE_X5Y149_C5Q;
  assign CLBLM_R_X11Y149_SLICE_X15Y149_A1 = CLBLM_R_X11Y151_SLICE_X14Y151_CO6;
  assign CLBLM_R_X11Y149_SLICE_X15Y149_A2 = CLBLM_L_X12Y147_SLICE_X16Y147_DO6;
  assign CLBLM_R_X11Y149_SLICE_X15Y149_A3 = CLBLM_R_X11Y147_SLICE_X15Y147_AO6;
  assign CLBLM_R_X11Y149_SLICE_X15Y149_A4 = CLBLM_R_X11Y149_SLICE_X15Y149_BO6;
  assign CLBLM_R_X11Y149_SLICE_X15Y149_A5 = CLBLM_L_X8Y146_SLICE_X10Y146_BO6;
  assign CLBLM_R_X11Y149_SLICE_X15Y149_A6 = CLBLM_L_X8Y149_SLICE_X10Y149_DO6;
  assign CLBLM_R_X11Y149_SLICE_X15Y149_B1 = CLBLL_L_X4Y150_SLICE_X4Y150_CQ;
  assign CLBLM_R_X11Y149_SLICE_X15Y149_B2 = CLBLM_R_X11Y144_SLICE_X14Y144_CO6;
  assign CLBLM_R_X11Y149_SLICE_X15Y149_B3 = CLBLM_L_X12Y146_SLICE_X16Y146_AO6;
  assign CLBLM_R_X11Y149_SLICE_X15Y149_B4 = CLBLM_L_X8Y152_SLICE_X10Y152_DQ;
  assign CLBLM_R_X11Y149_SLICE_X15Y149_B5 = CLBLM_L_X8Y151_SLICE_X11Y151_BO6;
  assign CLBLM_R_X11Y149_SLICE_X15Y149_B6 = CLBLM_R_X7Y148_SLICE_X8Y148_AO5;
  assign LIOI3_X0Y155_OLOGIC_X0Y156_D1 = CLBLM_R_X3Y152_SLICE_X3Y152_CQ;
  assign CLBLM_R_X11Y149_SLICE_X15Y149_C1 = CLBLM_L_X10Y145_SLICE_X13Y145_BO6;
  assign CLBLM_R_X11Y149_SLICE_X15Y149_C2 = CLBLM_R_X11Y149_SLICE_X14Y149_CO6;
  assign CLBLM_R_X11Y149_SLICE_X15Y149_C3 = CLBLM_R_X11Y152_SLICE_X15Y152_AQ;
  assign CLBLM_R_X11Y149_SLICE_X15Y149_C4 = CLBLM_R_X11Y148_SLICE_X15Y148_DO6;
  assign CLBLM_R_X11Y149_SLICE_X15Y149_C5 = RIOB33_X105Y131_IOB_X1Y132_I;
  assign CLBLL_L_X4Y152_SLICE_X4Y152_A1 = CLBLM_R_X3Y143_SLICE_X3Y143_BQ;
  assign CLBLL_L_X4Y152_SLICE_X4Y152_A2 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLL_L_X4Y152_SLICE_X4Y152_A3 = CLBLM_L_X10Y149_SLICE_X12Y149_BQ;
  assign CLBLL_L_X4Y152_SLICE_X4Y152_A4 = CLBLL_L_X4Y152_SLICE_X5Y152_BQ;
  assign CLBLL_L_X4Y152_SLICE_X4Y152_A5 = CLBLL_L_X4Y142_SLICE_X4Y142_AQ;
  assign CLBLL_L_X4Y152_SLICE_X4Y152_A6 = CLBLM_L_X8Y152_SLICE_X11Y152_BQ;
  assign CLBLM_R_X11Y149_SLICE_X15Y149_C6 = CLBLM_L_X12Y149_SLICE_X16Y149_CO6;
  assign LIOI3_X0Y155_OLOGIC_X0Y156_T1 = 1'b1;
  assign CLBLL_L_X4Y152_SLICE_X4Y152_B1 = CLBLL_L_X4Y147_SLICE_X4Y147_B5Q;
  assign CLBLL_L_X4Y152_SLICE_X4Y152_B2 = CLBLM_R_X3Y145_SLICE_X2Y145_DO6;
  assign CLBLL_L_X4Y152_SLICE_X4Y152_B3 = CLBLL_L_X4Y151_SLICE_X4Y151_B5Q;
  assign CLBLL_L_X4Y152_SLICE_X4Y152_B4 = CLBLL_L_X4Y152_SLICE_X5Y152_BQ;
  assign CLBLL_L_X4Y152_SLICE_X4Y152_B5 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLL_L_X4Y152_SLICE_X4Y152_B6 = 1'b1;
  assign CLBLM_R_X11Y149_SLICE_X15Y149_D1 = CLBLM_L_X10Y150_SLICE_X13Y150_BO5;
  assign CLBLM_R_X11Y149_SLICE_X15Y149_D2 = CLBLM_L_X12Y149_SLICE_X16Y149_DO6;
  assign CLBLM_R_X11Y149_SLICE_X15Y149_D3 = 1'b1;
  assign CLBLL_L_X4Y152_SLICE_X4Y152_C1 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLL_L_X4Y152_SLICE_X4Y152_C2 = CLBLM_R_X7Y152_SLICE_X8Y152_DQ;
  assign CLBLL_L_X4Y152_SLICE_X4Y152_C3 = CLBLL_L_X4Y152_SLICE_X4Y152_DQ;
  assign CLBLL_L_X4Y152_SLICE_X4Y152_C4 = CLBLL_L_X4Y152_SLICE_X4Y152_BQ;
  assign CLBLL_L_X4Y152_SLICE_X4Y152_C5 = CLBLM_R_X5Y153_SLICE_X6Y153_DQ;
  assign CLBLL_L_X4Y152_SLICE_X4Y152_C6 = 1'b1;
  assign CLBLM_R_X3Y143_SLICE_X2Y143_B2 = LIOB33_X0Y57_IOB_X0Y58_I;
  assign CLBLM_R_X11Y149_SLICE_X14Y149_A1 = CLBLM_L_X8Y150_SLICE_X10Y150_DO6;
  assign CLBLL_L_X4Y152_SLICE_X4Y152_CLK = CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O;
  assign CLBLM_R_X11Y149_SLICE_X14Y149_A2 = CLBLM_L_X12Y147_SLICE_X16Y147_DO6;
  assign CLBLM_R_X11Y149_SLICE_X14Y149_A3 = CLBLM_L_X10Y148_SLICE_X12Y148_DO6;
  assign CLBLM_R_X11Y149_SLICE_X14Y149_A4 = CLBLM_R_X11Y149_SLICE_X14Y149_BO6;
  assign CLBLM_R_X11Y149_SLICE_X14Y149_A5 = CLBLM_L_X8Y146_SLICE_X10Y146_DO6;
  assign CLBLM_R_X11Y149_SLICE_X14Y149_A6 = CLBLM_R_X11Y147_SLICE_X14Y147_CO6;
  assign CLBLL_L_X4Y152_SLICE_X4Y152_D1 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLL_L_X4Y152_SLICE_X4Y152_D2 = CLBLL_L_X4Y152_SLICE_X4Y152_CQ;
  assign CLBLL_L_X4Y152_SLICE_X4Y152_D3 = CLBLL_L_X4Y152_SLICE_X4Y152_DQ;
  assign CLBLL_L_X4Y152_SLICE_X4Y152_D4 = CLBLL_L_X4Y152_SLICE_X4Y152_BQ;
  assign CLBLL_L_X4Y152_SLICE_X4Y152_D5 = CLBLM_R_X5Y153_SLICE_X6Y153_DQ;
  assign CLBLL_L_X4Y152_SLICE_X4Y152_D6 = CLBLM_R_X5Y152_SLICE_X7Y152_A5Q;
  assign CLBLM_R_X11Y149_SLICE_X14Y149_B3 = CLBLM_R_X13Y149_SLICE_X18Y149_AO6;
  assign CLBLM_R_X11Y149_SLICE_X14Y149_B4 = CLBLM_L_X10Y149_SLICE_X13Y149_DO6;
  assign CLBLM_R_X11Y149_SLICE_X14Y149_B5 = CLBLM_L_X12Y149_SLICE_X17Y149_DO6;
  assign CLBLM_R_X11Y149_SLICE_X14Y149_B6 = CLBLM_R_X5Y146_SLICE_X7Y146_AQ;
  assign CLBLM_R_X11Y149_SLICE_X14Y149_C1 = CLBLM_L_X8Y149_SLICE_X11Y149_BO6;
  assign CLBLM_R_X11Y149_SLICE_X14Y149_C2 = CLBLM_L_X10Y147_SLICE_X13Y147_CO6;
  assign CLBLM_R_X11Y149_SLICE_X14Y149_C3 = CLBLM_R_X11Y148_SLICE_X14Y148_CO6;
  assign CLBLM_R_X11Y149_SLICE_X14Y149_C4 = CLBLM_L_X10Y149_SLICE_X12Y149_DO6;
  assign CLBLM_R_X11Y149_SLICE_X14Y149_C5 = CLBLM_L_X12Y147_SLICE_X16Y147_DO6;
  assign CLBLM_R_X11Y149_SLICE_X14Y149_C6 = CLBLM_R_X11Y148_SLICE_X14Y148_BO6;
  assign CLBLM_R_X11Y149_SLICE_X14Y149_D1 = CLBLM_L_X8Y149_SLICE_X11Y149_CO6;
  assign CLBLM_R_X11Y149_SLICE_X14Y149_D2 = CLBLM_R_X11Y150_SLICE_X14Y150_CO6;
  assign CLBLM_R_X11Y149_SLICE_X14Y149_D3 = CLBLM_R_X7Y150_SLICE_X9Y150_DO6;
  assign CLBLM_R_X11Y149_SLICE_X14Y149_D4 = CLBLM_L_X10Y149_SLICE_X13Y149_DO6;
  assign CLBLM_R_X11Y149_SLICE_X14Y149_D5 = CLBLM_L_X8Y150_SLICE_X10Y150_DO6;
  assign CLBLM_R_X11Y149_SLICE_X14Y149_D6 = 1'b1;
  assign RIOB33_SING_X105Y150_IOB_X1Y150_O = 1'b1;
  assign RIOI3_TBYTESRC_X105Y181_OLOGIC_X1Y182_D1 = CLBLM_R_X11Y146_SLICE_X14Y146_BO5;
  assign CLBLL_L_X4Y152_SLICE_X5Y152_A1 = CLBLL_L_X2Y150_SLICE_X1Y150_AQ;
  assign CLBLL_L_X4Y152_SLICE_X5Y152_A2 = CLBLM_R_X3Y152_SLICE_X3Y152_AQ;
  assign CLBLL_L_X4Y152_SLICE_X5Y152_A3 = CLBLL_L_X4Y152_SLICE_X5Y152_AQ;
  assign CLBLL_L_X4Y152_SLICE_X5Y152_A4 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLL_L_X4Y152_SLICE_X5Y152_A5 = CLBLL_L_X4Y144_SLICE_X4Y144_C5Q;
  assign CLBLL_L_X4Y152_SLICE_X5Y152_A6 = CLBLL_L_X4Y152_SLICE_X5Y152_CO6;
  assign CLBLL_L_X4Y152_SLICE_X5Y152_AX = CLBLL_L_X4Y152_SLICE_X5Y152_CO5;
  assign CLBLL_L_X4Y152_SLICE_X5Y152_B1 = CLBLM_L_X10Y153_SLICE_X13Y153_A5Q;
  assign CLBLL_L_X4Y152_SLICE_X5Y152_B2 = CLBLM_R_X3Y143_SLICE_X3Y143_BQ;
  assign CLBLL_L_X4Y152_SLICE_X5Y152_B3 = CLBLL_L_X4Y146_SLICE_X5Y146_DQ;
  assign CLBLL_L_X4Y152_SLICE_X5Y152_B4 = CLBLM_R_X5Y153_SLICE_X7Y153_BQ;
  assign CLBLL_L_X4Y152_SLICE_X5Y152_B5 = CLBLL_L_X4Y142_SLICE_X4Y142_AQ;
  assign CLBLL_L_X4Y152_SLICE_X5Y152_B6 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign RIOI3_TBYTESRC_X105Y181_OLOGIC_X1Y182_T1 = 1'b1;
  assign CLBLL_L_X4Y152_SLICE_X5Y152_C1 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLL_L_X4Y152_SLICE_X5Y152_C2 = CLBLM_R_X5Y152_SLICE_X6Y152_BQ;
  assign CLBLL_L_X4Y152_SLICE_X5Y152_C3 = CLBLL_L_X2Y150_SLICE_X1Y150_AQ;
  assign CLBLL_L_X4Y152_SLICE_X5Y152_C4 = CLBLL_L_X4Y152_SLICE_X5Y152_A5Q;
  assign CLBLL_L_X4Y152_SLICE_X5Y152_C5 = CLBLL_L_X4Y152_SLICE_X5Y152_DO6;
  assign CLBLL_L_X4Y152_SLICE_X5Y152_C6 = 1'b1;
  assign RIOI3_TBYTESRC_X105Y181_OLOGIC_X1Y181_D1 = CLBLM_L_X10Y154_SLICE_X12Y154_CO5;
  assign CLBLL_L_X4Y152_SLICE_X5Y152_CLK = CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O;
  assign CLBLL_L_X4Y152_SLICE_X5Y152_D1 = CLBLM_R_X5Y154_SLICE_X6Y154_AQ;
  assign CLBLL_L_X4Y152_SLICE_X5Y152_D2 = CLBLL_L_X4Y153_SLICE_X5Y153_AQ;
  assign CLBLL_L_X4Y152_SLICE_X5Y152_D3 = CLBLM_R_X7Y153_SLICE_X9Y153_AQ;
  assign CLBLL_L_X4Y152_SLICE_X5Y152_D4 = CLBLM_R_X3Y149_SLICE_X3Y149_AQ;
  assign CLBLL_L_X4Y152_SLICE_X5Y152_D5 = CLBLM_R_X3Y149_SLICE_X2Y149_AQ;
  assign CLBLL_L_X4Y152_SLICE_X5Y152_D6 = CLBLM_R_X5Y154_SLICE_X6Y154_BQ;
  assign RIOI3_TBYTESRC_X105Y181_OLOGIC_X1Y181_T1 = 1'b1;
  assign CLBLM_L_X8Y146_SLICE_X11Y146_A1 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_L_X8Y146_SLICE_X11Y146_A2 = CLBLM_L_X8Y146_SLICE_X11Y146_BQ;
  assign CLBLM_L_X8Y146_SLICE_X11Y146_A3 = CLBLM_L_X8Y146_SLICE_X11Y146_AQ;
  assign CLBLM_L_X8Y146_SLICE_X11Y146_A4 = 1'b1;
  assign CLBLM_L_X8Y146_SLICE_X11Y146_A5 = CLBLM_R_X7Y146_SLICE_X9Y146_AQ;
  assign CLBLM_L_X8Y146_SLICE_X11Y146_A6 = CLBLM_R_X11Y146_SLICE_X14Y146_DO6;
  assign CLBLM_L_X8Y146_SLICE_X11Y146_B1 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_L_X8Y146_SLICE_X11Y146_B2 = CLBLM_L_X8Y147_SLICE_X11Y147_C5Q;
  assign CLBLM_L_X8Y146_SLICE_X11Y146_B3 = CLBLM_R_X7Y146_SLICE_X8Y146_D5Q;
  assign CLBLM_L_X8Y146_SLICE_X11Y146_B4 = 1'b1;
  assign CLBLM_L_X8Y146_SLICE_X11Y146_B5 = CLBLM_R_X7Y153_SLICE_X9Y153_C5Q;
  assign CLBLM_L_X8Y146_SLICE_X11Y146_B6 = 1'b1;
  assign CLBLM_L_X8Y146_SLICE_X11Y146_C1 = CLBLM_L_X8Y146_SLICE_X11Y146_C5Q;
  assign CLBLM_L_X8Y146_SLICE_X11Y146_C2 = CLBLM_R_X3Y145_SLICE_X3Y145_BQ;
  assign CLBLM_L_X8Y146_SLICE_X11Y146_C3 = CLBLM_L_X8Y143_SLICE_X11Y143_AQ;
  assign CLBLM_L_X8Y146_SLICE_X11Y146_C4 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_L_X8Y146_SLICE_X11Y146_C5 = CLBLM_R_X13Y149_SLICE_X18Y149_AO6;
  assign CLBLM_L_X8Y146_SLICE_X11Y146_C6 = 1'b1;
  assign CLBLM_L_X8Y146_SLICE_X11Y146_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X8Y146_SLICE_X11Y146_D1 = CLBLM_L_X8Y148_SLICE_X11Y148_BQ;
  assign CLBLM_L_X8Y146_SLICE_X11Y146_D2 = CLBLM_R_X5Y152_SLICE_X6Y152_CQ;
  assign CLBLM_L_X8Y146_SLICE_X11Y146_D3 = CLBLL_L_X4Y142_SLICE_X5Y142_AQ;
  assign CLBLM_L_X8Y146_SLICE_X11Y146_D4 = CLBLM_L_X10Y146_SLICE_X13Y146_CQ;
  assign CLBLM_L_X8Y146_SLICE_X11Y146_D5 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_L_X8Y146_SLICE_X11Y146_D6 = 1'b1;
  assign LIOB33_X0Y151_IOB_X0Y151_O = CLBLL_L_X2Y146_SLICE_X0Y146_CQ;
  assign LIOB33_X0Y151_IOB_X0Y152_O = CLBLL_L_X4Y147_SLICE_X5Y147_C5Q;
  assign LIOI3_SING_X0Y199_OLOGIC_X0Y199_D1 = 1'b1;
  assign RIOB33_SING_X105Y199_IOB_X1Y199_O = CLBLM_R_X7Y153_SLICE_X8Y153_A5Q;
  assign CLBLM_L_X8Y146_SLICE_X10Y146_A1 = CLBLM_R_X7Y153_SLICE_X8Y153_A5Q;
  assign CLBLM_L_X8Y146_SLICE_X10Y146_A2 = CLBLM_R_X7Y149_SLICE_X8Y149_AQ;
  assign CLBLM_L_X8Y146_SLICE_X10Y146_A3 = CLBLM_R_X7Y146_SLICE_X9Y146_CO6;
  assign CLBLM_L_X8Y146_SLICE_X10Y146_A4 = CLBLL_L_X4Y148_SLICE_X4Y148_CQ;
  assign CLBLM_L_X8Y146_SLICE_X10Y146_A5 = CLBLM_R_X7Y144_SLICE_X9Y144_B5Q;
  assign CLBLM_L_X8Y146_SLICE_X10Y146_A6 = 1'b1;
  assign LIOI3_SING_X0Y199_OLOGIC_X0Y199_T1 = 1'b1;
  assign CLBLM_L_X8Y146_SLICE_X10Y146_AX = CLBLM_R_X5Y142_SLICE_X7Y142_A5Q;
  assign CLBLM_L_X8Y146_SLICE_X10Y146_B1 = CLBLM_R_X7Y144_SLICE_X8Y144_DQ;
  assign CLBLM_L_X8Y146_SLICE_X10Y146_B2 = CLBLL_L_X4Y142_SLICE_X5Y142_C5Q;
  assign CLBLM_L_X8Y146_SLICE_X10Y146_B3 = CLBLM_L_X8Y146_SLICE_X10Y146_AO5;
  assign CLBLM_L_X8Y146_SLICE_X10Y146_B4 = CLBLM_R_X7Y146_SLICE_X9Y146_DO6;
  assign CLBLM_L_X8Y146_SLICE_X10Y146_B5 = CLBLM_L_X8Y146_SLICE_X10Y146_CO6;
  assign CLBLM_L_X8Y146_SLICE_X10Y146_B6 = 1'b1;
  assign RIOI3_X105Y139_ILOGIC_X1Y140_D = RIOB33_X105Y139_IOB_X1Y140_I;
  assign RIOI3_X105Y139_ILOGIC_X1Y139_D = RIOB33_X105Y139_IOB_X1Y139_I;
  assign CLBLM_L_X8Y146_SLICE_X10Y146_BX = CLBLM_L_X8Y145_SLICE_X10Y145_A5Q;
  assign CLBLM_L_X8Y146_SLICE_X10Y146_C1 = CLBLM_L_X8Y144_SLICE_X10Y144_AQ;
  assign CLBLM_L_X8Y146_SLICE_X10Y146_C2 = CLBLM_L_X8Y146_SLICE_X10Y146_AO6;
  assign CLBLM_L_X8Y146_SLICE_X10Y146_C3 = CLBLM_R_X11Y146_SLICE_X14Y146_CO6;
  assign CLBLM_L_X8Y146_SLICE_X10Y146_C4 = CLBLM_L_X10Y148_SLICE_X12Y148_AO5;
  assign CLBLM_L_X8Y146_SLICE_X10Y146_C5 = CLBLM_R_X7Y148_SLICE_X9Y148_A5Q;
  assign CLBLM_L_X8Y146_SLICE_X10Y146_C6 = CLBLM_L_X10Y149_SLICE_X12Y149_BQ;
  assign CLBLM_L_X8Y146_SLICE_X10Y146_CE = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_L_X8Y146_SLICE_X10Y146_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X8Y146_SLICE_X10Y146_D1 = CLBLM_R_X5Y140_SLICE_X6Y140_A5Q;
  assign CLBLM_L_X8Y146_SLICE_X10Y146_D2 = CLBLM_R_X5Y150_SLICE_X7Y150_A5Q;
  assign CLBLM_L_X8Y146_SLICE_X10Y146_D3 = CLBLM_R_X11Y146_SLICE_X14Y146_CO6;
  assign CLBLM_L_X8Y146_SLICE_X10Y146_D4 = CLBLM_L_X8Y146_SLICE_X10Y146_AO5;
  assign CLBLM_L_X8Y146_SLICE_X10Y146_D5 = CLBLM_R_X5Y143_SLICE_X6Y143_CQ;
  assign CLBLM_L_X8Y146_SLICE_X10Y146_D6 = CLBLM_R_X7Y146_SLICE_X9Y146_DO6;
  assign CLBLM_R_X3Y144_SLICE_X3Y144_B1 = CLBLM_R_X5Y147_SLICE_X6Y147_B5Q;
  assign CLBLM_R_X3Y144_SLICE_X3Y144_B2 = CLBLM_R_X3Y144_SLICE_X2Y144_BO6;
  assign CLBLM_R_X11Y150_SLICE_X15Y150_A1 = CLBLM_R_X11Y150_SLICE_X15Y150_DO6;
  assign CLBLM_R_X11Y150_SLICE_X15Y150_A2 = CLBLM_L_X12Y149_SLICE_X17Y149_CO6;
  assign CLBLM_R_X11Y150_SLICE_X15Y150_A3 = CLBLM_R_X7Y153_SLICE_X9Y153_BQ;
  assign CLBLM_R_X11Y150_SLICE_X15Y150_A4 = CLBLM_L_X8Y150_SLICE_X11Y150_DO6;
  assign CLBLM_R_X11Y150_SLICE_X15Y150_A5 = CLBLM_R_X7Y143_SLICE_X9Y143_BQ;
  assign CLBLM_R_X11Y150_SLICE_X15Y150_A6 = CLBLM_L_X8Y150_SLICE_X10Y150_BO6;
  assign CLBLM_R_X11Y150_SLICE_X15Y150_B1 = CLBLM_R_X11Y150_SLICE_X15Y150_DO6;
  assign CLBLM_R_X11Y150_SLICE_X15Y150_B2 = CLBLM_L_X12Y149_SLICE_X17Y149_CO6;
  assign CLBLM_R_X11Y150_SLICE_X15Y150_B3 = CLBLM_R_X7Y153_SLICE_X9Y153_BQ;
  assign CLBLM_R_X3Y144_SLICE_X3Y144_B5 = CLBLM_R_X5Y143_SLICE_X6Y143_D5Q;
  assign CLBLM_R_X11Y150_SLICE_X15Y150_B4 = CLBLM_L_X8Y150_SLICE_X11Y150_DO6;
  assign CLBLM_R_X11Y150_SLICE_X15Y150_B5 = CLBLM_R_X7Y149_SLICE_X8Y149_CO6;
  assign CLBLM_R_X11Y150_SLICE_X15Y150_B6 = CLBLM_R_X11Y151_SLICE_X15Y151_BO6;
  assign CLBLL_L_X4Y153_SLICE_X4Y153_A1 = CLBLM_R_X5Y154_SLICE_X7Y154_AQ;
  assign CLBLL_L_X4Y153_SLICE_X4Y153_A2 = CLBLL_L_X4Y152_SLICE_X4Y152_BQ;
  assign CLBLL_L_X4Y153_SLICE_X4Y153_A3 = 1'b1;
  assign CLBLL_L_X4Y153_SLICE_X4Y153_A4 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLL_L_X4Y153_SLICE_X4Y153_A5 = CLBLM_R_X5Y150_SLICE_X6Y150_C5Q;
  assign CLBLL_L_X4Y153_SLICE_X4Y153_A6 = 1'b1;
  assign CLBLM_R_X11Y150_SLICE_X15Y150_C1 = CLBLM_L_X12Y150_SLICE_X16Y150_BO6;
  assign CLBLM_R_X11Y150_SLICE_X15Y150_C2 = CLBLM_R_X7Y150_SLICE_X8Y150_CO6;
  assign CLBLM_R_X11Y150_SLICE_X15Y150_C3 = CLBLM_L_X8Y149_SLICE_X10Y149_DO6;
  assign CLBLL_L_X4Y153_SLICE_X4Y153_B1 = CLBLM_L_X10Y152_SLICE_X13Y152_AQ;
  assign CLBLL_L_X4Y153_SLICE_X4Y153_B2 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLL_L_X4Y153_SLICE_X4Y153_B3 = CLBLM_L_X10Y153_SLICE_X13Y153_A5Q;
  assign CLBLL_L_X4Y153_SLICE_X4Y153_B4 = CLBLL_L_X4Y149_SLICE_X4Y149_CQ;
  assign CLBLL_L_X4Y153_SLICE_X4Y153_B5 = 1'b1;
  assign CLBLL_L_X4Y153_SLICE_X4Y153_B6 = 1'b1;
  assign CLBLM_R_X11Y150_SLICE_X15Y150_D1 = 1'b1;
  assign CLBLM_R_X11Y150_SLICE_X15Y150_D2 = CLBLM_R_X7Y151_SLICE_X8Y151_CQ;
  assign CLBLL_L_X4Y153_SLICE_X4Y153_C1 = CLBLL_L_X4Y142_SLICE_X4Y142_AQ;
  assign CLBLL_L_X4Y153_SLICE_X4Y153_C2 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLL_L_X4Y153_SLICE_X4Y153_C3 = RIOB33_X105Y131_IOB_X1Y131_I;
  assign CLBLL_L_X4Y153_SLICE_X4Y153_C4 = CLBLM_R_X5Y142_SLICE_X7Y142_CO6;
  assign CLBLL_L_X4Y153_SLICE_X4Y153_C5 = RIOB33_SING_X105Y100_IOB_X1Y100_I;
  assign CLBLL_L_X4Y153_SLICE_X4Y153_C6 = 1'b1;
  assign CLBLM_R_X11Y150_SLICE_X15Y150_D3 = CLBLM_L_X10Y148_SLICE_X12Y148_AO6;
  assign CLBLM_R_X11Y150_SLICE_X15Y150_D4 = CLBLM_R_X7Y152_SLICE_X8Y152_CQ;
  assign CLBLL_L_X4Y153_SLICE_X4Y153_CLK = CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O;
  assign CLBLM_R_X11Y150_SLICE_X14Y150_A1 = CLBLM_L_X10Y146_SLICE_X13Y146_DO6;
  assign CLBLM_R_X11Y150_SLICE_X14Y150_A2 = CLBLM_R_X11Y151_SLICE_X14Y151_BO6;
  assign CLBLM_R_X11Y150_SLICE_X14Y150_A3 = CLBLM_L_X12Y149_SLICE_X17Y149_BO5;
  assign CLBLM_R_X11Y150_SLICE_X14Y150_A4 = CLBLM_R_X7Y146_SLICE_X9Y146_BQ;
  assign CLBLM_R_X11Y150_SLICE_X14Y150_A5 = CLBLM_R_X11Y151_SLICE_X14Y151_AQ;
  assign CLBLL_L_X4Y153_SLICE_X4Y153_D1 = CLBLM_R_X5Y147_SLICE_X7Y147_AQ;
  assign CLBLL_L_X4Y153_SLICE_X4Y153_D2 = CLBLL_L_X4Y153_SLICE_X5Y153_A5Q;
  assign CLBLL_L_X4Y153_SLICE_X4Y153_D3 = CLBLM_R_X7Y145_SLICE_X8Y145_A5Q;
  assign CLBLL_L_X4Y153_SLICE_X4Y153_D4 = RIOB33_X105Y131_IOB_X1Y131_I;
  assign CLBLL_L_X4Y153_SLICE_X4Y153_D5 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLL_L_X4Y153_SLICE_X4Y153_D6 = 1'b1;
  assign CLBLM_R_X11Y150_SLICE_X14Y150_A6 = CLBLM_R_X11Y148_SLICE_X15Y148_AO6;
  assign CLBLM_R_X11Y150_SLICE_X14Y150_AX = CLBLM_L_X10Y150_SLICE_X13Y150_AQ;
  assign CLBLM_R_X11Y150_SLICE_X14Y150_B1 = CLBLM_R_X7Y152_SLICE_X8Y152_DQ;
  assign CLBLM_R_X11Y150_SLICE_X14Y150_B2 = CLBLM_R_X7Y146_SLICE_X8Y146_C5Q;
  assign CLBLM_R_X11Y150_SLICE_X14Y150_B3 = CLBLM_L_X10Y150_SLICE_X13Y150_BO6;
  assign CLBLM_R_X11Y150_SLICE_X14Y150_B4 = CLBLM_L_X8Y150_SLICE_X10Y150_BO6;
  assign CLBLM_R_X11Y150_SLICE_X14Y150_B5 = CLBLM_R_X11Y150_SLICE_X14Y150_AO6;
  assign CLBLM_R_X11Y150_SLICE_X14Y150_B6 = CLBLM_L_X10Y148_SLICE_X12Y148_AO6;
  assign CLBLM_R_X11Y150_SLICE_X14Y150_C1 = CLBLM_L_X12Y149_SLICE_X17Y149_BO5;
  assign CLBLM_R_X11Y150_SLICE_X14Y150_C2 = CLBLM_R_X5Y146_SLICE_X7Y146_AQ;
  assign CLBLM_R_X11Y150_SLICE_X14Y150_C3 = CLBLM_L_X10Y146_SLICE_X13Y146_DO6;
  assign CLBLM_R_X11Y150_SLICE_X14Y150_C4 = CLBLM_R_X13Y149_SLICE_X18Y149_AO6;
  assign CLBLM_R_X11Y150_SLICE_X14Y150_C5 = CLBLM_L_X8Y152_SLICE_X11Y152_CQ;
  assign CLBLM_R_X11Y150_SLICE_X14Y150_C6 = CLBLM_L_X12Y150_SLICE_X16Y150_CO6;
  assign CLBLM_R_X11Y150_SLICE_X14Y150_CE = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X11Y150_SLICE_X14Y150_CLK = CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O;
  assign CLBLM_R_X11Y150_SLICE_X14Y150_D1 = CLBLM_R_X7Y146_SLICE_X8Y146_C5Q;
  assign CLBLM_R_X11Y150_SLICE_X14Y150_D2 = CLBLM_R_X11Y147_SLICE_X15Y147_BO6;
  assign CLBLM_R_X11Y150_SLICE_X14Y150_D3 = CLBLM_R_X7Y152_SLICE_X8Y152_DQ;
  assign CLBLM_R_X11Y150_SLICE_X14Y150_D4 = CLBLM_R_X11Y144_SLICE_X14Y144_BO6;
  assign CLBLL_L_X4Y153_SLICE_X5Y153_A1 = CLBLL_L_X2Y150_SLICE_X1Y150_AQ;
  assign CLBLL_L_X4Y153_SLICE_X5Y153_A2 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLL_L_X4Y153_SLICE_X5Y153_A3 = CLBLL_L_X4Y153_SLICE_X5Y153_AQ;
  assign CLBLL_L_X4Y153_SLICE_X5Y153_A4 = CLBLL_L_X4Y153_SLICE_X5Y153_BO6;
  assign CLBLL_L_X4Y153_SLICE_X5Y153_A5 = CLBLL_L_X4Y148_SLICE_X5Y148_AQ;
  assign CLBLL_L_X4Y153_SLICE_X5Y153_A6 = 1'b1;
  assign CLBLM_R_X11Y150_SLICE_X14Y150_D5 = CLBLM_R_X7Y144_SLICE_X9Y144_B5Q;
  assign CLBLM_R_X11Y150_SLICE_X14Y150_D6 = CLBLM_R_X7Y153_SLICE_X8Y153_A5Q;
  assign CLBLL_L_X4Y153_SLICE_X5Y153_AX = CLBLL_L_X4Y153_SLICE_X4Y153_DO6;
  assign CLBLL_L_X4Y153_SLICE_X5Y153_B1 = CLBLM_R_X3Y149_SLICE_X2Y149_AQ;
  assign CLBLL_L_X4Y153_SLICE_X5Y153_B2 = CLBLM_R_X3Y149_SLICE_X3Y149_AQ;
  assign CLBLL_L_X4Y153_SLICE_X5Y153_B3 = CLBLM_R_X7Y153_SLICE_X9Y153_AQ;
  assign CLBLL_L_X4Y153_SLICE_X5Y153_B4 = CLBLM_R_X5Y154_SLICE_X6Y154_BQ;
  assign CLBLL_L_X4Y153_SLICE_X5Y153_B5 = CLBLM_R_X5Y154_SLICE_X6Y154_AQ;
  assign CLBLL_L_X4Y153_SLICE_X5Y153_B6 = 1'b1;
  assign CLBLL_L_X4Y153_SLICE_X5Y153_C1 = 1'b1;
  assign CLBLL_L_X4Y153_SLICE_X5Y153_C2 = 1'b1;
  assign CLBLL_L_X4Y153_SLICE_X5Y153_C3 = 1'b1;
  assign CLBLL_L_X4Y153_SLICE_X5Y153_C4 = 1'b1;
  assign CLBLL_L_X4Y153_SLICE_X5Y153_C5 = 1'b1;
  assign CLBLL_L_X4Y153_SLICE_X5Y153_C6 = 1'b1;
  assign CLBLL_L_X4Y153_SLICE_X5Y153_CLK = CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O;
  assign CLBLM_R_X3Y144_SLICE_X3Y144_D1 = CLBLL_L_X2Y146_SLICE_X1Y146_B5Q;
  assign CLBLM_R_X3Y144_SLICE_X3Y144_D2 = CLBLM_R_X5Y143_SLICE_X6Y143_D5Q;
  assign CLBLL_L_X4Y153_SLICE_X5Y153_D1 = 1'b1;
  assign CLBLL_L_X4Y153_SLICE_X5Y153_D2 = 1'b1;
  assign CLBLL_L_X4Y153_SLICE_X5Y153_D3 = 1'b1;
  assign CLBLL_L_X4Y153_SLICE_X5Y153_D4 = 1'b1;
  assign CLBLL_L_X4Y153_SLICE_X5Y153_D5 = 1'b1;
  assign CLBLL_L_X4Y153_SLICE_X5Y153_D6 = 1'b1;
  assign CLBLM_R_X3Y144_SLICE_X3Y144_D5 = CLBLM_R_X3Y144_SLICE_X3Y144_AQ;
  assign CLBLM_L_X8Y147_SLICE_X11Y147_A1 = CLBLM_R_X3Y148_SLICE_X3Y148_AQ;
  assign CLBLM_L_X8Y147_SLICE_X11Y147_A2 = CLBLM_R_X11Y146_SLICE_X14Y146_DO6;
  assign CLBLM_L_X8Y147_SLICE_X11Y147_A3 = CLBLM_L_X8Y147_SLICE_X11Y147_AQ;
  assign CLBLM_L_X8Y147_SLICE_X11Y147_A4 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_L_X8Y147_SLICE_X11Y147_A5 = CLBLM_R_X5Y151_SLICE_X6Y151_AQ;
  assign CLBLM_L_X8Y147_SLICE_X11Y147_A6 = 1'b1;
  assign CLBLM_R_X3Y144_SLICE_X2Y144_A3 = CLBLM_R_X3Y144_SLICE_X2Y144_AQ;
  assign LIOB33_X0Y153_IOB_X0Y154_O = CLBLM_R_X7Y153_SLICE_X9Y153_DQ;
  assign CLBLM_L_X8Y147_SLICE_X11Y147_B1 = CLBLM_L_X8Y148_SLICE_X10Y148_B5Q;
  assign CLBLM_L_X8Y147_SLICE_X11Y147_B2 = CLBLM_L_X8Y147_SLICE_X11Y147_BQ;
  assign CLBLM_L_X8Y147_SLICE_X11Y147_B3 = CLBLM_R_X7Y142_SLICE_X8Y142_C5Q;
  assign CLBLM_L_X8Y147_SLICE_X11Y147_B4 = CLBLM_R_X5Y146_SLICE_X7Y146_BQ;
  assign CLBLM_L_X8Y147_SLICE_X11Y147_B5 = CLBLM_R_X7Y152_SLICE_X8Y152_D5Q;
  assign CLBLM_L_X8Y147_SLICE_X11Y147_B6 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X3Y144_SLICE_X2Y144_A4 = CLBLM_R_X3Y144_SLICE_X2Y144_BO6;
  assign CLBLM_R_X3Y144_SLICE_X2Y144_A5 = CLBLM_R_X3Y144_SLICE_X3Y144_AQ;
  assign LIOB33_X0Y153_IOB_X0Y153_O = CLBLM_L_X8Y153_SLICE_X10Y153_A5Q;
  assign CLBLM_L_X8Y147_SLICE_X11Y147_C1 = CLBLM_L_X10Y153_SLICE_X13Y153_A5Q;
  assign CLBLM_L_X8Y147_SLICE_X11Y147_C2 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_L_X8Y147_SLICE_X11Y147_C3 = 1'b1;
  assign CLBLM_L_X8Y147_SLICE_X11Y147_C4 = CLBLM_L_X8Y145_SLICE_X10Y145_AQ;
  assign CLBLM_L_X8Y147_SLICE_X11Y147_C5 = CLBLM_R_X7Y153_SLICE_X9Y153_A5Q;
  assign CLBLM_L_X8Y147_SLICE_X11Y147_C6 = 1'b1;
  assign CLBLM_R_X3Y144_SLICE_X2Y144_A6 = 1'b1;
  assign CLBLM_L_X8Y147_SLICE_X11Y147_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X8Y147_SLICE_X11Y147_D1 = CLBLM_L_X10Y146_SLICE_X12Y146_BQ;
  assign CLBLM_L_X8Y147_SLICE_X11Y147_D2 = 1'b1;
  assign CLBLM_L_X8Y147_SLICE_X11Y147_D3 = CLBLM_L_X8Y147_SLICE_X11Y147_DQ;
  assign CLBLM_L_X8Y147_SLICE_X11Y147_D4 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_L_X8Y147_SLICE_X11Y147_D5 = CLBLM_R_X11Y148_SLICE_X15Y148_AO6;
  assign CLBLM_L_X8Y147_SLICE_X11Y147_D6 = CLBLL_L_X4Y144_SLICE_X5Y144_D5Q;
  assign CLBLM_L_X8Y147_SLICE_X10Y147_A1 = 1'b1;
  assign CLBLM_L_X8Y147_SLICE_X10Y147_A2 = CLBLM_R_X7Y149_SLICE_X9Y149_BQ;
  assign CLBLM_L_X8Y147_SLICE_X10Y147_A3 = CLBLM_L_X8Y147_SLICE_X10Y147_AQ;
  assign CLBLM_L_X8Y147_SLICE_X10Y147_A4 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_L_X8Y147_SLICE_X10Y147_A5 = CLBLM_L_X8Y145_SLICE_X11Y145_AQ;
  assign CLBLM_L_X8Y147_SLICE_X10Y147_A6 = CLBLM_R_X13Y149_SLICE_X18Y149_AO6;
  assign CLBLM_L_X8Y147_SLICE_X10Y147_B1 = CLBLM_L_X8Y147_SLICE_X11Y147_DQ;
  assign CLBLM_L_X8Y147_SLICE_X10Y147_B2 = 1'b1;
  assign CLBLM_L_X8Y147_SLICE_X10Y147_B3 = 1'b1;
  assign CLBLM_L_X8Y147_SLICE_X10Y147_B4 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_L_X8Y147_SLICE_X10Y147_B5 = CLBLM_R_X5Y143_SLICE_X6Y143_BQ;
  assign CLBLM_L_X8Y147_SLICE_X10Y147_B6 = CLBLM_R_X3Y147_SLICE_X3Y147_DO6;
  assign CLBLM_L_X10Y153_SLICE_X13Y153_C1 = CLBLM_R_X5Y152_SLICE_X6Y152_DQ;
  assign CLBLM_L_X8Y147_SLICE_X10Y147_C1 = RIOB33_X105Y111_IOB_X1Y112_I;
  assign CLBLM_L_X8Y147_SLICE_X10Y147_C2 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_L_X8Y147_SLICE_X10Y147_C3 = 1'b1;
  assign CLBLM_L_X8Y147_SLICE_X10Y147_C4 = CLBLM_L_X10Y146_SLICE_X12Y146_CQ;
  assign CLBLM_L_X8Y147_SLICE_X10Y147_C5 = CLBLM_L_X8Y151_SLICE_X10Y151_B5Q;
  assign CLBLM_L_X8Y147_SLICE_X10Y147_C6 = 1'b1;
  assign CLBLM_R_X3Y144_SLICE_X2Y144_B6 = 1'b1;
  assign CLBLM_L_X8Y147_SLICE_X10Y147_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X8Y147_SLICE_X10Y147_D1 = CLBLM_R_X7Y146_SLICE_X8Y146_B5Q;
  assign CLBLM_L_X8Y147_SLICE_X10Y147_D2 = CLBLM_L_X8Y147_SLICE_X10Y147_AQ;
  assign CLBLM_L_X8Y147_SLICE_X10Y147_D3 = 1'b1;
  assign CLBLM_L_X8Y147_SLICE_X10Y147_D4 = CLBLM_R_X7Y148_SLICE_X8Y148_AO5;
  assign CLBLM_L_X8Y147_SLICE_X10Y147_D5 = CLBLM_L_X8Y150_SLICE_X11Y150_BO5;
  assign CLBLM_L_X8Y147_SLICE_X10Y147_D6 = CLBLM_L_X8Y144_SLICE_X10Y144_DO6;
  assign CLBLM_L_X10Y153_SLICE_X13Y153_CLK = CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O;
  assign CLBLM_R_X11Y151_SLICE_X15Y151_A1 = 1'b1;
  assign CLBLM_R_X11Y151_SLICE_X15Y151_A2 = CLBLM_R_X5Y149_SLICE_X7Y149_D5Q;
  assign CLBLM_R_X11Y151_SLICE_X15Y151_A3 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X11Y151_SLICE_X15Y151_A4 = CLBLM_L_X12Y151_SLICE_X16Y151_AQ;
  assign CLBLM_R_X11Y151_SLICE_X15Y151_A5 = CLBLM_R_X11Y151_SLICE_X14Y151_AQ;
  assign CLBLM_R_X11Y151_SLICE_X15Y151_A6 = 1'b1;
  assign CLBLM_R_X11Y151_SLICE_X15Y151_B1 = CLBLL_L_X4Y148_SLICE_X4Y148_CQ;
  assign CLBLM_R_X11Y151_SLICE_X15Y151_B2 = CLBLM_R_X7Y153_SLICE_X8Y153_A5Q;
  assign CLBLM_R_X11Y151_SLICE_X15Y151_B3 = CLBLM_L_X12Y147_SLICE_X16Y147_DO6;
  assign CLBLM_R_X11Y151_SLICE_X15Y151_B4 = CLBLM_R_X7Y144_SLICE_X9Y144_B5Q;
  assign CLBLM_R_X11Y151_SLICE_X15Y151_B5 = CLBLM_R_X7Y149_SLICE_X8Y149_AQ;
  assign CLBLM_R_X11Y151_SLICE_X15Y151_B6 = CLBLM_R_X7Y143_SLICE_X9Y143_BQ;
  assign CLBLM_L_X10Y153_SLICE_X13Y153_D3 = CLBLM_L_X10Y152_SLICE_X13Y152_AQ;
  assign CLBLM_R_X7Y141_SLICE_X9Y141_A1 = CLBLM_R_X7Y141_SLICE_X9Y141_AQ;
  assign CLBLM_R_X7Y141_SLICE_X9Y141_A2 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X7Y141_SLICE_X9Y141_A3 = CLBLM_R_X7Y141_SLICE_X8Y141_AO6;
  assign CLBLM_R_X7Y141_SLICE_X9Y141_A4 = CLBLM_R_X7Y144_SLICE_X9Y144_BQ;
  assign CLBLM_R_X7Y141_SLICE_X9Y141_A5 = CLBLM_L_X8Y142_SLICE_X10Y142_DO6;
  assign CLBLM_R_X7Y141_SLICE_X9Y141_A6 = CLBLL_L_X4Y151_SLICE_X4Y151_CQ;
  assign CLBLM_L_X10Y153_SLICE_X13Y153_D4 = CLBLM_L_X8Y152_SLICE_X10Y152_CQ;
  assign CLBLM_R_X11Y151_SLICE_X15Y151_C1 = 1'b1;
  assign CLBLM_R_X11Y151_SLICE_X15Y151_C2 = 1'b1;
  assign CLBLM_R_X7Y141_SLICE_X9Y141_B1 = 1'b1;
  assign CLBLM_R_X7Y141_SLICE_X9Y141_B2 = 1'b1;
  assign CLBLM_R_X7Y141_SLICE_X9Y141_B3 = 1'b1;
  assign CLBLM_R_X7Y141_SLICE_X9Y141_B4 = 1'b1;
  assign CLBLM_R_X7Y141_SLICE_X9Y141_B5 = 1'b1;
  assign CLBLM_R_X7Y141_SLICE_X9Y141_B6 = 1'b1;
  assign CLBLM_R_X11Y151_SLICE_X15Y151_CLK = CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O;
  assign CLBLM_R_X11Y151_SLICE_X15Y151_D1 = 1'b1;
  assign CLBLM_R_X7Y141_SLICE_X9Y141_C1 = 1'b1;
  assign CLBLM_R_X7Y141_SLICE_X9Y141_C2 = 1'b1;
  assign CLBLM_R_X7Y141_SLICE_X9Y141_C3 = 1'b1;
  assign CLBLM_R_X7Y141_SLICE_X9Y141_C4 = 1'b1;
  assign CLBLM_R_X7Y141_SLICE_X9Y141_C5 = 1'b1;
  assign CLBLM_R_X7Y141_SLICE_X9Y141_C6 = 1'b1;
  assign CLBLM_R_X11Y151_SLICE_X15Y151_D3 = 1'b1;
  assign CLBLM_R_X11Y151_SLICE_X15Y151_D4 = 1'b1;
  assign CLBLM_R_X7Y141_SLICE_X9Y141_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X11Y151_SLICE_X14Y151_A1 = CLBLM_R_X7Y144_SLICE_X9Y144_AQ;
  assign CLBLM_R_X11Y151_SLICE_X14Y151_A2 = CLBLM_L_X12Y149_SLICE_X17Y149_CO6;
  assign CLBLM_R_X11Y151_SLICE_X14Y151_A3 = CLBLM_R_X11Y151_SLICE_X14Y151_AQ;
  assign CLBLM_R_X11Y151_SLICE_X14Y151_A4 = 1'b1;
  assign CLBLM_R_X11Y151_SLICE_X14Y151_A5 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X7Y141_SLICE_X9Y141_D1 = 1'b1;
  assign CLBLM_R_X7Y141_SLICE_X9Y141_D2 = 1'b1;
  assign CLBLM_R_X7Y141_SLICE_X9Y141_D3 = 1'b1;
  assign CLBLM_R_X7Y141_SLICE_X9Y141_D4 = 1'b1;
  assign CLBLM_R_X7Y141_SLICE_X9Y141_D5 = 1'b1;
  assign CLBLM_R_X7Y141_SLICE_X9Y141_D6 = 1'b1;
  assign CLBLM_R_X11Y151_SLICE_X14Y151_A6 = CLBLM_R_X7Y153_SLICE_X9Y153_DQ;
  assign CLBLM_R_X11Y151_SLICE_X14Y151_B1 = CLBLM_R_X11Y144_SLICE_X14Y144_BO6;
  assign CLBLM_R_X11Y151_SLICE_X14Y151_B2 = CLBLM_R_X7Y153_SLICE_X8Y153_A5Q;
  assign CLBLM_R_X11Y151_SLICE_X14Y151_B3 = CLBLM_R_X11Y151_SLICE_X15Y151_A5Q;
  assign CLBLM_R_X11Y151_SLICE_X14Y151_B4 = CLBLM_R_X11Y147_SLICE_X15Y147_BO6;
  assign CLBLM_R_X7Y141_SLICE_X8Y141_A1 = CLBLM_L_X8Y145_SLICE_X11Y145_DQ;
  assign CLBLM_R_X7Y141_SLICE_X8Y141_A2 = RIOB33_X105Y131_IOB_X1Y131_I;
  assign CLBLM_R_X7Y141_SLICE_X8Y141_A3 = RIOB33_X105Y101_IOB_X1Y102_I;
  assign CLBLM_R_X7Y141_SLICE_X8Y141_A4 = CLBLM_L_X10Y147_SLICE_X12Y147_CO6;
  assign CLBLM_R_X7Y141_SLICE_X8Y141_A5 = CLBLM_R_X3Y151_SLICE_X2Y151_AQ;
  assign CLBLM_R_X7Y141_SLICE_X8Y141_A6 = 1'b1;
  assign CLBLM_R_X11Y151_SLICE_X14Y151_C2 = CLBLM_R_X7Y150_SLICE_X8Y150_CO6;
  assign CLBLM_R_X11Y151_SLICE_X14Y151_C3 = CLBLM_L_X8Y150_SLICE_X10Y150_BO6;
  assign CLBLM_R_X11Y151_SLICE_X14Y151_C4 = CLBLM_R_X3Y150_SLICE_X3Y150_D5Q;
  assign CLBLM_R_X11Y151_SLICE_X14Y151_C5 = CLBLL_L_X4Y150_SLICE_X4Y150_A5Q;
  assign CLBLM_R_X7Y141_SLICE_X8Y141_B1 = 1'b1;
  assign CLBLM_R_X7Y141_SLICE_X8Y141_B2 = CLBLM_R_X7Y145_SLICE_X8Y145_AQ;
  assign CLBLM_R_X7Y141_SLICE_X8Y141_B3 = CLBLM_R_X3Y151_SLICE_X2Y151_AQ;
  assign CLBLM_R_X7Y141_SLICE_X8Y141_B4 = CLBLM_L_X10Y147_SLICE_X12Y147_CO6;
  assign CLBLM_R_X7Y141_SLICE_X8Y141_B5 = 1'b1;
  assign CLBLM_R_X7Y141_SLICE_X8Y141_B6 = RIOB33_SING_X105Y100_IOB_X1Y100_I;
  assign CLBLM_R_X11Y151_SLICE_X14Y151_CLK = CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O;
  assign CLBLM_R_X11Y151_SLICE_X14Y151_D1 = CLBLM_L_X10Y148_SLICE_X12Y148_AO6;
  assign CLBLM_R_X11Y151_SLICE_X14Y151_D2 = CLBLM_R_X3Y150_SLICE_X3Y150_D5Q;
  assign CLBLM_R_X7Y141_SLICE_X8Y141_C1 = 1'b1;
  assign CLBLM_R_X7Y141_SLICE_X8Y141_C2 = 1'b1;
  assign CLBLM_R_X7Y141_SLICE_X8Y141_C3 = 1'b1;
  assign CLBLM_R_X7Y141_SLICE_X8Y141_C4 = 1'b1;
  assign CLBLM_R_X7Y141_SLICE_X8Y141_C5 = 1'b1;
  assign CLBLM_R_X7Y141_SLICE_X8Y141_C6 = 1'b1;
  assign CLBLM_R_X11Y151_SLICE_X14Y151_D3 = CLBLL_L_X4Y150_SLICE_X4Y150_A5Q;
  assign CLBLM_R_X11Y151_SLICE_X14Y151_D4 = CLBLM_L_X8Y150_SLICE_X10Y150_BO6;
  assign CLBLM_R_X11Y151_SLICE_X14Y151_D5 = 1'b1;
  assign CLBLM_L_X10Y153_SLICE_X12Y153_A6 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X11Y151_SLICE_X14Y151_D6 = CLBLM_L_X10Y151_SLICE_X13Y151_DO6;
  assign CLBLM_R_X7Y141_SLICE_X8Y141_D1 = 1'b1;
  assign CLBLM_R_X7Y141_SLICE_X8Y141_D2 = 1'b1;
  assign CLBLM_R_X7Y141_SLICE_X8Y141_D3 = 1'b1;
  assign CLBLM_R_X7Y141_SLICE_X8Y141_D4 = 1'b1;
  assign CLBLM_R_X7Y141_SLICE_X8Y141_D5 = 1'b1;
  assign CLBLM_R_X7Y141_SLICE_X8Y141_D6 = 1'b1;
  assign CLBLM_L_X10Y153_SLICE_X12Y153_B1 = CLBLM_R_X7Y154_SLICE_X8Y154_DO6;
  assign LIOI3_X0Y159_OLOGIC_X0Y160_D1 = CLBLL_L_X2Y148_SLICE_X0Y148_AQ;
  assign LIOI3_X0Y159_OLOGIC_X0Y160_T1 = 1'b1;
  assign LIOI3_X0Y159_OLOGIC_X0Y159_D1 = CLBLL_L_X2Y146_SLICE_X0Y146_CQ;
  assign LIOI3_X0Y159_OLOGIC_X0Y159_T1 = 1'b1;
  assign LIOB33_X0Y155_IOB_X0Y156_O = CLBLM_R_X3Y152_SLICE_X3Y152_CQ;
  assign LIOB33_X0Y155_IOB_X0Y155_O = CLBLM_R_X5Y154_SLICE_X7Y154_AQ;
  assign CLBLM_L_X10Y153_SLICE_X12Y153_C1 = CLBLM_L_X10Y147_SLICE_X12Y147_AQ;
  assign CLBLM_L_X8Y148_SLICE_X11Y148_A1 = CLBLM_R_X7Y151_SLICE_X9Y151_A5Q;
  assign CLBLM_L_X8Y148_SLICE_X11Y148_A2 = CLBLM_R_X7Y147_SLICE_X9Y147_D5Q;
  assign CLBLM_L_X8Y148_SLICE_X11Y148_A3 = CLBLM_L_X8Y148_SLICE_X11Y148_AQ;
  assign CLBLM_L_X8Y148_SLICE_X11Y148_A4 = RIOB33_X105Y111_IOB_X1Y112_I;
  assign CLBLM_L_X8Y148_SLICE_X11Y148_A5 = CLBLM_L_X8Y147_SLICE_X10Y147_CQ;
  assign CLBLM_L_X8Y148_SLICE_X11Y148_A6 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_L_X8Y148_SLICE_X11Y148_B1 = CLBLM_R_X5Y153_SLICE_X6Y153_A5Q;
  assign CLBLM_L_X8Y148_SLICE_X11Y148_B2 = CLBLL_L_X4Y149_SLICE_X5Y149_C5Q;
  assign CLBLM_L_X8Y148_SLICE_X11Y148_B3 = CLBLM_L_X8Y147_SLICE_X11Y147_BQ;
  assign CLBLM_L_X8Y148_SLICE_X11Y148_B4 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_L_X8Y148_SLICE_X11Y148_B5 = CLBLM_L_X8Y145_SLICE_X11Y145_BQ;
  assign CLBLM_L_X8Y148_SLICE_X11Y148_B6 = 1'b1;
  assign CLBLM_L_X10Y153_SLICE_X12Y153_C4 = CLBLM_R_X5Y150_SLICE_X6Y150_B5Q;
  assign RIOI3_TBYTESRC_X105Y193_OLOGIC_X1Y194_D1 = CLBLM_L_X12Y151_SLICE_X16Y151_BO6;
  assign CLBLM_L_X8Y148_SLICE_X11Y148_C1 = CLBLM_R_X5Y149_SLICE_X6Y149_BQ;
  assign CLBLM_L_X8Y148_SLICE_X11Y148_C2 = CLBLM_L_X8Y147_SLICE_X11Y147_DQ;
  assign CLBLM_L_X8Y148_SLICE_X11Y148_C3 = CLBLM_L_X12Y149_SLICE_X17Y149_BO5;
  assign CLBLM_L_X8Y148_SLICE_X11Y148_C4 = CLBLM_L_X10Y151_SLICE_X13Y151_BO6;
  assign CLBLM_L_X8Y148_SLICE_X11Y148_C5 = CLBLM_R_X7Y143_SLICE_X8Y143_BQ;
  assign CLBLM_L_X8Y148_SLICE_X11Y148_C6 = CLBLM_L_X10Y148_SLICE_X12Y148_AO6;
  assign CLBLM_L_X8Y148_SLICE_X11Y148_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign RIOI3_TBYTESRC_X105Y193_OLOGIC_X1Y194_T1 = 1'b1;
  assign CLBLM_L_X8Y148_SLICE_X11Y148_D1 = 1'b1;
  assign CLBLM_L_X8Y148_SLICE_X11Y148_D2 = CLBLM_L_X10Y148_SLICE_X12Y148_BO6;
  assign CLBLM_L_X8Y148_SLICE_X11Y148_D3 = CLBLM_L_X8Y148_SLICE_X11Y148_BQ;
  assign CLBLM_L_X8Y148_SLICE_X11Y148_D4 = CLBLM_R_X7Y148_SLICE_X8Y148_AO5;
  assign CLBLM_L_X8Y148_SLICE_X11Y148_D5 = CLBLM_L_X8Y144_SLICE_X11Y144_CQ;
  assign CLBLM_L_X8Y148_SLICE_X11Y148_D6 = CLBLM_L_X8Y150_SLICE_X11Y150_BO6;
  assign CLBLM_L_X10Y153_SLICE_X12Y153_CLK = CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O;
  assign RIOI3_TBYTESRC_X105Y193_OLOGIC_X1Y193_D1 = CLBLM_L_X12Y151_SLICE_X16Y151_BO5;
  assign CLBLM_L_X8Y148_SLICE_X10Y148_A1 = CLBLM_L_X10Y146_SLICE_X12Y146_CQ;
  assign CLBLM_L_X8Y148_SLICE_X10Y148_A2 = CLBLM_R_X13Y149_SLICE_X18Y149_AO6;
  assign CLBLM_L_X8Y148_SLICE_X10Y148_A3 = CLBLM_L_X8Y148_SLICE_X10Y148_AQ;
  assign CLBLM_L_X8Y148_SLICE_X10Y148_A4 = 1'b1;
  assign CLBLM_L_X8Y148_SLICE_X10Y148_A5 = CLBLL_L_X2Y148_SLICE_X0Y148_AQ;
  assign CLBLM_L_X8Y148_SLICE_X10Y148_A6 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign RIOI3_TBYTESRC_X105Y193_OLOGIC_X1Y193_T1 = 1'b1;
  assign CLBLM_L_X8Y148_SLICE_X10Y148_B1 = CLBLM_R_X7Y148_SLICE_X9Y148_CQ;
  assign CLBLM_L_X8Y148_SLICE_X10Y148_B2 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_L_X8Y148_SLICE_X10Y148_B3 = CLBLM_L_X8Y147_SLICE_X10Y147_CQ;
  assign CLBLM_L_X8Y148_SLICE_X10Y148_B4 = CLBLM_R_X5Y152_SLICE_X6Y152_CQ;
  assign CLBLM_L_X8Y148_SLICE_X10Y148_B5 = CLBLM_R_X5Y146_SLICE_X6Y146_B5Q;
  assign CLBLM_L_X8Y148_SLICE_X10Y148_B6 = 1'b1;
  assign CLBLM_L_X8Y148_SLICE_X10Y148_C1 = CLBLM_R_X7Y148_SLICE_X9Y148_DO6;
  assign CLBLM_L_X8Y148_SLICE_X10Y148_C2 = CLBLM_L_X12Y146_SLICE_X16Y146_CO6;
  assign CLBLM_L_X8Y148_SLICE_X10Y148_C3 = CLBLL_L_X4Y148_SLICE_X4Y148_CQ;
  assign CLBLM_L_X8Y148_SLICE_X10Y148_C4 = CLBLM_R_X3Y146_SLICE_X2Y146_D5Q;
  assign CLBLM_L_X8Y148_SLICE_X10Y148_C5 = CLBLM_R_X3Y149_SLICE_X3Y149_DQ;
  assign CLBLM_L_X8Y148_SLICE_X10Y148_C6 = CLBLM_L_X8Y146_SLICE_X10Y146_AO5;
  assign CLBLM_L_X8Y148_SLICE_X10Y148_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X8Y148_SLICE_X10Y148_D1 = CLBLM_R_X5Y151_SLICE_X6Y151_AQ;
  assign CLBLM_L_X8Y148_SLICE_X10Y148_D2 = CLBLM_R_X7Y148_SLICE_X8Y148_AO5;
  assign CLBLM_L_X8Y148_SLICE_X10Y148_D3 = CLBLM_L_X8Y153_SLICE_X10Y153_DQ;
  assign CLBLM_L_X8Y148_SLICE_X10Y148_D4 = CLBLM_R_X7Y148_SLICE_X8Y148_AO6;
  assign CLBLM_L_X8Y148_SLICE_X10Y148_D5 = CLBLM_L_X8Y153_SLICE_X10Y153_D5Q;
  assign CLBLM_L_X8Y148_SLICE_X10Y148_D6 = CLBLM_L_X8Y150_SLICE_X11Y150_BO6;
  assign CLBLM_L_X10Y153_SLICE_X12Y153_D3 = RIOB33_X105Y131_IOB_X1Y131_I;
  assign CLBLM_L_X10Y153_SLICE_X12Y153_D4 = CLBLL_L_X4Y153_SLICE_X5Y153_A5Q;
  assign CLBLM_L_X10Y153_SLICE_X12Y153_D6 = CLBLM_R_X7Y145_SLICE_X8Y145_A5Q;
  assign CLBLM_R_X11Y152_SLICE_X15Y152_A1 = CLBLM_R_X11Y152_SLICE_X15Y152_CQ;
  assign CLBLM_R_X11Y152_SLICE_X15Y152_A2 = CLBLM_R_X11Y152_SLICE_X15Y152_BQ;
  assign CLBLM_R_X11Y152_SLICE_X15Y152_A3 = CLBLM_R_X11Y152_SLICE_X15Y152_A5Q;
  assign CLBLM_R_X11Y152_SLICE_X15Y152_A4 = CLBLM_L_X10Y151_SLICE_X13Y151_CO6;
  assign CLBLM_R_X11Y152_SLICE_X15Y152_A5 = CLBLM_R_X11Y152_SLICE_X15Y152_B5Q;
  assign CLBLM_R_X11Y152_SLICE_X15Y152_A6 = 1'b1;
  assign CLBLM_R_X11Y152_SLICE_X15Y152_B1 = CLBLM_R_X11Y152_SLICE_X15Y152_CQ;
  assign CLBLM_R_X11Y152_SLICE_X15Y152_B2 = CLBLM_R_X11Y152_SLICE_X15Y152_BQ;
  assign CLBLM_R_X11Y152_SLICE_X15Y152_B3 = CLBLM_R_X11Y152_SLICE_X15Y152_A5Q;
  assign CLBLM_R_X11Y152_SLICE_X15Y152_B4 = CLBLM_L_X10Y151_SLICE_X13Y151_CO6;
  assign CLBLM_R_X11Y152_SLICE_X15Y152_B5 = CLBLM_R_X11Y152_SLICE_X15Y152_B5Q;
  assign CLBLM_R_X11Y152_SLICE_X15Y152_B6 = 1'b1;
  assign CLBLM_R_X7Y142_SLICE_X9Y142_A1 = CLBLL_L_X4Y151_SLICE_X4Y151_BQ;
  assign CLBLM_R_X7Y142_SLICE_X9Y142_A2 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X7Y142_SLICE_X9Y142_A3 = CLBLM_R_X7Y142_SLICE_X9Y142_AQ;
  assign CLBLM_R_X7Y142_SLICE_X9Y142_A4 = CLBLL_L_X4Y143_SLICE_X5Y143_D5Q;
  assign CLBLM_R_X7Y142_SLICE_X9Y142_A5 = CLBLM_R_X3Y145_SLICE_X3Y145_D5Q;
  assign CLBLM_R_X7Y142_SLICE_X9Y142_A6 = CLBLM_R_X5Y145_SLICE_X6Y145_D5Q;
  assign CLBLM_R_X11Y152_SLICE_X15Y152_C1 = 1'b1;
  assign CLBLM_R_X11Y152_SLICE_X15Y152_C2 = CLBLM_R_X11Y152_SLICE_X15Y152_CQ;
  assign CLBLM_R_X11Y149_SLICE_X15Y149_D4 = CLBLM_R_X7Y148_SLICE_X8Y148_CO6;
  assign CLBLM_R_X7Y142_SLICE_X9Y142_B1 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X7Y142_SLICE_X9Y142_B2 = CLBLM_R_X7Y142_SLICE_X9Y142_BQ;
  assign CLBLM_R_X7Y142_SLICE_X9Y142_B3 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X7Y142_SLICE_X9Y142_B4 = CLBLM_R_X7Y146_SLICE_X8Y146_BQ;
  assign CLBLM_R_X7Y142_SLICE_X9Y142_B5 = 1'b1;
  assign CLBLM_R_X7Y142_SLICE_X9Y142_B6 = CLBLL_L_X4Y152_SLICE_X4Y152_B5Q;
  assign CLBLM_R_X11Y149_SLICE_X15Y149_D5 = CLBLM_R_X11Y150_SLICE_X14Y150_AO6;
  assign CLBLM_R_X11Y152_SLICE_X15Y152_CLK = CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O;
  assign CLBLM_R_X11Y149_SLICE_X15Y149_D6 = CLBLM_L_X8Y149_SLICE_X10Y149_AO6;
  assign CLBLM_R_X7Y142_SLICE_X9Y142_C1 = CLBLM_L_X10Y147_SLICE_X12Y147_CO6;
  assign CLBLM_R_X7Y142_SLICE_X9Y142_C2 = 1'b1;
  assign CLBLM_R_X7Y142_SLICE_X9Y142_C3 = CLBLM_R_X7Y145_SLICE_X8Y145_CQ;
  assign CLBLM_R_X7Y142_SLICE_X9Y142_C4 = 1'b1;
  assign CLBLM_R_X7Y142_SLICE_X9Y142_C5 = CLBLM_R_X7Y142_SLICE_X9Y142_DO6;
  assign CLBLM_R_X7Y142_SLICE_X9Y142_C6 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X11Y152_SLICE_X15Y152_D3 = 1'b1;
  assign CLBLM_R_X11Y152_SLICE_X15Y152_D4 = 1'b1;
  assign CLBLM_R_X7Y142_SLICE_X9Y142_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X11Y152_SLICE_X14Y152_A1 = CLBLM_L_X10Y153_SLICE_X13Y153_CQ;
  assign CLBLM_R_X11Y152_SLICE_X14Y152_A2 = CLBLM_L_X8Y152_SLICE_X10Y152_CQ;
  assign CLBLM_R_X11Y152_SLICE_X14Y152_A3 = CLBLM_R_X7Y146_SLICE_X8Y146_A5Q;
  assign CLBLM_R_X11Y152_SLICE_X14Y152_A4 = CLBLM_L_X10Y152_SLICE_X12Y152_AQ;
  assign CLBLM_R_X7Y142_SLICE_X9Y142_D1 = CLBLM_R_X3Y151_SLICE_X2Y151_AQ;
  assign CLBLM_R_X7Y142_SLICE_X9Y142_D2 = CLBLM_R_X7Y145_SLICE_X8Y145_AQ;
  assign CLBLM_R_X7Y142_SLICE_X9Y142_D3 = RIOB33_SING_X105Y100_IOB_X1Y100_I;
  assign CLBLM_R_X7Y142_SLICE_X9Y142_D4 = RIOB33_X105Y131_IOB_X1Y131_I;
  assign CLBLM_R_X7Y142_SLICE_X9Y142_D5 = 1'b1;
  assign CLBLM_R_X7Y142_SLICE_X9Y142_D6 = RIOB33_X105Y101_IOB_X1Y101_I;
  assign CLBLM_R_X11Y152_SLICE_X14Y152_A5 = CLBLM_R_X11Y153_SLICE_X14Y153_AQ;
  assign CLBLM_R_X11Y152_SLICE_X14Y152_A6 = CLBLM_R_X5Y147_SLICE_X6Y147_AQ;
  assign CLBLM_R_X11Y152_SLICE_X14Y152_B1 = 1'b1;
  assign CLBLM_R_X11Y152_SLICE_X14Y152_B2 = 1'b1;
  assign CLBLM_R_X11Y152_SLICE_X14Y152_B3 = 1'b1;
  assign CLBLM_R_X7Y142_SLICE_X8Y142_A1 = CLBLM_L_X8Y147_SLICE_X10Y147_C5Q;
  assign CLBLM_R_X7Y142_SLICE_X8Y142_A2 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X7Y142_SLICE_X8Y142_A3 = CLBLM_R_X7Y142_SLICE_X8Y142_AQ;
  assign CLBLM_R_X7Y142_SLICE_X8Y142_A4 = CLBLM_L_X10Y144_SLICE_X13Y144_CQ;
  assign CLBLM_R_X7Y142_SLICE_X8Y142_A5 = CLBLM_R_X5Y150_SLICE_X6Y150_AQ;
  assign CLBLM_R_X7Y142_SLICE_X8Y142_A6 = CLBLM_L_X8Y142_SLICE_X10Y142_BQ;
  assign CLBLM_R_X11Y152_SLICE_X14Y152_C1 = 1'b1;
  assign CLBLM_R_X11Y152_SLICE_X14Y152_C2 = 1'b1;
  assign CLBLM_R_X11Y152_SLICE_X14Y152_C3 = 1'b1;
  assign CLBLM_R_X7Y142_SLICE_X8Y142_B1 = 1'b1;
  assign CLBLM_R_X7Y142_SLICE_X8Y142_B2 = CLBLM_R_X7Y142_SLICE_X8Y142_BQ;
  assign CLBLM_R_X7Y142_SLICE_X8Y142_B3 = CLBLM_R_X7Y142_SLICE_X8Y142_AQ;
  assign CLBLM_R_X7Y142_SLICE_X8Y142_B4 = CLBLM_R_X13Y149_SLICE_X18Y149_AO6;
  assign CLBLM_R_X7Y142_SLICE_X8Y142_B5 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X7Y142_SLICE_X8Y142_B6 = CLBLM_R_X5Y143_SLICE_X6Y143_DQ;
  assign CLBLM_R_X11Y152_SLICE_X14Y152_D1 = 1'b1;
  assign CLBLM_R_X11Y152_SLICE_X14Y152_D2 = 1'b1;
  assign CLBLM_R_X11Y152_SLICE_X14Y152_D3 = 1'b1;
  assign CLBLM_R_X7Y142_SLICE_X8Y142_C1 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X7Y142_SLICE_X8Y142_C2 = CLBLM_R_X7Y152_SLICE_X8Y152_D5Q;
  assign CLBLM_R_X7Y142_SLICE_X8Y142_C3 = 1'b1;
  assign CLBLM_R_X7Y142_SLICE_X8Y142_C4 = CLBLM_R_X5Y145_SLICE_X6Y145_D5Q;
  assign CLBLM_R_X7Y142_SLICE_X8Y142_C5 = CLBLL_L_X4Y142_SLICE_X4Y142_A5Q;
  assign CLBLM_R_X7Y142_SLICE_X8Y142_C6 = 1'b1;
  assign CLBLM_R_X11Y152_SLICE_X14Y152_D4 = 1'b1;
  assign CLBLM_R_X11Y152_SLICE_X14Y152_D5 = 1'b1;
  assign CLBLM_R_X11Y152_SLICE_X14Y152_D6 = 1'b1;
  assign CLBLM_R_X7Y142_SLICE_X8Y142_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign LIOI3_X0Y155_OLOGIC_X0Y155_T1 = 1'b1;
  assign CLBLM_R_X7Y142_SLICE_X8Y142_D1 = CLBLM_R_X5Y147_SLICE_X7Y147_C5Q;
  assign CLBLM_R_X7Y142_SLICE_X8Y142_D2 = CLBLM_R_X7Y142_SLICE_X8Y142_CQ;
  assign CLBLM_R_X7Y142_SLICE_X8Y142_D3 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X7Y142_SLICE_X8Y142_D4 = CLBLL_L_X4Y149_SLICE_X5Y149_C5Q;
  assign CLBLM_R_X7Y142_SLICE_X8Y142_D5 = 1'b1;
  assign CLBLM_R_X7Y142_SLICE_X8Y142_D6 = 1'b1;
  assign CLBLM_R_X7Y151_SLICE_X9Y151_C1 = CLBLM_R_X7Y151_SLICE_X8Y151_AQ;
  assign CLBLM_R_X7Y151_SLICE_X9Y151_C2 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X7Y151_SLICE_X9Y151_C3 = CLBLM_R_X11Y151_SLICE_X15Y151_AQ;
  assign CLBLM_R_X7Y151_SLICE_X9Y151_C4 = CLBLM_R_X3Y150_SLICE_X3Y150_D5Q;
  assign CLBLM_R_X7Y151_SLICE_X9Y151_C5 = 1'b1;
  assign CLBLM_R_X11Y149_SLICE_X14Y149_B1 = CLBLM_R_X7Y150_SLICE_X9Y150_DO6;
  assign LIOB33_X0Y157_IOB_X0Y158_O = RIOB33_X105Y133_IOB_X1Y134_I;
  assign LIOB33_X0Y157_IOB_X0Y157_O = CLBLM_R_X3Y152_SLICE_X3Y152_BQ;
  assign CLBLM_R_X7Y151_SLICE_X9Y151_C6 = 1'b1;
  assign CLBLM_R_X11Y149_SLICE_X14Y149_B2 = CLBLM_L_X8Y149_SLICE_X11Y149_CO6;
  assign CLBLM_R_X7Y151_SLICE_X9Y151_CLK = CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O;
  assign CLBLM_R_X7Y151_SLICE_X9Y151_D1 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_L_X8Y149_SLICE_X11Y149_A1 = CLBLM_R_X7Y149_SLICE_X9Y149_B5Q;
  assign CLBLM_L_X8Y149_SLICE_X11Y149_A2 = RIOB33_SING_X105Y100_IOB_X1Y100_I;
  assign CLBLM_L_X8Y149_SLICE_X11Y149_A3 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_L_X8Y149_SLICE_X11Y149_A4 = CLBLM_L_X8Y146_SLICE_X11Y146_CQ;
  assign CLBLM_L_X8Y149_SLICE_X11Y149_A5 = CLBLL_L_X4Y148_SLICE_X4Y148_BQ;
  assign CLBLM_L_X8Y149_SLICE_X11Y149_A6 = 1'b1;
  assign CLBLM_R_X7Y151_SLICE_X9Y151_D2 = CLBLL_L_X4Y151_SLICE_X4Y151_AQ;
  assign CLBLM_L_X8Y149_SLICE_X11Y149_B1 = CLBLM_L_X8Y145_SLICE_X10Y145_DO6;
  assign CLBLM_L_X8Y149_SLICE_X11Y149_B2 = CLBLM_L_X8Y148_SLICE_X11Y148_DO6;
  assign CLBLM_L_X8Y149_SLICE_X11Y149_B3 = CLBLM_R_X11Y147_SLICE_X15Y147_DO6;
  assign CLBLM_L_X8Y149_SLICE_X11Y149_B4 = CLBLM_L_X8Y150_SLICE_X11Y150_CO6;
  assign CLBLM_L_X8Y149_SLICE_X11Y149_B5 = CLBLM_L_X8Y151_SLICE_X11Y151_DO6;
  assign CLBLM_L_X8Y149_SLICE_X11Y149_B6 = CLBLM_L_X12Y147_SLICE_X16Y147_DO6;
  assign CLBLM_R_X7Y151_SLICE_X9Y151_D3 = CLBLM_L_X10Y153_SLICE_X12Y153_AQ;
  assign CLBLM_R_X7Y151_SLICE_X9Y151_D4 = CLBLL_L_X2Y146_SLICE_X0Y146_DQ;
  assign CLBLM_L_X8Y149_SLICE_X11Y149_C1 = CLBLM_R_X5Y148_SLICE_X6Y148_AQ;
  assign CLBLM_L_X8Y149_SLICE_X11Y149_C2 = CLBLM_L_X8Y149_SLICE_X10Y149_CO6;
  assign CLBLM_L_X8Y149_SLICE_X11Y149_C3 = CLBLM_L_X10Y151_SLICE_X12Y151_CQ;
  assign CLBLM_L_X8Y149_SLICE_X11Y149_C4 = CLBLM_L_X10Y151_SLICE_X13Y151_BO5;
  assign CLBLM_L_X8Y149_SLICE_X11Y149_C5 = 1'b1;
  assign CLBLM_L_X8Y149_SLICE_X11Y149_C6 = CLBLM_L_X10Y151_SLICE_X13Y151_BO6;
  assign CLBLM_R_X7Y151_SLICE_X9Y151_D5 = CLBLM_R_X7Y149_SLICE_X9Y149_C5Q;
  assign CLBLM_R_X7Y151_SLICE_X9Y151_D6 = 1'b1;
  assign CLBLM_L_X8Y149_SLICE_X11Y149_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X8Y149_SLICE_X11Y149_D1 = CLBLM_L_X8Y143_SLICE_X10Y143_CQ;
  assign CLBLM_L_X8Y149_SLICE_X11Y149_D2 = 1'b1;
  assign CLBLM_L_X8Y149_SLICE_X11Y149_D3 = CLBLM_L_X8Y151_SLICE_X10Y151_DO6;
  assign CLBLM_L_X8Y149_SLICE_X11Y149_D4 = CLBLM_L_X8Y144_SLICE_X11Y144_DQ;
  assign CLBLM_L_X8Y149_SLICE_X11Y149_D5 = CLBLM_L_X12Y149_SLICE_X17Y149_BO5;
  assign CLBLM_L_X8Y149_SLICE_X11Y149_D6 = CLBLM_R_X11Y148_SLICE_X15Y148_AO6;
  assign CLBLM_L_X8Y149_SLICE_X10Y149_A1 = CLBLL_L_X4Y146_SLICE_X4Y146_CQ;
  assign CLBLM_L_X8Y149_SLICE_X10Y149_A2 = CLBLM_R_X5Y149_SLICE_X6Y149_C5Q;
  assign CLBLM_L_X8Y149_SLICE_X10Y149_A3 = CLBLM_L_X8Y150_SLICE_X10Y150_BO5;
  assign CLBLM_L_X8Y149_SLICE_X10Y149_A4 = CLBLM_L_X8Y149_SLICE_X10Y149_BO6;
  assign CLBLM_L_X8Y149_SLICE_X10Y149_A5 = CLBLL_L_X4Y143_SLICE_X5Y143_AQ;
  assign CLBLM_L_X8Y149_SLICE_X10Y149_A6 = CLBLM_L_X10Y150_SLICE_X12Y150_BO6;
  assign CLBLM_L_X8Y149_SLICE_X10Y149_AX = CLBLM_R_X5Y149_SLICE_X6Y149_BQ;
  assign CLBLM_L_X8Y149_SLICE_X10Y149_B1 = CLBLM_R_X7Y144_SLICE_X9Y144_B5Q;
  assign CLBLM_L_X8Y149_SLICE_X10Y149_B2 = CLBLM_R_X7Y153_SLICE_X8Y153_A5Q;
  assign CLBLM_L_X8Y149_SLICE_X10Y149_B3 = CLBLM_L_X12Y147_SLICE_X16Y147_DO6;
  assign CLBLM_L_X8Y149_SLICE_X10Y149_B4 = CLBLM_R_X7Y149_SLICE_X8Y149_AQ;
  assign CLBLM_L_X8Y149_SLICE_X10Y149_B5 = CLBLM_L_X10Y146_SLICE_X13Y146_DO6;
  assign CLBLM_L_X8Y149_SLICE_X10Y149_B6 = CLBLL_L_X4Y148_SLICE_X4Y148_CQ;
  assign CLBLM_L_X8Y149_SLICE_X10Y149_C1 = CLBLM_R_X11Y144_SLICE_X14Y144_BO6;
  assign CLBLM_L_X8Y149_SLICE_X10Y149_C2 = CLBLM_R_X7Y144_SLICE_X9Y144_B5Q;
  assign CLBLM_L_X8Y149_SLICE_X10Y149_C3 = CLBLM_R_X7Y153_SLICE_X8Y153_A5Q;
  assign CLBLM_L_X8Y149_SLICE_X10Y149_C4 = CLBLM_R_X5Y145_SLICE_X7Y145_A5Q;
  assign CLBLM_L_X8Y149_SLICE_X10Y149_C5 = CLBLM_R_X11Y147_SLICE_X15Y147_BO6;
  assign CLBLM_L_X8Y149_SLICE_X10Y149_C6 = CLBLM_R_X7Y151_SLICE_X8Y151_C5Q;
  assign CLBLM_L_X8Y149_SLICE_X10Y149_CE = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X7Y151_SLICE_X8Y151_A2 = CLBLM_R_X13Y149_SLICE_X18Y149_AO6;
  assign CLBLM_R_X7Y151_SLICE_X8Y151_A3 = CLBLM_R_X7Y151_SLICE_X8Y151_AQ;
  assign CLBLM_L_X8Y149_SLICE_X10Y149_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X7Y151_SLICE_X8Y151_A4 = CLBLM_R_X5Y144_SLICE_X7Y144_AQ;
  assign CLBLM_R_X7Y151_SLICE_X8Y151_A5 = 1'b1;
  assign CLBLM_L_X8Y149_SLICE_X10Y149_D1 = CLBLM_L_X8Y148_SLICE_X10Y148_AQ;
  assign CLBLM_L_X8Y149_SLICE_X10Y149_D2 = 1'b1;
  assign CLBLM_L_X8Y149_SLICE_X10Y149_D3 = CLBLL_L_X4Y150_SLICE_X4Y150_AQ;
  assign CLBLM_L_X8Y149_SLICE_X10Y149_D4 = CLBLM_L_X8Y150_SLICE_X10Y150_BO5;
  assign CLBLM_L_X8Y149_SLICE_X10Y149_D5 = CLBLM_L_X8Y150_SLICE_X11Y150_BO6;
  assign CLBLM_L_X8Y149_SLICE_X10Y149_D6 = CLBLM_R_X7Y149_SLICE_X9Y149_DO6;
  assign CLBLM_R_X7Y151_SLICE_X8Y151_A6 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X7Y151_SLICE_X8Y151_B1 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X7Y151_SLICE_X8Y151_B2 = CLBLM_R_X7Y151_SLICE_X8Y151_BQ;
  assign CLBLM_R_X11Y153_SLICE_X15Y153_A1 = CLBLM_R_X11Y153_SLICE_X14Y153_A5Q;
  assign CLBLM_R_X11Y153_SLICE_X15Y153_A2 = CLBLM_R_X11Y153_SLICE_X14Y153_BO6;
  assign CLBLM_R_X11Y153_SLICE_X15Y153_A3 = CLBLM_R_X11Y153_SLICE_X15Y153_AQ;
  assign CLBLM_R_X11Y153_SLICE_X15Y153_A4 = CLBLM_L_X8Y148_SLICE_X11Y148_B5Q;
  assign CLBLM_R_X7Y151_SLICE_X8Y151_B3 = CLBLM_R_X5Y151_SLICE_X6Y151_C5Q;
  assign CLBLM_R_X11Y153_SLICE_X15Y153_A5 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X11Y153_SLICE_X15Y153_A6 = CLBLM_R_X11Y153_SLICE_X15Y153_CO6;
  assign CLBLM_R_X7Y151_SLICE_X8Y151_B4 = CLBLM_R_X3Y145_SLICE_X3Y145_D5Q;
  assign CLBLM_R_X11Y153_SLICE_X15Y153_B1 = CLBLM_R_X11Y153_SLICE_X14Y153_A5Q;
  assign CLBLM_R_X11Y153_SLICE_X15Y153_B2 = CLBLM_R_X11Y153_SLICE_X14Y153_DO6;
  assign CLBLM_R_X11Y153_SLICE_X15Y153_B3 = CLBLM_L_X10Y153_SLICE_X13Y153_CQ;
  assign CLBLM_R_X11Y153_SLICE_X15Y153_B4 = CLBLM_R_X5Y147_SLICE_X6Y147_AQ;
  assign CLBLM_R_X7Y151_SLICE_X8Y151_B5 = CLBLL_L_X4Y150_SLICE_X5Y150_AQ;
  assign CLBLM_R_X11Y153_SLICE_X15Y153_B5 = CLBLM_R_X7Y146_SLICE_X8Y146_A5Q;
  assign CLBLM_R_X11Y153_SLICE_X15Y153_B6 = 1'b1;
  assign CLBLM_R_X7Y151_SLICE_X8Y151_B6 = CLBLL_L_X4Y151_SLICE_X4Y151_BQ;
  assign CLBLM_R_X7Y143_SLICE_X9Y143_A1 = CLBLM_R_X7Y151_SLICE_X9Y151_A5Q;
  assign CLBLM_R_X7Y143_SLICE_X9Y143_A2 = CLBLM_R_X7Y151_SLICE_X9Y151_CQ;
  assign CLBLM_R_X7Y143_SLICE_X9Y143_A3 = CLBLM_R_X7Y143_SLICE_X9Y143_AQ;
  assign CLBLM_R_X7Y143_SLICE_X9Y143_A4 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X7Y143_SLICE_X9Y143_A5 = CLBLM_L_X8Y149_SLICE_X11Y149_AQ;
  assign CLBLM_R_X7Y143_SLICE_X9Y143_A6 = 1'b1;
  assign CLBLM_R_X11Y153_SLICE_X15Y153_C1 = CLBLM_R_X7Y146_SLICE_X8Y146_A5Q;
  assign CLBLM_R_X11Y153_SLICE_X15Y153_C2 = CLBLM_R_X11Y153_SLICE_X14Y153_A5Q;
  assign CLBLM_R_X11Y153_SLICE_X15Y153_C3 = CLBLM_R_X11Y153_SLICE_X14Y153_DO6;
  assign CLBLM_R_X7Y143_SLICE_X9Y143_B1 = CLBLM_R_X7Y144_SLICE_X8Y144_BQ;
  assign CLBLM_R_X7Y143_SLICE_X9Y143_B2 = RIOB33_X105Y113_IOB_X1Y113_I;
  assign CLBLM_R_X7Y143_SLICE_X9Y143_B3 = CLBLM_R_X5Y143_SLICE_X7Y143_C5Q;
  assign CLBLM_R_X7Y143_SLICE_X9Y143_B4 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X7Y143_SLICE_X9Y143_B5 = CLBLM_L_X8Y144_SLICE_X10Y144_AQ;
  assign CLBLM_R_X7Y143_SLICE_X9Y143_B6 = 1'b1;
  assign CLBLM_R_X11Y153_SLICE_X15Y153_CLK = CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O;
  assign CLBLM_R_X11Y153_SLICE_X15Y153_D1 = 1'b1;
  assign CLBLM_R_X7Y143_SLICE_X9Y143_C1 = CLBLM_R_X11Y146_SLICE_X14Y146_BO6;
  assign CLBLM_R_X7Y143_SLICE_X9Y143_C2 = CLBLM_R_X7Y143_SLICE_X9Y143_CQ;
  assign CLBLM_R_X7Y143_SLICE_X9Y143_C3 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X7Y143_SLICE_X9Y143_C4 = CLBLL_L_X4Y151_SLICE_X4Y151_CQ;
  assign CLBLM_R_X7Y143_SLICE_X9Y143_C5 = CLBLM_R_X7Y143_SLICE_X9Y143_DO6;
  assign CLBLM_R_X7Y143_SLICE_X9Y143_C6 = CLBLL_L_X2Y146_SLICE_X1Y146_BQ;
  assign CLBLM_R_X11Y153_SLICE_X15Y153_D3 = CLBLM_R_X11Y153_SLICE_X14Y153_DO6;
  assign CLBLM_R_X11Y153_SLICE_X15Y153_D4 = 1'b1;
  assign CLBLM_R_X7Y143_SLICE_X9Y143_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X11Y153_SLICE_X14Y153_A1 = CLBLM_L_X10Y148_SLICE_X13Y148_C5Q;
  assign CLBLM_R_X11Y153_SLICE_X14Y153_A2 = CLBLM_R_X11Y153_SLICE_X15Y153_BO6;
  assign CLBLM_R_X11Y153_SLICE_X14Y153_A3 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X11Y153_SLICE_X14Y153_A4 = CLBLM_L_X8Y152_SLICE_X10Y152_C5Q;
  assign CLBLM_R_X11Y153_SLICE_X14Y153_A5 = CLBLM_R_X11Y153_SLICE_X14Y153_CO6;
  assign CLBLM_R_X7Y143_SLICE_X9Y143_D1 = 1'b1;
  assign CLBLM_R_X7Y143_SLICE_X9Y143_D2 = CLBLM_L_X8Y142_SLICE_X10Y142_CQ;
  assign CLBLM_R_X7Y143_SLICE_X9Y143_D3 = 1'b1;
  assign CLBLM_R_X7Y143_SLICE_X9Y143_D4 = CLBLM_R_X7Y141_SLICE_X9Y141_AQ;
  assign CLBLM_R_X7Y143_SLICE_X9Y143_D5 = 1'b1;
  assign CLBLM_R_X7Y143_SLICE_X9Y143_D6 = 1'b1;
  assign CLBLM_R_X7Y151_SLICE_X8Y151_C3 = CLBLM_R_X7Y155_SLICE_X8Y155_AQ;
  assign CLBLM_R_X11Y153_SLICE_X14Y153_A6 = 1'b1;
  assign CLBLM_R_X7Y151_SLICE_X8Y151_C4 = CLBLM_R_X3Y146_SLICE_X2Y146_D5Q;
  assign CLBLM_R_X11Y153_SLICE_X14Y153_B1 = CLBLM_L_X8Y152_SLICE_X10Y152_CQ;
  assign CLBLM_R_X11Y153_SLICE_X14Y153_B2 = CLBLM_L_X10Y152_SLICE_X13Y152_BQ;
  assign CLBLM_R_X7Y143_SLICE_X8Y143_A1 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X7Y143_SLICE_X8Y143_A2 = CLBLM_L_X8Y149_SLICE_X11Y149_AQ;
  assign CLBLM_R_X7Y143_SLICE_X8Y143_A3 = CLBLM_R_X7Y143_SLICE_X8Y143_AQ;
  assign CLBLM_R_X7Y143_SLICE_X8Y143_A4 = CLBLM_L_X10Y146_SLICE_X12Y146_D5Q;
  assign CLBLM_R_X7Y143_SLICE_X8Y143_A5 = CLBLL_L_X4Y147_SLICE_X5Y147_B5Q;
  assign CLBLM_R_X7Y143_SLICE_X8Y143_A6 = CLBLM_R_X7Y143_SLICE_X8Y143_CO6;
  assign CLBLM_R_X7Y151_SLICE_X8Y151_C5 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X7Y151_SLICE_X8Y151_C6 = 1'b1;
  assign CLBLM_R_X11Y153_SLICE_X14Y153_C1 = CLBLM_R_X7Y146_SLICE_X8Y146_A5Q;
  assign CLBLM_R_X7Y143_SLICE_X8Y143_B1 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X7Y143_SLICE_X8Y143_B2 = CLBLM_R_X7Y143_SLICE_X8Y143_BQ;
  assign CLBLM_R_X7Y143_SLICE_X8Y143_B3 = CLBLM_R_X3Y143_SLICE_X3Y143_AQ;
  assign CLBLM_R_X7Y143_SLICE_X8Y143_B4 = CLBLM_L_X12Y149_SLICE_X17Y149_CO6;
  assign CLBLM_R_X7Y143_SLICE_X8Y143_B5 = 1'b1;
  assign CLBLM_R_X7Y143_SLICE_X8Y143_B6 = CLBLM_R_X7Y144_SLICE_X8Y144_CQ;
  assign CLBLM_R_X11Y153_SLICE_X14Y153_D1 = CLBLM_L_X10Y152_SLICE_X13Y152_AQ;
  assign CLBLM_R_X11Y153_SLICE_X14Y153_D2 = CLBLM_L_X10Y152_SLICE_X13Y152_BQ;
  assign CLBLM_R_X11Y153_SLICE_X14Y153_D3 = CLBLM_R_X11Y153_SLICE_X14Y153_AQ;
  assign CLBLM_R_X7Y143_SLICE_X8Y143_C1 = CLBLM_R_X7Y143_SLICE_X9Y143_AQ;
  assign CLBLM_R_X7Y143_SLICE_X8Y143_C2 = CLBLM_L_X10Y143_SLICE_X12Y143_BQ;
  assign CLBLM_R_X7Y143_SLICE_X8Y143_C3 = CLBLM_L_X10Y144_SLICE_X13Y144_DQ;
  assign CLBLM_R_X7Y143_SLICE_X8Y143_C4 = CLBLM_L_X8Y143_SLICE_X10Y143_BQ;
  assign CLBLM_R_X7Y143_SLICE_X8Y143_C5 = CLBLM_R_X7Y144_SLICE_X8Y144_AQ;
  assign CLBLM_R_X7Y143_SLICE_X8Y143_C6 = 1'b1;
  assign CLBLM_R_X11Y153_SLICE_X14Y153_D4 = CLBLM_L_X10Y152_SLICE_X12Y152_AQ;
  assign CLBLM_R_X11Y153_SLICE_X14Y153_D5 = 1'b1;
  assign CLBLM_R_X11Y153_SLICE_X14Y153_D6 = CLBLM_L_X8Y152_SLICE_X10Y152_CQ;
  assign CLBLM_R_X7Y143_SLICE_X8Y143_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign LIOB33_X0Y159_IOB_X0Y160_O = CLBLL_L_X2Y148_SLICE_X0Y148_AQ;
  assign CLBLM_R_X7Y143_SLICE_X8Y143_D1 = CLBLM_R_X7Y143_SLICE_X9Y143_AQ;
  assign CLBLM_R_X7Y143_SLICE_X8Y143_D2 = CLBLM_R_X7Y143_SLICE_X8Y143_AQ;
  assign CLBLM_R_X7Y143_SLICE_X8Y143_D3 = CLBLM_L_X10Y144_SLICE_X13Y144_DQ;
  assign CLBLM_R_X7Y143_SLICE_X8Y143_D4 = CLBLM_R_X7Y144_SLICE_X8Y144_AQ;
  assign CLBLM_R_X7Y143_SLICE_X8Y143_D5 = CLBLM_L_X10Y143_SLICE_X12Y143_BQ;
  assign CLBLM_R_X7Y143_SLICE_X8Y143_D6 = CLBLM_L_X8Y143_SLICE_X10Y143_BQ;
  assign LIOB33_X0Y159_IOB_X0Y159_O = CLBLL_L_X2Y146_SLICE_X0Y146_CQ;
  assign CLBLM_R_X5Y153_SLICE_X6Y153_A5 = CLBLM_R_X7Y152_SLICE_X8Y152_BQ;
  assign CLBLM_R_X5Y153_SLICE_X6Y153_A6 = 1'b1;
  assign CLBLM_R_X7Y151_SLICE_X8Y151_D3 = CLBLM_L_X10Y151_SLICE_X13Y151_A5Q;
  assign CLBLM_R_X7Y151_SLICE_X8Y151_D4 = CLBLM_L_X8Y152_SLICE_X10Y152_A5Q;
  assign CLBLM_R_X7Y151_SLICE_X8Y151_D5 = 1'b1;
  assign CLBLM_R_X7Y151_SLICE_X8Y151_D6 = 1'b1;
  assign CLBLM_L_X8Y145_SLICE_X10Y145_A3 = CLBLM_R_X3Y145_SLICE_X3Y145_BQ;
  assign CLBLM_R_X5Y153_SLICE_X6Y153_B1 = CLBLM_R_X5Y153_SLICE_X6Y153_CQ;
  assign CLBLM_L_X8Y145_SLICE_X10Y145_A4 = CLBLL_L_X4Y146_SLICE_X5Y146_AQ;
  assign CLBLM_R_X5Y153_SLICE_X6Y153_B2 = CLBLM_R_X5Y153_SLICE_X7Y153_CQ;
  assign CLBLM_L_X8Y145_SLICE_X10Y145_A5 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_L_X8Y145_SLICE_X10Y145_A6 = 1'b1;
  assign CLBLM_L_X8Y150_SLICE_X11Y150_A1 = CLBLM_R_X7Y148_SLICE_X9Y148_CQ;
  assign CLBLM_L_X8Y150_SLICE_X11Y150_A2 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_L_X8Y150_SLICE_X11Y150_A3 = CLBLM_L_X8Y150_SLICE_X11Y150_AQ;
  assign CLBLM_L_X8Y150_SLICE_X11Y150_A4 = CLBLM_R_X3Y145_SLICE_X3Y145_D5Q;
  assign CLBLM_L_X8Y150_SLICE_X11Y150_A5 = CLBLM_R_X11Y151_SLICE_X15Y151_AQ;
  assign CLBLM_L_X8Y150_SLICE_X11Y150_A6 = CLBLL_L_X4Y151_SLICE_X4Y151_BQ;
  assign CLBLM_L_X8Y150_SLICE_X11Y150_B1 = CLBLM_R_X7Y153_SLICE_X8Y153_A5Q;
  assign CLBLM_L_X8Y150_SLICE_X11Y150_B2 = CLBLM_R_X7Y144_SLICE_X9Y144_B5Q;
  assign CLBLM_L_X8Y150_SLICE_X11Y150_B3 = CLBLM_R_X7Y149_SLICE_X8Y149_AQ;
  assign CLBLM_L_X8Y150_SLICE_X11Y150_B4 = CLBLM_L_X12Y147_SLICE_X16Y147_DO6;
  assign CLBLM_L_X8Y150_SLICE_X11Y150_B5 = CLBLL_L_X4Y148_SLICE_X4Y148_CQ;
  assign CLBLM_L_X8Y150_SLICE_X11Y150_B6 = 1'b1;
  assign CLBLM_L_X8Y150_SLICE_X11Y150_C1 = CLBLL_L_X2Y148_SLICE_X0Y148_AQ;
  assign CLBLM_L_X8Y150_SLICE_X11Y150_C2 = CLBLM_R_X7Y142_SLICE_X8Y142_D5Q;
  assign CLBLM_L_X8Y150_SLICE_X11Y150_C3 = CLBLM_L_X10Y151_SLICE_X13Y151_BO5;
  assign CLBLM_L_X8Y150_SLICE_X11Y150_C4 = CLBLM_L_X10Y150_SLICE_X12Y150_BO5;
  assign CLBLM_L_X8Y150_SLICE_X11Y150_C5 = CLBLM_L_X8Y143_SLICE_X11Y143_CQ;
  assign CLBLM_L_X8Y150_SLICE_X11Y150_C6 = CLBLM_L_X12Y149_SLICE_X17Y149_BO5;
  assign CLBLM_L_X8Y150_SLICE_X11Y150_CLK = CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O;
  assign CLBLM_L_X8Y150_SLICE_X11Y150_D1 = CLBLM_R_X7Y150_SLICE_X9Y150_CO6;
  assign CLBLM_L_X8Y150_SLICE_X11Y150_D2 = CLBLM_R_X11Y148_SLICE_X15Y148_AO6;
  assign CLBLM_L_X8Y150_SLICE_X11Y150_D3 = CLBLM_L_X10Y151_SLICE_X13Y151_BO5;
  assign CLBLM_L_X8Y150_SLICE_X11Y150_D4 = 1'b1;
  assign CLBLM_L_X8Y150_SLICE_X11Y150_D5 = CLBLM_L_X8Y146_SLICE_X10Y146_AQ;
  assign CLBLM_L_X8Y150_SLICE_X11Y150_D6 = CLBLM_L_X8Y152_SLICE_X11Y152_BQ;
  assign CLBLM_L_X8Y150_SLICE_X10Y150_A1 = CLBLM_L_X10Y146_SLICE_X12Y146_BQ;
  assign CLBLM_L_X8Y150_SLICE_X10Y150_A2 = CLBLM_R_X13Y149_SLICE_X18Y149_AO6;
  assign CLBLM_L_X8Y150_SLICE_X10Y150_A3 = CLBLM_L_X8Y150_SLICE_X10Y150_AQ;
  assign CLBLM_L_X8Y150_SLICE_X10Y150_A4 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_L_X8Y150_SLICE_X10Y150_A5 = 1'b1;
  assign CLBLM_L_X8Y150_SLICE_X10Y150_A6 = CLBLM_R_X7Y151_SLICE_X9Y151_AQ;
  assign LIOI3_X0Y161_OLOGIC_X0Y162_D1 = CLBLM_L_X10Y144_SLICE_X12Y144_BO6;
  assign CLBLM_L_X8Y150_SLICE_X10Y150_B1 = CLBLM_R_X7Y153_SLICE_X8Y153_A5Q;
  assign CLBLM_L_X8Y150_SLICE_X10Y150_B2 = CLBLL_L_X4Y148_SLICE_X4Y148_CQ;
  assign CLBLM_L_X8Y150_SLICE_X10Y150_B3 = CLBLM_R_X7Y149_SLICE_X8Y149_AQ;
  assign CLBLM_L_X8Y150_SLICE_X10Y150_B4 = CLBLM_R_X7Y144_SLICE_X9Y144_B5Q;
  assign CLBLM_L_X8Y150_SLICE_X10Y150_B5 = CLBLM_L_X12Y147_SLICE_X16Y147_DO6;
  assign CLBLM_L_X8Y150_SLICE_X10Y150_B6 = 1'b1;
  assign LIOI3_X0Y161_OLOGIC_X0Y162_T1 = 1'b1;
  assign CLBLM_L_X8Y150_SLICE_X10Y150_C1 = CLBLM_R_X7Y144_SLICE_X9Y144_B5Q;
  assign CLBLM_L_X8Y150_SLICE_X10Y150_C2 = 1'b1;
  assign CLBLM_L_X8Y150_SLICE_X10Y150_C3 = CLBLM_L_X8Y153_SLICE_X10Y153_B5Q;
  assign CLBLM_L_X8Y150_SLICE_X10Y150_C4 = CLBLL_L_X4Y145_SLICE_X4Y145_CQ;
  assign CLBLM_L_X8Y150_SLICE_X10Y150_C5 = CLBLM_R_X7Y153_SLICE_X8Y153_A5Q;
  assign CLBLM_L_X8Y150_SLICE_X10Y150_C6 = CLBLM_R_X11Y144_SLICE_X14Y144_AO6;
  assign LIOI3_X0Y101_OLOGIC_X0Y102_D1 = CLBLM_R_X5Y141_SLICE_X6Y141_DQ;
  assign LIOI3_X0Y161_OLOGIC_X0Y161_D1 = CLBLM_R_X5Y152_SLICE_X7Y152_DQ;
  assign CLBLM_L_X8Y150_SLICE_X10Y150_CLK = CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O;
  assign LIOI3_X0Y101_OLOGIC_X0Y102_T1 = 1'b1;
  assign CLBLM_L_X8Y150_SLICE_X10Y150_D1 = CLBLM_L_X8Y150_SLICE_X10Y150_CO6;
  assign CLBLM_L_X8Y150_SLICE_X10Y150_D2 = CLBLM_L_X8Y153_SLICE_X10Y153_BQ;
  assign CLBLM_L_X8Y150_SLICE_X10Y150_D3 = CLBLM_L_X8Y150_SLICE_X11Y150_BO5;
  assign CLBLM_L_X8Y150_SLICE_X10Y150_D4 = CLBLM_R_X7Y148_SLICE_X8Y148_AO5;
  assign CLBLM_L_X8Y150_SLICE_X10Y150_D5 = 1'b1;
  assign CLBLM_L_X8Y150_SLICE_X10Y150_D6 = CLBLM_L_X8Y150_SLICE_X10Y150_AQ;
  assign LIOI3_X0Y161_OLOGIC_X0Y161_T1 = 1'b1;
  assign LIOI3_X0Y101_OLOGIC_X0Y101_D1 = CLBLM_L_X8Y145_SLICE_X11Y145_C5Q;
  assign LIOI3_TBYTETERM_X0Y63_OLOGIC_X0Y64_D1 = CLBLM_R_X7Y141_SLICE_X8Y141_AO5;
  assign LIOI3_X0Y101_OLOGIC_X0Y101_T1 = 1'b1;
  assign LIOI3_TBYTETERM_X0Y63_OLOGIC_X0Y64_T1 = 1'b1;
  assign CLBLM_R_X7Y144_SLICE_X9Y144_A1 = CLBLM_R_X7Y144_SLICE_X9Y144_AQ;
  assign CLBLM_R_X7Y144_SLICE_X9Y144_A2 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X7Y144_SLICE_X9Y144_A3 = CLBLM_R_X3Y145_SLICE_X3Y145_D5Q;
  assign CLBLM_R_X7Y144_SLICE_X9Y144_A4 = CLBLM_R_X5Y144_SLICE_X6Y144_D5Q;
  assign CLBLM_R_X7Y144_SLICE_X9Y144_A5 = CLBLM_L_X10Y144_SLICE_X13Y144_C5Q;
  assign CLBLM_R_X7Y144_SLICE_X9Y144_A6 = CLBLL_L_X4Y151_SLICE_X4Y151_BQ;
  assign CLBLM_R_X7Y144_SLICE_X9Y144_AX = CLBLM_L_X8Y144_SLICE_X10Y144_BO5;
  assign CLBLM_R_X7Y144_SLICE_X9Y144_B1 = CLBLL_L_X4Y146_SLICE_X4Y146_BQ;
  assign CLBLM_R_X7Y144_SLICE_X9Y144_B2 = 1'b1;
  assign CLBLM_R_X7Y144_SLICE_X9Y144_B3 = CLBLM_L_X8Y143_SLICE_X10Y143_AQ;
  assign CLBLM_R_X7Y144_SLICE_X9Y144_B4 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X7Y144_SLICE_X9Y144_B5 = CLBLM_L_X12Y151_SLICE_X16Y151_AQ;
  assign CLBLM_R_X7Y144_SLICE_X9Y144_B6 = 1'b1;
  assign CLBLM_R_X7Y144_SLICE_X9Y144_C1 = CLBLM_R_X5Y142_SLICE_X6Y142_D5Q;
  assign CLBLM_R_X7Y144_SLICE_X9Y144_C2 = CLBLL_L_X4Y148_SLICE_X4Y148_CQ;
  assign CLBLM_R_X7Y144_SLICE_X9Y144_C3 = CLBLM_R_X7Y149_SLICE_X8Y149_AQ;
  assign CLBLM_R_X7Y144_SLICE_X9Y144_C4 = CLBLL_L_X4Y147_SLICE_X4Y147_CQ;
  assign CLBLM_R_X7Y144_SLICE_X9Y144_C5 = CLBLM_R_X7Y151_SLICE_X8Y151_D5Q;
  assign CLBLM_R_X7Y144_SLICE_X9Y144_C6 = CLBLM_L_X10Y146_SLICE_X12Y146_DQ;
  assign CLBLM_R_X7Y144_SLICE_X9Y144_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X7Y144_SLICE_X9Y144_D1 = CLBLM_R_X5Y146_SLICE_X7Y146_C5Q;
  assign CLBLM_R_X7Y144_SLICE_X9Y144_D2 = CLBLM_R_X7Y153_SLICE_X8Y153_A5Q;
  assign CLBLM_R_X7Y144_SLICE_X9Y144_D3 = 1'b1;
  assign CLBLM_R_X7Y144_SLICE_X9Y144_D4 = CLBLM_R_X7Y144_SLICE_X9Y144_CO6;
  assign CLBLM_R_X7Y144_SLICE_X9Y144_D5 = CLBLM_R_X7Y144_SLICE_X9Y144_B5Q;
  assign CLBLM_R_X7Y144_SLICE_X9Y144_D6 = CLBLM_R_X5Y148_SLICE_X6Y148_BQ;
  assign CLBLM_R_X7Y144_SLICE_X8Y144_A1 = CLBLM_L_X8Y149_SLICE_X11Y149_AQ;
  assign CLBLM_R_X7Y144_SLICE_X8Y144_A2 = CLBLM_R_X5Y145_SLICE_X6Y145_C5Q;
  assign CLBLM_R_X7Y144_SLICE_X8Y144_A3 = CLBLM_R_X7Y144_SLICE_X8Y144_AQ;
  assign CLBLM_R_X7Y144_SLICE_X8Y144_A4 = CLBLM_R_X5Y152_SLICE_X6Y152_CQ;
  assign CLBLM_R_X7Y144_SLICE_X8Y144_A5 = CLBLM_R_X7Y143_SLICE_X8Y143_CO5;
  assign CLBLM_R_X7Y144_SLICE_X8Y144_A6 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X7Y152_SLICE_X8Y152_C5 = 1'b1;
  assign LIOB33_X0Y161_IOB_X0Y161_O = CLBLM_R_X5Y152_SLICE_X7Y152_DQ;
  assign LIOB33_X0Y161_IOB_X0Y162_O = CLBLM_L_X10Y144_SLICE_X12Y144_BO6;
  assign CLBLM_R_X7Y144_SLICE_X8Y144_B1 = CLBLM_R_X3Y146_SLICE_X2Y146_D5Q;
  assign CLBLM_R_X7Y144_SLICE_X8Y144_B2 = 1'b1;
  assign CLBLM_R_X7Y144_SLICE_X8Y144_B3 = CLBLM_R_X7Y144_SLICE_X8Y144_AQ;
  assign CLBLM_R_X7Y144_SLICE_X8Y144_B4 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X7Y144_SLICE_X8Y144_B5 = CLBLL_L_X4Y147_SLICE_X5Y147_AQ;
  assign CLBLM_R_X7Y144_SLICE_X8Y144_B6 = 1'b1;
  assign CLBLM_R_X7Y144_SLICE_X8Y144_C1 = 1'b1;
  assign CLBLM_R_X7Y144_SLICE_X8Y144_C2 = CLBLL_L_X4Y142_SLICE_X5Y142_CQ;
  assign CLBLM_R_X7Y144_SLICE_X8Y144_C3 = CLBLM_R_X7Y144_SLICE_X9Y144_B5Q;
  assign CLBLM_R_X7Y144_SLICE_X8Y144_C4 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X7Y144_SLICE_X8Y144_C5 = CLBLM_R_X11Y149_SLICE_X15Y149_CO6;
  assign CLBLM_R_X7Y144_SLICE_X8Y144_C6 = 1'b1;
  assign CLBLM_R_X7Y144_SLICE_X8Y144_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X7Y144_SLICE_X8Y144_D1 = 1'b1;
  assign CLBLM_R_X7Y144_SLICE_X8Y144_D2 = CLBLM_L_X10Y149_SLICE_X12Y149_BQ;
  assign CLBLM_R_X7Y144_SLICE_X8Y144_D3 = CLBLM_R_X5Y142_SLICE_X6Y142_BQ;
  assign CLBLM_R_X7Y144_SLICE_X8Y144_D4 = CLBLM_L_X10Y147_SLICE_X12Y147_BQ;
  assign CLBLM_R_X7Y144_SLICE_X8Y144_D5 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X7Y144_SLICE_X8Y144_D6 = 1'b1;
  assign RIOI3_X105Y145_ILOGIC_X1Y146_D = RIOB33_X105Y145_IOB_X1Y146_I;
  assign RIOI3_X105Y145_ILOGIC_X1Y145_D = RIOB33_X105Y145_IOB_X1Y145_I;
  assign LIOI3_TBYTETERM_X0Y63_ILOGIC_X0Y63_D = LIOB33_X0Y63_IOB_X0Y63_I;
  assign CLBLM_L_X8Y151_SLICE_X11Y151_A1 = CLBLM_R_X3Y145_SLICE_X3Y145_D5Q;
  assign CLBLM_L_X8Y151_SLICE_X11Y151_A2 = CLBLL_L_X4Y151_SLICE_X4Y151_BQ;
  assign CLBLM_L_X8Y151_SLICE_X11Y151_A3 = CLBLM_L_X8Y151_SLICE_X11Y151_AQ;
  assign CLBLM_L_X8Y151_SLICE_X11Y151_A4 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_L_X8Y151_SLICE_X11Y151_A5 = CLBLL_L_X4Y151_SLICE_X4Y151_A5Q;
  assign CLBLM_L_X8Y151_SLICE_X11Y151_A6 = CLBLM_L_X8Y152_SLICE_X11Y152_DQ;
  assign CLBLM_R_X7Y152_SLICE_X8Y152_C6 = CLBLM_R_X7Y152_SLICE_X8Y152_AQ;
  assign CLBLM_L_X8Y151_SLICE_X11Y151_B1 = CLBLM_R_X7Y152_SLICE_X9Y152_B5Q;
  assign CLBLM_L_X8Y151_SLICE_X11Y151_B2 = CLBLM_L_X8Y150_SLICE_X11Y150_BO5;
  assign CLBLM_L_X8Y151_SLICE_X11Y151_B3 = CLBLM_L_X10Y151_SLICE_X13Y151_BO6;
  assign CLBLM_L_X8Y151_SLICE_X11Y151_B4 = CLBLM_L_X10Y150_SLICE_X12Y150_BO5;
  assign CLBLM_L_X8Y151_SLICE_X11Y151_B5 = CLBLM_R_X5Y153_SLICE_X7Y153_CQ;
  assign CLBLM_L_X8Y151_SLICE_X11Y151_B6 = CLBLM_L_X10Y152_SLICE_X12Y152_CQ;
  assign CLBLM_L_X8Y151_SLICE_X11Y151_C1 = CLBLM_R_X7Y153_SLICE_X8Y153_A5Q;
  assign CLBLM_L_X8Y151_SLICE_X11Y151_C2 = CLBLM_R_X3Y148_SLICE_X3Y148_CQ;
  assign CLBLM_L_X8Y151_SLICE_X11Y151_C3 = CLBLM_R_X7Y149_SLICE_X8Y149_AQ;
  assign CLBLM_L_X8Y151_SLICE_X11Y151_C4 = CLBLL_L_X4Y148_SLICE_X4Y148_CQ;
  assign CLBLM_L_X8Y151_SLICE_X11Y151_C5 = CLBLM_L_X12Y147_SLICE_X16Y147_DO6;
  assign CLBLM_L_X8Y151_SLICE_X11Y151_C6 = CLBLM_R_X7Y144_SLICE_X9Y144_B5Q;
  assign CLBLM_L_X8Y151_SLICE_X11Y151_CLK = CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O;
  assign CLBLM_L_X8Y151_SLICE_X11Y151_D1 = CLBLM_R_X5Y146_SLICE_X6Y146_BQ;
  assign CLBLM_L_X8Y151_SLICE_X11Y151_D2 = CLBLM_L_X10Y151_SLICE_X13Y151_BO6;
  assign CLBLM_L_X8Y151_SLICE_X11Y151_D3 = CLBLM_L_X10Y152_SLICE_X13Y152_CQ;
  assign CLBLM_L_X8Y151_SLICE_X11Y151_D4 = CLBLM_L_X8Y151_SLICE_X11Y151_CO6;
  assign CLBLM_L_X8Y151_SLICE_X11Y151_D5 = CLBLM_L_X10Y146_SLICE_X13Y146_DO6;
  assign CLBLM_L_X8Y151_SLICE_X11Y151_D6 = CLBLM_L_X10Y148_SLICE_X12Y148_AO6;
  assign CLBLM_L_X8Y151_SLICE_X10Y151_A1 = CLBLM_R_X7Y152_SLICE_X9Y152_BQ;
  assign CLBLM_L_X8Y151_SLICE_X10Y151_A2 = CLBLM_L_X8Y153_SLICE_X10Y153_C5Q;
  assign CLBLM_L_X8Y151_SLICE_X10Y151_A3 = CLBLM_L_X8Y151_SLICE_X10Y151_AQ;
  assign CLBLM_L_X8Y151_SLICE_X10Y151_A4 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_L_X8Y151_SLICE_X10Y151_A5 = CLBLL_L_X4Y143_SLICE_X4Y143_BQ;
  assign CLBLM_L_X8Y151_SLICE_X10Y151_A6 = 1'b1;
  assign CLBLM_L_X8Y151_SLICE_X10Y151_B1 = CLBLM_R_X7Y152_SLICE_X9Y152_B5Q;
  assign CLBLM_L_X8Y151_SLICE_X10Y151_B2 = 1'b1;
  assign CLBLM_L_X8Y151_SLICE_X10Y151_B3 = CLBLM_L_X10Y152_SLICE_X13Y152_BQ;
  assign CLBLM_L_X8Y151_SLICE_X10Y151_B4 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_L_X8Y151_SLICE_X10Y151_B5 = CLBLL_L_X4Y149_SLICE_X4Y149_B5Q;
  assign CLBLM_L_X8Y151_SLICE_X10Y151_B6 = 1'b1;
  assign CLBLM_L_X8Y151_SLICE_X10Y151_C1 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_L_X8Y151_SLICE_X10Y151_C2 = CLBLM_L_X8Y151_SLICE_X10Y151_CQ;
  assign CLBLM_L_X8Y151_SLICE_X10Y151_C3 = CLBLM_L_X8Y152_SLICE_X11Y152_DQ;
  assign CLBLM_L_X8Y151_SLICE_X10Y151_C4 = CLBLM_R_X7Y152_SLICE_X9Y152_C5Q;
  assign CLBLM_L_X8Y151_SLICE_X10Y151_C5 = CLBLM_R_X5Y145_SLICE_X6Y145_AQ;
  assign CLBLM_L_X8Y151_SLICE_X10Y151_C6 = 1'b1;
  assign CLBLM_L_X8Y151_SLICE_X10Y151_CLK = CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O;
  assign CLBLM_L_X8Y151_SLICE_X10Y151_D1 = CLBLM_R_X11Y146_SLICE_X15Y146_BO6;
  assign CLBLM_L_X8Y151_SLICE_X10Y151_D2 = CLBLM_R_X7Y153_SLICE_X8Y153_DQ;
  assign CLBLM_L_X8Y151_SLICE_X10Y151_D3 = CLBLM_L_X12Y147_SLICE_X16Y147_DO6;
  assign CLBLM_L_X8Y151_SLICE_X10Y151_D4 = CLBLM_L_X8Y152_SLICE_X11Y152_DQ;
  assign CLBLM_L_X8Y151_SLICE_X10Y151_D5 = CLBLM_R_X7Y149_SLICE_X8Y149_AQ;
  assign CLBLM_L_X8Y151_SLICE_X10Y151_D6 = CLBLL_L_X4Y148_SLICE_X4Y148_CQ;
  assign CLBLM_R_X7Y145_SLICE_X9Y145_A1 = CLBLM_R_X7Y144_SLICE_X9Y144_B5Q;
  assign CLBLM_R_X7Y145_SLICE_X9Y145_A2 = CLBLM_R_X7Y146_SLICE_X9Y146_CO5;
  assign CLBLM_R_X7Y145_SLICE_X9Y145_A3 = CLBLM_R_X7Y147_SLICE_X9Y147_DQ;
  assign CLBLM_R_X7Y145_SLICE_X9Y145_A4 = CLBLM_R_X5Y141_SLICE_X6Y141_B5Q;
  assign CLBLM_R_X7Y145_SLICE_X9Y145_A5 = CLBLM_R_X7Y144_SLICE_X9Y144_CO6;
  assign CLBLM_R_X7Y145_SLICE_X9Y145_A6 = CLBLM_R_X7Y153_SLICE_X8Y153_A5Q;
  assign CLBLM_R_X7Y145_SLICE_X9Y145_B1 = CLBLM_R_X7Y144_SLICE_X9Y144_B5Q;
  assign CLBLM_R_X7Y145_SLICE_X9Y145_B2 = CLBLM_R_X7Y146_SLICE_X9Y146_CO5;
  assign CLBLM_R_X7Y145_SLICE_X9Y145_B3 = CLBLM_R_X3Y148_SLICE_X3Y148_BQ;
  assign CLBLM_R_X7Y145_SLICE_X9Y145_B4 = CLBLM_R_X7Y146_SLICE_X8Y146_BQ;
  assign CLBLM_R_X7Y145_SLICE_X9Y145_B5 = CLBLM_R_X7Y144_SLICE_X9Y144_CO6;
  assign CLBLM_R_X7Y145_SLICE_X9Y145_B6 = CLBLM_R_X7Y153_SLICE_X8Y153_A5Q;
  assign CLBLM_R_X7Y145_SLICE_X9Y145_C1 = CLBLM_R_X7Y144_SLICE_X9Y144_CO6;
  assign CLBLM_R_X7Y145_SLICE_X9Y145_C2 = CLBLM_R_X5Y142_SLICE_X7Y142_A5Q;
  assign CLBLM_R_X7Y145_SLICE_X9Y145_C3 = CLBLM_R_X7Y144_SLICE_X9Y144_B5Q;
  assign CLBLM_R_X7Y145_SLICE_X9Y145_C4 = CLBLM_R_X7Y153_SLICE_X8Y153_A5Q;
  assign CLBLM_R_X7Y145_SLICE_X9Y145_C5 = CLBLM_R_X5Y147_SLICE_X7Y147_B5Q;
  assign CLBLM_R_X7Y145_SLICE_X9Y145_C6 = CLBLM_R_X7Y146_SLICE_X9Y146_CO5;
  assign LIOB33_X0Y163_IOB_X0Y163_O = CLBLM_R_X5Y152_SLICE_X7Y152_DO6;
  assign LIOB33_X0Y163_IOB_X0Y164_O = RIOB33_X105Y101_IOB_X1Y102_I;
  assign CLBLM_R_X7Y145_SLICE_X9Y145_D1 = CLBLM_R_X7Y144_SLICE_X9Y144_CO6;
  assign CLBLM_R_X7Y145_SLICE_X9Y145_D2 = CLBLM_R_X7Y146_SLICE_X9Y146_CO5;
  assign CLBLM_R_X7Y145_SLICE_X9Y145_D3 = CLBLM_R_X7Y144_SLICE_X9Y144_B5Q;
  assign CLBLM_R_X7Y145_SLICE_X9Y145_D4 = CLBLM_R_X7Y153_SLICE_X8Y153_A5Q;
  assign CLBLM_R_X7Y145_SLICE_X9Y145_D5 = CLBLM_R_X7Y145_SLICE_X8Y145_BQ;
  assign CLBLM_R_X7Y145_SLICE_X9Y145_D6 = CLBLM_R_X3Y148_SLICE_X3Y148_C5Q;
  assign CLBLM_R_X7Y145_SLICE_X8Y145_A1 = CLBLM_R_X7Y145_SLICE_X8Y145_B5Q;
  assign CLBLM_R_X7Y145_SLICE_X8Y145_A2 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X7Y145_SLICE_X8Y145_A3 = CLBLL_L_X4Y153_SLICE_X5Y153_A5Q;
  assign CLBLM_R_X7Y145_SLICE_X8Y145_A4 = CLBLM_L_X8Y154_SLICE_X10Y154_BO5;
  assign CLBLM_R_X7Y145_SLICE_X8Y145_A5 = CLBLL_L_X4Y143_SLICE_X5Y143_D5Q;
  assign CLBLM_R_X7Y145_SLICE_X8Y145_A6 = 1'b1;
  assign CLBLL_L_X2Y144_SLICE_X0Y144_A1 = 1'b1;
  assign CLBLL_L_X2Y144_SLICE_X0Y144_A2 = 1'b1;
  assign CLBLL_L_X2Y144_SLICE_X0Y144_A3 = 1'b1;
  assign CLBLL_L_X2Y144_SLICE_X0Y144_A4 = 1'b1;
  assign CLBLL_L_X2Y144_SLICE_X0Y144_A5 = 1'b1;
  assign CLBLL_L_X2Y144_SLICE_X0Y144_A6 = 1'b1;
  assign CLBLM_R_X7Y145_SLICE_X8Y145_B1 = CLBLM_R_X7Y146_SLICE_X8Y146_DQ;
  assign CLBLM_L_X12Y152_SLICE_X17Y152_C1 = 1'b1;
  assign CLBLL_L_X2Y144_SLICE_X0Y144_B1 = 1'b1;
  assign CLBLL_L_X2Y144_SLICE_X0Y144_B2 = 1'b1;
  assign CLBLL_L_X2Y144_SLICE_X0Y144_B3 = 1'b1;
  assign CLBLL_L_X2Y144_SLICE_X0Y144_B4 = 1'b1;
  assign CLBLL_L_X2Y144_SLICE_X0Y144_B5 = 1'b1;
  assign CLBLL_L_X2Y144_SLICE_X0Y144_B6 = 1'b1;
  assign CLBLM_R_X7Y145_SLICE_X8Y145_C2 = CLBLL_L_X4Y142_SLICE_X4Y142_CQ;
  assign CLBLM_R_X7Y145_SLICE_X8Y145_C3 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X7Y145_SLICE_X8Y145_C4 = CLBLM_R_X5Y152_SLICE_X6Y152_DQ;
  assign CLBLL_L_X2Y144_SLICE_X0Y144_C1 = 1'b1;
  assign CLBLL_L_X2Y144_SLICE_X0Y144_C2 = 1'b1;
  assign CLBLL_L_X2Y144_SLICE_X0Y144_C3 = 1'b1;
  assign CLBLL_L_X2Y144_SLICE_X0Y144_C4 = 1'b1;
  assign CLBLL_L_X2Y144_SLICE_X0Y144_C5 = 1'b1;
  assign CLBLL_L_X2Y144_SLICE_X0Y144_C6 = 1'b1;
  assign CLBLM_R_X7Y145_SLICE_X8Y145_C5 = CLBLM_R_X5Y147_SLICE_X7Y147_B5Q;
  assign CLBLM_R_X7Y145_SLICE_X8Y145_C6 = 1'b1;
  assign CLBLM_R_X7Y145_SLICE_X8Y145_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X7Y145_SLICE_X8Y145_D1 = CLBLM_R_X5Y145_SLICE_X6Y145_D5Q;
  assign CLBLM_R_X7Y145_SLICE_X8Y145_D2 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X7Y145_SLICE_X8Y145_D3 = CLBLM_R_X5Y150_SLICE_X7Y150_A5Q;
  assign CLBLL_L_X2Y144_SLICE_X0Y144_D1 = 1'b1;
  assign CLBLL_L_X2Y144_SLICE_X0Y144_D2 = 1'b1;
  assign CLBLL_L_X2Y144_SLICE_X0Y144_D3 = 1'b1;
  assign CLBLL_L_X2Y144_SLICE_X0Y144_D4 = 1'b1;
  assign CLBLL_L_X2Y144_SLICE_X0Y144_D5 = 1'b1;
  assign CLBLL_L_X2Y144_SLICE_X0Y144_D6 = 1'b1;
  assign CLBLM_R_X7Y145_SLICE_X8Y145_D4 = CLBLM_R_X7Y144_SLICE_X9Y144_A5Q;
  assign CLBLM_R_X7Y145_SLICE_X8Y145_D5 = CLBLM_R_X5Y153_SLICE_X6Y153_D5Q;
  assign CLBLM_R_X7Y145_SLICE_X8Y145_D6 = 1'b1;
  assign CLBLL_L_X2Y144_SLICE_X1Y144_A1 = CLBLM_R_X3Y145_SLICE_X3Y145_CQ;
  assign CLBLL_L_X2Y144_SLICE_X1Y144_A2 = CLBLL_L_X2Y146_SLICE_X1Y146_B5Q;
  assign CLBLL_L_X2Y144_SLICE_X1Y144_A3 = 1'b1;
  assign CLBLL_L_X2Y144_SLICE_X1Y144_A4 = CLBLM_R_X3Y144_SLICE_X3Y144_AQ;
  assign CLBLL_L_X2Y144_SLICE_X1Y144_A5 = CLBLL_L_X2Y146_SLICE_X0Y146_DQ;
  assign CLBLL_L_X2Y144_SLICE_X1Y144_A6 = CLBLM_R_X5Y143_SLICE_X6Y143_D5Q;
  assign CLBLL_L_X2Y144_SLICE_X1Y144_B1 = 1'b1;
  assign CLBLL_L_X2Y144_SLICE_X1Y144_B2 = 1'b1;
  assign CLBLL_L_X2Y144_SLICE_X1Y144_B3 = 1'b1;
  assign CLBLL_L_X2Y144_SLICE_X1Y144_B4 = 1'b1;
  assign CLBLL_L_X2Y144_SLICE_X1Y144_B5 = 1'b1;
  assign CLBLL_L_X2Y144_SLICE_X1Y144_B6 = 1'b1;
  assign CLBLL_L_X2Y144_SLICE_X1Y144_C1 = 1'b1;
  assign CLBLL_L_X2Y144_SLICE_X1Y144_C2 = 1'b1;
  assign CLBLL_L_X2Y144_SLICE_X1Y144_C3 = 1'b1;
  assign CLBLL_L_X2Y144_SLICE_X1Y144_C4 = 1'b1;
  assign CLBLL_L_X2Y144_SLICE_X1Y144_C5 = 1'b1;
  assign CLBLL_L_X2Y144_SLICE_X1Y144_C6 = 1'b1;
  assign CLBLM_L_X12Y152_SLICE_X17Y152_D3 = 1'b1;
  assign CLBLM_L_X12Y152_SLICE_X17Y152_D4 = 1'b1;
  assign CLBLM_L_X12Y152_SLICE_X17Y152_D5 = 1'b1;
  assign CLBLL_L_X2Y144_SLICE_X1Y144_D1 = 1'b1;
  assign CLBLL_L_X2Y144_SLICE_X1Y144_D2 = 1'b1;
  assign CLBLL_L_X2Y144_SLICE_X1Y144_D3 = 1'b1;
  assign CLBLL_L_X2Y144_SLICE_X1Y144_D4 = 1'b1;
  assign CLBLL_L_X2Y144_SLICE_X1Y144_D5 = 1'b1;
  assign CLBLL_L_X2Y144_SLICE_X1Y144_D6 = 1'b1;
  assign CLBLM_L_X12Y152_SLICE_X17Y152_D6 = 1'b1;
  assign LIOI3_TBYTETERM_X0Y137_OLOGIC_X0Y137_T1 = 1'b1;
  assign CLBLM_L_X8Y152_SLICE_X11Y152_A1 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_L_X8Y152_SLICE_X11Y152_A2 = CLBLM_R_X11Y150_SLICE_X14Y150_AQ;
  assign CLBLM_L_X8Y152_SLICE_X11Y152_A3 = CLBLM_L_X8Y152_SLICE_X11Y152_AQ;
  assign CLBLM_L_X8Y152_SLICE_X11Y152_A4 = CLBLM_R_X7Y142_SLICE_X8Y142_C5Q;
  assign CLBLM_L_X8Y152_SLICE_X11Y152_A5 = CLBLM_R_X7Y152_SLICE_X8Y152_D5Q;
  assign CLBLM_L_X8Y152_SLICE_X11Y152_A6 = CLBLM_L_X8Y151_SLICE_X10Y151_A5Q;
  assign CLBLM_L_X8Y152_SLICE_X11Y152_B1 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_L_X8Y152_SLICE_X11Y152_B2 = CLBLM_L_X8Y152_SLICE_X11Y152_BQ;
  assign CLBLM_L_X8Y152_SLICE_X11Y152_B3 = CLBLM_R_X5Y150_SLICE_X7Y150_AQ;
  assign CLBLM_L_X8Y152_SLICE_X11Y152_B4 = CLBLL_L_X4Y147_SLICE_X5Y147_CQ;
  assign CLBLM_L_X8Y152_SLICE_X11Y152_B5 = CLBLM_R_X11Y153_SLICE_X15Y153_AQ;
  assign CLBLM_L_X8Y152_SLICE_X11Y152_B6 = CLBLL_L_X4Y142_SLICE_X5Y142_DQ;
  assign CLBLM_L_X8Y152_SLICE_X11Y152_C1 = CLBLM_L_X12Y149_SLICE_X17Y149_CO6;
  assign CLBLM_L_X8Y152_SLICE_X11Y152_C2 = CLBLM_L_X8Y152_SLICE_X11Y152_CQ;
  assign CLBLM_L_X8Y152_SLICE_X11Y152_C3 = CLBLM_R_X5Y153_SLICE_X6Y153_B5Q;
  assign CLBLM_L_X8Y152_SLICE_X11Y152_C4 = CLBLM_L_X8Y153_SLICE_X11Y153_BQ;
  assign CLBLM_L_X8Y152_SLICE_X11Y152_C5 = 1'b1;
  assign CLBLM_L_X8Y152_SLICE_X11Y152_C6 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_L_X8Y152_SLICE_X11Y152_CLK = CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O;
  assign CLBLM_L_X8Y152_SLICE_X11Y152_D1 = 1'b1;
  assign CLBLM_L_X8Y152_SLICE_X11Y152_D2 = CLBLM_L_X8Y152_SLICE_X11Y152_CQ;
  assign CLBLM_L_X8Y152_SLICE_X11Y152_D3 = CLBLM_R_X7Y146_SLICE_X8Y146_C5Q;
  assign CLBLM_L_X8Y152_SLICE_X11Y152_D4 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_L_X8Y152_SLICE_X11Y152_D5 = CLBLM_L_X10Y151_SLICE_X13Y151_AQ;
  assign CLBLM_L_X8Y152_SLICE_X11Y152_D6 = 1'b1;
  assign CLBLM_L_X8Y152_SLICE_X10Y152_A1 = CLBLM_R_X11Y153_SLICE_X14Y153_AQ;
  assign CLBLM_L_X8Y152_SLICE_X10Y152_A2 = CLBLM_L_X8Y152_SLICE_X10Y152_BQ;
  assign CLBLM_L_X8Y152_SLICE_X10Y152_A3 = CLBLM_L_X8Y152_SLICE_X10Y152_AQ;
  assign CLBLM_L_X8Y152_SLICE_X10Y152_A4 = RIOB33_X105Y131_IOB_X1Y131_I;
  assign CLBLM_L_X8Y152_SLICE_X10Y152_A5 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_L_X8Y152_SLICE_X10Y152_A6 = CLBLM_R_X7Y152_SLICE_X9Y152_AQ;
  assign CLBLM_L_X12Y152_SLICE_X16Y152_A4 = CLBLM_L_X8Y144_SLICE_X10Y144_BQ;
  assign CLBLM_L_X12Y152_SLICE_X16Y152_A5 = CLBLM_R_X11Y148_SLICE_X14Y148_BO6;
  assign CLBLM_L_X8Y152_SLICE_X10Y152_AX = CLBLM_L_X8Y154_SLICE_X10Y154_BO6;
  assign CLBLM_L_X8Y152_SLICE_X10Y152_B1 = CLBLM_R_X7Y148_SLICE_X9Y148_C5Q;
  assign CLBLM_L_X8Y152_SLICE_X10Y152_B2 = CLBLM_L_X8Y152_SLICE_X10Y152_BQ;
  assign CLBLM_L_X8Y152_SLICE_X10Y152_B3 = 1'b1;
  assign CLBLM_L_X8Y152_SLICE_X10Y152_B4 = RIOB33_X105Y131_IOB_X1Y131_I;
  assign CLBLM_L_X8Y152_SLICE_X10Y152_B5 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_L_X8Y152_SLICE_X10Y152_B6 = CLBLM_R_X7Y152_SLICE_X9Y152_AQ;
  assign CLBLM_L_X8Y152_SLICE_X10Y152_C1 = CLBLM_L_X8Y142_SLICE_X10Y142_A5Q;
  assign CLBLM_L_X8Y152_SLICE_X10Y152_C2 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_L_X8Y152_SLICE_X10Y152_C3 = CLBLM_R_X5Y153_SLICE_X7Y153_AQ;
  assign CLBLM_L_X8Y152_SLICE_X10Y152_C4 = CLBLM_L_X8Y151_SLICE_X10Y151_A5Q;
  assign CLBLM_L_X8Y152_SLICE_X10Y152_C5 = CLBLM_L_X10Y152_SLICE_X12Y152_DO6;
  assign CLBLM_L_X8Y152_SLICE_X10Y152_C6 = 1'b1;
  assign CLBLM_L_X8Y152_SLICE_X10Y152_CLK = CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O;
  assign CLBLM_L_X10Y154_SLICE_X13Y154_C3 = CLBLM_L_X10Y154_SLICE_X12Y154_BQ;
  assign CLBLM_L_X8Y152_SLICE_X10Y152_D1 = CLBLM_R_X7Y152_SLICE_X8Y152_B5Q;
  assign CLBLM_L_X8Y152_SLICE_X10Y152_D2 = CLBLM_R_X7Y152_SLICE_X9Y152_BQ;
  assign CLBLM_L_X8Y152_SLICE_X10Y152_D3 = CLBLM_L_X8Y152_SLICE_X10Y152_DQ;
  assign CLBLM_L_X8Y152_SLICE_X10Y152_D4 = CLBLM_R_X7Y152_SLICE_X8Y152_D5Q;
  assign CLBLM_L_X8Y152_SLICE_X10Y152_D5 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_L_X8Y152_SLICE_X10Y152_D6 = CLBLM_R_X7Y142_SLICE_X8Y142_C5Q;
  assign CLBLM_L_X10Y154_SLICE_X13Y154_CLK = CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O;
  assign LIOB33_X0Y165_IOB_X0Y166_O = RIOB33_SING_X105Y100_IOB_X1Y100_I;
  assign LIOB33_X0Y165_IOB_X0Y165_O = LIOB33_X0Y57_IOB_X0Y57_I;
  assign CLBLM_L_X12Y152_SLICE_X16Y152_C1 = 1'b1;
  assign CLBLM_R_X7Y146_SLICE_X9Y146_A1 = CLBLM_R_X7Y143_SLICE_X9Y143_B5Q;
  assign CLBLM_R_X7Y146_SLICE_X9Y146_A2 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X7Y146_SLICE_X9Y146_A3 = CLBLM_R_X7Y146_SLICE_X9Y146_AQ;
  assign CLBLM_R_X7Y146_SLICE_X9Y146_A4 = CLBLM_R_X5Y148_SLICE_X7Y148_C5Q;
  assign CLBLM_R_X7Y146_SLICE_X9Y146_A5 = CLBLM_L_X10Y145_SLICE_X12Y145_AQ;
  assign CLBLM_R_X7Y146_SLICE_X9Y146_A6 = CLBLM_R_X5Y142_SLICE_X7Y142_BQ;
  assign CLBLM_L_X10Y154_SLICE_X13Y154_D3 = CLBLM_L_X10Y155_SLICE_X13Y155_AO6;
  assign CLBLM_R_X7Y146_SLICE_X9Y146_B1 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X7Y146_SLICE_X9Y146_B2 = CLBLM_R_X7Y146_SLICE_X9Y146_BQ;
  assign CLBLM_R_X7Y146_SLICE_X9Y146_B3 = CLBLL_L_X4Y142_SLICE_X5Y142_DQ;
  assign CLBLM_L_X10Y154_SLICE_X13Y154_D4 = CLBLM_R_X7Y146_SLICE_X8Y146_A5Q;
  assign CLBLM_R_X7Y146_SLICE_X9Y146_B4 = CLBLM_R_X5Y152_SLICE_X7Y152_BQ;
  assign CLBLM_R_X7Y146_SLICE_X9Y146_B5 = CLBLM_R_X7Y144_SLICE_X8Y144_BQ;
  assign CLBLM_R_X7Y146_SLICE_X9Y146_B6 = CLBLL_L_X4Y147_SLICE_X5Y147_CQ;
  assign CLBLM_R_X7Y146_SLICE_X9Y146_C1 = CLBLM_R_X7Y149_SLICE_X8Y149_AQ;
  assign CLBLM_R_X7Y146_SLICE_X9Y146_C2 = CLBLM_L_X10Y146_SLICE_X12Y146_DQ;
  assign CLBLM_R_X7Y146_SLICE_X9Y146_C3 = CLBLM_R_X7Y151_SLICE_X8Y151_D5Q;
  assign CLBLM_R_X7Y146_SLICE_X9Y146_C4 = CLBLL_L_X4Y147_SLICE_X4Y147_CQ;
  assign CLBLM_R_X7Y146_SLICE_X9Y146_C5 = CLBLM_R_X5Y142_SLICE_X6Y142_D5Q;
  assign CLBLM_R_X7Y146_SLICE_X9Y146_C6 = 1'b1;
  assign LIOI3_X0Y165_OLOGIC_X0Y166_D1 = RIOB33_SING_X105Y100_IOB_X1Y100_I;
  assign CLBLM_R_X7Y146_SLICE_X9Y146_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign LIOI3_X0Y165_OLOGIC_X0Y166_T1 = 1'b1;
  assign CLBLM_R_X7Y146_SLICE_X9Y146_D1 = CLBLM_R_X7Y149_SLICE_X8Y149_AQ;
  assign CLBLM_R_X7Y146_SLICE_X9Y146_D2 = CLBLM_L_X10Y146_SLICE_X12Y146_DQ;
  assign CLBLM_R_X7Y146_SLICE_X9Y146_D3 = CLBLM_R_X7Y151_SLICE_X8Y151_D5Q;
  assign CLBLM_R_X7Y146_SLICE_X9Y146_D4 = CLBLL_L_X4Y147_SLICE_X4Y147_CQ;
  assign CLBLM_R_X7Y146_SLICE_X9Y146_D5 = CLBLM_R_X5Y142_SLICE_X6Y142_D5Q;
  assign CLBLM_R_X7Y146_SLICE_X9Y146_D6 = CLBLM_R_X11Y146_SLICE_X15Y146_BO6;
  assign LIOI3_X0Y103_OLOGIC_X0Y104_D1 = CLBLM_R_X3Y145_SLICE_X2Y145_C5Q;
  assign LIOI3_X0Y145_OLOGIC_X0Y146_D1 = CLBLM_R_X3Y143_SLICE_X3Y143_DO6;
  assign LIOI3_X0Y165_OLOGIC_X0Y165_D1 = LIOB33_X0Y57_IOB_X0Y57_I;
  assign CLBLM_R_X7Y146_SLICE_X8Y146_A1 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X7Y146_SLICE_X8Y146_A2 = CLBLM_R_X3Y147_SLICE_X2Y147_CQ;
  assign CLBLL_L_X2Y145_SLICE_X0Y145_A1 = CLBLM_R_X5Y142_SLICE_X6Y142_D5Q;
  assign CLBLL_L_X2Y145_SLICE_X0Y145_A2 = CLBLL_L_X2Y146_SLICE_X0Y146_BQ;
  assign CLBLL_L_X2Y145_SLICE_X0Y145_A3 = CLBLL_L_X2Y145_SLICE_X0Y145_AQ;
  assign CLBLL_L_X2Y145_SLICE_X0Y145_A4 = CLBLL_L_X2Y146_SLICE_X0Y146_AQ;
  assign CLBLL_L_X2Y145_SLICE_X0Y145_A5 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLL_L_X2Y145_SLICE_X0Y145_A6 = CLBLM_R_X3Y146_SLICE_X2Y146_CQ;
  assign CLBLM_R_X7Y146_SLICE_X8Y146_A3 = CLBLM_R_X3Y146_SLICE_X2Y146_C5Q;
  assign CLBLM_R_X7Y146_SLICE_X8Y146_A4 = CLBLM_L_X8Y150_SLICE_X10Y150_AQ;
  assign CLBLM_R_X7Y146_SLICE_X8Y146_A5 = CLBLM_R_X7Y142_SLICE_X8Y142_AQ;
  assign CLBLL_L_X2Y145_SLICE_X0Y145_B1 = 1'b1;
  assign CLBLL_L_X2Y145_SLICE_X0Y145_B2 = CLBLL_L_X2Y146_SLICE_X0Y146_BQ;
  assign CLBLL_L_X2Y145_SLICE_X0Y145_B3 = CLBLL_L_X2Y145_SLICE_X0Y145_AQ;
  assign CLBLL_L_X2Y145_SLICE_X0Y145_B4 = CLBLL_L_X2Y146_SLICE_X0Y146_AQ;
  assign CLBLL_L_X2Y145_SLICE_X0Y145_B5 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLL_L_X2Y145_SLICE_X0Y145_B6 = CLBLM_R_X5Y144_SLICE_X7Y144_B5Q;
  assign CLBLM_R_X7Y146_SLICE_X8Y146_B1 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X7Y146_SLICE_X8Y146_B2 = CLBLM_R_X7Y142_SLICE_X8Y142_BQ;
  assign CLBLL_L_X2Y145_SLICE_X0Y145_C1 = 1'b1;
  assign CLBLL_L_X2Y145_SLICE_X0Y145_C2 = 1'b1;
  assign CLBLL_L_X2Y145_SLICE_X0Y145_C3 = 1'b1;
  assign CLBLL_L_X2Y145_SLICE_X0Y145_C4 = 1'b1;
  assign CLBLL_L_X2Y145_SLICE_X0Y145_C5 = 1'b1;
  assign CLBLL_L_X2Y145_SLICE_X0Y145_C6 = 1'b1;
  assign CLBLM_R_X7Y146_SLICE_X8Y146_C1 = CLBLM_R_X7Y147_SLICE_X8Y147_AQ;
  assign CLBLL_L_X2Y145_SLICE_X0Y145_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X7Y146_SLICE_X8Y146_C2 = CLBLM_R_X5Y146_SLICE_X7Y146_CQ;
  assign CLBLM_R_X7Y146_SLICE_X8Y146_C3 = CLBLL_L_X4Y153_SLICE_X4Y153_AQ;
  assign CLBLM_R_X7Y146_SLICE_X8Y146_C4 = CLBLM_R_X5Y140_SLICE_X6Y140_A5Q;
  assign CLBLM_R_X7Y146_SLICE_X8Y146_C5 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X7Y146_SLICE_X8Y146_C6 = 1'b1;
  assign CLBLL_L_X2Y145_SLICE_X0Y145_D1 = 1'b1;
  assign CLBLL_L_X2Y145_SLICE_X0Y145_D2 = 1'b1;
  assign CLBLL_L_X2Y145_SLICE_X0Y145_D3 = 1'b1;
  assign CLBLL_L_X2Y145_SLICE_X0Y145_D4 = 1'b1;
  assign CLBLL_L_X2Y145_SLICE_X0Y145_D5 = 1'b1;
  assign CLBLL_L_X2Y145_SLICE_X0Y145_D6 = 1'b1;
  assign CLBLM_L_X10Y154_SLICE_X12Y154_A6 = CLBLM_L_X10Y154_SLICE_X13Y154_DO6;
  assign CLBLM_R_X7Y146_SLICE_X8Y146_D1 = CLBLM_R_X7Y153_SLICE_X9Y153_A5Q;
  assign CLBLM_R_X7Y146_SLICE_X8Y146_D2 = CLBLM_R_X5Y145_SLICE_X7Y145_A5Q;
  assign CLBLM_R_X7Y146_SLICE_X8Y146_D3 = CLBLM_R_X7Y145_SLICE_X8Y145_A5Q;
  assign CLBLM_R_X7Y146_SLICE_X8Y146_D4 = CLBLM_R_X5Y147_SLICE_X6Y147_B5Q;
  assign CLBLM_R_X7Y146_SLICE_X8Y146_D5 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X7Y146_SLICE_X8Y146_D6 = 1'b1;
  assign LIOI3_X0Y145_OLOGIC_X0Y146_T1 = 1'b1;
  assign CLBLL_L_X2Y145_SLICE_X1Y145_A1 = CLBLL_L_X2Y146_SLICE_X1Y146_DO6;
  assign CLBLL_L_X2Y145_SLICE_X1Y145_A2 = CLBLM_R_X3Y146_SLICE_X2Y146_BQ;
  assign CLBLL_L_X2Y145_SLICE_X1Y145_A3 = CLBLL_L_X2Y145_SLICE_X1Y145_AQ;
  assign CLBLL_L_X2Y145_SLICE_X1Y145_A4 = CLBLL_L_X4Y143_SLICE_X4Y143_D5Q;
  assign CLBLL_L_X2Y145_SLICE_X1Y145_A5 = CLBLM_R_X5Y143_SLICE_X6Y143_C5Q;
  assign CLBLL_L_X2Y145_SLICE_X1Y145_A6 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLL_L_X2Y145_SLICE_X1Y145_B1 = CLBLL_L_X2Y145_SLICE_X1Y145_DO6;
  assign CLBLL_L_X2Y145_SLICE_X1Y145_B2 = CLBLL_L_X2Y146_SLICE_X0Y146_AQ;
  assign CLBLL_L_X2Y145_SLICE_X1Y145_B3 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLL_L_X2Y145_SLICE_X1Y145_B4 = CLBLL_L_X4Y143_SLICE_X4Y143_D5Q;
  assign CLBLL_L_X2Y145_SLICE_X1Y145_B5 = CLBLL_L_X2Y145_SLICE_X1Y145_BQ;
  assign CLBLL_L_X2Y145_SLICE_X1Y145_B6 = 1'b1;
  assign CLBLL_L_X2Y145_SLICE_X1Y145_C1 = CLBLL_L_X4Y143_SLICE_X4Y143_D5Q;
  assign CLBLL_L_X2Y145_SLICE_X1Y145_C2 = CLBLL_L_X2Y145_SLICE_X1Y145_CQ;
  assign CLBLL_L_X2Y145_SLICE_X1Y145_C3 = CLBLL_L_X4Y145_SLICE_X4Y145_C5Q;
  assign CLBLL_L_X2Y145_SLICE_X1Y145_C4 = CLBLL_L_X2Y146_SLICE_X1Y146_CO6;
  assign CLBLL_L_X2Y145_SLICE_X1Y145_C5 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLL_L_X2Y145_SLICE_X1Y145_C6 = CLBLL_L_X2Y145_SLICE_X1Y145_DO5;
  assign CLBLL_L_X2Y145_SLICE_X1Y145_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLL_L_X2Y145_SLICE_X1Y145_D1 = CLBLL_L_X2Y145_SLICE_X1Y145_BQ;
  assign CLBLL_L_X2Y145_SLICE_X1Y145_D2 = CLBLL_L_X2Y145_SLICE_X1Y145_CQ;
  assign CLBLL_L_X2Y145_SLICE_X1Y145_D3 = CLBLL_L_X2Y146_SLICE_X1Y146_DO6;
  assign CLBLL_L_X2Y145_SLICE_X1Y145_D4 = CLBLL_L_X2Y145_SLICE_X1Y145_AQ;
  assign CLBLL_L_X2Y145_SLICE_X1Y145_D5 = CLBLM_R_X3Y146_SLICE_X2Y146_BQ;
  assign CLBLL_L_X2Y145_SLICE_X1Y145_D6 = 1'b1;
  assign CLBLM_L_X10Y154_SLICE_X12Y154_BX = CLBLM_L_X10Y154_SLICE_X12Y154_DO6;
  assign LIOI3_X0Y145_OLOGIC_X0Y145_D1 = CLBLM_R_X3Y148_SLICE_X3Y148_DO6;
  assign CLBLM_L_X8Y153_SLICE_X11Y153_A1 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_L_X8Y153_SLICE_X11Y153_A2 = CLBLM_R_X11Y153_SLICE_X14Y153_A5Q;
  assign CLBLM_L_X8Y153_SLICE_X11Y153_A3 = CLBLM_L_X8Y153_SLICE_X11Y153_AQ;
  assign CLBLM_L_X8Y153_SLICE_X11Y153_A4 = CLBLM_L_X10Y153_SLICE_X12Y153_CO5;
  assign CLBLM_L_X8Y153_SLICE_X11Y153_A5 = CLBLM_L_X8Y154_SLICE_X11Y154_AQ;
  assign CLBLM_L_X8Y153_SLICE_X11Y153_A6 = CLBLM_R_X5Y150_SLICE_X6Y150_B5Q;
  assign CLBLM_L_X10Y154_SLICE_X12Y154_C1 = CLBLM_L_X10Y155_SLICE_X13Y155_BO6;
  assign CLBLM_L_X8Y153_SLICE_X11Y153_B1 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_L_X8Y153_SLICE_X11Y153_B2 = CLBLM_L_X8Y153_SLICE_X11Y153_BQ;
  assign CLBLM_L_X8Y153_SLICE_X11Y153_B3 = CLBLM_R_X3Y145_SLICE_X3Y145_D5Q;
  assign CLBLM_L_X8Y153_SLICE_X11Y153_B4 = CLBLM_L_X10Y154_SLICE_X12Y154_A5Q;
  assign CLBLM_L_X8Y153_SLICE_X11Y153_B5 = CLBLL_L_X4Y151_SLICE_X4Y151_BQ;
  assign CLBLM_L_X8Y153_SLICE_X11Y153_B6 = CLBLM_L_X8Y153_SLICE_X10Y153_CQ;
  assign CLBLM_L_X10Y154_SLICE_X12Y154_C2 = CLBLM_L_X10Y155_SLICE_X13Y155_CO6;
  assign CLBLM_L_X10Y154_SLICE_X12Y154_C3 = CLBLM_R_X3Y150_SLICE_X2Y150_BQ;
  assign CLBLM_L_X8Y153_SLICE_X11Y153_C1 = CLBLM_R_X7Y153_SLICE_X9Y153_C5Q;
  assign CLBLM_L_X8Y153_SLICE_X11Y153_C2 = CLBLM_L_X10Y153_SLICE_X12Y153_BQ;
  assign CLBLM_L_X8Y153_SLICE_X11Y153_C3 = CLBLM_R_X7Y154_SLICE_X8Y154_DO6;
  assign CLBLM_L_X8Y153_SLICE_X11Y153_C4 = CLBLM_L_X10Y153_SLICE_X12Y153_AQ;
  assign CLBLM_L_X8Y153_SLICE_X11Y153_C5 = CLBLM_L_X8Y146_SLICE_X11Y146_BQ;
  assign CLBLM_L_X8Y153_SLICE_X11Y153_C6 = CLBLM_R_X7Y151_SLICE_X9Y151_D5Q;
  assign CLBLM_L_X8Y153_SLICE_X11Y153_CLK = CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O;
  assign CLBLM_L_X8Y153_SLICE_X11Y153_D1 = CLBLM_R_X7Y145_SLICE_X8Y145_A5Q;
  assign CLBLM_L_X8Y153_SLICE_X11Y153_D2 = CLBLL_L_X4Y153_SLICE_X5Y153_A5Q;
  assign CLBLM_L_X8Y153_SLICE_X11Y153_D3 = 1'b1;
  assign CLBLM_L_X8Y153_SLICE_X11Y153_D4 = 1'b1;
  assign CLBLM_L_X8Y153_SLICE_X11Y153_D5 = CLBLM_L_X8Y145_SLICE_X11Y145_DQ;
  assign CLBLM_L_X8Y153_SLICE_X11Y153_D6 = RIOB33_X105Y131_IOB_X1Y131_I;
  assign CLBLM_L_X8Y153_SLICE_X10Y153_A1 = CLBLM_R_X7Y155_SLICE_X8Y155_A5Q;
  assign CLBLM_L_X8Y153_SLICE_X10Y153_A2 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_L_X8Y153_SLICE_X10Y153_A3 = CLBLM_R_X5Y153_SLICE_X7Y153_DO6;
  assign CLBLM_L_X8Y153_SLICE_X10Y153_A4 = CLBLM_L_X10Y152_SLICE_X12Y152_BQ;
  assign CLBLM_L_X8Y153_SLICE_X10Y153_A5 = CLBLM_L_X10Y147_SLICE_X13Y147_AQ;
  assign CLBLM_L_X8Y153_SLICE_X10Y153_A6 = 1'b1;
  assign LIOI3_X0Y145_OLOGIC_X0Y145_T1 = 1'b1;
  assign CLBLM_L_X8Y153_SLICE_X10Y153_B1 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_L_X8Y153_SLICE_X10Y153_B2 = CLBLM_L_X8Y153_SLICE_X10Y153_A5Q;
  assign CLBLM_L_X8Y153_SLICE_X10Y153_B3 = 1'b1;
  assign CLBLM_L_X8Y153_SLICE_X10Y153_B4 = CLBLM_R_X7Y152_SLICE_X9Y152_CQ;
  assign CLBLM_L_X8Y153_SLICE_X10Y153_B5 = CLBLM_L_X10Y153_SLICE_X13Y153_A5Q;
  assign CLBLM_L_X8Y153_SLICE_X10Y153_B6 = 1'b1;
  assign CLBLM_L_X8Y153_SLICE_X10Y153_C1 = CLBLM_R_X3Y150_SLICE_X2Y150_D5Q;
  assign CLBLM_L_X8Y153_SLICE_X10Y153_C2 = CLBLL_L_X4Y143_SLICE_X4Y143_AQ;
  assign CLBLM_L_X8Y153_SLICE_X10Y153_C3 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_L_X8Y153_SLICE_X10Y153_C4 = CLBLM_R_X7Y153_SLICE_X9Y153_BQ;
  assign CLBLM_L_X8Y153_SLICE_X10Y153_C5 = CLBLM_L_X8Y153_SLICE_X10Y153_B5Q;
  assign CLBLM_L_X8Y153_SLICE_X10Y153_C6 = 1'b1;
  assign CLBLM_L_X8Y153_SLICE_X10Y153_CLK = CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O;
  assign CLBLM_L_X8Y153_SLICE_X10Y153_D1 = 1'b1;
  assign CLBLM_L_X8Y153_SLICE_X10Y153_D2 = CLBLM_L_X10Y151_SLICE_X13Y151_A5Q;
  assign CLBLM_L_X8Y153_SLICE_X10Y153_D3 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_L_X8Y153_SLICE_X10Y153_D4 = CLBLM_L_X10Y145_SLICE_X12Y145_BQ;
  assign CLBLM_L_X8Y153_SLICE_X10Y153_D5 = CLBLM_R_X3Y149_SLICE_X3Y149_AQ;
  assign CLBLM_L_X8Y153_SLICE_X10Y153_D6 = 1'b1;
  assign CLBLM_R_X11Y150_SLICE_X15Y150_C4 = 1'b1;
  assign RIOI3_X105Y147_ILOGIC_X1Y148_D = RIOB33_X105Y147_IOB_X1Y148_I;
  assign CLBLM_R_X11Y150_SLICE_X15Y150_C5 = CLBLM_R_X11Y151_SLICE_X14Y151_DO6;
  assign CLBLM_L_X10Y154_SLICE_X12Y154_D3 = RIOB33_SING_X105Y100_IOB_X1Y100_I;
  assign RIOI3_X105Y147_ILOGIC_X1Y147_D = RIOB33_X105Y147_IOB_X1Y147_I;
  assign CLBLM_R_X11Y150_SLICE_X15Y150_C6 = CLBLM_L_X8Y151_SLICE_X11Y151_BO6;
  assign CLBLM_L_X10Y154_SLICE_X12Y154_D4 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign LIOB33_X0Y167_IOB_X0Y168_O = RIOB33_X105Y101_IOB_X1Y101_I;
  assign LIOB33_X0Y167_IOB_X0Y167_O = RIOB33_X105Y105_IOB_X1Y106_I;
  assign CLBLM_L_X10Y154_SLICE_X12Y154_D6 = 1'b1;
  assign CLBLM_R_X7Y147_SLICE_X9Y147_A1 = CLBLM_R_X3Y145_SLICE_X3Y145_BQ;
  assign CLBLM_R_X7Y147_SLICE_X9Y147_A2 = CLBLM_R_X7Y146_SLICE_X8Y146_B5Q;
  assign CLBLM_R_X7Y147_SLICE_X9Y147_A3 = CLBLM_R_X3Y146_SLICE_X2Y146_D5Q;
  assign CLBLM_R_X7Y147_SLICE_X9Y147_A4 = CLBLM_R_X3Y149_SLICE_X2Y149_BQ;
  assign CLBLM_R_X7Y147_SLICE_X9Y147_A5 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X7Y147_SLICE_X9Y147_A6 = 1'b1;
  assign CLBLM_R_X7Y147_SLICE_X9Y147_B1 = CLBLL_L_X4Y151_SLICE_X4Y151_BQ;
  assign CLBLM_R_X7Y147_SLICE_X9Y147_B2 = CLBLM_R_X7Y147_SLICE_X9Y147_BQ;
  assign CLBLM_R_X7Y147_SLICE_X9Y147_B3 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X7Y147_SLICE_X9Y147_B4 = CLBLM_L_X8Y147_SLICE_X10Y147_C5Q;
  assign CLBLM_R_X7Y147_SLICE_X9Y147_B5 = CLBLM_L_X10Y144_SLICE_X13Y144_CQ;
  assign CLBLM_R_X7Y147_SLICE_X9Y147_B6 = CLBLM_R_X7Y147_SLICE_X9Y147_A5Q;
  assign CLBLM_R_X7Y147_SLICE_X9Y147_C1 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X7Y147_SLICE_X9Y147_C2 = CLBLM_R_X5Y145_SLICE_X6Y145_CQ;
  assign CLBLM_R_X7Y147_SLICE_X9Y147_C3 = CLBLM_R_X7Y146_SLICE_X9Y146_BQ;
  assign CLBLM_R_X7Y147_SLICE_X9Y147_C4 = CLBLM_L_X8Y146_SLICE_X11Y146_AQ;
  assign CLBLM_R_X7Y147_SLICE_X9Y147_C5 = CLBLL_L_X4Y150_SLICE_X4Y150_B5Q;
  assign CLBLM_R_X7Y147_SLICE_X9Y147_C6 = 1'b1;
  assign CLBLM_R_X11Y150_SLICE_X15Y150_D5 = CLBLM_L_X12Y149_SLICE_X17Y149_BO5;
  assign CLBLM_R_X7Y147_SLICE_X9Y147_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X11Y150_SLICE_X15Y150_D6 = 1'b1;
  assign CLBLM_R_X7Y147_SLICE_X9Y147_D1 = CLBLM_L_X8Y147_SLICE_X10Y147_AQ;
  assign CLBLM_R_X7Y147_SLICE_X9Y147_D2 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X7Y147_SLICE_X9Y147_D3 = CLBLM_L_X10Y151_SLICE_X13Y151_AQ;
  assign CLBLM_R_X7Y147_SLICE_X9Y147_D4 = CLBLL_L_X4Y149_SLICE_X5Y149_AQ;
  assign CLBLM_R_X7Y147_SLICE_X9Y147_D5 = 1'b1;
  assign CLBLM_R_X7Y147_SLICE_X9Y147_D6 = 1'b1;
  assign CLBLL_L_X2Y146_SLICE_X0Y146_A1 = CLBLL_L_X4Y146_SLICE_X4Y146_B5Q;
  assign CLBLL_L_X2Y146_SLICE_X0Y146_A2 = CLBLL_L_X2Y146_SLICE_X0Y146_BQ;
  assign CLBLL_L_X2Y146_SLICE_X0Y146_A3 = CLBLL_L_X2Y146_SLICE_X0Y146_AQ;
  assign CLBLL_L_X2Y146_SLICE_X0Y146_A4 = CLBLM_R_X3Y146_SLICE_X2Y146_CQ;
  assign CLBLL_L_X2Y146_SLICE_X0Y146_A5 = CLBLL_L_X2Y145_SLICE_X0Y145_AQ;
  assign CLBLL_L_X2Y146_SLICE_X0Y146_A6 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X7Y147_SLICE_X8Y147_A1 = CLBLM_R_X7Y145_SLICE_X8Y145_DQ;
  assign CLBLM_R_X7Y147_SLICE_X8Y147_A2 = CLBLM_L_X8Y145_SLICE_X10Y145_A5Q;
  assign CLBLM_R_X7Y147_SLICE_X8Y147_A3 = CLBLM_R_X7Y147_SLICE_X9Y147_C5Q;
  assign CLBLL_L_X2Y146_SLICE_X0Y146_B1 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLL_L_X2Y146_SLICE_X0Y146_B2 = CLBLL_L_X2Y146_SLICE_X0Y146_BQ;
  assign CLBLL_L_X2Y146_SLICE_X0Y146_B3 = CLBLL_L_X2Y146_SLICE_X0Y146_AQ;
  assign CLBLL_L_X2Y146_SLICE_X0Y146_B4 = CLBLM_R_X3Y146_SLICE_X2Y146_CQ;
  assign CLBLL_L_X2Y146_SLICE_X0Y146_B5 = CLBLL_L_X2Y145_SLICE_X0Y145_AQ;
  assign CLBLL_L_X2Y146_SLICE_X0Y146_B6 = CLBLM_R_X3Y147_SLICE_X2Y147_BQ;
  assign CLBLM_R_X7Y147_SLICE_X8Y147_A5 = CLBLM_R_X7Y145_SLICE_X8Y145_CQ;
  assign CLBLM_R_X7Y147_SLICE_X8Y147_A6 = CLBLM_R_X3Y150_SLICE_X3Y150_DQ;
  assign CLBLM_L_X10Y144_SLICE_X13Y144_A5 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLL_L_X2Y146_SLICE_X0Y146_C1 = CLBLL_L_X2Y145_SLICE_X0Y145_AQ;
  assign CLBLL_L_X2Y146_SLICE_X0Y146_C2 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLL_L_X2Y146_SLICE_X0Y146_C3 = CLBLL_L_X2Y146_SLICE_X0Y146_AQ;
  assign CLBLL_L_X2Y146_SLICE_X0Y146_C4 = CLBLL_L_X2Y146_SLICE_X0Y146_BQ;
  assign CLBLL_L_X2Y146_SLICE_X0Y146_C5 = 1'b1;
  assign CLBLL_L_X2Y146_SLICE_X0Y146_C6 = CLBLL_L_X4Y149_SLICE_X4Y149_D5Q;
  assign CLBLM_R_X7Y147_SLICE_X8Y147_B4 = CLBLM_R_X7Y153_SLICE_X8Y153_A5Q;
  assign CLBLM_R_X7Y147_SLICE_X8Y147_B5 = CLBLM_R_X7Y144_SLICE_X9Y144_B5Q;
  assign CLBLL_L_X2Y146_SLICE_X0Y146_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X7Y147_SLICE_X8Y147_C1 = CLBLM_R_X7Y144_SLICE_X9Y144_B5Q;
  assign CLBLM_R_X7Y147_SLICE_X8Y147_C2 = CLBLM_R_X7Y153_SLICE_X8Y153_A5Q;
  assign CLBLM_R_X7Y147_SLICE_X8Y147_C3 = CLBLM_R_X7Y144_SLICE_X8Y144_B5Q;
  assign CLBLM_R_X7Y147_SLICE_X8Y147_C4 = 1'b1;
  assign CLBLL_L_X2Y146_SLICE_X0Y146_D1 = CLBLM_R_X3Y144_SLICE_X3Y144_AQ;
  assign CLBLL_L_X2Y146_SLICE_X0Y146_D2 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLL_L_X2Y146_SLICE_X0Y146_D3 = CLBLL_L_X2Y146_SLICE_X1Y146_B5Q;
  assign CLBLL_L_X2Y146_SLICE_X0Y146_D4 = CLBLM_R_X3Y145_SLICE_X3Y145_CQ;
  assign CLBLL_L_X2Y146_SLICE_X0Y146_D5 = CLBLM_R_X5Y153_SLICE_X6Y153_B5Q;
  assign CLBLL_L_X2Y146_SLICE_X0Y146_D6 = CLBLM_R_X5Y145_SLICE_X6Y145_BQ;
  assign CLBLM_L_X10Y144_SLICE_X13Y144_AX = CLBLM_L_X10Y144_SLICE_X12Y144_BO5;
  assign CLBLM_R_X7Y147_SLICE_X8Y147_D1 = CLBLM_R_X7Y147_SLICE_X8Y147_CO6;
  assign CLBLM_R_X7Y147_SLICE_X8Y147_D2 = CLBLM_R_X11Y147_SLICE_X14Y147_AO6;
  assign CLBLM_R_X7Y147_SLICE_X8Y147_D3 = CLBLM_L_X8Y150_SLICE_X11Y150_BO6;
  assign CLBLM_R_X7Y147_SLICE_X8Y147_D4 = CLBLM_R_X5Y145_SLICE_X6Y145_CQ;
  assign CLBLM_R_X7Y147_SLICE_X8Y147_D5 = 1'b1;
  assign CLBLM_R_X7Y147_SLICE_X8Y147_D6 = CLBLM_R_X7Y142_SLICE_X8Y142_BQ;
  assign CLBLM_L_X10Y144_SLICE_X13Y144_B2 = CLBLM_L_X10Y144_SLICE_X13Y144_BQ;
  assign RIOI3_X105Y123_ILOGIC_X1Y123_D = RIOB33_X105Y123_IOB_X1Y123_I;
  assign CLBLL_L_X2Y146_SLICE_X1Y146_A1 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLL_L_X2Y146_SLICE_X1Y146_A2 = CLBLL_L_X4Y143_SLICE_X4Y143_D5Q;
  assign CLBLL_L_X2Y146_SLICE_X1Y146_A3 = CLBLL_L_X2Y146_SLICE_X1Y146_AQ;
  assign CLBLL_L_X2Y146_SLICE_X1Y146_A4 = CLBLM_L_X8Y144_SLICE_X11Y144_BQ;
  assign CLBLL_L_X2Y146_SLICE_X1Y146_A5 = 1'b1;
  assign CLBLL_L_X2Y146_SLICE_X1Y146_A6 = CLBLL_L_X4Y149_SLICE_X5Y149_CQ;
  assign CLBLM_R_X7Y152_SLICE_X9Y152_C4 = CLBLM_L_X8Y153_SLICE_X10Y153_BQ;
  assign CLBLM_R_X7Y152_SLICE_X9Y152_C5 = CLBLM_R_X7Y146_SLICE_X8Y146_C5Q;
  assign CLBLL_L_X2Y146_SLICE_X1Y146_B1 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLL_L_X2Y146_SLICE_X1Y146_B2 = CLBLM_R_X5Y150_SLICE_X6Y150_AQ;
  assign CLBLL_L_X2Y146_SLICE_X1Y146_B3 = CLBLL_L_X4Y147_SLICE_X4Y147_CQ;
  assign CLBLL_L_X2Y146_SLICE_X1Y146_B4 = CLBLM_R_X3Y144_SLICE_X2Y144_CO6;
  assign CLBLL_L_X2Y146_SLICE_X1Y146_B5 = CLBLL_L_X2Y148_SLICE_X1Y148_AO6;
  assign CLBLL_L_X2Y146_SLICE_X1Y146_B6 = 1'b1;
  assign CLBLM_R_X7Y152_SLICE_X9Y152_C6 = 1'b1;
  assign CLBLL_L_X2Y146_SLICE_X1Y146_C1 = CLBLL_L_X2Y146_SLICE_X1Y146_AQ;
  assign CLBLL_L_X2Y146_SLICE_X1Y146_C2 = CLBLM_R_X3Y149_SLICE_X2Y149_BQ;
  assign CLBLL_L_X2Y146_SLICE_X1Y146_C3 = CLBLL_L_X4Y149_SLICE_X4Y149_AQ;
  assign CLBLL_L_X2Y146_SLICE_X1Y146_C4 = CLBLL_L_X4Y149_SLICE_X5Y149_CQ;
  assign CLBLL_L_X2Y146_SLICE_X1Y146_C5 = CLBLM_R_X3Y147_SLICE_X2Y147_CQ;
  assign CLBLL_L_X2Y146_SLICE_X1Y146_C6 = 1'b1;
  assign CLBLL_L_X2Y146_SLICE_X1Y146_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLL_L_X2Y146_SLICE_X1Y146_D1 = CLBLL_L_X2Y145_SLICE_X1Y145_CQ;
  assign CLBLL_L_X2Y146_SLICE_X1Y146_D2 = CLBLL_L_X4Y149_SLICE_X5Y149_CQ;
  assign CLBLL_L_X2Y146_SLICE_X1Y146_D3 = CLBLL_L_X4Y149_SLICE_X4Y149_AQ;
  assign CLBLL_L_X2Y146_SLICE_X1Y146_D4 = CLBLM_R_X3Y147_SLICE_X2Y147_CQ;
  assign CLBLL_L_X2Y146_SLICE_X1Y146_D5 = CLBLL_L_X2Y146_SLICE_X1Y146_AQ;
  assign CLBLL_L_X2Y146_SLICE_X1Y146_D6 = CLBLM_R_X3Y149_SLICE_X2Y149_BQ;
  assign CLBLM_L_X8Y154_SLICE_X11Y154_A1 = CLBLM_L_X10Y153_SLICE_X12Y153_A5Q;
  assign CLBLM_L_X8Y154_SLICE_X11Y154_A2 = CLBLM_L_X10Y155_SLICE_X12Y155_AQ;
  assign CLBLM_L_X8Y154_SLICE_X11Y154_A3 = CLBLM_L_X8Y154_SLICE_X11Y154_AQ;
  assign CLBLM_L_X8Y154_SLICE_X11Y154_A4 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_L_X8Y154_SLICE_X11Y154_A5 = CLBLM_R_X5Y152_SLICE_X6Y152_BQ;
  assign CLBLM_L_X8Y154_SLICE_X11Y154_A6 = CLBLM_R_X5Y150_SLICE_X6Y150_B5Q;
  assign CLBLM_L_X8Y154_SLICE_X11Y154_B1 = 1'b1;
  assign CLBLM_L_X8Y154_SLICE_X11Y154_B2 = 1'b1;
  assign CLBLM_L_X8Y154_SLICE_X11Y154_B3 = 1'b1;
  assign CLBLM_L_X8Y154_SLICE_X11Y154_B4 = 1'b1;
  assign CLBLM_L_X8Y154_SLICE_X11Y154_B5 = 1'b1;
  assign CLBLM_L_X8Y154_SLICE_X11Y154_B6 = 1'b1;
  assign CLBLM_R_X7Y152_SLICE_X9Y152_D2 = CLBLM_R_X7Y152_SLICE_X9Y152_AQ;
  assign CLBLM_R_X7Y152_SLICE_X9Y152_D3 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_L_X8Y154_SLICE_X11Y154_C1 = 1'b1;
  assign CLBLM_L_X8Y154_SLICE_X11Y154_C2 = 1'b1;
  assign CLBLM_L_X8Y154_SLICE_X11Y154_C3 = 1'b1;
  assign CLBLM_L_X8Y154_SLICE_X11Y154_C4 = 1'b1;
  assign CLBLM_L_X8Y154_SLICE_X11Y154_C5 = 1'b1;
  assign CLBLM_L_X8Y154_SLICE_X11Y154_C6 = 1'b1;
  assign CLBLM_L_X8Y154_SLICE_X11Y154_CLK = CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O;
  assign CLBLM_R_X7Y152_SLICE_X9Y152_D5 = CLBLM_L_X8Y152_SLICE_X10Y152_AQ;
  assign CLBLM_R_X7Y152_SLICE_X9Y152_D6 = 1'b1;
  assign CLBLM_L_X8Y154_SLICE_X11Y154_D1 = 1'b1;
  assign CLBLM_L_X8Y154_SLICE_X11Y154_D2 = 1'b1;
  assign CLBLM_L_X8Y154_SLICE_X11Y154_D3 = 1'b1;
  assign CLBLM_L_X8Y154_SLICE_X11Y154_D4 = 1'b1;
  assign CLBLM_L_X8Y154_SLICE_X11Y154_D5 = 1'b1;
  assign CLBLM_L_X8Y154_SLICE_X11Y154_D6 = 1'b1;
  assign CLBLM_L_X8Y154_SLICE_X10Y154_A1 = CLBLM_R_X7Y155_SLICE_X8Y155_BO5;
  assign CLBLM_L_X8Y154_SLICE_X10Y154_A2 = CLBLM_L_X10Y154_SLICE_X13Y154_AQ;
  assign CLBLM_L_X8Y154_SLICE_X10Y154_A3 = CLBLM_L_X8Y154_SLICE_X10Y154_AQ;
  assign CLBLM_L_X8Y154_SLICE_X10Y154_A4 = CLBLM_R_X7Y154_SLICE_X8Y154_AQ;
  assign CLBLM_L_X8Y154_SLICE_X10Y154_A5 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_L_X8Y154_SLICE_X10Y154_A6 = CLBLM_R_X5Y150_SLICE_X6Y150_B5Q;
  assign CLBLM_L_X8Y154_SLICE_X10Y154_B1 = CLBLM_L_X10Y154_SLICE_X12Y154_B5Q;
  assign CLBLM_L_X8Y154_SLICE_X10Y154_B2 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_L_X8Y154_SLICE_X10Y154_B3 = CLBLM_R_X5Y142_SLICE_X7Y142_CO6;
  assign CLBLM_L_X8Y154_SLICE_X10Y154_B4 = CLBLM_L_X8Y153_SLICE_X10Y153_B5Q;
  assign CLBLM_L_X8Y154_SLICE_X10Y154_B5 = RIOB33_X105Y131_IOB_X1Y131_I;
  assign CLBLM_L_X8Y154_SLICE_X10Y154_B6 = 1'b1;
  assign CLBLM_L_X8Y154_SLICE_X10Y154_C1 = 1'b1;
  assign CLBLM_L_X8Y154_SLICE_X10Y154_C2 = 1'b1;
  assign CLBLM_L_X8Y154_SLICE_X10Y154_C3 = 1'b1;
  assign CLBLM_L_X8Y154_SLICE_X10Y154_C4 = 1'b1;
  assign CLBLM_L_X8Y154_SLICE_X10Y154_C5 = 1'b1;
  assign CLBLM_L_X8Y154_SLICE_X10Y154_C6 = 1'b1;
  assign LIOB33_X0Y169_IOB_X0Y170_O = RIOB33_X105Y117_IOB_X1Y118_I;
  assign LIOB33_X0Y169_IOB_X0Y169_O = RIOB33_X105Y117_IOB_X1Y117_I;
  assign CLBLM_L_X8Y154_SLICE_X10Y154_CLK = CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O;
  assign CLBLM_L_X8Y154_SLICE_X10Y154_D1 = 1'b1;
  assign CLBLM_L_X8Y154_SLICE_X10Y154_D2 = 1'b1;
  assign CLBLM_L_X8Y154_SLICE_X10Y154_D3 = 1'b1;
  assign CLBLM_L_X8Y154_SLICE_X10Y154_D4 = 1'b1;
  assign CLBLM_L_X8Y154_SLICE_X10Y154_D5 = 1'b1;
  assign CLBLM_L_X8Y154_SLICE_X10Y154_D6 = 1'b1;
  assign RIOI3_X105Y123_ILOGIC_X1Y124_D = RIOB33_X105Y123_IOB_X1Y124_I;
  assign CLBLM_R_X7Y148_SLICE_X9Y148_A1 = 1'b1;
  assign CLBLM_R_X7Y148_SLICE_X9Y148_A2 = CLBLM_R_X3Y148_SLICE_X3Y148_BQ;
  assign CLBLM_R_X7Y148_SLICE_X9Y148_A3 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X7Y148_SLICE_X9Y148_A4 = CLBLM_L_X8Y143_SLICE_X10Y143_CQ;
  assign CLBLM_R_X7Y148_SLICE_X9Y148_A5 = CLBLM_L_X10Y149_SLICE_X12Y149_BQ;
  assign CLBLM_R_X7Y148_SLICE_X9Y148_A6 = 1'b1;
  assign CLBLM_R_X7Y152_SLICE_X8Y152_B5 = CLBLM_L_X8Y146_SLICE_X10Y146_BQ;
  assign CLBLM_R_X7Y152_SLICE_X8Y152_B6 = 1'b1;
  assign CLBLM_R_X7Y148_SLICE_X9Y148_B1 = 1'b1;
  assign CLBLM_R_X7Y148_SLICE_X9Y148_B2 = CLBLM_R_X7Y148_SLICE_X9Y148_BQ;
  assign CLBLM_R_X7Y148_SLICE_X9Y148_B3 = CLBLM_R_X5Y143_SLICE_X7Y143_BQ;
  assign CLBLM_R_X7Y148_SLICE_X9Y148_B4 = CLBLM_L_X12Y149_SLICE_X17Y149_CO6;
  assign CLBLM_R_X7Y148_SLICE_X9Y148_B5 = CLBLM_L_X8Y148_SLICE_X10Y148_AQ;
  assign CLBLM_R_X7Y148_SLICE_X9Y148_B6 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X7Y148_SLICE_X9Y148_C1 = CLBLM_L_X8Y148_SLICE_X10Y148_BQ;
  assign CLBLM_R_X7Y148_SLICE_X9Y148_C2 = CLBLM_R_X3Y151_SLICE_X3Y151_BQ;
  assign CLBLM_R_X7Y148_SLICE_X9Y148_C3 = CLBLM_R_X5Y152_SLICE_X6Y152_CQ;
  assign CLBLM_R_X7Y148_SLICE_X9Y148_C4 = CLBLM_R_X7Y151_SLICE_X9Y151_CQ;
  assign CLBLM_R_X7Y148_SLICE_X9Y148_C5 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X7Y148_SLICE_X9Y148_C6 = 1'b1;
  assign CLBLM_R_X7Y148_SLICE_X9Y148_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X7Y148_SLICE_X9Y148_D1 = CLBLM_R_X11Y146_SLICE_X15Y146_BO6;
  assign CLBLM_R_X7Y148_SLICE_X9Y148_D2 = CLBLM_R_X7Y146_SLICE_X9Y146_CO6;
  assign CLBLM_R_X7Y148_SLICE_X9Y148_D3 = CLBLM_R_X5Y146_SLICE_X7Y146_D5Q;
  assign CLBLM_R_X7Y148_SLICE_X9Y148_D4 = CLBLM_R_X7Y149_SLICE_X8Y149_AQ;
  assign CLBLM_R_X7Y148_SLICE_X9Y148_D5 = CLBLM_R_X5Y144_SLICE_X7Y144_B5Q;
  assign CLBLL_L_X2Y147_SLICE_X0Y147_A1 = 1'b1;
  assign CLBLL_L_X2Y147_SLICE_X0Y147_A2 = 1'b1;
  assign CLBLL_L_X2Y147_SLICE_X0Y147_A3 = 1'b1;
  assign CLBLL_L_X2Y147_SLICE_X0Y147_A4 = 1'b1;
  assign CLBLL_L_X2Y147_SLICE_X0Y147_A5 = 1'b1;
  assign CLBLL_L_X2Y147_SLICE_X0Y147_A6 = 1'b1;
  assign CLBLM_R_X7Y148_SLICE_X9Y148_D6 = CLBLL_L_X4Y148_SLICE_X4Y148_CQ;
  assign CLBLM_R_X7Y148_SLICE_X8Y148_A1 = CLBLM_R_X7Y144_SLICE_X9Y144_B5Q;
  assign CLBLL_L_X2Y147_SLICE_X0Y147_B1 = 1'b1;
  assign CLBLL_L_X2Y147_SLICE_X0Y147_B2 = 1'b1;
  assign CLBLL_L_X2Y147_SLICE_X0Y147_B3 = 1'b1;
  assign CLBLL_L_X2Y147_SLICE_X0Y147_B4 = 1'b1;
  assign CLBLL_L_X2Y147_SLICE_X0Y147_B5 = 1'b1;
  assign CLBLL_L_X2Y147_SLICE_X0Y147_B6 = 1'b1;
  assign CLBLM_R_X7Y148_SLICE_X8Y148_A2 = CLBLL_L_X4Y148_SLICE_X4Y148_CQ;
  assign CLBLM_R_X7Y148_SLICE_X8Y148_A3 = CLBLM_L_X12Y147_SLICE_X16Y147_DO6;
  assign CLBLM_R_X7Y148_SLICE_X8Y148_A4 = CLBLM_R_X7Y153_SLICE_X8Y153_A5Q;
  assign CLBLL_L_X2Y147_SLICE_X0Y147_C1 = 1'b1;
  assign CLBLL_L_X2Y147_SLICE_X0Y147_C2 = 1'b1;
  assign CLBLL_L_X2Y147_SLICE_X0Y147_C3 = 1'b1;
  assign CLBLL_L_X2Y147_SLICE_X0Y147_C4 = 1'b1;
  assign CLBLL_L_X2Y147_SLICE_X0Y147_C5 = 1'b1;
  assign CLBLL_L_X2Y147_SLICE_X0Y147_C6 = 1'b1;
  assign CLBLM_R_X7Y148_SLICE_X8Y148_AX = CLBLM_R_X7Y147_SLICE_X9Y147_AQ;
  assign CLBLM_R_X7Y148_SLICE_X8Y148_B1 = CLBLM_R_X7Y144_SLICE_X9Y144_B5Q;
  assign CLBLM_R_X7Y148_SLICE_X8Y148_B2 = CLBLM_R_X11Y144_SLICE_X14Y144_CO6;
  assign CLBLM_R_X7Y148_SLICE_X8Y148_B3 = CLBLM_R_X5Y149_SLICE_X7Y149_BQ;
  assign CLBLM_R_X7Y148_SLICE_X8Y148_B4 = CLBLM_R_X7Y153_SLICE_X8Y153_A5Q;
  assign CLBLM_R_X7Y148_SLICE_X8Y148_B5 = CLBLM_L_X8Y146_SLICE_X11Y146_C5Q;
  assign CLBLM_R_X7Y148_SLICE_X8Y148_B6 = CLBLM_L_X10Y146_SLICE_X13Y146_DO6;
  assign CLBLL_L_X2Y147_SLICE_X0Y147_D1 = 1'b1;
  assign CLBLL_L_X2Y147_SLICE_X0Y147_D2 = 1'b1;
  assign CLBLL_L_X2Y147_SLICE_X0Y147_D3 = 1'b1;
  assign CLBLL_L_X2Y147_SLICE_X0Y147_D4 = 1'b1;
  assign CLBLL_L_X2Y147_SLICE_X0Y147_D5 = 1'b1;
  assign CLBLL_L_X2Y147_SLICE_X0Y147_D6 = 1'b1;
  assign CLBLM_R_X7Y148_SLICE_X8Y148_C3 = CLBLM_L_X8Y150_SLICE_X11Y150_BO6;
  assign CLBLM_R_X7Y148_SLICE_X8Y148_C4 = 1'b1;
  assign CLBLM_R_X7Y148_SLICE_X8Y148_C6 = CLBLM_R_X7Y148_SLICE_X8Y148_BO6;
  assign CLBLM_R_X7Y148_SLICE_X8Y148_CE = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X7Y148_SLICE_X8Y148_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X7Y148_SLICE_X8Y148_D1 = CLBLM_R_X3Y149_SLICE_X3Y149_AQ;
  assign CLBLM_R_X7Y148_SLICE_X8Y148_D2 = CLBLM_R_X5Y144_SLICE_X7Y144_B5Q;
  assign CLBLM_R_X7Y148_SLICE_X8Y148_D3 = CLBLL_L_X4Y152_SLICE_X5Y152_A5Q;
  assign CLBLM_R_X7Y148_SLICE_X8Y148_D4 = 1'b1;
  assign CLBLM_R_X7Y148_SLICE_X8Y148_D5 = 1'b1;
  assign CLBLM_R_X7Y148_SLICE_X8Y148_D6 = CLBLM_R_X7Y144_SLICE_X9Y144_BQ;
  assign CLBLL_L_X2Y147_SLICE_X1Y147_A1 = 1'b1;
  assign CLBLL_L_X2Y147_SLICE_X1Y147_A2 = CLBLM_R_X5Y147_SLICE_X7Y147_BQ;
  assign CLBLL_L_X2Y147_SLICE_X1Y147_A3 = 1'b1;
  assign CLBLL_L_X2Y147_SLICE_X1Y147_A4 = 1'b1;
  assign CLBLL_L_X2Y147_SLICE_X1Y147_A5 = 1'b1;
  assign CLBLL_L_X2Y147_SLICE_X1Y147_A6 = CLBLL_L_X4Y147_SLICE_X4Y147_C5Q;
  assign CLBLM_R_X5Y154_SLICE_X6Y154_A3 = CLBLL_L_X4Y153_SLICE_X5Y153_BO5;
  assign CLBLL_L_X2Y147_SLICE_X1Y147_B1 = 1'b1;
  assign CLBLL_L_X2Y147_SLICE_X1Y147_B2 = 1'b1;
  assign CLBLL_L_X2Y147_SLICE_X1Y147_B3 = 1'b1;
  assign CLBLL_L_X2Y147_SLICE_X1Y147_B4 = 1'b1;
  assign CLBLL_L_X2Y147_SLICE_X1Y147_B5 = 1'b1;
  assign CLBLL_L_X2Y147_SLICE_X1Y147_B6 = 1'b1;
  assign CLBLM_R_X5Y154_SLICE_X6Y154_A5 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLL_L_X2Y147_SLICE_X1Y147_C1 = 1'b1;
  assign CLBLL_L_X2Y147_SLICE_X1Y147_C2 = 1'b1;
  assign CLBLL_L_X2Y147_SLICE_X1Y147_C3 = 1'b1;
  assign CLBLL_L_X2Y147_SLICE_X1Y147_C4 = 1'b1;
  assign CLBLL_L_X2Y147_SLICE_X1Y147_C5 = 1'b1;
  assign CLBLL_L_X2Y147_SLICE_X1Y147_C6 = 1'b1;
  assign LIOI3_X0Y167_OLOGIC_X0Y168_D1 = RIOB33_X105Y101_IOB_X1Y101_I;
  assign LIOB33_X0Y179_IOB_X0Y180_O = RIOB33_X105Y127_IOB_X1Y127_I;
  assign CLBLL_L_X2Y147_SLICE_X1Y147_D1 = 1'b1;
  assign CLBLL_L_X2Y147_SLICE_X1Y147_D2 = 1'b1;
  assign CLBLL_L_X2Y147_SLICE_X1Y147_D3 = 1'b1;
  assign CLBLL_L_X2Y147_SLICE_X1Y147_D4 = 1'b1;
  assign CLBLL_L_X2Y147_SLICE_X1Y147_D5 = 1'b1;
  assign CLBLL_L_X2Y147_SLICE_X1Y147_D6 = 1'b1;
  assign LIOB33_X0Y179_IOB_X0Y179_O = RIOB33_X105Y125_IOB_X1Y126_I;
  assign LIOI3_X0Y105_OLOGIC_X0Y106_D1 = CLBLM_R_X3Y146_SLICE_X3Y146_BQ;
  assign LIOI3_X0Y167_OLOGIC_X0Y168_T1 = 1'b1;
  assign LIOI3_X0Y167_OLOGIC_X0Y167_D1 = RIOB33_X105Y105_IOB_X1Y106_I;
  assign LIOI3_X0Y105_OLOGIC_X0Y106_T1 = 1'b1;
  assign RIOI3_X105Y151_OLOGIC_X1Y152_D1 = 1'b1;
  assign LIOI3_X0Y167_OLOGIC_X0Y167_T1 = 1'b1;
  assign LIOI3_X0Y105_OLOGIC_X0Y105_D1 = CLBLL_L_X4Y150_SLICE_X4Y150_C5Q;
  assign RIOI3_X105Y151_OLOGIC_X1Y152_T1 = 1'b1;
  assign LIOI3_TBYTETERM_X0Y113_OLOGIC_X0Y114_D1 = CLBLM_L_X8Y142_SLICE_X10Y142_A5Q;
  assign LIOI3_X0Y105_OLOGIC_X0Y105_T1 = 1'b1;
  assign RIOI3_X105Y151_OLOGIC_X1Y151_D1 = 1'b1;
  assign LIOI3_TBYTETERM_X0Y113_OLOGIC_X0Y114_T1 = 1'b1;
  assign RIOI3_X105Y151_OLOGIC_X1Y151_T1 = 1'b1;
  assign LIOI3_TBYTETERM_X0Y113_OLOGIC_X0Y113_D1 = CLBLM_R_X3Y147_SLICE_X3Y147_C5Q;
  assign LIOB33_X0Y171_IOB_X0Y172_O = RIOB33_X105Y119_IOB_X1Y120_I;
  assign LIOB33_X0Y171_IOB_X0Y171_O = RIOB33_X105Y119_IOB_X1Y119_I;
  assign LIOI3_TBYTETERM_X0Y113_OLOGIC_X0Y113_T1 = 1'b1;
  assign CLBLM_R_X7Y149_SLICE_X9Y149_A1 = CLBLM_R_X7Y149_SLICE_X9Y149_B5Q;
  assign CLBLM_R_X7Y149_SLICE_X9Y149_A2 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X7Y149_SLICE_X9Y149_A3 = CLBLM_L_X8Y148_SLICE_X11Y148_AQ;
  assign CLBLM_R_X7Y149_SLICE_X9Y149_A4 = CLBLM_L_X8Y153_SLICE_X10Y153_AQ;
  assign CLBLM_R_X7Y149_SLICE_X9Y149_A5 = CLBLM_R_X7Y149_SLICE_X9Y149_C5Q;
  assign CLBLM_R_X7Y149_SLICE_X9Y149_A6 = 1'b1;
  assign CLBLM_R_X7Y150_SLICE_X9Y150_D5 = 1'b1;
  assign CLBLM_R_X7Y149_SLICE_X9Y149_B1 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X7Y149_SLICE_X9Y149_B2 = CLBLM_R_X7Y146_SLICE_X8Y146_B5Q;
  assign CLBLM_R_X7Y149_SLICE_X9Y149_B3 = CLBLL_L_X4Y150_SLICE_X5Y150_AQ;
  assign CLBLM_R_X7Y149_SLICE_X9Y149_B4 = CLBLL_L_X4Y149_SLICE_X5Y149_DQ;
  assign CLBLM_R_X7Y149_SLICE_X9Y149_B5 = CLBLM_L_X12Y151_SLICE_X16Y151_AQ;
  assign CLBLM_R_X7Y149_SLICE_X9Y149_B6 = 1'b1;
  assign CLBLM_R_X7Y149_SLICE_X9Y149_C1 = CLBLM_R_X7Y151_SLICE_X9Y151_C5Q;
  assign CLBLM_R_X7Y149_SLICE_X9Y149_C2 = CLBLM_L_X10Y151_SLICE_X13Y151_AQ;
  assign CLBLM_R_X7Y149_SLICE_X9Y149_C3 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X7Y149_SLICE_X9Y149_C4 = CLBLM_R_X7Y149_SLICE_X9Y149_AQ;
  assign CLBLM_R_X7Y149_SLICE_X9Y149_C5 = 1'b1;
  assign CLBLM_R_X7Y149_SLICE_X9Y149_C6 = 1'b1;
  assign CLBLM_R_X7Y149_SLICE_X9Y149_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X7Y150_SLICE_X9Y150_D6 = CLBLM_L_X8Y150_SLICE_X11Y150_BO6;
  assign CLBLL_L_X2Y148_SLICE_X0Y148_A1 = 1'b1;
  assign CLBLL_L_X2Y148_SLICE_X0Y148_A2 = 1'b1;
  assign CLBLL_L_X2Y148_SLICE_X0Y148_A3 = 1'b1;
  assign CLBLL_L_X2Y148_SLICE_X0Y148_A4 = 1'b1;
  assign CLBLL_L_X2Y148_SLICE_X0Y148_A5 = 1'b1;
  assign CLBLL_L_X2Y148_SLICE_X0Y148_A6 = 1'b1;
  assign CLBLM_R_X7Y149_SLICE_X9Y149_D1 = CLBLM_R_X7Y148_SLICE_X9Y148_AQ;
  assign CLBLM_R_X7Y149_SLICE_X9Y149_D2 = CLBLM_R_X7Y153_SLICE_X8Y153_AQ;
  assign CLBLL_L_X2Y148_SLICE_X0Y148_AX = CLBLM_R_X3Y145_SLICE_X3Y145_CQ;
  assign CLBLM_R_X7Y149_SLICE_X9Y149_D3 = CLBLM_R_X11Y144_SLICE_X14Y144_AO6;
  assign CLBLL_L_X2Y148_SLICE_X0Y148_B1 = 1'b1;
  assign CLBLL_L_X2Y148_SLICE_X0Y148_B2 = 1'b1;
  assign CLBLL_L_X2Y148_SLICE_X0Y148_B3 = 1'b1;
  assign CLBLL_L_X2Y148_SLICE_X0Y148_B4 = 1'b1;
  assign CLBLL_L_X2Y148_SLICE_X0Y148_B5 = 1'b1;
  assign CLBLL_L_X2Y148_SLICE_X0Y148_B6 = 1'b1;
  assign CLBLM_R_X7Y149_SLICE_X8Y149_A1 = CLBLM_R_X5Y152_SLICE_X7Y152_B5Q;
  assign CLBLM_R_X7Y149_SLICE_X8Y149_A2 = CLBLM_L_X8Y149_SLICE_X10Y149_AQ;
  assign CLBLM_R_X7Y149_SLICE_X8Y149_A3 = 1'b1;
  assign CLBLL_L_X2Y148_SLICE_X0Y148_C1 = 1'b1;
  assign CLBLL_L_X2Y148_SLICE_X0Y148_C2 = 1'b1;
  assign CLBLL_L_X2Y148_SLICE_X0Y148_C3 = 1'b1;
  assign CLBLL_L_X2Y148_SLICE_X0Y148_C4 = 1'b1;
  assign CLBLL_L_X2Y148_SLICE_X0Y148_C5 = 1'b1;
  assign CLBLL_L_X2Y148_SLICE_X0Y148_C6 = 1'b1;
  assign CLBLL_L_X2Y148_SLICE_X0Y148_CE = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X7Y149_SLICE_X8Y149_A6 = 1'b1;
  assign CLBLL_L_X2Y148_SLICE_X0Y148_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X7Y149_SLICE_X8Y149_B1 = CLBLM_R_X11Y144_SLICE_X14Y144_AO6;
  assign CLBLM_R_X7Y149_SLICE_X8Y149_B2 = CLBLM_R_X5Y142_SLICE_X6Y142_CQ;
  assign CLBLM_R_X7Y149_SLICE_X8Y149_B3 = CLBLM_R_X7Y144_SLICE_X9Y144_B5Q;
  assign CLBLM_R_X7Y149_SLICE_X8Y149_B4 = CLBLM_R_X11Y144_SLICE_X14Y144_CO6;
  assign CLBLL_L_X2Y148_SLICE_X0Y148_D1 = 1'b1;
  assign CLBLL_L_X2Y148_SLICE_X0Y148_D2 = 1'b1;
  assign CLBLL_L_X2Y148_SLICE_X0Y148_D3 = 1'b1;
  assign CLBLL_L_X2Y148_SLICE_X0Y148_D4 = 1'b1;
  assign CLBLL_L_X2Y148_SLICE_X0Y148_D5 = 1'b1;
  assign CLBLL_L_X2Y148_SLICE_X0Y148_D6 = 1'b1;
  assign CLBLM_R_X7Y149_SLICE_X8Y149_C1 = CLBLM_L_X10Y146_SLICE_X13Y146_DO6;
  assign CLBLM_R_X7Y149_SLICE_X8Y149_C2 = CLBLM_R_X3Y149_SLICE_X3Y149_D5Q;
  assign CLBLM_R_X7Y149_SLICE_X8Y149_C3 = CLBLM_R_X7Y147_SLICE_X8Y147_BO6;
  assign CLBLM_R_X7Y149_SLICE_X8Y149_C4 = CLBLM_L_X10Y150_SLICE_X12Y150_BO6;
  assign CLBLM_R_X7Y149_SLICE_X8Y149_C5 = CLBLM_R_X7Y148_SLICE_X8Y148_AO6;
  assign CLBLM_R_X7Y149_SLICE_X8Y149_C6 = CLBLM_R_X5Y149_SLICE_X7Y149_D5Q;
  assign CLBLM_R_X7Y149_SLICE_X8Y149_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X7Y149_SLICE_X8Y149_D1 = CLBLM_R_X7Y148_SLICE_X8Y148_AO5;
  assign CLBLM_R_X7Y149_SLICE_X8Y149_D2 = CLBLL_L_X4Y151_SLICE_X5Y151_AQ;
  assign CLBLM_R_X7Y149_SLICE_X8Y149_D3 = CLBLM_R_X13Y149_SLICE_X18Y149_AO6;
  assign CLBLM_R_X7Y149_SLICE_X8Y149_D4 = CLBLM_R_X7Y149_SLICE_X8Y149_A5Q;
  assign CLBLM_R_X7Y149_SLICE_X8Y149_D5 = 1'b1;
  assign CLBLM_R_X7Y149_SLICE_X8Y149_D6 = CLBLM_R_X7Y149_SLICE_X8Y149_BO6;
  assign CLBLL_L_X2Y148_SLICE_X1Y148_A1 = LIOB33_X0Y55_IOB_X0Y55_I;
  assign CLBLL_L_X2Y148_SLICE_X1Y148_A2 = CLBLM_R_X3Y148_SLICE_X2Y148_BQ;
  assign CLBLL_L_X2Y148_SLICE_X1Y148_A3 = CLBLL_L_X4Y149_SLICE_X4Y149_D5Q;
  assign CLBLL_L_X2Y148_SLICE_X1Y148_A4 = CLBLL_L_X2Y146_SLICE_X1Y146_BQ;
  assign CLBLL_L_X2Y148_SLICE_X1Y148_A5 = CLBLM_R_X3Y149_SLICE_X2Y149_DQ;
  assign CLBLL_L_X2Y148_SLICE_X1Y148_A6 = CLBLL_L_X4Y149_SLICE_X4Y149_DQ;
  assign CLBLL_L_X2Y148_SLICE_X1Y148_B1 = LIOB33_X0Y55_IOB_X0Y55_I;
  assign CLBLL_L_X2Y148_SLICE_X1Y148_B2 = CLBLM_R_X3Y148_SLICE_X2Y148_BQ;
  assign CLBLL_L_X2Y148_SLICE_X1Y148_B3 = CLBLL_L_X4Y149_SLICE_X4Y149_D5Q;
  assign CLBLL_L_X2Y148_SLICE_X1Y148_B4 = CLBLL_L_X2Y146_SLICE_X1Y146_BQ;
  assign CLBLL_L_X2Y148_SLICE_X1Y148_B5 = CLBLM_R_X3Y149_SLICE_X2Y149_DQ;
  assign CLBLL_L_X2Y148_SLICE_X1Y148_B6 = CLBLL_L_X4Y149_SLICE_X4Y149_DQ;
  assign CLBLL_L_X2Y148_SLICE_X1Y148_C1 = CLBLL_L_X2Y146_SLICE_X1Y146_B5Q;
  assign CLBLL_L_X2Y148_SLICE_X1Y148_C2 = CLBLL_L_X4Y148_SLICE_X5Y148_BQ;
  assign CLBLL_L_X2Y148_SLICE_X1Y148_C3 = 1'b1;
  assign CLBLL_L_X2Y148_SLICE_X1Y148_C4 = CLBLM_R_X3Y145_SLICE_X3Y145_CQ;
  assign CLBLL_L_X2Y148_SLICE_X1Y148_C5 = CLBLM_R_X3Y144_SLICE_X3Y144_AQ;
  assign CLBLL_L_X2Y148_SLICE_X1Y148_C6 = CLBLM_R_X5Y145_SLICE_X7Y145_CO6;
  assign CLBLL_L_X2Y148_SLICE_X1Y148_D1 = 1'b1;
  assign CLBLL_L_X2Y148_SLICE_X1Y148_D2 = 1'b1;
  assign CLBLL_L_X2Y148_SLICE_X1Y148_D3 = 1'b1;
  assign CLBLL_L_X2Y148_SLICE_X1Y148_D4 = 1'b1;
  assign CLBLL_L_X2Y148_SLICE_X1Y148_D5 = 1'b1;
  assign CLBLL_L_X2Y148_SLICE_X1Y148_D6 = 1'b1;
  assign LIOB33_X0Y173_IOB_X0Y174_O = RIOB33_X105Y121_IOB_X1Y122_I;
  assign LIOB33_X0Y173_IOB_X0Y173_O = RIOB33_X105Y121_IOB_X1Y121_I;
  assign CLBLM_R_X7Y150_SLICE_X9Y150_A1 = CLBLM_R_X7Y153_SLICE_X8Y153_A5Q;
  assign CLBLM_R_X7Y150_SLICE_X9Y150_A2 = CLBLM_R_X3Y150_SLICE_X2Y150_D5Q;
  assign CLBLM_R_X7Y150_SLICE_X9Y150_A3 = CLBLM_R_X11Y144_SLICE_X14Y144_AO6;
  assign CLBLM_R_X7Y150_SLICE_X9Y150_A4 = CLBLM_R_X11Y144_SLICE_X14Y144_CO6;
  assign CLBLM_R_X7Y150_SLICE_X9Y150_A5 = CLBLM_R_X5Y151_SLICE_X6Y151_BQ;
  assign CLBLM_R_X7Y150_SLICE_X9Y150_A6 = CLBLM_R_X7Y144_SLICE_X9Y144_B5Q;
  assign CLBLM_R_X7Y152_SLICE_X8Y152_C4 = CLBLM_L_X12Y149_SLICE_X17Y149_CO6;
  assign CLBLM_R_X7Y150_SLICE_X9Y150_B1 = CLBLM_R_X3Y149_SLICE_X2Y149_C5Q;
  assign CLBLM_R_X7Y150_SLICE_X9Y150_B2 = CLBLM_L_X8Y150_SLICE_X10Y150_BO6;
  assign CLBLM_R_X7Y150_SLICE_X9Y150_B3 = CLBLM_R_X7Y148_SLICE_X8Y148_AO6;
  assign CLBLM_R_X7Y150_SLICE_X9Y150_B4 = CLBLM_R_X7Y149_SLICE_X9Y149_C5Q;
  assign CLBLM_R_X7Y150_SLICE_X9Y150_B5 = CLBLM_R_X7Y150_SLICE_X9Y150_AO6;
  assign CLBLM_R_X7Y150_SLICE_X9Y150_B6 = CLBLM_L_X10Y146_SLICE_X13Y146_DO6;
  assign CLBLM_R_X5Y140_SLICE_X7Y140_A1 = 1'b1;
  assign CLBLM_R_X5Y140_SLICE_X7Y140_A2 = 1'b1;
  assign CLBLM_R_X5Y140_SLICE_X7Y140_A3 = 1'b1;
  assign CLBLM_R_X5Y140_SLICE_X7Y140_A4 = 1'b1;
  assign CLBLM_R_X5Y140_SLICE_X7Y140_A5 = 1'b1;
  assign CLBLM_R_X5Y140_SLICE_X7Y140_A6 = 1'b1;
  assign CLBLM_R_X7Y150_SLICE_X9Y150_C1 = CLBLM_R_X11Y146_SLICE_X15Y146_BO6;
  assign CLBLM_R_X7Y150_SLICE_X9Y150_C2 = CLBLL_L_X4Y148_SLICE_X4Y148_CQ;
  assign CLBLM_R_X7Y150_SLICE_X9Y150_C3 = CLBLM_R_X5Y142_SLICE_X6Y142_DQ;
  assign CLBLM_R_X5Y140_SLICE_X7Y140_B1 = 1'b1;
  assign CLBLM_R_X5Y140_SLICE_X7Y140_B2 = 1'b1;
  assign CLBLM_R_X5Y140_SLICE_X7Y140_B3 = 1'b1;
  assign CLBLM_R_X5Y140_SLICE_X7Y140_B4 = 1'b1;
  assign CLBLM_R_X5Y140_SLICE_X7Y140_B5 = 1'b1;
  assign CLBLM_R_X5Y140_SLICE_X7Y140_B6 = 1'b1;
  assign CLBLM_R_X7Y150_SLICE_X9Y150_D1 = CLBLM_R_X7Y151_SLICE_X8Y151_AQ;
  assign CLBLM_R_X7Y150_SLICE_X9Y150_D2 = CLBLL_L_X4Y153_SLICE_X4Y153_B5Q;
  assign CLBLM_R_X5Y140_SLICE_X7Y140_C1 = 1'b1;
  assign CLBLM_R_X5Y140_SLICE_X7Y140_C2 = 1'b1;
  assign CLBLM_R_X5Y140_SLICE_X7Y140_C3 = 1'b1;
  assign CLBLM_R_X5Y140_SLICE_X7Y140_C4 = 1'b1;
  assign CLBLM_R_X5Y140_SLICE_X7Y140_C5 = 1'b1;
  assign CLBLM_R_X5Y140_SLICE_X7Y140_C6 = 1'b1;
  assign CLBLM_R_X7Y150_SLICE_X9Y150_D3 = 1'b1;
  assign CLBLM_R_X7Y150_SLICE_X9Y150_D4 = CLBLM_L_X8Y150_SLICE_X10Y150_BO5;
  assign CLBLM_R_X7Y150_SLICE_X8Y150_A1 = CLBLM_R_X7Y150_SLICE_X8Y150_BO5;
  assign CLBLM_R_X7Y150_SLICE_X8Y150_A2 = CLBLM_L_X10Y151_SLICE_X12Y151_AQ;
  assign CLBLM_R_X7Y150_SLICE_X8Y150_A3 = CLBLM_R_X7Y150_SLICE_X8Y150_AQ;
  assign CLBLM_R_X7Y150_SLICE_X8Y150_A4 = CLBLM_R_X7Y146_SLICE_X8Y146_D5Q;
  assign CLBLM_R_X7Y150_SLICE_X8Y150_A5 = CLBLM_L_X8Y149_SLICE_X11Y149_AQ;
  assign CLBLM_R_X7Y150_SLICE_X8Y150_A6 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X5Y140_SLICE_X7Y140_D1 = 1'b1;
  assign CLBLM_R_X5Y140_SLICE_X7Y140_D2 = 1'b1;
  assign CLBLM_R_X5Y140_SLICE_X7Y140_D3 = 1'b1;
  assign CLBLM_R_X5Y140_SLICE_X7Y140_D4 = 1'b1;
  assign CLBLM_R_X5Y140_SLICE_X7Y140_D5 = 1'b1;
  assign CLBLM_R_X5Y140_SLICE_X7Y140_D6 = 1'b1;
  assign CLBLM_R_X7Y150_SLICE_X8Y150_B1 = 1'b1;
  assign CLBLM_R_X7Y150_SLICE_X8Y150_B2 = CLBLM_R_X5Y143_SLICE_X7Y143_AQ;
  assign CLBLM_R_X7Y150_SLICE_X8Y150_B3 = CLBLM_R_X7Y150_SLICE_X8Y150_AQ;
  assign CLBLM_R_X7Y150_SLICE_X8Y150_B4 = 1'b1;
  assign CLBLM_R_X7Y150_SLICE_X8Y150_B5 = CLBLM_R_X7Y143_SLICE_X8Y143_DO6;
  assign CLBLM_R_X5Y140_SLICE_X6Y140_A1 = CLBLM_R_X5Y140_SLICE_X6Y140_CQ;
  assign CLBLM_R_X5Y140_SLICE_X6Y140_A2 = CLBLL_L_X4Y140_SLICE_X4Y140_CO6;
  assign CLBLM_R_X5Y140_SLICE_X6Y140_A3 = CLBLM_R_X5Y140_SLICE_X6Y140_AQ;
  assign CLBLM_R_X5Y140_SLICE_X6Y140_A4 = CLBLL_L_X4Y140_SLICE_X4Y140_AQ;
  assign CLBLM_R_X5Y140_SLICE_X6Y140_A5 = CLBLM_R_X5Y144_SLICE_X6Y144_DQ;
  assign CLBLM_R_X5Y140_SLICE_X6Y140_A6 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X7Y150_SLICE_X8Y150_C1 = CLBLM_R_X7Y153_SLICE_X8Y153_CQ;
  assign CLBLM_R_X7Y150_SLICE_X8Y150_C2 = CLBLM_R_X11Y148_SLICE_X15Y148_AO6;
  assign CLBLM_R_X5Y140_SLICE_X6Y140_AX = CLBLM_R_X5Y140_SLICE_X6Y140_DO6;
  assign CLBLM_R_X7Y150_SLICE_X8Y150_C3 = CLBLM_R_X7Y149_SLICE_X9Y149_A5Q;
  assign CLBLM_R_X5Y140_SLICE_X6Y140_B1 = CLBLL_L_X4Y140_SLICE_X4Y140_CO6;
  assign CLBLM_R_X5Y140_SLICE_X6Y140_B2 = CLBLM_R_X5Y140_SLICE_X6Y140_BQ;
  assign CLBLM_R_X5Y140_SLICE_X6Y140_B3 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X5Y140_SLICE_X6Y140_B4 = CLBLM_R_X5Y140_SLICE_X6Y140_DO5;
  assign CLBLM_R_X5Y140_SLICE_X6Y140_B5 = 1'b1;
  assign CLBLM_R_X5Y140_SLICE_X6Y140_B6 = CLBLM_R_X5Y142_SLICE_X6Y142_CQ;
  assign CLBLM_L_X12Y153_SLICE_X17Y153_C3 = 1'b1;
  assign CLBLM_R_X7Y150_SLICE_X8Y150_CLK = CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O;
  assign CLBLM_R_X7Y150_SLICE_X8Y150_D1 = CLBLM_R_X11Y147_SLICE_X15Y147_BO6;
  assign CLBLM_R_X5Y140_SLICE_X6Y140_C1 = CLBLL_L_X4Y140_SLICE_X4Y140_AQ;
  assign CLBLM_R_X5Y140_SLICE_X6Y140_C2 = CLBLM_R_X5Y140_SLICE_X6Y140_CQ;
  assign CLBLM_R_X5Y140_SLICE_X6Y140_C3 = CLBLM_R_X7Y147_SLICE_X9Y147_DQ;
  assign CLBLM_R_X5Y140_SLICE_X6Y140_C4 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X5Y140_SLICE_X6Y140_C5 = CLBLL_L_X4Y140_SLICE_X4Y140_CO6;
  assign CLBLM_R_X5Y140_SLICE_X6Y140_C6 = 1'b1;
  assign CLBLM_R_X7Y150_SLICE_X8Y150_D2 = CLBLM_R_X7Y153_SLICE_X8Y153_A5Q;
  assign CLBLM_R_X7Y150_SLICE_X8Y150_D3 = CLBLM_R_X11Y144_SLICE_X14Y144_BO6;
  assign CLBLM_R_X7Y150_SLICE_X8Y150_D4 = CLBLM_R_X7Y144_SLICE_X9Y144_B5Q;
  assign CLBLM_R_X5Y140_SLICE_X6Y140_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X7Y150_SLICE_X8Y150_D6 = CLBLM_R_X3Y151_SLICE_X2Y151_AQ;
  assign CLBLM_R_X5Y140_SLICE_X6Y140_D1 = CLBLL_L_X4Y140_SLICE_X4Y140_AQ;
  assign CLBLM_R_X5Y140_SLICE_X6Y140_D2 = CLBLM_R_X5Y141_SLICE_X6Y141_BQ;
  assign CLBLM_R_X5Y140_SLICE_X6Y140_D3 = CLBLM_R_X5Y140_SLICE_X6Y140_AQ;
  assign CLBLM_R_X5Y140_SLICE_X6Y140_D4 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X5Y140_SLICE_X6Y140_D5 = CLBLM_R_X5Y140_SLICE_X6Y140_CQ;
  assign CLBLM_R_X5Y140_SLICE_X6Y140_D6 = 1'b1;
  assign LIOB33_X0Y175_IOB_X0Y176_O = RIOB33_X105Y115_IOB_X1Y116_I;
  assign LIOB33_X0Y175_IOB_X0Y175_O = RIOB33_X105Y123_IOB_X1Y123_I;
  assign CLBLM_L_X12Y153_SLICE_X17Y153_D6 = 1'b1;
  assign CLBLM_R_X11Y146_SLICE_X14Y146_C2 = CLBLM_R_X7Y144_SLICE_X9Y144_B5Q;
  assign CLBLM_L_X12Y153_SLICE_X16Y153_A6 = 1'b1;
  assign LIOI3_X0Y171_OLOGIC_X0Y172_D1 = RIOB33_X105Y119_IOB_X1Y120_I;
  assign RIOI3_SING_X105Y100_ILOGIC_X1Y100_D = RIOB33_SING_X105Y100_IOB_X1Y100_I;
  assign CLBLM_L_X10Y155_SLICE_X13Y155_C3 = CLBLM_R_X5Y147_SLICE_X6Y147_AQ;
  assign LIOI3_X0Y171_OLOGIC_X0Y172_T1 = 1'b1;
  assign LIOI3_X0Y109_OLOGIC_X0Y110_D1 = CLBLM_R_X5Y145_SLICE_X7Y145_AQ;
  assign LIOI3_X0Y171_OLOGIC_X0Y171_D1 = RIOB33_X105Y119_IOB_X1Y119_I;
  assign LIOI3_X0Y109_OLOGIC_X0Y110_T1 = 1'b1;
  assign RIOI3_X105Y153_OLOGIC_X1Y154_D1 = 1'b1;
  assign LIOI3_X0Y171_OLOGIC_X0Y171_T1 = 1'b1;
  assign LIOI3_X0Y109_OLOGIC_X0Y109_D1 = CLBLM_R_X5Y141_SLICE_X6Y141_BQ;
  assign RIOI3_X105Y153_OLOGIC_X1Y154_T1 = 1'b1;
  assign LIOI3_TBYTETERM_X0Y137_OLOGIC_X0Y138_D1 = CLBLM_R_X3Y148_SLICE_X2Y148_A5Q;
  assign LIOI3_X0Y109_OLOGIC_X0Y109_T1 = 1'b1;
  assign CLBLM_R_X11Y146_SLICE_X14Y146_C5 = CLBLM_R_X7Y146_SLICE_X9Y146_CO6;
  assign RIOI3_X105Y153_OLOGIC_X1Y153_D1 = 1'b1;
  assign LIOI3_TBYTETERM_X0Y137_OLOGIC_X0Y138_T1 = 1'b1;
  assign CLBLM_R_X7Y151_SLICE_X9Y151_A1 = CLBLM_R_X7Y142_SLICE_X8Y142_C5Q;
  assign CLBLM_R_X7Y151_SLICE_X9Y151_A2 = CLBLM_R_X7Y152_SLICE_X8Y152_D5Q;
  assign CLBLM_R_X7Y151_SLICE_X9Y151_A3 = CLBLM_R_X7Y151_SLICE_X9Y151_AQ;
  assign CLBLM_R_X7Y151_SLICE_X9Y151_A4 = CLBLL_L_X4Y151_SLICE_X4Y151_C5Q;
  assign CLBLM_R_X7Y151_SLICE_X9Y151_A5 = CLBLM_L_X8Y153_SLICE_X10Y153_AQ;
  assign CLBLM_R_X7Y151_SLICE_X9Y151_A6 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign RIOI3_X105Y153_OLOGIC_X1Y153_T1 = 1'b1;
  assign LIOI3_TBYTETERM_X0Y137_OLOGIC_X0Y137_D1 = CLBLM_R_X5Y153_SLICE_X6Y153_B5Q;
  assign CLBLM_R_X7Y151_SLICE_X9Y151_AX = CLBLM_R_X7Y152_SLICE_X9Y152_DO5;
  assign CLBLM_L_X12Y153_SLICE_X16Y153_C1 = 1'b1;
  assign CLBLM_R_X7Y151_SLICE_X9Y151_B1 = CLBLM_L_X8Y149_SLICE_X11Y149_AQ;
  assign CLBLM_R_X7Y151_SLICE_X9Y151_B2 = CLBLM_R_X7Y152_SLICE_X9Y152_C5Q;
  assign CLBLM_R_X7Y151_SLICE_X9Y151_B3 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X7Y151_SLICE_X9Y151_B4 = CLBLM_R_X7Y150_SLICE_X8Y150_BO6;
  assign CLBLM_R_X7Y151_SLICE_X9Y151_B5 = CLBLM_R_X7Y151_SLICE_X9Y151_BQ;
  assign CLBLM_R_X7Y151_SLICE_X9Y151_B6 = CLBLM_L_X10Y153_SLICE_X13Y153_CQ;
  assign CLBLM_L_X10Y155_SLICE_X13Y155_D3 = 1'b1;
  assign CLBLM_R_X5Y141_SLICE_X7Y141_A1 = 1'b1;
  assign CLBLM_R_X5Y141_SLICE_X7Y141_A2 = 1'b1;
  assign CLBLM_R_X5Y141_SLICE_X7Y141_A3 = 1'b1;
  assign CLBLM_R_X5Y141_SLICE_X7Y141_A4 = 1'b1;
  assign CLBLM_R_X5Y141_SLICE_X7Y141_A5 = 1'b1;
  assign CLBLL_L_X2Y150_SLICE_X0Y150_A1 = 1'b1;
  assign CLBLL_L_X2Y150_SLICE_X0Y150_A2 = 1'b1;
  assign CLBLL_L_X2Y150_SLICE_X0Y150_A3 = 1'b1;
  assign CLBLL_L_X2Y150_SLICE_X0Y150_A4 = 1'b1;
  assign CLBLL_L_X2Y150_SLICE_X0Y150_A5 = 1'b1;
  assign CLBLL_L_X2Y150_SLICE_X0Y150_A6 = 1'b1;
  assign CLBLM_L_X12Y153_SLICE_X16Y153_C5 = 1'b1;
  assign CLBLM_R_X5Y141_SLICE_X7Y141_A6 = 1'b1;
  assign CLBLM_R_X5Y141_SLICE_X7Y141_B4 = 1'b1;
  assign CLBLL_L_X2Y150_SLICE_X0Y150_B1 = 1'b1;
  assign CLBLL_L_X2Y150_SLICE_X0Y150_B2 = 1'b1;
  assign CLBLL_L_X2Y150_SLICE_X0Y150_B3 = 1'b1;
  assign CLBLL_L_X2Y150_SLICE_X0Y150_B4 = 1'b1;
  assign CLBLL_L_X2Y150_SLICE_X0Y150_B5 = 1'b1;
  assign CLBLL_L_X2Y150_SLICE_X0Y150_B6 = 1'b1;
  assign CLBLM_R_X5Y141_SLICE_X7Y141_B6 = 1'b1;
  assign CLBLM_R_X5Y141_SLICE_X7Y141_B5 = 1'b1;
  assign CLBLM_R_X5Y141_SLICE_X7Y141_C4 = 1'b1;
  assign CLBLL_L_X2Y150_SLICE_X0Y150_C1 = 1'b1;
  assign CLBLL_L_X2Y150_SLICE_X0Y150_C2 = 1'b1;
  assign CLBLL_L_X2Y150_SLICE_X0Y150_C3 = 1'b1;
  assign CLBLL_L_X2Y150_SLICE_X0Y150_C4 = 1'b1;
  assign CLBLL_L_X2Y150_SLICE_X0Y150_C5 = 1'b1;
  assign CLBLL_L_X2Y150_SLICE_X0Y150_C6 = 1'b1;
  assign CLBLM_R_X5Y141_SLICE_X7Y141_C5 = 1'b1;
  assign CLBLM_R_X5Y141_SLICE_X7Y141_C6 = 1'b1;
  assign CLBLM_R_X7Y151_SLICE_X8Y151_A1 = CLBLM_R_X5Y147_SLICE_X7Y147_AQ;
  assign CLBLM_R_X5Y141_SLICE_X7Y141_D1 = 1'b1;
  assign CLBLM_R_X5Y141_SLICE_X7Y141_D2 = 1'b1;
  assign CLBLM_R_X5Y141_SLICE_X7Y141_D3 = 1'b1;
  assign CLBLM_R_X5Y141_SLICE_X7Y141_D4 = 1'b1;
  assign CLBLL_L_X2Y150_SLICE_X0Y150_D1 = 1'b1;
  assign CLBLL_L_X2Y150_SLICE_X0Y150_D2 = 1'b1;
  assign CLBLL_L_X2Y150_SLICE_X0Y150_D3 = 1'b1;
  assign CLBLL_L_X2Y150_SLICE_X0Y150_D4 = 1'b1;
  assign CLBLL_L_X2Y150_SLICE_X0Y150_D5 = 1'b1;
  assign CLBLL_L_X2Y150_SLICE_X0Y150_D6 = 1'b1;
  assign CLBLM_R_X5Y141_SLICE_X7Y141_D5 = 1'b1;
  assign CLBLM_R_X5Y141_SLICE_X7Y141_D6 = 1'b1;
  assign CLBLM_R_X5Y141_SLICE_X6Y141_A1 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X5Y141_SLICE_X6Y141_A2 = CLBLM_R_X5Y141_SLICE_X6Y141_DQ;
  assign CLBLM_R_X5Y141_SLICE_X6Y141_A3 = CLBLM_R_X5Y141_SLICE_X6Y141_AQ;
  assign CLBLM_R_X5Y141_SLICE_X6Y141_A4 = 1'b1;
  assign CLBLM_R_X5Y141_SLICE_X6Y141_A5 = CLBLM_R_X5Y142_SLICE_X6Y142_AQ;
  assign CLBLM_R_X5Y141_SLICE_X6Y141_A6 = CLBLM_R_X11Y146_SLICE_X14Y146_DO6;
  assign CLBLM_R_X7Y151_SLICE_X8Y151_C1 = CLBLM_R_X3Y147_SLICE_X3Y147_AQ;
  assign CLBLM_R_X7Y151_SLICE_X8Y151_C2 = CLBLL_L_X4Y151_SLICE_X5Y151_BQ;
  assign CLBLM_R_X5Y141_SLICE_X6Y141_B1 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X5Y141_SLICE_X6Y141_B2 = CLBLM_R_X5Y145_SLICE_X7Y145_AQ;
  assign CLBLM_R_X5Y141_SLICE_X6Y141_B3 = CLBLM_R_X5Y140_SLICE_X6Y140_CQ;
  assign CLBLM_R_X5Y141_SLICE_X6Y141_B4 = CLBLM_L_X8Y144_SLICE_X10Y144_BQ;
  assign CLBLM_R_X5Y141_SLICE_X6Y141_B5 = 1'b1;
  assign CLBLM_R_X5Y141_SLICE_X6Y141_B6 = 1'b1;
  assign CLBLM_R_X7Y151_SLICE_X8Y151_CLK = CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O;
  assign CLBLM_R_X7Y151_SLICE_X8Y151_D1 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X7Y151_SLICE_X8Y151_D2 = CLBLM_R_X5Y149_SLICE_X7Y149_BQ;
  assign CLBLM_R_X5Y141_SLICE_X6Y141_C1 = 1'b1;
  assign CLBLM_R_X5Y141_SLICE_X6Y141_C2 = CLBLM_R_X5Y141_SLICE_X6Y141_D5Q;
  assign CLBLM_R_X5Y141_SLICE_X6Y141_C3 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X5Y141_SLICE_X6Y141_C4 = CLBLM_L_X8Y151_SLICE_X10Y151_B5Q;
  assign CLBLM_R_X5Y141_SLICE_X6Y141_C5 = CLBLM_L_X10Y145_SLICE_X12Y145_AQ;
  assign CLBLL_L_X2Y150_SLICE_X1Y150_A1 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLL_L_X2Y150_SLICE_X1Y150_A2 = CLBLL_L_X4Y146_SLICE_X5Y146_BQ;
  assign CLBLL_L_X2Y150_SLICE_X1Y150_A3 = 1'b1;
  assign CLBLL_L_X2Y150_SLICE_X1Y150_A4 = CLBLL_L_X4Y150_SLICE_X4Y150_DO6;
  assign CLBLL_L_X2Y150_SLICE_X1Y150_A5 = 1'b1;
  assign CLBLL_L_X2Y150_SLICE_X1Y150_A6 = CLBLM_R_X5Y153_SLICE_X6Y153_DQ;
  assign CLBLM_R_X5Y141_SLICE_X6Y141_C6 = 1'b1;
  assign CLBLM_R_X5Y141_SLICE_X6Y141_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLL_L_X2Y150_SLICE_X1Y150_B1 = 1'b1;
  assign CLBLL_L_X2Y150_SLICE_X1Y150_B2 = 1'b1;
  assign CLBLL_L_X2Y150_SLICE_X1Y150_B3 = 1'b1;
  assign CLBLL_L_X2Y150_SLICE_X1Y150_B4 = 1'b1;
  assign CLBLM_R_X5Y141_SLICE_X6Y141_D4 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X5Y141_SLICE_X6Y141_D5 = RIOB33_X105Y123_IOB_X1Y123_I;
  assign CLBLM_R_X5Y141_SLICE_X6Y141_D6 = 1'b1;
  assign CLBLL_L_X2Y150_SLICE_X1Y150_B5 = 1'b1;
  assign CLBLL_L_X2Y150_SLICE_X1Y150_B6 = 1'b1;
  assign CLBLM_R_X5Y141_SLICE_X6Y141_D1 = RIOB33_X105Y107_IOB_X1Y108_I;
  assign CLBLM_R_X5Y141_SLICE_X6Y141_D2 = CLBLM_R_X5Y141_SLICE_X6Y141_AQ;
  assign CLBLM_R_X5Y141_SLICE_X6Y141_D3 = CLBLM_L_X8Y146_SLICE_X11Y146_DQ;
  assign CLBLL_L_X2Y150_SLICE_X1Y150_C1 = 1'b1;
  assign CLBLL_L_X2Y150_SLICE_X1Y150_C2 = 1'b1;
  assign CLBLL_L_X2Y150_SLICE_X1Y150_C3 = 1'b1;
  assign CLBLL_L_X2Y150_SLICE_X1Y150_C4 = 1'b1;
  assign CLBLL_L_X2Y150_SLICE_X1Y150_C5 = 1'b1;
  assign CLBLL_L_X2Y150_SLICE_X1Y150_C6 = 1'b1;
  assign CLBLL_L_X2Y150_SLICE_X1Y150_CLK = CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O;
  assign LIOB33_X0Y177_IOB_X0Y177_O = RIOB33_X105Y123_IOB_X1Y124_I;
  assign LIOB33_X0Y177_IOB_X0Y178_O = RIOB33_X105Y125_IOB_X1Y125_I;
  assign CLBLL_L_X2Y150_SLICE_X1Y150_D1 = 1'b1;
  assign CLBLL_L_X2Y150_SLICE_X1Y150_D2 = 1'b1;
  assign CLBLL_L_X2Y150_SLICE_X1Y150_D3 = 1'b1;
  assign CLBLL_L_X2Y150_SLICE_X1Y150_D4 = 1'b1;
  assign CLBLL_L_X2Y150_SLICE_X1Y150_D5 = 1'b1;
  assign CLBLL_L_X2Y150_SLICE_X1Y150_D6 = 1'b1;
  assign CLBLM_L_X10Y155_SLICE_X12Y155_B3 = CLBLM_R_X11Y153_SLICE_X15Y153_DO6;
  assign CLBLM_L_X10Y155_SLICE_X12Y155_B4 = CLBLM_L_X10Y153_SLICE_X13Y153_CQ;
  assign CLBLM_L_X10Y155_SLICE_X12Y155_C6 = 1'b1;
  assign CLBLM_R_X11Y151_SLICE_X15Y151_C3 = 1'b1;
  assign CLBLM_R_X11Y151_SLICE_X15Y151_C4 = 1'b1;
  assign CLBLM_R_X11Y151_SLICE_X15Y151_C5 = 1'b1;
  assign CLBLM_R_X11Y151_SLICE_X15Y151_C6 = 1'b1;
  assign RIOI3_SING_X105Y149_ILOGIC_X1Y149_D = RIOB33_SING_X105Y149_IOB_X1Y149_I;
  assign CLBLM_R_X7Y152_SLICE_X9Y152_A1 = CLBLM_L_X8Y152_SLICE_X10Y152_AQ;
  assign CLBLM_R_X7Y152_SLICE_X9Y152_A2 = CLBLL_L_X4Y151_SLICE_X4Y151_C5Q;
  assign CLBLM_R_X7Y152_SLICE_X9Y152_A3 = CLBLM_R_X7Y152_SLICE_X9Y152_AQ;
  assign CLBLM_R_X7Y152_SLICE_X9Y152_A4 = RIOB33_X105Y131_IOB_X1Y131_I;
  assign CLBLM_R_X7Y152_SLICE_X9Y152_A5 = CLBLM_L_X8Y152_SLICE_X10Y152_BQ;
  assign CLBLM_R_X7Y152_SLICE_X9Y152_A6 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X7Y152_SLICE_X9Y152_B1 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X7Y152_SLICE_X9Y152_B2 = 1'b1;
  assign CLBLM_R_X7Y152_SLICE_X9Y152_B3 = CLBLM_R_X5Y152_SLICE_X7Y152_AQ;
  assign CLBLM_R_X7Y152_SLICE_X9Y152_B4 = CLBLM_L_X10Y149_SLICE_X12Y149_BQ;
  assign CLBLM_R_X7Y152_SLICE_X9Y152_B5 = CLBLM_R_X7Y142_SLICE_X8Y142_D5Q;
  assign CLBLM_R_X7Y152_SLICE_X9Y152_B6 = 1'b1;
  assign CLBLM_R_X11Y151_SLICE_X15Y151_D2 = 1'b1;
  assign CLBLM_R_X5Y142_SLICE_X7Y142_A1 = CLBLM_R_X5Y142_SLICE_X7Y142_AQ;
  assign CLBLM_R_X5Y142_SLICE_X7Y142_A2 = CLBLM_R_X7Y143_SLICE_X9Y143_CQ;
  assign CLBLM_R_X5Y142_SLICE_X7Y142_A3 = CLBLL_L_X4Y149_SLICE_X5Y149_C5Q;
  assign CLBLM_R_X5Y142_SLICE_X7Y142_A4 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X5Y142_SLICE_X7Y142_A5 = CLBLM_R_X5Y147_SLICE_X6Y147_C5Q;
  assign CLBLM_R_X5Y142_SLICE_X7Y142_A6 = 1'b1;
  assign CLBLM_R_X7Y152_SLICE_X9Y152_C1 = CLBLL_L_X4Y143_SLICE_X4Y143_BQ;
  assign CLBLM_R_X7Y152_SLICE_X9Y152_C2 = CLBLM_R_X7Y152_SLICE_X9Y152_AQ;
  assign CLBLM_R_X7Y152_SLICE_X9Y152_C3 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X5Y142_SLICE_X7Y142_B1 = CLBLL_L_X4Y143_SLICE_X4Y143_DQ;
  assign CLBLM_R_X5Y142_SLICE_X7Y142_B2 = CLBLM_R_X5Y141_SLICE_X6Y141_BQ;
  assign CLBLM_R_X5Y142_SLICE_X7Y142_B3 = 1'b1;
  assign CLBLM_R_X5Y142_SLICE_X7Y142_B4 = CLBLL_L_X4Y142_SLICE_X5Y142_C5Q;
  assign CLBLM_R_X5Y142_SLICE_X7Y142_B5 = 1'b1;
  assign CLBLM_R_X5Y142_SLICE_X7Y142_B6 = CLBLM_R_X5Y140_SLICE_X6Y140_A5Q;
  assign CLBLM_R_X7Y152_SLICE_X9Y152_CLK = CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O;
  assign CLBLM_R_X5Y142_SLICE_X7Y142_BX = CLBLM_R_X5Y141_SLICE_X6Y141_CO6;
  assign CLBLM_R_X7Y152_SLICE_X9Y152_D1 = CLBLM_L_X8Y152_SLICE_X10Y152_BQ;
  assign CLBLM_R_X5Y142_SLICE_X7Y142_C1 = CLBLM_R_X5Y147_SLICE_X6Y147_C5Q;
  assign CLBLM_R_X5Y142_SLICE_X7Y142_C2 = CLBLM_R_X5Y144_SLICE_X7Y144_DO6;
  assign CLBLM_R_X5Y142_SLICE_X7Y142_C3 = 1'b1;
  assign CLBLM_R_X5Y142_SLICE_X7Y142_C4 = LIOB33_X0Y61_IOB_X0Y61_I;
  assign CLBLM_R_X5Y142_SLICE_X7Y142_C5 = CLBLM_R_X5Y142_SLICE_X7Y142_AQ;
  assign CLBLM_R_X5Y142_SLICE_X7Y142_C6 = 1'b1;
  assign CLBLM_R_X7Y152_SLICE_X9Y152_D4 = CLBLL_L_X4Y145_SLICE_X5Y145_C5Q;
  assign CLBLM_R_X5Y142_SLICE_X7Y142_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X7Y152_SLICE_X8Y152_A1 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X7Y152_SLICE_X8Y152_A2 = CLBLL_L_X4Y151_SLICE_X4Y151_BQ;
  assign CLBLM_R_X7Y152_SLICE_X8Y152_A3 = CLBLM_R_X3Y145_SLICE_X3Y145_D5Q;
  assign CLBLM_R_X7Y152_SLICE_X8Y152_A4 = CLBLM_R_X7Y152_SLICE_X8Y152_AQ;
  assign CLBLM_R_X7Y152_SLICE_X8Y152_A5 = CLBLM_R_X5Y151_SLICE_X7Y151_BQ;
  assign CLBLM_R_X5Y142_SLICE_X7Y142_D1 = 1'b1;
  assign CLBLM_R_X5Y142_SLICE_X7Y142_D2 = 1'b1;
  assign CLBLM_R_X5Y142_SLICE_X7Y142_D3 = 1'b1;
  assign CLBLM_R_X5Y142_SLICE_X7Y142_D4 = 1'b1;
  assign CLBLM_R_X5Y142_SLICE_X7Y142_D5 = 1'b1;
  assign CLBLM_R_X5Y142_SLICE_X7Y142_D6 = 1'b1;
  assign CLBLM_R_X7Y152_SLICE_X8Y152_A6 = CLBLM_R_X3Y151_SLICE_X3Y151_CQ;
  assign CLBLM_R_X7Y152_SLICE_X8Y152_B1 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X7Y152_SLICE_X8Y152_B2 = CLBLM_R_X3Y151_SLICE_X3Y151_CQ;
  assign CLBLM_R_X7Y152_SLICE_X8Y152_B3 = CLBLL_L_X4Y150_SLICE_X4Y150_AQ;
  assign CLBLM_R_X7Y152_SLICE_X8Y152_B4 = CLBLL_L_X4Y152_SLICE_X4Y152_B5Q;
  assign CLBLM_R_X5Y142_SLICE_X6Y142_A1 = CLBLM_L_X8Y143_SLICE_X11Y143_DQ;
  assign CLBLM_R_X5Y142_SLICE_X6Y142_A2 = CLBLM_R_X3Y151_SLICE_X3Y151_AQ;
  assign CLBLM_R_X5Y142_SLICE_X6Y142_A3 = CLBLM_R_X5Y142_SLICE_X6Y142_AQ;
  assign CLBLM_R_X5Y142_SLICE_X6Y142_A4 = CLBLM_R_X5Y142_SLICE_X7Y142_BQ;
  assign CLBLM_R_X5Y142_SLICE_X6Y142_A5 = CLBLM_L_X10Y145_SLICE_X12Y145_AQ;
  assign CLBLM_R_X5Y142_SLICE_X6Y142_A6 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X7Y152_SLICE_X8Y152_C1 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X7Y152_SLICE_X8Y152_C2 = CLBLM_R_X7Y152_SLICE_X8Y152_CQ;
  assign CLBLM_R_X7Y152_SLICE_X8Y152_C3 = CLBLM_R_X7Y153_SLICE_X8Y153_BQ;
  assign CLBLM_R_X5Y142_SLICE_X6Y142_B1 = CLBLL_L_X2Y146_SLICE_X0Y146_CQ;
  assign CLBLM_R_X5Y142_SLICE_X6Y142_B2 = CLBLM_R_X5Y142_SLICE_X6Y142_BQ;
  assign CLBLM_R_X5Y142_SLICE_X6Y142_B3 = 1'b1;
  assign CLBLM_R_X5Y142_SLICE_X6Y142_B4 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X5Y142_SLICE_X6Y142_B5 = CLBLL_L_X4Y142_SLICE_X5Y142_BQ;
  assign CLBLM_R_X5Y142_SLICE_X6Y142_B6 = CLBLM_R_X13Y149_SLICE_X18Y149_AO6;
  assign CLBLM_R_X7Y152_SLICE_X8Y152_CLK = CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O;
  assign CLBLM_R_X7Y152_SLICE_X8Y152_D1 = CLBLM_L_X12Y151_SLICE_X16Y151_AQ;
  assign CLBLM_R_X7Y152_SLICE_X8Y152_D2 = RIOB33_X105Y111_IOB_X1Y112_I;
  assign CLBLM_R_X5Y142_SLICE_X6Y142_C1 = CLBLM_R_X5Y143_SLICE_X6Y143_AQ;
  assign CLBLM_R_X5Y142_SLICE_X6Y142_C2 = CLBLM_R_X5Y142_SLICE_X6Y142_CQ;
  assign CLBLM_R_X5Y142_SLICE_X6Y142_C3 = CLBLM_R_X13Y149_SLICE_X18Y149_AO6;
  assign CLBLM_R_X5Y142_SLICE_X6Y142_C4 = CLBLM_R_X7Y151_SLICE_X8Y151_C5Q;
  assign CLBLM_R_X5Y142_SLICE_X6Y142_C5 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X5Y142_SLICE_X6Y142_C6 = 1'b1;
  assign CLBLM_R_X7Y152_SLICE_X8Y152_D3 = CLBLM_R_X3Y152_SLICE_X3Y152_BQ;
  assign CLBLM_R_X7Y152_SLICE_X8Y152_D4 = CLBLM_R_X7Y152_SLICE_X8Y152_AQ;
  assign CLBLM_R_X7Y152_SLICE_X8Y152_D5 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X5Y142_SLICE_X6Y142_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X7Y152_SLICE_X8Y152_D6 = 1'b1;
  assign CLBLM_R_X5Y142_SLICE_X6Y142_D1 = CLBLM_R_X3Y142_SLICE_X2Y142_AQ;
  assign CLBLM_R_X5Y142_SLICE_X6Y142_D2 = 1'b1;
  assign CLBLM_R_X5Y142_SLICE_X6Y142_D3 = CLBLM_L_X8Y143_SLICE_X11Y143_DQ;
  assign CLBLM_R_X5Y142_SLICE_X6Y142_D4 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X5Y142_SLICE_X6Y142_D5 = CLBLM_R_X3Y146_SLICE_X2Y146_D5Q;
  assign CLBLM_R_X5Y142_SLICE_X6Y142_D6 = 1'b1;
  assign CLBLM_R_X7Y153_SLICE_X9Y153_C4 = CLBLL_L_X4Y145_SLICE_X5Y145_BQ;
  assign CLBLM_R_X7Y153_SLICE_X9Y153_C5 = CLBLM_R_X7Y149_SLICE_X9Y149_BQ;
  assign CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_I0 = LIOB33_X0Y77_IOB_X0Y78_I;
  assign CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_I1 = 1'b1;
  assign CLBLM_R_X7Y153_SLICE_X9Y153_C6 = 1'b1;
  assign CLBLM_R_X11Y151_SLICE_X14Y151_B5 = CLBLM_R_X11Y151_SLICE_X15Y151_AQ;
  assign CLBLM_R_X11Y151_SLICE_X14Y151_B6 = CLBLM_R_X7Y144_SLICE_X9Y144_B5Q;
  assign CLBLM_R_X11Y151_SLICE_X14Y151_C1 = CLBLM_L_X10Y148_SLICE_X12Y148_AO6;
  assign CLBLM_R_X7Y153_SLICE_X9Y153_D2 = CLBLM_R_X7Y152_SLICE_X9Y152_B5Q;
  assign CLBLM_R_X7Y153_SLICE_X9Y153_D5 = 1'b1;
  assign CLBLM_R_X7Y153_SLICE_X9Y153_D6 = 1'b1;
  assign CLBLM_R_X11Y151_SLICE_X14Y151_C6 = CLBLM_L_X10Y151_SLICE_X13Y151_DO6;
  assign RIOI3_X105Y197_OLOGIC_X1Y198_D1 = CLBLM_L_X12Y150_SLICE_X16Y150_AO5;
  assign RIOI3_SING_X105Y150_OLOGIC_X1Y150_D1 = 1'b1;
  assign RIOI3_SING_X105Y150_OLOGIC_X1Y150_T1 = 1'b1;
  assign RIOI3_X105Y197_OLOGIC_X1Y198_T1 = 1'b1;
  assign LIOB33_X0Y181_IOB_X0Y182_O = RIOB33_X105Y129_IOB_X1Y129_I;
  assign LIOB33_X0Y181_IOB_X0Y181_O = RIOB33_X105Y127_IOB_X1Y128_I;
  assign CLBLM_R_X7Y153_SLICE_X9Y153_A1 = CLBLM_L_X10Y151_SLICE_X13Y151_A5Q;
  assign CLBLM_R_X7Y153_SLICE_X9Y153_A2 = CLBLM_L_X8Y152_SLICE_X10Y152_CQ;
  assign CLBLM_R_X7Y153_SLICE_X9Y153_A3 = CLBLM_R_X7Y153_SLICE_X9Y153_AQ;
  assign CLBLM_R_X7Y153_SLICE_X9Y153_A4 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X7Y153_SLICE_X9Y153_A5 = CLBLL_L_X2Y150_SLICE_X1Y150_AQ;
  assign CLBLM_R_X7Y153_SLICE_X9Y153_A6 = 1'b1;
  assign CLBLM_R_X7Y153_SLICE_X9Y153_B1 = CLBLM_R_X7Y147_SLICE_X9Y147_CQ;
  assign CLBLM_R_X7Y153_SLICE_X9Y153_B2 = CLBLM_R_X7Y153_SLICE_X9Y153_BQ;
  assign CLBLM_R_X7Y153_SLICE_X9Y153_B3 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X7Y153_SLICE_X9Y153_B4 = CLBLM_R_X3Y145_SLICE_X3Y145_D5Q;
  assign CLBLM_R_X7Y153_SLICE_X8Y153_B5 = CLBLL_L_X4Y142_SLICE_X5Y142_DQ;
  assign CLBLM_R_X7Y153_SLICE_X9Y153_B5 = CLBLM_R_X5Y147_SLICE_X6Y147_AQ;
  assign CLBLM_R_X7Y153_SLICE_X9Y153_B6 = CLBLL_L_X4Y151_SLICE_X4Y151_BQ;
  assign CLBLM_R_X7Y153_SLICE_X8Y153_B6 = CLBLM_R_X7Y153_SLICE_X8Y153_BQ;
  assign CLBLM_R_X5Y143_SLICE_X7Y143_A1 = CLBLM_R_X5Y143_SLICE_X6Y143_DQ;
  assign CLBLM_R_X5Y143_SLICE_X7Y143_A2 = CLBLM_L_X8Y149_SLICE_X11Y149_AQ;
  assign CLBLM_R_X5Y143_SLICE_X7Y143_A3 = CLBLM_R_X5Y143_SLICE_X7Y143_AQ;
  assign CLBLM_R_X5Y143_SLICE_X7Y143_A4 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X5Y143_SLICE_X7Y143_A5 = CLBLM_R_X5Y142_SLICE_X6Y142_AQ;
  assign CLBLM_R_X5Y143_SLICE_X7Y143_A6 = CLBLM_R_X7Y143_SLICE_X8Y143_DO6;
  assign CLBLM_R_X7Y153_SLICE_X9Y153_C1 = CLBLM_R_X7Y151_SLICE_X9Y151_D5Q;
  assign CLBLM_R_X7Y153_SLICE_X9Y153_C2 = CLBLM_R_X7Y154_SLICE_X8Y154_AQ;
  assign CLBLM_R_X7Y153_SLICE_X9Y153_C3 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X5Y143_SLICE_X7Y143_B1 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X5Y143_SLICE_X7Y143_B2 = CLBLM_R_X5Y143_SLICE_X7Y143_BQ;
  assign CLBLM_R_X5Y143_SLICE_X7Y143_B3 = CLBLM_R_X3Y145_SLICE_X3Y145_D5Q;
  assign CLBLM_R_X5Y143_SLICE_X7Y143_B4 = CLBLM_R_X7Y145_SLICE_X8Y145_C5Q;
  assign CLBLM_R_X5Y143_SLICE_X7Y143_B5 = CLBLM_R_X3Y151_SLICE_X3Y151_BQ;
  assign CLBLM_R_X5Y143_SLICE_X7Y143_B6 = CLBLL_L_X4Y151_SLICE_X4Y151_BQ;
  assign CLBLM_R_X7Y153_SLICE_X9Y153_CLK = CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O;
  assign CLBLM_R_X7Y153_SLICE_X9Y153_D1 = CLBLM_R_X5Y153_SLICE_X6Y153_AQ;
  assign CLBLM_R_X5Y143_SLICE_X7Y143_C1 = CLBLM_R_X3Y151_SLICE_X3Y151_BQ;
  assign CLBLM_R_X5Y143_SLICE_X7Y143_C2 = CLBLM_R_X5Y143_SLICE_X7Y143_CQ;
  assign CLBLM_R_X5Y143_SLICE_X7Y143_C3 = CLBLM_R_X5Y151_SLICE_X7Y151_AQ;
  assign CLBLM_R_X5Y143_SLICE_X7Y143_C4 = CLBLL_L_X4Y144_SLICE_X5Y144_CQ;
  assign CLBLM_R_X5Y143_SLICE_X7Y143_C5 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X5Y143_SLICE_X7Y143_C6 = 1'b1;
  assign CLBLM_R_X7Y153_SLICE_X9Y153_D3 = CLBLM_R_X7Y143_SLICE_X9Y143_BQ;
  assign CLBLM_R_X7Y153_SLICE_X9Y153_D4 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X5Y143_SLICE_X7Y143_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X7Y153_SLICE_X8Y153_A1 = 1'b1;
  assign CLBLM_R_X7Y153_SLICE_X8Y153_A2 = CLBLM_L_X10Y149_SLICE_X12Y149_BQ;
  assign CLBLM_R_X7Y153_SLICE_X8Y153_A3 = CLBLM_R_X7Y148_SLICE_X8Y148_AQ;
  assign CLBLM_R_X7Y153_SLICE_X8Y153_A4 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X7Y153_SLICE_X8Y153_A5 = CLBLM_R_X3Y153_SLICE_X2Y153_AQ;
  assign CLBLM_R_X5Y143_SLICE_X7Y143_D1 = CLBLM_R_X5Y145_SLICE_X7Y145_AQ;
  assign CLBLM_R_X5Y143_SLICE_X7Y143_D2 = CLBLL_L_X4Y142_SLICE_X5Y142_CQ;
  assign CLBLM_R_X5Y143_SLICE_X7Y143_D3 = 1'b1;
  assign CLBLM_R_X5Y143_SLICE_X7Y143_D4 = CLBLM_R_X5Y141_SLICE_X6Y141_B5Q;
  assign CLBLM_R_X5Y143_SLICE_X7Y143_D5 = CLBLM_R_X7Y144_SLICE_X8Y144_CQ;
  assign CLBLM_R_X5Y143_SLICE_X7Y143_D6 = CLBLM_R_X5Y142_SLICE_X7Y142_BO6;
  assign CLBLM_R_X7Y153_SLICE_X8Y153_A6 = 1'b1;
  assign CLBLM_R_X7Y153_SLICE_X8Y153_B1 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X7Y153_SLICE_X8Y153_B2 = CLBLL_L_X4Y147_SLICE_X5Y147_CQ;
  assign CLBLM_R_X7Y153_SLICE_X8Y153_B3 = CLBLM_L_X8Y153_SLICE_X11Y153_BQ;
  assign CLBLM_R_X7Y153_SLICE_X8Y153_B4 = CLBLM_R_X5Y147_SLICE_X6Y147_BQ;
  assign CLBLM_R_X5Y143_SLICE_X6Y143_A1 = CLBLM_R_X3Y151_SLICE_X2Y151_AQ;
  assign CLBLM_R_X5Y143_SLICE_X6Y143_A2 = CLBLM_R_X7Y142_SLICE_X8Y142_C5Q;
  assign CLBLM_R_X5Y143_SLICE_X6Y143_A3 = CLBLM_R_X5Y143_SLICE_X6Y143_AQ;
  assign CLBLM_R_X5Y143_SLICE_X6Y143_A4 = CLBLM_R_X7Y152_SLICE_X8Y152_D5Q;
  assign CLBLM_R_X5Y143_SLICE_X6Y143_A5 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X5Y143_SLICE_X6Y143_A6 = CLBLL_L_X4Y143_SLICE_X5Y143_DQ;
  assign CLBLM_R_X7Y153_SLICE_X8Y153_C1 = CLBLL_L_X4Y142_SLICE_X5Y142_DQ;
  assign CLBLM_R_X7Y153_SLICE_X8Y153_C2 = CLBLM_R_X7Y153_SLICE_X8Y153_CQ;
  assign CLBLM_R_X7Y153_SLICE_X8Y153_C3 = CLBLM_L_X10Y148_SLICE_X13Y148_C5Q;
  assign CLBLM_R_X5Y143_SLICE_X6Y143_B1 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X5Y143_SLICE_X6Y143_B2 = CLBLL_L_X2Y145_SLICE_X1Y145_DO5;
  assign CLBLM_R_X5Y143_SLICE_X6Y143_B3 = CLBLM_R_X7Y143_SLICE_X8Y143_AQ;
  assign CLBLM_R_X5Y143_SLICE_X6Y143_B4 = 1'b1;
  assign CLBLM_R_X5Y143_SLICE_X6Y143_B5 = CLBLL_L_X2Y146_SLICE_X1Y146_CO5;
  assign CLBLM_R_X5Y143_SLICE_X6Y143_B6 = 1'b1;
  assign CLBLM_R_X7Y153_SLICE_X8Y153_CLK = CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O;
  assign CLBLM_R_X7Y153_SLICE_X8Y153_D1 = 1'b1;
  assign CLBLM_R_X7Y153_SLICE_X8Y153_D2 = CLBLM_R_X7Y147_SLICE_X9Y147_C5Q;
  assign CLBLM_R_X5Y143_SLICE_X6Y143_C1 = RIOB33_X105Y111_IOB_X1Y111_I;
  assign CLBLM_R_X5Y143_SLICE_X6Y143_C2 = CLBLM_R_X5Y143_SLICE_X6Y143_CQ;
  assign CLBLM_R_X5Y143_SLICE_X6Y143_C3 = CLBLM_R_X5Y143_SLICE_X6Y143_D5Q;
  assign CLBLM_R_X5Y143_SLICE_X6Y143_C4 = CLBLM_L_X8Y143_SLICE_X10Y143_BQ;
  assign CLBLM_R_X5Y143_SLICE_X6Y143_C5 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X5Y143_SLICE_X6Y143_C6 = 1'b1;
  assign CLBLM_R_X7Y153_SLICE_X8Y153_D3 = CLBLM_R_X7Y153_SLICE_X8Y153_DQ;
  assign CLBLM_R_X7Y153_SLICE_X8Y153_D4 = CLBLM_R_X7Y153_SLICE_X8Y153_BQ;
  assign CLBLM_R_X7Y153_SLICE_X8Y153_D5 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X5Y143_SLICE_X6Y143_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X7Y153_SLICE_X8Y153_D6 = CLBLM_R_X11Y148_SLICE_X15Y148_AO6;
  assign LIOI3_X0Y111_OLOGIC_X0Y111_T1 = 1'b1;
  assign LIOI3_TBYTETERM_X0Y163_OLOGIC_X0Y164_D1 = RIOB33_X105Y101_IOB_X1Y102_I;
  assign RIOI3_X105Y155_OLOGIC_X1Y155_D1 = 1'b1;
  assign CLBLM_R_X5Y143_SLICE_X6Y143_D1 = CLBLM_R_X5Y153_SLICE_X6Y153_B5Q;
  assign CLBLM_R_X5Y143_SLICE_X6Y143_D2 = CLBLM_R_X5Y143_SLICE_X6Y143_AQ;
  assign CLBLM_R_X5Y143_SLICE_X6Y143_D3 = CLBLM_R_X3Y144_SLICE_X2Y144_AQ;
  assign CLBLM_R_X5Y143_SLICE_X6Y143_D4 = CLBLM_R_X7Y142_SLICE_X8Y142_D5Q;
  assign CLBLM_R_X5Y143_SLICE_X6Y143_D5 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X5Y143_SLICE_X6Y143_D6 = 1'b1;
  assign LIOI3_TBYTETERM_X0Y163_OLOGIC_X0Y164_T1 = 1'b1;
  assign RIOI3_X105Y155_OLOGIC_X1Y155_T1 = 1'b1;
  assign LIOI3_TBYTETERM_X0Y163_OLOGIC_X0Y163_D1 = CLBLM_R_X5Y152_SLICE_X7Y152_DO6;
  assign LIOI3_TBYTETERM_X0Y163_OLOGIC_X0Y163_T1 = 1'b1;
  assign CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_CE0 = 1'b1;
  assign CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_CE1 = 1'b1;
  assign CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_IGNORE0 = 1'b1;
  assign CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_IGNORE1 = 1'b1;
  assign CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_S0 = 1'b1;
  assign CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_S1 = 1'b1;
  assign LIOB33_X0Y63_IOB_X0Y64_O = CLBLM_R_X7Y141_SLICE_X8Y141_AO5;
  assign LIOI3_X0Y51_ILOGIC_X0Y52_D = LIOB33_X0Y51_IOB_X0Y52_I;
  assign LIOI3_X0Y51_ILOGIC_X0Y51_D = LIOB33_X0Y51_IOB_X0Y51_I;
  assign RIOI3_SING_X105Y199_OLOGIC_X1Y199_D1 = CLBLM_R_X7Y153_SLICE_X8Y153_A5Q;
  assign RIOB33_X105Y151_IOB_X1Y152_O = 1'b1;
  assign RIOB33_X105Y151_IOB_X1Y151_O = 1'b1;
  assign RIOI3_SING_X105Y199_OLOGIC_X1Y199_T1 = 1'b1;
  assign CLBLM_R_X7Y154_SLICE_X9Y154_A1 = CLBLL_L_X4Y143_SLICE_X4Y143_AQ;
  assign CLBLM_R_X7Y154_SLICE_X9Y154_A2 = 1'b1;
  assign CLBLM_R_X7Y154_SLICE_X9Y154_A3 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X7Y154_SLICE_X9Y154_A4 = CLBLM_R_X7Y154_SLICE_X9Y154_AQ;
  assign CLBLM_R_X7Y154_SLICE_X9Y154_A5 = CLBLM_R_X5Y150_SLICE_X6Y150_B5Q;
  assign CLBLM_R_X7Y154_SLICE_X9Y154_A6 = CLBLM_R_X7Y154_SLICE_X9Y154_CO6;
  assign LIOI3_TBYTESRC_X0Y57_ILOGIC_X0Y58_D = LIOB33_X0Y57_IOB_X0Y58_I;
  assign LIOI3_TBYTESRC_X0Y57_ILOGIC_X0Y57_D = LIOB33_X0Y57_IOB_X0Y57_I;
  assign CLBLM_R_X7Y154_SLICE_X9Y154_B1 = 1'b1;
  assign CLBLM_R_X7Y154_SLICE_X9Y154_B2 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X7Y154_SLICE_X9Y154_B3 = CLBLL_L_X4Y149_SLICE_X4Y149_AQ;
  assign CLBLM_R_X7Y154_SLICE_X9Y154_B4 = CLBLM_R_X5Y150_SLICE_X6Y150_B5Q;
  assign CLBLM_R_X7Y154_SLICE_X9Y154_B5 = CLBLM_R_X7Y154_SLICE_X9Y154_CO5;
  assign CLBLM_R_X7Y154_SLICE_X9Y154_B6 = CLBLM_R_X7Y154_SLICE_X9Y154_BQ;
  assign CLBLM_R_X5Y144_SLICE_X7Y144_A1 = 1'b1;
  assign CLBLM_R_X5Y144_SLICE_X7Y144_A2 = CLBLL_L_X4Y150_SLICE_X4Y150_C5Q;
  assign CLBLM_R_X5Y144_SLICE_X7Y144_A3 = CLBLM_R_X5Y144_SLICE_X7Y144_AQ;
  assign CLBLM_R_X5Y144_SLICE_X7Y144_A4 = CLBLM_R_X11Y146_SLICE_X14Y146_DO6;
  assign CLBLM_R_X5Y144_SLICE_X7Y144_A5 = CLBLM_R_X3Y150_SLICE_X2Y150_AQ;
  assign CLBLM_R_X5Y144_SLICE_X7Y144_A6 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X7Y154_SLICE_X9Y154_C1 = CLBLM_R_X5Y152_SLICE_X6Y152_BQ;
  assign CLBLM_R_X7Y154_SLICE_X9Y154_C2 = CLBLM_L_X10Y153_SLICE_X12Y153_A5Q;
  assign CLBLM_R_X7Y154_SLICE_X9Y154_C3 = CLBLM_L_X8Y154_SLICE_X11Y154_AQ;
  assign CLBLM_R_X5Y144_SLICE_X7Y144_B1 = 1'b1;
  assign CLBLM_R_X5Y144_SLICE_X7Y144_B2 = CLBLM_R_X3Y146_SLICE_X2Y146_D5Q;
  assign CLBLM_R_X5Y144_SLICE_X7Y144_B3 = CLBLM_R_X5Y151_SLICE_X7Y151_B5Q;
  assign CLBLM_R_X5Y144_SLICE_X7Y144_B4 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X5Y144_SLICE_X7Y144_B5 = CLBLM_R_X5Y144_SLICE_X7Y144_C5Q;
  assign CLBLM_R_X5Y144_SLICE_X7Y144_B6 = 1'b1;
  assign CLBLM_R_X7Y154_SLICE_X9Y154_CLK = CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O;
  assign CLBLM_R_X7Y154_SLICE_X9Y154_D1 = CLBLM_L_X8Y154_SLICE_X11Y154_AQ;
  assign CLBLM_R_X5Y144_SLICE_X7Y144_C1 = CLBLM_R_X5Y143_SLICE_X7Y143_C5Q;
  assign CLBLM_R_X5Y144_SLICE_X7Y144_C2 = 1'b1;
  assign CLBLM_R_X5Y144_SLICE_X7Y144_C3 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X5Y144_SLICE_X7Y144_C4 = CLBLM_R_X7Y144_SLICE_X8Y144_C5Q;
  assign CLBLM_R_X5Y144_SLICE_X7Y144_C5 = CLBLM_L_X8Y145_SLICE_X11Y145_DQ;
  assign CLBLM_R_X5Y144_SLICE_X7Y144_C6 = 1'b1;
  assign CLBLM_R_X7Y154_SLICE_X9Y154_D3 = CLBLM_R_X7Y154_SLICE_X9Y154_BQ;
  assign CLBLM_R_X7Y154_SLICE_X9Y154_D4 = CLBLM_L_X8Y153_SLICE_X11Y153_AQ;
  assign CLBLM_R_X5Y144_SLICE_X7Y144_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X7Y154_SLICE_X8Y154_A1 = CLBLM_R_X7Y148_SLICE_X9Y148_A5Q;
  assign CLBLM_R_X7Y154_SLICE_X8Y154_A2 = CLBLM_R_X5Y150_SLICE_X6Y150_B5Q;
  assign CLBLM_R_X7Y154_SLICE_X8Y154_A3 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X7Y154_SLICE_X8Y154_A5 = 1'b1;
  assign CLBLM_R_X7Y154_SLICE_X8Y154_A6 = CLBLM_R_X7Y155_SLICE_X8Y155_BO5;
  assign CLBLM_R_X5Y144_SLICE_X7Y144_D1 = CLBLM_R_X5Y144_SLICE_X7Y144_C5Q;
  assign CLBLM_R_X5Y144_SLICE_X7Y144_D2 = CLBLL_L_X4Y148_SLICE_X5Y148_B5Q;
  assign CLBLM_R_X5Y144_SLICE_X7Y144_D3 = CLBLM_L_X8Y142_SLICE_X10Y142_A5Q;
  assign CLBLM_R_X5Y144_SLICE_X7Y144_D4 = 1'b1;
  assign CLBLM_R_X5Y144_SLICE_X7Y144_D5 = CLBLM_L_X8Y152_SLICE_X10Y152_C5Q;
  assign CLBLM_R_X5Y144_SLICE_X7Y144_D6 = 1'b1;
  assign CLBLM_R_X7Y154_SLICE_X8Y154_B1 = CLBLM_R_X5Y152_SLICE_X7Y152_C5Q;
  assign CLBLM_R_X7Y154_SLICE_X8Y154_B2 = CLBLM_R_X7Y154_SLICE_X8Y154_BQ;
  assign CLBLM_R_X7Y154_SLICE_X8Y154_B3 = CLBLM_R_X5Y150_SLICE_X6Y150_B5Q;
  assign CLBLM_R_X7Y154_SLICE_X8Y154_B4 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X7Y154_SLICE_X8Y154_B5 = CLBLM_R_X7Y154_SLICE_X8Y154_CO5;
  assign CLBLM_R_X5Y144_SLICE_X6Y144_A1 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X5Y144_SLICE_X6Y144_A2 = CLBLM_R_X5Y152_SLICE_X6Y152_AQ;
  assign CLBLM_R_X5Y144_SLICE_X6Y144_A3 = CLBLM_R_X5Y144_SLICE_X6Y144_AQ;
  assign CLBLM_R_X5Y144_SLICE_X6Y144_A4 = CLBLM_R_X7Y144_SLICE_X8Y144_D5Q;
  assign CLBLM_R_X5Y144_SLICE_X6Y144_A5 = 1'b1;
  assign CLBLM_R_X5Y144_SLICE_X6Y144_A6 = CLBLM_R_X11Y146_SLICE_X14Y146_DO6;
  assign CLBLM_R_X7Y154_SLICE_X8Y154_C1 = CLBLM_R_X5Y152_SLICE_X6Y152_BQ;
  assign CLBLM_R_X7Y154_SLICE_X8Y154_C2 = CLBLM_R_X7Y154_SLICE_X8Y154_AQ;
  assign CLBLM_R_X7Y154_SLICE_X8Y154_C3 = CLBLM_L_X8Y154_SLICE_X10Y154_AQ;
  assign CLBLM_R_X5Y144_SLICE_X6Y144_B1 = CLBLM_R_X13Y149_SLICE_X18Y149_AO6;
  assign CLBLM_R_X5Y144_SLICE_X6Y144_B2 = CLBLM_R_X5Y144_SLICE_X6Y144_BQ;
  assign CLBLM_R_X5Y144_SLICE_X6Y144_B3 = CLBLL_L_X4Y145_SLICE_X4Y145_AQ;
  assign CLBLM_R_X5Y144_SLICE_X6Y144_B4 = CLBLM_L_X8Y150_SLICE_X11Y150_AQ;
  assign CLBLM_R_X5Y144_SLICE_X6Y144_B5 = 1'b1;
  assign CLBLM_R_X5Y144_SLICE_X6Y144_B6 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X7Y154_SLICE_X8Y154_CLK = CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O;
  assign CLBLM_R_X7Y154_SLICE_X8Y154_D1 = CLBLM_R_X7Y155_SLICE_X8Y155_AQ;
  assign CLBLM_R_X7Y154_SLICE_X8Y154_D2 = CLBLM_L_X8Y154_SLICE_X10Y154_AQ;
  assign CLBLM_R_X5Y144_SLICE_X6Y144_C1 = 1'b1;
  assign CLBLM_R_X5Y144_SLICE_X6Y144_C2 = CLBLM_R_X5Y145_SLICE_X6Y145_D5Q;
  assign CLBLM_R_X5Y144_SLICE_X6Y144_C3 = CLBLL_L_X4Y143_SLICE_X4Y143_BQ;
  assign CLBLM_R_X5Y144_SLICE_X6Y144_C4 = CLBLL_L_X4Y145_SLICE_X4Y145_DO5;
  assign CLBLM_R_X5Y144_SLICE_X6Y144_C5 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X5Y144_SLICE_X6Y144_C6 = CLBLM_R_X5Y144_SLICE_X6Y144_D5Q;
  assign CLBLM_R_X7Y154_SLICE_X8Y154_D3 = CLBLM_R_X7Y154_SLICE_X9Y154_DO6;
  assign CLBLM_R_X7Y154_SLICE_X8Y154_D4 = CLBLM_R_X7Y154_SLICE_X8Y154_BQ;
  assign CLBLM_R_X7Y154_SLICE_X8Y154_D5 = 1'b1;
  assign CLBLM_R_X5Y144_SLICE_X6Y144_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X7Y154_SLICE_X8Y154_D6 = CLBLM_R_X7Y154_SLICE_X8Y154_AQ;
  assign CLBLM_R_X5Y144_SLICE_X6Y144_D1 = CLBLM_R_X5Y144_SLICE_X6Y144_BQ;
  assign CLBLM_R_X5Y144_SLICE_X6Y144_D2 = CLBLL_L_X4Y144_SLICE_X4Y144_BQ;
  assign CLBLM_R_X5Y144_SLICE_X6Y144_D3 = CLBLM_R_X5Y145_SLICE_X6Y145_D5Q;
  assign CLBLM_R_X5Y144_SLICE_X6Y144_D4 = CLBLL_L_X4Y144_SLICE_X4Y144_D5Q;
  assign CLBLM_R_X5Y144_SLICE_X6Y144_D5 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X5Y144_SLICE_X6Y144_D6 = 1'b1;
  assign LIOB33_X0Y65_IOB_X0Y66_O = CLBLL_L_X4Y151_SLICE_X4Y151_CQ;
  assign LIOB33_X0Y65_IOB_X0Y65_O = CLBLM_R_X7Y141_SLICE_X8Y141_BO6;
  assign RIOB33_X105Y153_IOB_X1Y154_O = 1'b1;
  assign RIOB33_X105Y153_IOB_X1Y153_O = 1'b1;
  assign LIOB33_X0Y185_IOB_X0Y186_O = RIOB33_X105Y119_IOB_X1Y120_I;
  assign LIOB33_X0Y185_IOB_X0Y185_O = RIOB33_X105Y133_IOB_X1Y133_I;
  assign CLBLM_R_X7Y155_SLICE_X9Y155_A1 = 1'b1;
  assign CLBLM_R_X7Y155_SLICE_X9Y155_A2 = 1'b1;
  assign CLBLM_R_X3Y147_SLICE_X3Y147_B1 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X7Y155_SLICE_X9Y155_A3 = 1'b1;
  assign CLBLM_R_X7Y155_SLICE_X9Y155_A4 = 1'b1;
  assign CLBLM_R_X7Y155_SLICE_X9Y155_A5 = 1'b1;
  assign CLBLM_R_X7Y155_SLICE_X9Y155_A6 = 1'b1;
  assign CLBLM_R_X3Y147_SLICE_X3Y147_B2 = CLBLM_R_X3Y147_SLICE_X3Y147_BQ;
  assign CLBLM_R_X7Y155_SLICE_X9Y155_B1 = 1'b1;
  assign CLBLM_R_X7Y155_SLICE_X9Y155_B2 = 1'b1;
  assign CLBLM_R_X3Y147_SLICE_X3Y147_B3 = RIOB33_X105Y119_IOB_X1Y119_I;
  assign CLBLM_R_X7Y155_SLICE_X9Y155_B3 = 1'b1;
  assign CLBLM_R_X7Y155_SLICE_X9Y155_B4 = 1'b1;
  assign CLBLM_R_X7Y155_SLICE_X9Y155_B5 = 1'b1;
  assign CLBLM_R_X7Y155_SLICE_X9Y155_B6 = 1'b1;
  assign CLBLM_R_X5Y145_SLICE_X7Y145_A1 = CLBLM_R_X5Y147_SLICE_X7Y147_CQ;
  assign CLBLM_R_X5Y145_SLICE_X7Y145_A2 = CLBLM_R_X3Y145_SLICE_X2Y145_B5Q;
  assign CLBLM_R_X5Y145_SLICE_X7Y145_A3 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X5Y145_SLICE_X7Y145_A4 = 1'b1;
  assign CLBLM_R_X5Y145_SLICE_X7Y145_A5 = CLBLM_L_X10Y153_SLICE_X13Y153_A5Q;
  assign CLBLM_R_X5Y145_SLICE_X7Y145_A6 = 1'b1;
  assign CLBLM_R_X7Y155_SLICE_X9Y155_C1 = 1'b1;
  assign CLBLM_R_X7Y155_SLICE_X9Y155_C2 = 1'b1;
  assign CLBLM_R_X7Y155_SLICE_X9Y155_C3 = 1'b1;
  assign CLBLM_R_X5Y145_SLICE_X7Y145_B1 = CLBLM_L_X8Y144_SLICE_X10Y144_AO5;
  assign CLBLM_R_X5Y145_SLICE_X7Y145_B2 = CLBLL_L_X4Y147_SLICE_X4Y147_D5Q;
  assign CLBLM_R_X5Y145_SLICE_X7Y145_B3 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X5Y145_SLICE_X7Y145_B4 = CLBLM_L_X10Y144_SLICE_X12Y144_AO6;
  assign CLBLM_R_X5Y145_SLICE_X7Y145_B5 = CLBLM_L_X10Y151_SLICE_X12Y151_CQ;
  assign CLBLM_R_X5Y145_SLICE_X7Y145_B6 = 1'b1;
  assign CLBLM_R_X7Y155_SLICE_X9Y155_D1 = 1'b1;
  assign CLBLM_R_X7Y155_SLICE_X9Y155_D2 = 1'b1;
  assign CLBLM_R_X5Y145_SLICE_X7Y145_C1 = CLBLM_R_X3Y147_SLICE_X3Y147_C5Q;
  assign CLBLM_R_X5Y145_SLICE_X7Y145_C2 = CLBLM_R_X3Y148_SLICE_X3Y148_BQ;
  assign CLBLM_R_X5Y145_SLICE_X7Y145_C3 = CLBLL_L_X4Y146_SLICE_X4Y146_C5Q;
  assign CLBLM_R_X5Y145_SLICE_X7Y145_C4 = CLBLM_R_X5Y143_SLICE_X7Y143_DO6;
  assign CLBLM_R_X5Y145_SLICE_X7Y145_C5 = CLBLM_R_X5Y145_SLICE_X7Y145_DO6;
  assign CLBLM_R_X5Y145_SLICE_X7Y145_C6 = CLBLM_R_X5Y147_SLICE_X7Y147_B5Q;
  assign CLBLM_R_X7Y155_SLICE_X9Y155_D3 = 1'b1;
  assign CLBLM_R_X7Y155_SLICE_X9Y155_D4 = 1'b1;
  assign CLBLM_R_X5Y145_SLICE_X7Y145_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X7Y155_SLICE_X8Y155_A1 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X7Y155_SLICE_X8Y155_A2 = CLBLM_R_X7Y154_SLICE_X9Y154_CO6;
  assign CLBLM_R_X7Y155_SLICE_X8Y155_A3 = CLBLM_R_X7Y155_SLICE_X8Y155_AQ;
  assign CLBLM_R_X7Y155_SLICE_X8Y155_A4 = CLBLL_L_X4Y140_SLICE_X4Y140_A5Q;
  assign CLBLM_R_X7Y155_SLICE_X8Y155_A5 = CLBLM_R_X7Y154_SLICE_X9Y154_AQ;
  assign CLBLM_R_X5Y145_SLICE_X7Y145_D1 = 1'b1;
  assign CLBLM_R_X5Y145_SLICE_X7Y145_D2 = CLBLM_R_X7Y145_SLICE_X8Y145_BQ;
  assign CLBLM_R_X5Y145_SLICE_X7Y145_D3 = CLBLM_R_X7Y146_SLICE_X8Y146_DQ;
  assign CLBLM_R_X5Y145_SLICE_X7Y145_D4 = CLBLM_R_X5Y146_SLICE_X7Y146_D5Q;
  assign CLBLM_R_X5Y145_SLICE_X7Y145_D5 = CLBLM_R_X3Y145_SLICE_X2Y145_B5Q;
  assign CLBLM_R_X5Y145_SLICE_X7Y145_D6 = 1'b1;
  assign CLBLM_R_X7Y155_SLICE_X8Y155_A6 = CLBLM_R_X5Y150_SLICE_X6Y150_B5Q;
  assign CLBLM_R_X7Y155_SLICE_X8Y155_AX = CLBLM_R_X7Y155_SLICE_X8Y155_BO6;
  assign CLBLM_R_X7Y155_SLICE_X8Y155_B1 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X7Y155_SLICE_X8Y155_B2 = CLBLM_R_X7Y154_SLICE_X9Y154_CO6;
  assign CLBLM_R_X7Y155_SLICE_X8Y155_B3 = CLBLM_R_X7Y155_SLICE_X8Y155_AQ;
  assign CLBLM_R_X7Y155_SLICE_X8Y155_B4 = CLBLL_L_X4Y153_SLICE_X4Y153_BQ;
  assign CLBLM_R_X5Y145_SLICE_X6Y145_A1 = RIOB33_X105Y109_IOB_X1Y109_I;
  assign CLBLM_R_X5Y145_SLICE_X6Y145_A2 = CLBLM_R_X5Y147_SLICE_X7Y147_C5Q;
  assign CLBLM_R_X5Y145_SLICE_X6Y145_A3 = CLBLM_R_X5Y145_SLICE_X6Y145_AQ;
  assign CLBLM_R_X5Y145_SLICE_X6Y145_A4 = CLBLL_L_X2Y146_SLICE_X0Y146_BQ;
  assign CLBLM_R_X5Y145_SLICE_X6Y145_A5 = CLBLM_R_X7Y151_SLICE_X9Y151_A5Q;
  assign CLBLM_R_X5Y145_SLICE_X6Y145_A6 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X7Y155_SLICE_X8Y155_C1 = 1'b1;
  assign CLBLM_R_X7Y155_SLICE_X8Y155_C2 = 1'b1;
  assign CLBLM_R_X7Y155_SLICE_X8Y155_C3 = 1'b1;
  assign CLBLM_R_X5Y145_SLICE_X6Y145_B1 = CLBLL_L_X4Y145_SLICE_X5Y145_CQ;
  assign CLBLM_R_X5Y145_SLICE_X6Y145_B2 = CLBLL_L_X4Y151_SLICE_X4Y151_AQ;
  assign CLBLM_R_X5Y145_SLICE_X6Y145_B3 = CLBLM_R_X5Y145_SLICE_X6Y145_AQ;
  assign CLBLM_R_X5Y145_SLICE_X6Y145_B4 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X5Y145_SLICE_X6Y145_B5 = CLBLM_R_X7Y149_SLICE_X8Y149_A5Q;
  assign CLBLM_R_X5Y145_SLICE_X6Y145_B6 = 1'b1;
  assign CLBLM_R_X7Y155_SLICE_X8Y155_CLK = CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O;
  assign CLBLM_R_X7Y155_SLICE_X8Y155_D1 = 1'b1;
  assign CLBLM_R_X7Y155_SLICE_X8Y155_D2 = 1'b1;
  assign CLBLM_R_X5Y145_SLICE_X6Y145_C1 = CLBLM_L_X8Y142_SLICE_X10Y142_A5Q;
  assign CLBLM_R_X5Y145_SLICE_X6Y145_C2 = CLBLM_R_X3Y146_SLICE_X2Y146_D5Q;
  assign CLBLM_R_X5Y145_SLICE_X6Y145_C3 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X5Y145_SLICE_X6Y145_C4 = CLBLM_R_X5Y142_SLICE_X6Y142_DQ;
  assign CLBLM_R_X5Y145_SLICE_X6Y145_C5 = 1'b1;
  assign CLBLM_R_X5Y145_SLICE_X6Y145_C6 = 1'b1;
  assign CLBLM_R_X7Y155_SLICE_X8Y155_D3 = 1'b1;
  assign CLBLM_R_X7Y155_SLICE_X8Y155_D4 = 1'b1;
  assign CLBLM_R_X7Y155_SLICE_X8Y155_D5 = 1'b1;
  assign CLBLM_R_X5Y145_SLICE_X6Y145_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X7Y155_SLICE_X8Y155_D6 = 1'b1;
  assign CLBLM_R_X5Y145_SLICE_X6Y145_D1 = CLBLM_R_X3Y145_SLICE_X2Y145_CQ;
  assign CLBLM_R_X5Y145_SLICE_X6Y145_D2 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X5Y145_SLICE_X6Y145_D3 = CLBLM_R_X3Y151_SLICE_X3Y151_AQ;
  assign CLBLM_R_X5Y145_SLICE_X6Y145_D4 = CLBLM_R_X5Y149_SLICE_X7Y149_CQ;
  assign CLBLM_R_X5Y145_SLICE_X6Y145_D5 = CLBLM_R_X5Y145_SLICE_X6Y145_D5Q;
  assign CLBLM_R_X5Y145_SLICE_X6Y145_D6 = 1'b1;
  assign LIOI3_X0Y175_OLOGIC_X0Y176_D1 = RIOB33_X105Y115_IOB_X1Y116_I;
  assign LIOI3_X0Y175_OLOGIC_X0Y176_T1 = 1'b1;
  assign LIOI3_X0Y115_OLOGIC_X0Y116_D1 = CLBLM_R_X7Y143_SLICE_X9Y143_B5Q;
  assign LIOI3_X0Y175_OLOGIC_X0Y175_D1 = RIOB33_X105Y123_IOB_X1Y123_I;
  assign LIOI3_X0Y115_OLOGIC_X0Y116_T1 = 1'b1;
  assign RIOI3_X105Y159_OLOGIC_X1Y160_D1 = 1'b1;
  assign LIOI3_X0Y175_OLOGIC_X0Y175_T1 = 1'b1;
  assign LIOI3_X0Y115_OLOGIC_X0Y115_D1 = CLBLM_R_X5Y147_SLICE_X6Y147_C5Q;
  assign RIOI3_X105Y159_OLOGIC_X1Y160_T1 = 1'b1;
  assign LIOI3_TBYTETERM_X0Y187_OLOGIC_X0Y188_D1 = CLBLM_R_X5Y147_SLICE_X6Y147_AQ;
  assign LIOI3_X0Y115_OLOGIC_X0Y115_T1 = 1'b1;
  assign RIOI3_X105Y159_OLOGIC_X1Y159_D1 = 1'b1;
  assign LIOI3_TBYTETERM_X0Y187_OLOGIC_X0Y188_T1 = 1'b1;
  assign RIOI3_X105Y159_OLOGIC_X1Y159_T1 = 1'b1;
  assign RIOB33_X105Y155_IOB_X1Y156_O = 1'b1;
  assign RIOB33_X105Y155_IOB_X1Y155_O = 1'b1;
  assign LIOI3_TBYTETERM_X0Y187_OLOGIC_X0Y187_D1 = CLBLM_L_X8Y145_SLICE_X11Y145_DQ;
  assign LIOI3_TBYTETERM_X0Y187_OLOGIC_X0Y187_T1 = 1'b1;
  assign LIOB33_X0Y187_IOB_X0Y188_O = CLBLM_R_X5Y147_SLICE_X6Y147_AQ;
  assign LIOB33_X0Y187_IOB_X0Y187_O = CLBLM_L_X8Y145_SLICE_X11Y145_DQ;
  assign CLBLM_R_X5Y146_SLICE_X7Y146_A1 = CLBLL_L_X4Y146_SLICE_X4Y146_BQ;
  assign CLBLM_R_X5Y146_SLICE_X7Y146_A2 = CLBLM_R_X7Y152_SLICE_X8Y152_D5Q;
  assign CLBLM_R_X5Y146_SLICE_X7Y146_A3 = CLBLM_R_X5Y146_SLICE_X7Y146_AQ;
  assign CLBLM_R_X5Y146_SLICE_X7Y146_A4 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X5Y146_SLICE_X7Y146_A5 = CLBLL_L_X2Y145_SLICE_X1Y145_AQ;
  assign CLBLM_R_X5Y146_SLICE_X7Y146_A6 = CLBLM_R_X7Y142_SLICE_X8Y142_C5Q;
  assign CLBLM_R_X5Y146_SLICE_X7Y146_B1 = 1'b1;
  assign CLBLM_R_X5Y146_SLICE_X7Y146_B2 = CLBLM_R_X5Y145_SLICE_X6Y145_D5Q;
  assign CLBLM_R_X5Y146_SLICE_X7Y146_B3 = CLBLL_L_X4Y145_SLICE_X4Y145_DO5;
  assign CLBLM_R_X5Y146_SLICE_X7Y146_B4 = CLBLM_L_X8Y148_SLICE_X11Y148_BQ;
  assign CLBLM_R_X5Y146_SLICE_X7Y146_B5 = CLBLL_L_X4Y143_SLICE_X4Y143_BQ;
  assign CLBLM_R_X5Y146_SLICE_X7Y146_B6 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X5Y146_SLICE_X7Y146_C1 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X5Y146_SLICE_X7Y146_C2 = CLBLM_L_X12Y151_SLICE_X16Y151_AQ;
  assign CLBLM_R_X5Y146_SLICE_X7Y146_C3 = CLBLM_R_X3Y146_SLICE_X2Y146_AQ;
  assign CLBLM_R_X5Y146_SLICE_X7Y146_C4 = 1'b1;
  assign CLBLM_R_X5Y146_SLICE_X7Y146_C5 = CLBLM_R_X5Y145_SLICE_X7Y145_BQ;
  assign CLBLM_R_X5Y146_SLICE_X7Y146_C6 = 1'b1;
  assign CLBLM_R_X5Y146_SLICE_X7Y146_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X5Y146_SLICE_X7Y146_D1 = CLBLM_L_X8Y154_SLICE_X11Y154_AQ;
  assign CLBLM_R_X5Y146_SLICE_X7Y146_D2 = CLBLM_L_X8Y152_SLICE_X10Y152_DQ;
  assign CLBLM_R_X5Y146_SLICE_X7Y146_D3 = CLBLM_R_X3Y145_SLICE_X2Y145_B5Q;
  assign CLBLM_R_X5Y146_SLICE_X7Y146_D4 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X5Y146_SLICE_X7Y146_D5 = CLBLM_R_X5Y149_SLICE_X6Y149_B5Q;
  assign CLBLM_R_X5Y146_SLICE_X7Y146_D6 = 1'b1;
  assign CLBLM_R_X5Y146_SLICE_X6Y146_A1 = 1'b1;
  assign CLBLM_R_X5Y146_SLICE_X6Y146_A2 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X5Y146_SLICE_X6Y146_A3 = CLBLM_R_X5Y146_SLICE_X6Y146_AQ;
  assign CLBLM_R_X5Y146_SLICE_X6Y146_A4 = CLBLM_R_X5Y147_SLICE_X6Y147_BQ;
  assign CLBLM_R_X5Y146_SLICE_X6Y146_A5 = CLBLL_L_X4Y144_SLICE_X5Y144_AQ;
  assign CLBLM_R_X5Y146_SLICE_X6Y146_A6 = CLBLM_R_X11Y148_SLICE_X15Y148_AO6;
  assign CLBLM_R_X5Y146_SLICE_X6Y146_B1 = 1'b1;
  assign CLBLM_R_X5Y146_SLICE_X6Y146_B2 = CLBLM_R_X3Y146_SLICE_X3Y146_BQ;
  assign CLBLM_R_X5Y146_SLICE_X6Y146_B3 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X5Y146_SLICE_X6Y146_B4 = CLBLM_R_X7Y149_SLICE_X8Y149_A5Q;
  assign CLBLM_R_X5Y146_SLICE_X6Y146_B5 = CLBLL_L_X4Y149_SLICE_X5Y149_C5Q;
  assign CLBLM_R_X5Y146_SLICE_X6Y146_B6 = 1'b1;
  assign LIOI3_X0Y53_ILOGIC_X0Y54_D = LIOB33_X0Y53_IOB_X0Y54_I;
  assign LIOI3_X0Y53_ILOGIC_X0Y53_D = LIOB33_X0Y53_IOB_X0Y53_I;
  assign CLBLM_R_X5Y146_SLICE_X6Y146_C1 = CLBLL_L_X2Y145_SLICE_X1Y145_AQ;
  assign CLBLM_R_X5Y146_SLICE_X6Y146_C2 = CLBLM_R_X3Y149_SLICE_X2Y149_BQ;
  assign CLBLM_R_X5Y146_SLICE_X6Y146_C3 = 1'b1;
  assign CLBLM_R_X5Y146_SLICE_X6Y146_C4 = 1'b1;
  assign CLBLM_R_X5Y146_SLICE_X6Y146_C5 = CLBLM_R_X7Y147_SLICE_X9Y147_DQ;
  assign CLBLM_R_X5Y146_SLICE_X6Y146_C6 = CLBLM_R_X5Y142_SLICE_X7Y142_A5Q;
  assign CLBLM_R_X5Y146_SLICE_X6Y146_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X5Y146_SLICE_X6Y146_D1 = 1'b1;
  assign CLBLM_R_X5Y146_SLICE_X6Y146_D2 = 1'b1;
  assign CLBLM_R_X5Y146_SLICE_X6Y146_D3 = CLBLM_R_X3Y147_SLICE_X2Y147_BQ;
  assign CLBLM_R_X5Y146_SLICE_X6Y146_D4 = CLBLL_L_X4Y144_SLICE_X4Y144_DQ;
  assign CLBLM_R_X5Y146_SLICE_X6Y146_D5 = CLBLM_R_X3Y145_SLICE_X3Y145_C5Q;
  assign CLBLM_R_X5Y146_SLICE_X6Y146_D6 = CLBLM_R_X3Y147_SLICE_X2Y147_AQ;
  assign RIOB33_X105Y157_IOB_X1Y158_O = 1'b1;
  assign RIOB33_X105Y157_IOB_X1Y157_O = 1'b1;
  assign LIOB33_X0Y189_IOB_X0Y190_O = CLBLM_L_X10Y154_SLICE_X12Y154_CO5;
  assign LIOB33_X0Y189_IOB_X0Y189_O = CLBLM_L_X8Y147_SLICE_X10Y147_BQ;
  assign CLBLM_R_X11Y152_SLICE_X15Y152_C3 = 1'b1;
  assign CLBLM_R_X11Y152_SLICE_X15Y152_C4 = CLBLM_L_X10Y151_SLICE_X13Y151_CO6;
  assign CLBLM_R_X11Y152_SLICE_X15Y152_C5 = 1'b1;
  assign CLBLM_R_X11Y152_SLICE_X15Y152_C6 = 1'b1;
  assign LIOI3_X0Y61_ILOGIC_X0Y62_D = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X5Y147_SLICE_X7Y147_A1 = CLBLM_R_X5Y149_SLICE_X7Y149_DQ;
  assign CLBLM_R_X5Y147_SLICE_X7Y147_A2 = CLBLM_L_X8Y147_SLICE_X10Y147_C5Q;
  assign CLBLM_R_X5Y147_SLICE_X7Y147_A3 = CLBLM_R_X5Y147_SLICE_X7Y147_AQ;
  assign CLBLM_R_X5Y147_SLICE_X7Y147_A4 = CLBLM_L_X10Y144_SLICE_X13Y144_CQ;
  assign CLBLM_R_X5Y147_SLICE_X7Y147_A5 = CLBLM_R_X5Y148_SLICE_X7Y148_C5Q;
  assign CLBLM_R_X5Y147_SLICE_X7Y147_A6 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X11Y152_SLICE_X15Y152_D1 = 1'b1;
  assign CLBLM_R_X11Y152_SLICE_X15Y152_D2 = 1'b1;
  assign CLBLM_R_X5Y147_SLICE_X7Y147_B1 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X5Y147_SLICE_X7Y147_B2 = CLBLM_R_X7Y154_SLICE_X8Y154_BQ;
  assign CLBLM_R_X5Y147_SLICE_X7Y147_B3 = RIOB33_X105Y123_IOB_X1Y124_I;
  assign CLBLM_R_X5Y147_SLICE_X7Y147_B4 = CLBLM_R_X7Y147_SLICE_X9Y147_CQ;
  assign CLBLM_R_X5Y147_SLICE_X7Y147_B5 = CLBLM_R_X3Y147_SLICE_X3Y147_C5Q;
  assign CLBLM_R_X5Y147_SLICE_X7Y147_B6 = 1'b1;
  assign CLBLM_R_X5Y147_SLICE_X7Y147_C1 = CLBLM_R_X7Y151_SLICE_X9Y151_DQ;
  assign CLBLM_R_X5Y147_SLICE_X7Y147_C2 = CLBLM_R_X5Y145_SLICE_X6Y145_D5Q;
  assign CLBLM_R_X5Y147_SLICE_X7Y147_C3 = RIOB33_X105Y109_IOB_X1Y109_I;
  assign CLBLM_R_X5Y147_SLICE_X7Y147_C4 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X5Y147_SLICE_X7Y147_C5 = CLBLM_L_X10Y153_SLICE_X12Y153_A5Q;
  assign CLBLM_R_X5Y147_SLICE_X7Y147_C6 = 1'b1;
  assign CLBLM_R_X11Y152_SLICE_X15Y152_D5 = 1'b1;
  assign CLBLM_R_X5Y147_SLICE_X7Y147_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X11Y152_SLICE_X15Y152_D6 = 1'b1;
  assign CLBLM_R_X5Y147_SLICE_X7Y147_D1 = CLBLM_R_X7Y151_SLICE_X9Y151_DQ;
  assign CLBLM_R_X5Y147_SLICE_X7Y147_D2 = CLBLM_R_X7Y147_SLICE_X8Y147_AO6;
  assign CLBLM_R_X5Y147_SLICE_X7Y147_D3 = CLBLM_R_X7Y153_SLICE_X9Y153_CQ;
  assign CLBLM_R_X5Y147_SLICE_X7Y147_D4 = CLBLM_R_X3Y148_SLICE_X2Y148_DO6;
  assign CLBLM_R_X5Y147_SLICE_X7Y147_D5 = 1'b1;
  assign CLBLM_R_X5Y147_SLICE_X7Y147_D6 = CLBLM_L_X8Y148_SLICE_X10Y148_BQ;
  assign CLBLM_R_X5Y147_SLICE_X6Y147_A1 = CLBLL_L_X4Y150_SLICE_X4Y150_DO6;
  assign CLBLM_R_X5Y147_SLICE_X6Y147_A2 = CLBLL_L_X4Y146_SLICE_X5Y146_BQ;
  assign CLBLM_R_X5Y147_SLICE_X6Y147_A3 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X5Y147_SLICE_X6Y147_A4 = CLBLL_L_X2Y150_SLICE_X1Y150_AQ;
  assign CLBLM_R_X5Y147_SLICE_X6Y147_A5 = CLBLM_R_X5Y146_SLICE_X7Y146_BQ;
  assign CLBLM_R_X5Y147_SLICE_X6Y147_A6 = CLBLM_L_X8Y147_SLICE_X11Y147_CQ;
  assign CLBLM_R_X5Y147_SLICE_X6Y147_B1 = CLBLM_R_X5Y153_SLICE_X6Y153_B5Q;
  assign CLBLM_R_X5Y147_SLICE_X6Y147_B2 = CLBLM_R_X7Y144_SLICE_X8Y144_B5Q;
  assign CLBLM_R_X5Y147_SLICE_X6Y147_B3 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X5Y147_SLICE_X6Y147_B4 = CLBLM_R_X3Y150_SLICE_X3Y150_BQ;
  assign CLBLM_R_X5Y147_SLICE_X6Y147_B5 = CLBLL_L_X4Y151_SLICE_X4Y151_AQ;
  assign CLBLM_R_X5Y147_SLICE_X6Y147_B6 = 1'b1;
  assign CLBLM_R_X5Y147_SLICE_X6Y147_C1 = CLBLL_L_X4Y143_SLICE_X4Y143_BQ;
  assign CLBLM_R_X5Y147_SLICE_X6Y147_C2 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X5Y147_SLICE_X6Y147_C3 = CLBLM_R_X7Y153_SLICE_X8Y153_AQ;
  assign CLBLM_R_X5Y147_SLICE_X6Y147_C4 = CLBLL_L_X4Y151_SLICE_X4Y151_CQ;
  assign CLBLM_R_X5Y147_SLICE_X6Y147_C5 = CLBLM_L_X8Y154_SLICE_X10Y154_BO5;
  assign CLBLM_R_X5Y147_SLICE_X6Y147_C6 = 1'b1;
  assign CLBLM_R_X5Y147_SLICE_X6Y147_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X5Y147_SLICE_X6Y147_D1 = CLBLM_R_X3Y147_SLICE_X2Y147_AQ;
  assign CLBLM_R_X5Y147_SLICE_X6Y147_D2 = CLBLM_R_X7Y144_SLICE_X8Y144_D5Q;
  assign CLBLM_R_X5Y147_SLICE_X6Y147_D3 = 1'b1;
  assign CLBLM_R_X5Y147_SLICE_X6Y147_D4 = CLBLM_R_X5Y145_SLICE_X7Y145_A5Q;
  assign CLBLM_R_X5Y147_SLICE_X6Y147_D5 = 1'b1;
  assign CLBLM_R_X5Y147_SLICE_X6Y147_D6 = CLBLM_R_X3Y147_SLICE_X2Y147_BQ;
  assign CLBLM_L_X10Y146_SLICE_X13Y146_B1 = CLBLM_L_X10Y148_SLICE_X13Y148_CQ;
  assign CLBLM_L_X10Y146_SLICE_X13Y146_B2 = CLBLM_L_X10Y146_SLICE_X13Y146_BQ;
  assign CLBLM_L_X10Y146_SLICE_X13Y146_B3 = CLBLM_L_X8Y146_SLICE_X11Y146_CQ;
  assign CLBLM_L_X10Y146_SLICE_X13Y146_B4 = CLBLM_L_X10Y145_SLICE_X12Y145_AQ;
  assign CLBLM_L_X10Y146_SLICE_X13Y146_B5 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_L_X10Y146_SLICE_X13Y146_B6 = CLBLM_R_X5Y142_SLICE_X7Y142_BQ;
  assign CLBLM_R_X7Y154_SLICE_X9Y154_C4 = CLBLM_R_X7Y154_SLICE_X9Y154_BQ;
  assign CLBLM_R_X7Y154_SLICE_X9Y154_C5 = CLBLM_L_X8Y153_SLICE_X11Y153_AQ;
  assign CLBLM_R_X7Y154_SLICE_X9Y154_C6 = 1'b1;
  assign CLBLM_R_X11Y152_SLICE_X14Y152_B4 = 1'b1;
  assign CLBLM_L_X10Y146_SLICE_X13Y146_C1 = CLBLM_L_X10Y145_SLICE_X12Y145_AQ;
  assign CLBLM_R_X11Y152_SLICE_X14Y152_B5 = 1'b1;
  assign LIOB33_X0Y183_IOB_X0Y184_O = RIOB33_X105Y131_IOB_X1Y132_I;
  assign CLBLM_L_X10Y146_SLICE_X13Y146_C2 = CLBLM_L_X10Y146_SLICE_X13Y146_CQ;
  assign CLBLM_R_X11Y152_SLICE_X14Y152_B6 = 1'b1;
  assign LIOB33_X0Y183_IOB_X0Y183_O = RIOB33_X105Y129_IOB_X1Y130_I;
  assign RIOB33_X105Y159_IOB_X1Y159_O = 1'b1;
  assign RIOB33_X105Y159_IOB_X1Y160_O = 1'b1;
  assign CLBLM_L_X10Y146_SLICE_X13Y146_C3 = CLBLM_R_X5Y142_SLICE_X7Y142_BQ;
  assign CLBLM_L_X10Y146_SLICE_X13Y146_C4 = CLBLM_L_X10Y146_SLICE_X13Y146_BQ;
  assign CLBLM_L_X10Y146_SLICE_X13Y146_C5 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_L_X10Y146_SLICE_X13Y146_C6 = CLBLL_L_X4Y144_SLICE_X5Y144_D5Q;
  assign CLBLM_R_X7Y154_SLICE_X9Y154_D2 = CLBLM_R_X7Y154_SLICE_X9Y154_AQ;
  assign CLBLM_R_X11Y152_SLICE_X14Y152_C4 = 1'b1;
  assign CLBLM_R_X7Y154_SLICE_X9Y154_D5 = 1'b1;
  assign CLBLM_R_X11Y152_SLICE_X14Y152_C5 = 1'b1;
  assign LIOB33_X0Y191_IOB_X0Y191_O = CLBLL_L_X2Y148_SLICE_X1Y148_CO6;
  assign LIOB33_X0Y191_IOB_X0Y192_O = CLBLL_L_X4Y153_SLICE_X4Y153_DO5;
  assign CLBLM_R_X7Y154_SLICE_X9Y154_D6 = CLBLM_L_X10Y153_SLICE_X12Y153_A5Q;
  assign CLBLM_R_X11Y152_SLICE_X14Y152_C6 = 1'b1;
  assign LIOI3_X0Y177_OLOGIC_X0Y178_D1 = RIOB33_X105Y125_IOB_X1Y125_I;
  assign CLBLM_R_X7Y154_SLICE_X8Y154_A4 = CLBLM_R_X7Y154_SLICE_X8Y154_AQ;
  assign LIOI3_X0Y177_OLOGIC_X0Y178_T1 = 1'b1;
  assign LIOI3_X0Y117_OLOGIC_X0Y118_D1 = CLBLM_R_X7Y142_SLICE_X9Y142_BQ;
  assign LIOI3_X0Y177_OLOGIC_X0Y177_D1 = RIOB33_X105Y123_IOB_X1Y124_I;
  assign LIOI3_X0Y117_OLOGIC_X0Y118_T1 = 1'b1;
  assign RIOI3_X105Y161_OLOGIC_X1Y162_D1 = CLBLM_R_X7Y153_SLICE_X9Y153_C5Q;
  assign LIOI3_X0Y177_OLOGIC_X0Y177_T1 = 1'b1;
  assign LIOI3_X0Y117_OLOGIC_X0Y117_D1 = CLBLM_L_X10Y143_SLICE_X13Y143_C5Q;
  assign RIOI3_X105Y161_OLOGIC_X1Y162_T1 = 1'b1;
  assign CLBLM_L_X10Y146_SLICE_X12Y146_A6 = CLBLL_L_X4Y147_SLICE_X5Y147_CQ;
  assign LIOI3_X0Y117_OLOGIC_X0Y117_T1 = 1'b1;
  assign RIOI3_X105Y161_OLOGIC_X1Y161_D1 = CLBLM_L_X10Y154_SLICE_X12Y154_DO5;
  assign CLBLM_R_X5Y148_SLICE_X7Y148_A1 = CLBLM_R_X5Y147_SLICE_X7Y147_CQ;
  assign CLBLM_R_X5Y148_SLICE_X7Y148_A2 = CLBLL_L_X4Y142_SLICE_X5Y142_DQ;
  assign CLBLM_R_X5Y148_SLICE_X7Y148_A3 = CLBLM_R_X5Y148_SLICE_X7Y148_AQ;
  assign CLBLM_R_X5Y148_SLICE_X7Y148_A4 = CLBLL_L_X4Y147_SLICE_X5Y147_CQ;
  assign CLBLM_R_X5Y148_SLICE_X7Y148_A5 = CLBLM_R_X3Y148_SLICE_X3Y148_CQ;
  assign CLBLM_R_X5Y148_SLICE_X7Y148_A6 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X7Y154_SLICE_X8Y154_B6 = CLBLM_R_X7Y154_SLICE_X8Y154_CO6;
  assign CLBLM_R_X5Y148_SLICE_X7Y148_B1 = CLBLM_R_X11Y148_SLICE_X15Y148_AO6;
  assign CLBLM_R_X5Y148_SLICE_X7Y148_B2 = CLBLM_R_X5Y148_SLICE_X7Y148_BQ;
  assign CLBLM_R_X5Y148_SLICE_X7Y148_B3 = 1'b1;
  assign CLBLM_R_X5Y148_SLICE_X7Y148_B4 = CLBLM_R_X5Y148_SLICE_X7Y148_AQ;
  assign CLBLM_R_X5Y148_SLICE_X7Y148_B5 = CLBLM_R_X5Y146_SLICE_X7Y146_D5Q;
  assign CLBLM_R_X5Y148_SLICE_X7Y148_B6 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign RIOI3_X105Y161_OLOGIC_X1Y161_T1 = 1'b1;
  assign CLBLM_R_X5Y148_SLICE_X7Y148_C1 = CLBLL_L_X4Y143_SLICE_X4Y143_BQ;
  assign CLBLM_R_X5Y148_SLICE_X7Y148_C2 = CLBLM_R_X5Y148_SLICE_X7Y148_AQ;
  assign CLBLM_R_X5Y148_SLICE_X7Y148_C3 = CLBLL_L_X4Y150_SLICE_X4Y150_CQ;
  assign CLBLM_R_X5Y148_SLICE_X7Y148_C4 = CLBLM_R_X7Y143_SLICE_X8Y143_BQ;
  assign CLBLM_R_X5Y148_SLICE_X7Y148_C5 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X5Y148_SLICE_X7Y148_C6 = 1'b1;
  assign CLBLM_R_X5Y148_SLICE_X7Y148_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X5Y148_SLICE_X7Y148_D1 = CLBLM_R_X5Y154_SLICE_X6Y154_AQ;
  assign CLBLM_R_X5Y148_SLICE_X7Y148_D2 = CLBLM_R_X5Y154_SLICE_X6Y154_BQ;
  assign CLBLM_R_X5Y148_SLICE_X7Y148_D3 = 1'b1;
  assign CLBLM_R_X5Y148_SLICE_X7Y148_D4 = CLBLM_R_X7Y148_SLICE_X9Y148_A5Q;
  assign CLBLM_R_X5Y148_SLICE_X7Y148_D5 = 1'b1;
  assign CLBLM_R_X5Y148_SLICE_X7Y148_D6 = CLBLM_L_X8Y147_SLICE_X11Y147_CQ;
  assign CLBLM_R_X5Y148_SLICE_X6Y148_A1 = CLBLM_R_X7Y150_SLICE_X8Y150_AQ;
  assign CLBLM_R_X5Y148_SLICE_X6Y148_A2 = CLBLM_R_X7Y151_SLICE_X9Y151_BQ;
  assign CLBLM_R_X5Y148_SLICE_X6Y148_A3 = CLBLM_R_X7Y143_SLICE_X8Y143_DO6;
  assign CLBLM_R_X5Y148_SLICE_X6Y148_A4 = CLBLM_R_X5Y149_SLICE_X6Y149_AQ;
  assign CLBLM_R_X5Y148_SLICE_X6Y148_A5 = CLBLM_R_X5Y143_SLICE_X7Y143_AQ;
  assign CLBLM_R_X5Y148_SLICE_X6Y148_A6 = 1'b1;
  assign CLBLM_R_X7Y154_SLICE_X8Y154_C4 = CLBLM_R_X7Y155_SLICE_X8Y155_BO5;
  assign CLBLM_R_X5Y148_SLICE_X6Y148_AX = CLBLL_L_X4Y151_SLICE_X5Y151_CQ;
  assign CLBLM_R_X5Y148_SLICE_X6Y148_B1 = CLBLM_R_X5Y146_SLICE_X6Y146_DO6;
  assign CLBLM_R_X5Y148_SLICE_X6Y148_B2 = CLBLM_R_X5Y148_SLICE_X7Y148_DO6;
  assign CLBLM_R_X5Y148_SLICE_X6Y148_B3 = CLBLM_R_X7Y142_SLICE_X8Y142_DQ;
  assign CLBLM_R_X5Y148_SLICE_X6Y148_B4 = CLBLM_R_X7Y148_SLICE_X8Y148_DO6;
  assign CLBLM_R_X5Y148_SLICE_X6Y148_B5 = CLBLL_L_X4Y152_SLICE_X5Y152_AQ;
  assign CLBLM_R_X5Y148_SLICE_X6Y148_B6 = CLBLM_R_X5Y149_SLICE_X6Y149_DO6;
  assign CLBLM_R_X7Y154_SLICE_X8Y154_C5 = CLBLM_R_X7Y154_SLICE_X8Y154_DO6;
  assign CLBLM_R_X7Y154_SLICE_X8Y154_C6 = 1'b1;
  assign CLBLM_R_X5Y148_SLICE_X6Y148_BX = CLBLL_L_X4Y147_SLICE_X5Y147_CQ;
  assign CLBLM_R_X5Y148_SLICE_X6Y148_C1 = CLBLM_R_X7Y151_SLICE_X9Y151_BQ;
  assign CLBLM_R_X5Y148_SLICE_X6Y148_C2 = CLBLM_R_X5Y149_SLICE_X6Y149_AQ;
  assign CLBLM_R_X5Y148_SLICE_X6Y148_C3 = CLBLM_R_X5Y143_SLICE_X7Y143_AQ;
  assign CLBLM_R_X5Y148_SLICE_X6Y148_C4 = CLBLM_R_X7Y143_SLICE_X8Y143_DO6;
  assign CLBLM_R_X5Y148_SLICE_X6Y148_C5 = CLBLM_R_X7Y150_SLICE_X8Y150_AQ;
  assign CLBLM_R_X5Y148_SLICE_X6Y148_C6 = CLBLL_L_X4Y147_SLICE_X5Y147_AQ;
  assign CLBLM_R_X5Y148_SLICE_X6Y148_CE = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X5Y148_SLICE_X6Y148_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X5Y148_SLICE_X6Y148_CX = CLBLM_R_X5Y149_SLICE_X7Y149_C5Q;
  assign CLBLM_R_X5Y148_SLICE_X6Y148_D1 = 1'b1;
  assign CLBLM_R_X5Y148_SLICE_X6Y148_D2 = CLBLM_R_X7Y153_SLICE_X8Y153_CQ;
  assign CLBLM_R_X5Y148_SLICE_X6Y148_D3 = CLBLM_R_X3Y150_SLICE_X3Y150_A5Q;
  assign CLBLM_R_X5Y148_SLICE_X6Y148_D4 = CLBLM_R_X3Y144_SLICE_X3Y144_AQ;
  assign CLBLM_R_X5Y148_SLICE_X6Y148_D5 = CLBLM_L_X10Y148_SLICE_X13Y148_C5Q;
  assign CLBLM_R_X5Y148_SLICE_X6Y148_D6 = CLBLL_L_X4Y146_SLICE_X5Y146_AO5;
  assign RIOB33_X105Y161_IOB_X1Y162_O = CLBLM_R_X7Y153_SLICE_X9Y153_C5Q;
  assign RIOB33_X105Y161_IOB_X1Y161_O = CLBLM_L_X10Y154_SLICE_X12Y154_DO5;
  assign LIOB33_X0Y193_IOB_X0Y194_O = RIOB33_X105Y103_IOB_X1Y103_I;
  assign LIOB33_X0Y193_IOB_X0Y193_O = CLBLL_L_X2Y166_SLICE_X0Y166_AO6;
  assign CLBLM_L_X10Y155_SLICE_X13Y155_D4 = 1'b1;
  assign LIOI3_X0Y55_ILOGIC_X0Y56_D = LIOB33_X0Y55_IOB_X0Y56_I;
  assign LIOI3_X0Y55_ILOGIC_X0Y55_D = LIOB33_X0Y55_IOB_X0Y55_I;
  assign RIOI3_X105Y101_ILOGIC_X1Y102_D = RIOB33_X105Y101_IOB_X1Y102_I;
  assign RIOI3_X105Y101_ILOGIC_X1Y101_D = RIOB33_X105Y101_IOB_X1Y101_I;
  assign CLBLM_L_X12Y153_SLICE_X16Y153_C3 = 1'b1;
  assign CLBLM_R_X5Y149_SLICE_X7Y149_A1 = CLBLL_L_X4Y151_SLICE_X4Y151_B5Q;
  assign CLBLM_R_X5Y149_SLICE_X7Y149_A2 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X5Y149_SLICE_X7Y149_A3 = CLBLM_R_X7Y151_SLICE_X9Y151_A5Q;
  assign CLBLM_R_X5Y149_SLICE_X7Y149_A4 = CLBLM_L_X10Y149_SLICE_X12Y149_A5Q;
  assign CLBLM_R_X5Y149_SLICE_X7Y149_A5 = RIOB33_X105Y107_IOB_X1Y107_I;
  assign CLBLM_R_X5Y149_SLICE_X7Y149_A6 = CLBLM_R_X5Y149_SLICE_X7Y149_AQ;
  assign CLBLM_R_X5Y149_SLICE_X7Y149_B1 = CLBLM_R_X3Y144_SLICE_X3Y144_AQ;
  assign CLBLM_R_X5Y149_SLICE_X7Y149_B2 = CLBLM_R_X5Y149_SLICE_X7Y149_BQ;
  assign CLBLM_R_X5Y149_SLICE_X7Y149_B3 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X5Y149_SLICE_X7Y149_B4 = CLBLM_R_X7Y152_SLICE_X8Y152_D5Q;
  assign CLBLM_R_X5Y149_SLICE_X7Y149_B5 = CLBLM_R_X7Y142_SLICE_X8Y142_C5Q;
  assign CLBLM_R_X5Y149_SLICE_X7Y149_B6 = CLBLM_R_X5Y152_SLICE_X7Y152_B5Q;
  assign CLBLM_R_X5Y149_SLICE_X7Y149_C1 = CLBLM_L_X10Y153_SLICE_X13Y153_A5Q;
  assign CLBLM_R_X5Y149_SLICE_X7Y149_C2 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X5Y149_SLICE_X7Y149_C3 = CLBLM_R_X3Y151_SLICE_X3Y151_BQ;
  assign CLBLM_R_X5Y149_SLICE_X7Y149_C4 = CLBLM_R_X7Y149_SLICE_X9Y149_CQ;
  assign CLBLM_R_X5Y149_SLICE_X7Y149_C5 = CLBLM_R_X7Y144_SLICE_X9Y144_AQ;
  assign CLBLM_R_X5Y149_SLICE_X7Y149_C6 = 1'b1;
  assign CLBLM_R_X5Y149_SLICE_X7Y149_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X5Y149_SLICE_X7Y149_D1 = CLBLM_R_X5Y150_SLICE_X6Y150_A5Q;
  assign CLBLM_R_X5Y149_SLICE_X7Y149_D2 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X5Y149_SLICE_X7Y149_D3 = 1'b1;
  assign CLBLM_R_X5Y149_SLICE_X7Y149_D4 = CLBLL_L_X4Y149_SLICE_X4Y149_AQ;
  assign CLBLM_R_X5Y149_SLICE_X7Y149_D5 = CLBLM_R_X5Y149_SLICE_X7Y149_AQ;
  assign CLBLM_R_X5Y149_SLICE_X7Y149_D6 = 1'b1;
  assign CLBLM_R_X5Y149_SLICE_X6Y149_A1 = CLBLM_L_X8Y149_SLICE_X11Y149_AQ;
  assign CLBLM_R_X5Y149_SLICE_X6Y149_A2 = CLBLM_R_X7Y151_SLICE_X9Y151_C5Q;
  assign CLBLM_R_X5Y149_SLICE_X6Y149_A3 = CLBLM_R_X5Y149_SLICE_X6Y149_AQ;
  assign CLBLM_R_X5Y149_SLICE_X6Y149_A4 = CLBLL_L_X4Y145_SLICE_X5Y145_C5Q;
  assign CLBLM_R_X5Y149_SLICE_X6Y149_A5 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X5Y149_SLICE_X6Y149_A6 = CLBLM_R_X5Y148_SLICE_X6Y148_AO5;
  assign CLBLM_R_X5Y149_SLICE_X6Y149_B1 = CLBLM_L_X10Y149_SLICE_X13Y149_AQ;
  assign CLBLM_R_X5Y149_SLICE_X6Y149_B2 = CLBLL_L_X4Y148_SLICE_X5Y148_BQ;
  assign CLBLM_R_X5Y149_SLICE_X6Y149_B3 = 1'b1;
  assign CLBLM_R_X5Y149_SLICE_X6Y149_B4 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X5Y149_SLICE_X6Y149_B5 = CLBLM_R_X5Y148_SLICE_X6Y148_AQ;
  assign CLBLM_R_X5Y149_SLICE_X6Y149_B6 = 1'b1;
  assign CLBLM_R_X5Y149_SLICE_X6Y149_C1 = CLBLL_L_X4Y148_SLICE_X4Y148_C5Q;
  assign CLBLM_R_X5Y149_SLICE_X6Y149_C2 = CLBLM_L_X8Y151_SLICE_X10Y151_AQ;
  assign CLBLM_R_X5Y149_SLICE_X6Y149_C3 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X5Y149_SLICE_X6Y149_C4 = CLBLL_L_X4Y143_SLICE_X5Y143_DQ;
  assign CLBLM_R_X5Y149_SLICE_X6Y149_C5 = CLBLM_L_X8Y145_SLICE_X11Y145_DQ;
  assign CLBLM_R_X5Y149_SLICE_X6Y149_C6 = 1'b1;
  assign CLBLM_R_X5Y149_SLICE_X6Y149_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X5Y149_SLICE_X6Y149_D1 = CLBLM_R_X3Y149_SLICE_X2Y149_AQ;
  assign CLBLM_R_X5Y149_SLICE_X6Y149_D2 = CLBLL_L_X4Y153_SLICE_X5Y153_AQ;
  assign CLBLM_R_X5Y149_SLICE_X6Y149_D3 = 1'b1;
  assign CLBLM_R_X5Y149_SLICE_X6Y149_D4 = CLBLM_L_X8Y152_SLICE_X11Y152_D5Q;
  assign CLBLM_R_X5Y149_SLICE_X6Y149_D5 = CLBLM_L_X8Y144_SLICE_X11Y144_BQ;
  assign CLBLM_R_X5Y149_SLICE_X6Y149_D6 = CLBLM_R_X3Y152_SLICE_X3Y152_AQ;
  assign RIOB33_X105Y163_IOB_X1Y163_O = CLBLM_R_X7Y151_SLICE_X9Y151_D5Q;
  assign RIOB33_X105Y163_IOB_X1Y164_O = CLBLM_L_X10Y153_SLICE_X12Y153_AQ;
  assign LIOB33_X0Y195_IOB_X0Y196_O = CLBLM_R_X3Y148_SLICE_X3Y148_DO5;
  assign LIOB33_X0Y195_IOB_X0Y195_O = CLBLM_R_X3Y151_SLICE_X2Y151_AO5;
  assign LIOI3_X0Y111_OLOGIC_X0Y112_D1 = CLBLL_L_X4Y146_SLICE_X4Y146_C5Q;
  assign LIOI3_X0Y111_OLOGIC_X0Y112_T1 = 1'b1;
  assign CLBLM_L_X10Y155_SLICE_X12Y155_A6 = CLBLM_R_X5Y146_SLICE_X7Y146_CQ;
  assign LIOI3_X0Y111_OLOGIC_X0Y111_D1 = CLBLM_R_X3Y145_SLICE_X2Y145_B5Q;
  assign CLBLM_R_X5Y150_SLICE_X7Y150_A1 = CLBLL_L_X4Y150_SLICE_X4Y150_B5Q;
  assign CLBLM_R_X5Y150_SLICE_X7Y150_A2 = CLBLM_R_X5Y149_SLICE_X7Y149_DQ;
  assign CLBLM_R_X5Y150_SLICE_X7Y150_A3 = CLBLM_R_X5Y150_SLICE_X7Y150_AQ;
  assign CLBLM_R_X5Y150_SLICE_X7Y150_A4 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X5Y150_SLICE_X7Y150_A5 = CLBLM_L_X10Y153_SLICE_X13Y153_A5Q;
  assign CLBLM_R_X5Y150_SLICE_X7Y150_A6 = 1'b1;
  assign CLBLM_R_X5Y150_SLICE_X7Y150_B1 = CLBLL_L_X4Y152_SLICE_X5Y152_A5Q;
  assign CLBLM_R_X5Y150_SLICE_X7Y150_B2 = CLBLM_R_X5Y151_SLICE_X7Y151_DO6;
  assign CLBLM_R_X5Y150_SLICE_X7Y150_B3 = CLBLM_R_X5Y147_SLICE_X6Y147_DO6;
  assign CLBLM_R_X5Y150_SLICE_X7Y150_B4 = CLBLM_R_X5Y150_SLICE_X7Y150_DO6;
  assign CLBLM_R_X5Y150_SLICE_X7Y150_B5 = CLBLM_R_X5Y146_SLICE_X6Y146_BQ;
  assign CLBLM_R_X5Y150_SLICE_X7Y150_B6 = CLBLM_R_X5Y150_SLICE_X7Y150_CO6;
  assign CLBLM_R_X5Y150_SLICE_X7Y150_C1 = CLBLM_R_X5Y154_SLICE_X6Y154_AQ;
  assign CLBLM_R_X5Y150_SLICE_X7Y150_C2 = CLBLM_R_X5Y154_SLICE_X6Y154_BQ;
  assign CLBLM_R_X5Y150_SLICE_X7Y150_C3 = CLBLM_R_X7Y151_SLICE_X8Y151_CQ;
  assign CLBLM_R_X5Y150_SLICE_X7Y150_C4 = CLBLL_L_X4Y153_SLICE_X5Y153_AQ;
  assign CLBLM_R_X5Y150_SLICE_X7Y150_C5 = CLBLM_R_X7Y147_SLICE_X9Y147_D5Q;
  assign CLBLM_R_X5Y150_SLICE_X7Y150_C6 = CLBLM_R_X5Y149_SLICE_X6Y149_BQ;
  assign CLBLM_R_X5Y150_SLICE_X7Y150_CLK = CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O;
  assign CLBLM_L_X12Y153_SLICE_X16Y153_D4 = 1'b1;
  assign CLBLM_R_X5Y150_SLICE_X7Y150_D1 = 1'b1;
  assign CLBLM_R_X5Y150_SLICE_X7Y150_D2 = CLBLM_R_X7Y153_SLICE_X9Y153_AQ;
  assign CLBLM_R_X5Y150_SLICE_X7Y150_D3 = CLBLM_R_X3Y149_SLICE_X3Y149_AQ;
  assign CLBLM_R_X5Y150_SLICE_X7Y150_D4 = CLBLM_R_X5Y149_SLICE_X7Y149_CQ;
  assign CLBLM_R_X5Y150_SLICE_X7Y150_D5 = CLBLM_R_X7Y152_SLICE_X8Y152_DQ;
  assign CLBLM_R_X5Y150_SLICE_X7Y150_D6 = 1'b1;
  assign CLBLM_R_X5Y150_SLICE_X6Y150_A1 = CLBLM_L_X8Y153_SLICE_X10Y153_DQ;
  assign CLBLM_R_X5Y150_SLICE_X6Y150_A2 = CLBLM_R_X5Y150_SLICE_X6Y150_BQ;
  assign CLBLM_R_X5Y150_SLICE_X6Y150_A3 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X5Y150_SLICE_X6Y150_A4 = CLBLL_L_X2Y145_SLICE_X1Y145_CQ;
  assign CLBLM_R_X5Y150_SLICE_X6Y150_A5 = CLBLM_R_X5Y152_SLICE_X6Y152_DQ;
  assign CLBLM_R_X5Y150_SLICE_X6Y150_A6 = 1'b1;
  assign LIOI3_X0Y179_OLOGIC_X0Y180_D1 = RIOB33_X105Y127_IOB_X1Y127_I;
  assign RIOB33_X105Y165_IOB_X1Y165_O = CLBLM_L_X12Y152_SLICE_X16Y152_AO6;
  assign CLBLM_R_X5Y150_SLICE_X6Y150_B1 = CLBLM_R_X5Y150_SLICE_X6Y150_CQ;
  assign CLBLM_R_X5Y150_SLICE_X6Y150_B2 = CLBLM_L_X8Y153_SLICE_X10Y153_BQ;
  assign CLBLM_R_X5Y150_SLICE_X6Y150_B3 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X5Y150_SLICE_X6Y150_B4 = CLBLL_L_X4Y143_SLICE_X4Y143_AQ;
  assign CLBLM_R_X5Y150_SLICE_X6Y150_B5 = CLBLM_R_X3Y142_SLICE_X3Y142_AQ;
  assign CLBLM_R_X5Y150_SLICE_X6Y150_B6 = 1'b1;
  assign RIOB33_X105Y165_IOB_X1Y166_O = CLBLM_L_X8Y153_SLICE_X10Y153_A5Q;
  assign LIOI3_X0Y179_OLOGIC_X0Y180_T1 = 1'b1;
  assign CLBLM_R_X5Y150_SLICE_X6Y150_C1 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X5Y150_SLICE_X6Y150_C2 = CLBLM_R_X5Y144_SLICE_X6Y144_CQ;
  assign CLBLM_R_X5Y150_SLICE_X6Y150_C3 = CLBLM_L_X10Y144_SLICE_X13Y144_A5Q;
  assign CLBLM_R_X5Y150_SLICE_X6Y150_C4 = CLBLL_L_X4Y150_SLICE_X4Y150_DO6;
  assign CLBLM_R_X5Y150_SLICE_X6Y150_C5 = CLBLM_R_X5Y152_SLICE_X6Y152_B5Q;
  assign CLBLM_R_X5Y150_SLICE_X6Y150_C6 = 1'b1;
  assign LIOI3_X0Y121_OLOGIC_X0Y122_D1 = CLBLL_L_X4Y144_SLICE_X5Y144_CQ;
  assign CLBLM_R_X5Y150_SLICE_X6Y150_CLK = CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O;
  assign LIOI3_X0Y179_OLOGIC_X0Y179_D1 = RIOB33_X105Y125_IOB_X1Y126_I;
  assign LIOI3_X0Y121_OLOGIC_X0Y122_T1 = 1'b1;
  assign CLBLM_R_X5Y150_SLICE_X6Y150_D1 = CLBLM_R_X5Y150_SLICE_X6Y150_BQ;
  assign CLBLM_R_X5Y150_SLICE_X6Y150_D2 = CLBLM_R_X5Y151_SLICE_X7Y151_B5Q;
  assign CLBLM_R_X5Y150_SLICE_X6Y150_D3 = CLBLM_R_X5Y151_SLICE_X6Y151_DO6;
  assign CLBLM_R_X5Y150_SLICE_X6Y150_D4 = CLBLM_R_X5Y150_SLICE_X6Y150_A5Q;
  assign CLBLM_R_X5Y150_SLICE_X6Y150_D5 = CLBLM_R_X5Y145_SLICE_X6Y145_BQ;
  assign CLBLM_R_X5Y150_SLICE_X6Y150_D6 = CLBLM_L_X8Y146_SLICE_X11Y146_DQ;
  assign LIOI3_X0Y179_OLOGIC_X0Y179_T1 = 1'b1;
  assign RIOI3_X105Y165_OLOGIC_X1Y166_D1 = CLBLM_L_X8Y153_SLICE_X10Y153_A5Q;
  assign LIOI3_X0Y121_OLOGIC_X0Y121_D1 = CLBLM_L_X8Y147_SLICE_X10Y147_C5Q;
  assign RIOI3_X105Y165_OLOGIC_X1Y166_T1 = 1'b1;
  assign LIOB33_X0Y197_IOB_X0Y198_O = 1'b1;
  assign LIOB33_X0Y197_IOB_X0Y197_O = CLBLL_L_X4Y153_SLICE_X4Y153_CO5;
  assign LIOI3_X0Y121_OLOGIC_X0Y121_T1 = 1'b1;
  assign RIOI3_X105Y165_OLOGIC_X1Y165_D1 = CLBLM_L_X12Y152_SLICE_X16Y152_AO6;
  assign RIOI3_X105Y165_OLOGIC_X1Y165_T1 = 1'b1;
  assign LIOI3_X0Y173_OLOGIC_X0Y174_D1 = RIOB33_X105Y121_IOB_X1Y122_I;
  assign LIOI3_X0Y59_ILOGIC_X0Y60_D = LIOB33_X0Y59_IOB_X0Y60_I;
  assign LIOI3_X0Y59_ILOGIC_X0Y59_D = LIOB33_X0Y59_IOB_X0Y59_I;
  assign RIOI3_X105Y103_ILOGIC_X1Y104_D = RIOB33_X105Y103_IOB_X1Y104_I;
  assign RIOI3_X105Y103_ILOGIC_X1Y103_D = RIOB33_X105Y103_IOB_X1Y103_I;
  assign CLBLM_R_X5Y151_SLICE_X7Y151_A1 = CLBLM_L_X8Y149_SLICE_X11Y149_AQ;
  assign CLBLM_R_X5Y151_SLICE_X7Y151_A2 = CLBLM_R_X7Y145_SLICE_X8Y145_BQ;
  assign CLBLM_R_X5Y151_SLICE_X7Y151_A3 = CLBLM_R_X5Y151_SLICE_X7Y151_AQ;
  assign CLBLM_R_X5Y151_SLICE_X7Y151_A4 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X5Y151_SLICE_X7Y151_A5 = CLBLM_R_X5Y148_SLICE_X6Y148_CO6;
  assign CLBLM_R_X5Y151_SLICE_X7Y151_A6 = CLBLL_L_X4Y151_SLICE_X5Y151_D5Q;
  assign CLBLM_R_X5Y151_SLICE_X7Y151_B1 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X5Y151_SLICE_X7Y151_B2 = CLBLL_L_X4Y151_SLICE_X5Y151_CQ;
  assign CLBLM_R_X5Y151_SLICE_X7Y151_B3 = CLBLL_L_X4Y151_SLICE_X4Y151_A5Q;
  assign CLBLM_R_X5Y151_SLICE_X7Y151_B4 = CLBLM_R_X7Y144_SLICE_X8Y144_B5Q;
  assign CLBLM_R_X5Y151_SLICE_X7Y151_B5 = CLBLM_L_X10Y154_SLICE_X12Y154_AQ;
  assign CLBLM_R_X5Y151_SLICE_X7Y151_B6 = 1'b1;
  assign CLBLM_R_X5Y151_SLICE_X7Y151_C1 = CLBLM_R_X5Y148_SLICE_X7Y148_CQ;
  assign CLBLM_R_X5Y151_SLICE_X7Y151_C2 = CLBLM_R_X5Y144_SLICE_X6Y144_DQ;
  assign CLBLM_R_X5Y151_SLICE_X7Y151_C3 = CLBLL_L_X4Y151_SLICE_X5Y151_B5Q;
  assign CLBLM_R_X5Y151_SLICE_X7Y151_C4 = 1'b1;
  assign CLBLM_R_X5Y151_SLICE_X7Y151_C5 = CLBLM_R_X7Y147_SLICE_X9Y147_AQ;
  assign CLBLM_R_X5Y151_SLICE_X7Y151_C6 = 1'b1;
  assign LIOI3_X0Y173_OLOGIC_X0Y174_T1 = 1'b1;
  assign RIOB33_X105Y167_IOB_X1Y167_O = CLBLM_R_X7Y153_SLICE_X9Y153_DQ;
  assign CLBLM_R_X5Y151_SLICE_X7Y151_CLK = CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O;
  assign RIOB33_X105Y167_IOB_X1Y168_O = CLBLM_R_X5Y154_SLICE_X7Y154_AQ;
  assign CLBLM_R_X5Y151_SLICE_X7Y151_D1 = 1'b1;
  assign CLBLM_R_X5Y151_SLICE_X7Y151_D2 = CLBLM_R_X11Y151_SLICE_X15Y151_A5Q;
  assign CLBLM_R_X5Y151_SLICE_X7Y151_D3 = CLBLM_R_X7Y151_SLICE_X8Y151_DQ;
  assign CLBLM_R_X5Y151_SLICE_X7Y151_D4 = 1'b1;
  assign CLBLM_R_X5Y151_SLICE_X7Y151_D5 = CLBLL_L_X4Y152_SLICE_X5Y152_AQ;
  assign CLBLM_R_X5Y151_SLICE_X7Y151_D6 = CLBLM_R_X3Y152_SLICE_X3Y152_AQ;
  assign CLBLM_R_X5Y151_SLICE_X6Y151_A1 = CLBLM_R_X13Y149_SLICE_X18Y149_AO6;
  assign CLBLM_R_X5Y151_SLICE_X6Y151_A2 = 1'b1;
  assign CLBLM_R_X5Y151_SLICE_X6Y151_A3 = CLBLL_L_X4Y151_SLICE_X5Y151_D5Q;
  assign CLBLM_R_X5Y151_SLICE_X6Y151_A4 = CLBLM_R_X5Y151_SLICE_X6Y151_AQ;
  assign CLBLM_R_X5Y151_SLICE_X6Y151_A5 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X5Y151_SLICE_X6Y151_A6 = CLBLL_L_X4Y145_SLICE_X5Y145_AQ;
  assign CLBLM_R_X5Y151_SLICE_X6Y151_B1 = CLBLM_R_X13Y149_SLICE_X18Y149_AO6;
  assign CLBLM_R_X5Y151_SLICE_X6Y151_B2 = CLBLM_R_X5Y151_SLICE_X6Y151_BQ;
  assign CLBLM_R_X5Y151_SLICE_X6Y151_B3 = CLBLM_R_X7Y147_SLICE_X9Y147_BQ;
  assign CLBLM_R_X5Y151_SLICE_X6Y151_B4 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X5Y151_SLICE_X6Y151_B5 = CLBLL_L_X2Y146_SLICE_X1Y146_B5Q;
  assign CLBLM_R_X5Y151_SLICE_X6Y151_B6 = 1'b1;
  assign CLBLM_R_X5Y151_SLICE_X6Y151_C1 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X5Y151_SLICE_X6Y151_C2 = CLBLM_R_X5Y146_SLICE_X6Y146_B5Q;
  assign CLBLM_R_X5Y151_SLICE_X6Y151_C3 = CLBLL_L_X4Y153_SLICE_X4Y153_B5Q;
  assign CLBLM_R_X5Y151_SLICE_X6Y151_C4 = CLBLM_R_X3Y151_SLICE_X3Y151_AQ;
  assign CLBLM_R_X5Y151_SLICE_X6Y151_C5 = CLBLM_L_X10Y152_SLICE_X12Y152_CQ;
  assign CLBLM_R_X5Y151_SLICE_X6Y151_C6 = 1'b1;
  assign CLBLM_R_X5Y151_SLICE_X6Y151_CLK = CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O;
  assign LIOI3_X0Y173_OLOGIC_X0Y173_D1 = RIOB33_X105Y121_IOB_X1Y121_I;
  assign CLBLM_R_X5Y151_SLICE_X6Y151_D1 = CLBLM_R_X5Y149_SLICE_X7Y149_C5Q;
  assign CLBLM_R_X5Y151_SLICE_X6Y151_D2 = CLBLM_R_X5Y151_SLICE_X6Y151_CQ;
  assign CLBLM_R_X5Y151_SLICE_X6Y151_D3 = CLBLL_L_X4Y144_SLICE_X4Y144_B5Q;
  assign CLBLM_R_X5Y151_SLICE_X6Y151_D4 = 1'b1;
  assign CLBLM_R_X5Y151_SLICE_X6Y151_D5 = 1'b1;
  assign CLBLM_R_X5Y151_SLICE_X6Y151_D6 = CLBLM_R_X7Y152_SLICE_X8Y152_BQ;
  assign LIOI3_X0Y173_OLOGIC_X0Y173_T1 = 1'b1;
  assign CLBLM_R_X11Y153_SLICE_X15Y153_C4 = CLBLM_R_X5Y147_SLICE_X6Y147_AQ;
  assign CLBLM_R_X11Y153_SLICE_X15Y153_C5 = CLBLM_L_X10Y153_SLICE_X13Y153_CQ;
  assign CLBLM_R_X11Y153_SLICE_X15Y153_C6 = CLBLM_R_X11Y153_SLICE_X15Y153_AQ;
  assign RIOB33_X105Y169_IOB_X1Y170_O = CLBLM_R_X3Y152_SLICE_X3Y152_BQ;
  assign RIOB33_X105Y169_IOB_X1Y169_O = CLBLM_R_X3Y152_SLICE_X3Y152_CQ;
  assign CLBLM_R_X5Y152_SLICE_X7Y152_A1 = CLBLL_L_X4Y146_SLICE_X4Y146_C5Q;
  assign CLBLM_R_X5Y152_SLICE_X7Y152_A2 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X5Y152_SLICE_X7Y152_A3 = CLBLM_R_X7Y151_SLICE_X8Y151_D5Q;
  assign CLBLM_R_X5Y152_SLICE_X7Y152_A4 = CLBLM_R_X5Y149_SLICE_X6Y149_CQ;
  assign CLBLM_R_X5Y152_SLICE_X7Y152_A5 = CLBLM_R_X7Y146_SLICE_X8Y146_A5Q;
  assign CLBLM_R_X5Y152_SLICE_X7Y152_A6 = 1'b1;
  assign CLBLM_R_X5Y152_SLICE_X7Y152_B1 = CLBLM_R_X5Y151_SLICE_X6Y151_CQ;
  assign CLBLM_R_X5Y152_SLICE_X7Y152_B2 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X5Y152_SLICE_X7Y152_B3 = 1'b1;
  assign CLBLM_R_X5Y152_SLICE_X7Y152_B4 = CLBLL_L_X4Y145_SLICE_X5Y145_BQ;
  assign CLBLM_R_X5Y152_SLICE_X7Y152_B5 = CLBLM_R_X7Y155_SLICE_X8Y155_A5Q;
  assign CLBLM_R_X5Y152_SLICE_X7Y152_B6 = 1'b1;
  assign CLBLM_R_X11Y153_SLICE_X15Y153_D2 = CLBLM_R_X11Y153_SLICE_X14Y153_A5Q;
  assign CLBLM_R_X3Y142_SLICE_X3Y142_A1 = CLBLM_R_X7Y142_SLICE_X9Y142_BQ;
  assign CLBLM_R_X3Y142_SLICE_X3Y142_A2 = 1'b1;
  assign CLBLM_R_X3Y142_SLICE_X3Y142_A3 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X3Y142_SLICE_X3Y142_A4 = CLBLM_R_X3Y142_SLICE_X3Y142_AQ;
  assign CLBLM_R_X3Y142_SLICE_X3Y142_A5 = CLBLM_R_X5Y147_SLICE_X6Y147_AQ;
  assign CLBLM_R_X3Y142_SLICE_X3Y142_A6 = CLBLM_L_X10Y144_SLICE_X12Y144_AO6;
  assign CLBLM_R_X5Y152_SLICE_X7Y152_C1 = CLBLM_L_X8Y152_SLICE_X10Y152_BQ;
  assign CLBLM_R_X5Y152_SLICE_X7Y152_C2 = CLBLM_R_X5Y151_SLICE_X7Y151_BQ;
  assign CLBLM_R_X5Y152_SLICE_X7Y152_C3 = CLBLM_R_X5Y152_SLICE_X6Y152_CQ;
  assign CLBLM_R_X3Y142_SLICE_X3Y142_B1 = CLBLM_R_X7Y146_SLICE_X8Y146_DQ;
  assign CLBLM_R_X3Y142_SLICE_X3Y142_B2 = 1'b1;
  assign CLBLM_R_X3Y142_SLICE_X3Y142_B3 = CLBLM_R_X3Y147_SLICE_X3Y147_C5Q;
  assign CLBLM_R_X3Y142_SLICE_X3Y142_B4 = CLBLL_L_X4Y142_SLICE_X5Y142_CQ;
  assign CLBLM_R_X3Y142_SLICE_X3Y142_B5 = CLBLM_R_X5Y141_SLICE_X6Y141_BQ;
  assign CLBLM_R_X3Y142_SLICE_X3Y142_B6 = CLBLM_R_X3Y142_SLICE_X3Y142_CO6;
  assign CLBLM_R_X5Y152_SLICE_X7Y152_CLK = CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O;
  assign CLBLM_R_X5Y152_SLICE_X7Y152_D5 = CLBLM_R_X5Y150_SLICE_X6Y150_DO6;
  assign CLBLM_R_X5Y152_SLICE_X7Y152_D6 = 1'b1;
  assign CLBLM_R_X3Y142_SLICE_X3Y142_C1 = 1'b1;
  assign CLBLM_R_X3Y142_SLICE_X3Y142_C2 = CLBLM_R_X5Y145_SLICE_X7Y145_AQ;
  assign CLBLM_R_X3Y142_SLICE_X3Y142_C3 = CLBLL_L_X4Y143_SLICE_X4Y143_DQ;
  assign CLBLM_R_X3Y142_SLICE_X3Y142_C4 = 1'b1;
  assign CLBLM_R_X3Y142_SLICE_X3Y142_C5 = CLBLM_R_X3Y145_SLICE_X2Y145_B5Q;
  assign CLBLM_R_X3Y142_SLICE_X3Y142_C6 = CLBLL_L_X4Y146_SLICE_X4Y146_C5Q;
  assign CLBLM_R_X5Y152_SLICE_X7Y152_D4 = CLBLM_R_X7Y153_SLICE_X9Y153_DQ;
  assign CLBLM_R_X5Y152_SLICE_X6Y152_A1 = CLBLM_L_X8Y153_SLICE_X11Y153_AQ;
  assign CLBLM_R_X5Y152_SLICE_X6Y152_A2 = CLBLM_L_X10Y145_SLICE_X12Y145_AQ;
  assign CLBLM_R_X5Y152_SLICE_X6Y152_A3 = CLBLM_R_X5Y152_SLICE_X6Y152_AQ;
  assign CLBLM_R_X5Y152_SLICE_X6Y152_A4 = CLBLM_R_X5Y142_SLICE_X7Y142_BQ;
  assign CLBLM_R_X3Y142_SLICE_X3Y142_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X5Y152_SLICE_X6Y152_A5 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X3Y142_SLICE_X3Y142_D1 = 1'b1;
  assign CLBLM_R_X3Y142_SLICE_X3Y142_D2 = 1'b1;
  assign CLBLM_R_X3Y142_SLICE_X3Y142_D3 = 1'b1;
  assign CLBLM_R_X3Y142_SLICE_X3Y142_D4 = 1'b1;
  assign CLBLM_R_X3Y142_SLICE_X3Y142_D5 = 1'b1;
  assign CLBLM_R_X3Y142_SLICE_X3Y142_D6 = 1'b1;
  assign CLBLM_R_X5Y152_SLICE_X6Y152_A6 = CLBLM_R_X5Y152_SLICE_X7Y152_CQ;
  assign CLBLM_R_X5Y152_SLICE_X6Y152_B1 = CLBLL_L_X4Y152_SLICE_X5Y152_A5Q;
  assign CLBLM_R_X5Y152_SLICE_X6Y152_B2 = CLBLL_L_X4Y144_SLICE_X4Y144_C5Q;
  assign CLBLM_R_X5Y152_SLICE_X6Y152_B3 = CLBLM_R_X7Y153_SLICE_X8Y153_DQ;
  assign CLBLM_R_X5Y152_SLICE_X6Y152_B4 = CLBLM_R_X5Y144_SLICE_X7Y144_CQ;
  assign CLBLM_R_X3Y142_SLICE_X2Y142_A1 = CLBLM_R_X3Y142_SLICE_X2Y142_BO5;
  assign CLBLM_R_X5Y152_SLICE_X6Y152_C1 = CLBLM_R_X7Y147_SLICE_X9Y147_BQ;
  assign CLBLM_R_X5Y152_SLICE_X6Y152_C2 = CLBLM_R_X5Y152_SLICE_X6Y152_CQ;
  assign CLBLM_R_X5Y152_SLICE_X6Y152_C3 = 1'b1;
  assign CLBLM_R_X5Y152_SLICE_X6Y152_C4 = CLBLM_R_X3Y145_SLICE_X2Y145_CQ;
  assign CLBLM_R_X5Y152_SLICE_X6Y152_C5 = CLBLL_L_X4Y148_SLICE_X4Y148_DO6;
  assign CLBLM_R_X5Y152_SLICE_X6Y152_C6 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X3Y142_SLICE_X2Y142_A2 = CLBLM_R_X3Y143_SLICE_X3Y143_AQ;
  assign CLBLM_R_X3Y142_SLICE_X2Y142_A3 = CLBLM_R_X3Y142_SLICE_X2Y142_AQ;
  assign CLBLM_R_X3Y142_SLICE_X2Y142_A4 = CLBLM_R_X3Y142_SLICE_X2Y142_BO6;
  assign CLBLM_R_X5Y152_SLICE_X6Y152_CLK = CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O;
  assign CLBLM_R_X3Y142_SLICE_X2Y142_A5 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X3Y142_SLICE_X2Y142_B3 = CLBLM_R_X3Y142_SLICE_X2Y142_AQ;
  assign CLBLM_R_X3Y142_SLICE_X2Y142_A6 = CLBLM_L_X10Y144_SLICE_X12Y144_AO6;
  assign CLBLM_R_X3Y142_SLICE_X2Y142_B5 = CLBLM_R_X5Y147_SLICE_X6Y147_AQ;
  assign CLBLM_R_X3Y142_SLICE_X2Y142_B6 = 1'b1;
  assign CLBLM_R_X5Y152_SLICE_X6Y152_D1 = CLBLM_R_X5Y152_SLICE_X7Y152_AQ;
  assign CLBLM_R_X5Y152_SLICE_X6Y152_D2 = CLBLM_R_X5Y152_SLICE_X6Y152_CQ;
  assign CLBLM_R_X5Y152_SLICE_X6Y152_D3 = CLBLM_R_X5Y152_SLICE_X6Y152_DQ;
  assign CLBLM_R_X5Y152_SLICE_X6Y152_D4 = CLBLM_R_X3Y145_SLICE_X2Y145_CQ;
  assign CLBLM_R_X5Y152_SLICE_X6Y152_D5 = CLBLL_L_X4Y148_SLICE_X4Y148_DO6;
  assign CLBLM_R_X5Y152_SLICE_X6Y152_D6 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X3Y142_SLICE_X2Y142_C2 = 1'b1;
  assign CLBLM_R_X3Y142_SLICE_X2Y142_C3 = 1'b1;
  assign CLBLM_R_X3Y142_SLICE_X2Y142_C4 = 1'b1;
  assign CLBLM_R_X3Y142_SLICE_X2Y142_C1 = 1'b1;
  assign CLBLM_R_X3Y142_SLICE_X2Y142_C5 = 1'b1;
  assign CLBLM_R_X3Y142_SLICE_X2Y142_C6 = 1'b1;
  assign CLBLM_R_X3Y142_SLICE_X2Y142_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X3Y142_SLICE_X2Y142_D1 = 1'b1;
  assign CLBLM_R_X3Y142_SLICE_X2Y142_D2 = 1'b1;
  assign CLBLM_R_X3Y142_SLICE_X2Y142_D3 = 1'b1;
  assign CLBLM_R_X3Y142_SLICE_X2Y142_D4 = 1'b1;
  assign CLBLM_R_X3Y142_SLICE_X2Y142_D5 = 1'b1;
  assign CLBLM_R_X3Y142_SLICE_X2Y142_D6 = 1'b1;
  assign CLBLM_L_X10Y147_SLICE_X13Y147_B3 = CLBLM_R_X7Y151_SLICE_X8Y151_D5Q;
  assign CLBLM_L_X10Y147_SLICE_X13Y147_B4 = CLBLL_L_X4Y147_SLICE_X4Y147_CQ;
  assign CLBLM_R_X7Y155_SLICE_X9Y155_C4 = 1'b1;
  assign CLBLM_R_X7Y155_SLICE_X9Y155_C5 = 1'b1;
  assign CLBLM_R_X7Y155_SLICE_X9Y155_C6 = 1'b1;
  assign CLBLM_R_X11Y153_SLICE_X14Y153_B3 = CLBLM_R_X11Y153_SLICE_X14Y153_AQ;
  assign CLBLM_R_X11Y153_SLICE_X14Y153_B4 = CLBLM_L_X10Y152_SLICE_X12Y152_AQ;
  assign CLBLM_R_X11Y153_SLICE_X14Y153_B5 = CLBLM_L_X10Y152_SLICE_X13Y152_AQ;
  assign CLBLM_R_X11Y153_SLICE_X14Y153_B6 = CLBLM_R_X11Y153_SLICE_X15Y153_BO5;
  assign LIOI3_X0Y183_OLOGIC_X0Y184_D1 = RIOB33_X105Y131_IOB_X1Y132_I;
  assign LIOI3_X0Y183_OLOGIC_X0Y184_T1 = 1'b1;
  assign LIOI3_X0Y123_OLOGIC_X0Y124_D1 = CLBLL_L_X4Y151_SLICE_X4Y151_CQ;
  assign CLBLM_R_X11Y153_SLICE_X14Y153_C2 = CLBLM_R_X11Y153_SLICE_X14Y153_AQ;
  assign LIOI3_X0Y183_OLOGIC_X0Y183_D1 = RIOB33_X105Y129_IOB_X1Y130_I;
  assign LIOI3_X0Y123_OLOGIC_X0Y124_T1 = 1'b1;
  assign CLBLM_R_X11Y153_SLICE_X14Y153_C3 = CLBLM_R_X5Y147_SLICE_X6Y147_AQ;
  assign RIOI3_X105Y167_OLOGIC_X1Y168_D1 = CLBLM_R_X5Y154_SLICE_X7Y154_AQ;
  assign CLBLM_R_X11Y153_SLICE_X14Y153_C4 = CLBLM_L_X10Y152_SLICE_X12Y152_AQ;
  assign LIOI3_X0Y183_OLOGIC_X0Y183_T1 = 1'b1;
  assign CLBLM_R_X7Y155_SLICE_X9Y155_D5 = 1'b1;
  assign CLBLM_R_X11Y153_SLICE_X14Y153_C5 = CLBLM_L_X10Y153_SLICE_X13Y153_CQ;
  assign LIOI3_X0Y123_OLOGIC_X0Y123_D1 = CLBLL_L_X2Y146_SLICE_X0Y146_CQ;
  assign CLBLM_R_X7Y155_SLICE_X9Y155_D6 = 1'b1;
  assign CLBLM_R_X11Y153_SLICE_X14Y153_C6 = CLBLM_L_X8Y152_SLICE_X10Y152_CQ;
  assign RIOI3_X105Y167_OLOGIC_X1Y168_T1 = 1'b1;
  assign LIOI3_X0Y123_OLOGIC_X0Y123_T1 = 1'b1;
  assign RIOI3_X105Y167_OLOGIC_X1Y167_D1 = CLBLM_R_X7Y153_SLICE_X9Y153_DQ;
  assign CLBLM_R_X11Y153_SLICE_X14Y153_CLK = CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O;
  assign LIOI3_TBYTESRC_X0Y107_OLOGIC_X0Y108_D1 = CLBLL_L_X4Y143_SLICE_X4Y143_DQ;
  assign RIOI3_X105Y167_OLOGIC_X1Y167_T1 = 1'b1;
  assign LIOI3_TBYTESRC_X0Y107_OLOGIC_X0Y108_T1 = 1'b1;
  assign LIOI3_TBYTESRC_X0Y107_OLOGIC_X0Y107_D1 = CLBLM_R_X7Y146_SLICE_X8Y146_DQ;
  assign LIOI3_TBYTESRC_X0Y107_OLOGIC_X0Y107_T1 = 1'b1;
  assign RIOB33_X105Y171_IOB_X1Y172_O = CLBLL_L_X2Y148_SLICE_X0Y148_AQ;
  assign RIOB33_X105Y171_IOB_X1Y171_O = CLBLM_L_X8Y153_SLICE_X11Y153_DO6;
  assign CLBLM_R_X5Y153_SLICE_X7Y153_A1 = CLBLM_R_X5Y153_SLICE_X7Y153_AQ;
  assign CLBLM_R_X5Y153_SLICE_X7Y153_A2 = CLBLM_R_X7Y153_SLICE_X9Y153_D5Q;
  assign CLBLM_R_X5Y153_SLICE_X7Y153_A3 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X5Y153_SLICE_X7Y153_A4 = CLBLM_R_X5Y153_SLICE_X7Y153_DO5;
  assign CLBLM_R_X5Y153_SLICE_X7Y153_A5 = CLBLL_L_X4Y147_SLICE_X4Y147_B5Q;
  assign CLBLM_R_X5Y153_SLICE_X7Y153_A6 = CLBLM_L_X8Y149_SLICE_X11Y149_AQ;
  assign CLBLM_R_X5Y153_SLICE_X7Y153_B1 = CLBLM_R_X7Y152_SLICE_X9Y152_CQ;
  assign CLBLM_R_X5Y153_SLICE_X7Y153_B2 = CLBLM_R_X5Y153_SLICE_X7Y153_BQ;
  assign CLBLM_R_X5Y153_SLICE_X7Y153_B3 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X5Y153_SLICE_X7Y153_B4 = CLBLL_L_X4Y147_SLICE_X5Y147_CQ;
  assign CLBLM_R_X5Y153_SLICE_X7Y153_B5 = CLBLL_L_X4Y153_SLICE_X4Y153_A5Q;
  assign CLBLM_R_X5Y153_SLICE_X7Y153_B6 = CLBLL_L_X4Y142_SLICE_X5Y142_DQ;
  assign CLBLM_R_X7Y155_SLICE_X8Y155_B5 = CLBLM_R_X7Y154_SLICE_X9Y154_AQ;
  assign CLBLM_R_X7Y155_SLICE_X8Y155_B6 = 1'b1;
  assign CLBLM_R_X5Y153_SLICE_X7Y153_C1 = CLBLM_L_X12Y151_SLICE_X16Y151_AQ;
  assign CLBLM_R_X5Y153_SLICE_X7Y153_C2 = CLBLM_R_X11Y148_SLICE_X15Y148_AO6;
  assign CLBLM_R_X5Y153_SLICE_X7Y153_C3 = 1'b1;
  assign CLBLM_R_X5Y153_SLICE_X7Y153_C4 = CLBLM_R_X5Y153_SLICE_X7Y153_BQ;
  assign CLBLM_R_X5Y153_SLICE_X7Y153_C5 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X5Y153_SLICE_X7Y153_C6 = CLBLM_R_X5Y153_SLICE_X7Y153_CQ;
  assign CLBLM_R_X3Y143_SLICE_X3Y143_A1 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X3Y143_SLICE_X3Y143_A2 = CLBLM_R_X3Y147_SLICE_X3Y147_BQ;
  assign CLBLM_R_X5Y153_SLICE_X7Y153_CLK = CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O;
  assign CLBLM_R_X3Y143_SLICE_X3Y143_A3 = CLBLM_R_X3Y143_SLICE_X3Y143_AQ;
  assign CLBLM_R_X3Y143_SLICE_X3Y143_A4 = CLBLL_L_X4Y151_SLICE_X4Y151_BQ;
  assign CLBLM_R_X3Y143_SLICE_X3Y143_A5 = CLBLM_R_X3Y145_SLICE_X3Y145_D5Q;
  assign CLBLM_R_X3Y143_SLICE_X3Y143_A6 = CLBLL_L_X4Y143_SLICE_X4Y143_D5Q;
  assign CLBLM_R_X5Y153_SLICE_X7Y153_D1 = CLBLM_R_X5Y148_SLICE_X6Y148_CO6;
  assign CLBLM_R_X5Y153_SLICE_X7Y153_D2 = CLBLM_L_X8Y153_SLICE_X10Y153_A5Q;
  assign CLBLM_R_X5Y153_SLICE_X7Y153_D3 = CLBLM_R_X5Y151_SLICE_X7Y151_AQ;
  assign CLBLM_R_X5Y153_SLICE_X7Y153_D4 = CLBLM_L_X8Y149_SLICE_X11Y149_AQ;
  assign CLBLM_R_X5Y153_SLICE_X7Y153_D5 = CLBLM_R_X5Y153_SLICE_X7Y153_AQ;
  assign CLBLM_R_X5Y153_SLICE_X7Y153_D6 = 1'b1;
  assign CLBLM_R_X3Y143_SLICE_X3Y143_B3 = CLBLM_R_X5Y141_SLICE_X6Y141_BQ;
  assign CLBLM_R_X3Y143_SLICE_X3Y143_B4 = 1'b1;
  assign CLBLM_R_X3Y143_SLICE_X3Y143_B6 = CLBLL_L_X4Y143_SLICE_X5Y143_B5Q;
  assign CLBLM_R_X3Y143_SLICE_X3Y143_C1 = CLBLM_R_X3Y151_SLICE_X3Y151_AQ;
  assign CLBLM_R_X3Y143_SLICE_X3Y143_C2 = LIOB33_X0Y57_IOB_X0Y58_I;
  assign CLBLM_R_X3Y143_SLICE_X3Y143_C3 = CLBLM_R_X5Y146_SLICE_X6Y146_AQ;
  assign CLBLM_R_X5Y153_SLICE_X6Y153_A2 = CLBLM_R_X5Y153_SLICE_X6Y153_BQ;
  assign CLBLM_R_X5Y153_SLICE_X6Y153_A3 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X5Y153_SLICE_X6Y153_A4 = CLBLL_L_X4Y148_SLICE_X5Y148_AQ;
  assign CLBLM_R_X3Y143_SLICE_X3Y143_C4 = CLBLM_R_X3Y143_SLICE_X3Y143_CQ;
  assign CLBLM_R_X3Y143_SLICE_X3Y143_C5 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X3Y143_SLICE_X3Y143_C6 = 1'b1;
  assign CLBLM_R_X3Y143_SLICE_X3Y143_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X5Y153_SLICE_X6Y153_A1 = 1'b1;
  assign CLBLM_R_X3Y143_SLICE_X3Y143_D1 = CLBLL_L_X4Y143_SLICE_X4Y143_C5Q;
  assign CLBLM_R_X3Y143_SLICE_X3Y143_D2 = CLBLL_L_X4Y144_SLICE_X4Y144_CQ;
  assign CLBLM_R_X3Y143_SLICE_X3Y143_D3 = 1'b1;
  assign CLBLM_R_X5Y153_SLICE_X6Y153_B3 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X5Y153_SLICE_X6Y153_B4 = RIOB33_X105Y131_IOB_X1Y131_I;
  assign CLBLM_R_X5Y153_SLICE_X6Y153_B5 = CLBLM_R_X3Y151_SLICE_X2Y151_AQ;
  assign CLBLM_R_X5Y153_SLICE_X6Y153_B6 = 1'b1;
  assign CLBLM_R_X3Y143_SLICE_X3Y143_D4 = 1'b1;
  assign CLBLM_R_X3Y143_SLICE_X3Y143_D5 = 1'b1;
  assign CLBLM_R_X3Y143_SLICE_X3Y143_D6 = 1'b1;
  assign CLBLM_R_X5Y153_SLICE_X6Y153_C1 = CLBLM_R_X3Y153_SLICE_X2Y153_AQ;
  assign CLBLM_R_X5Y153_SLICE_X6Y153_C2 = CLBLM_R_X3Y147_SLICE_X2Y147_CQ;
  assign CLBLM_R_X5Y153_SLICE_X6Y153_C3 = CLBLM_L_X8Y144_SLICE_X10Y144_AQ;
  assign CLBLM_R_X5Y153_SLICE_X6Y153_C4 = RIOB33_X105Y105_IOB_X1Y106_I;
  assign CLBLM_R_X5Y153_SLICE_X6Y153_C5 = 1'b1;
  assign CLBLM_R_X5Y153_SLICE_X6Y153_C6 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X3Y143_SLICE_X2Y143_A1 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X3Y143_SLICE_X2Y143_A2 = CLBLM_L_X8Y144_SLICE_X11Y144_B5Q;
  assign CLBLM_R_X3Y143_SLICE_X2Y143_A3 = CLBLM_R_X3Y143_SLICE_X2Y143_AQ;
  assign CLBLM_R_X5Y153_SLICE_X6Y153_CLK = CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O;
  assign CLBLM_R_X3Y143_SLICE_X2Y143_AX = CLBLM_R_X3Y143_SLICE_X2Y143_BO6;
  assign CLBLM_R_X3Y143_SLICE_X2Y143_B3 = CLBLL_L_X4Y145_SLICE_X4Y145_AQ;
  assign CLBLM_R_X3Y143_SLICE_X2Y143_B4 = CLBLM_R_X3Y143_SLICE_X3Y143_CQ;
  assign CLBLM_R_X3Y143_SLICE_X2Y143_B5 = CLBLM_R_X3Y143_SLICE_X2Y143_A5Q;
  assign CLBLM_R_X3Y143_SLICE_X2Y143_B1 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X5Y153_SLICE_X6Y153_D1 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X5Y153_SLICE_X6Y153_D2 = 1'b1;
  assign CLBLM_R_X5Y153_SLICE_X6Y153_D3 = CLBLM_L_X8Y153_SLICE_X10Y153_DQ;
  assign CLBLM_R_X5Y153_SLICE_X6Y153_D4 = CLBLM_L_X8Y144_SLICE_X11Y144_AQ;
  assign CLBLM_R_X5Y153_SLICE_X6Y153_D5 = CLBLL_L_X4Y153_SLICE_X4Y153_A5Q;
  assign CLBLM_R_X5Y153_SLICE_X6Y153_D6 = 1'b1;
  assign CLBLM_R_X3Y143_SLICE_X2Y143_B6 = 1'b1;
  assign CLBLM_R_X3Y143_SLICE_X2Y143_C1 = CLBLL_L_X4Y142_SLICE_X4Y142_BQ;
  assign CLBLM_R_X3Y143_SLICE_X2Y143_C6 = 1'b1;
  assign CLBLM_R_X3Y143_SLICE_X2Y143_C2 = CLBLM_R_X3Y142_SLICE_X3Y142_AQ;
  assign CLBLM_R_X3Y143_SLICE_X2Y143_C3 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X3Y143_SLICE_X2Y143_C4 = CLBLM_R_X5Y144_SLICE_X6Y144_AQ;
  assign CLBLM_R_X3Y143_SLICE_X2Y143_C5 = CLBLM_R_X5Y147_SLICE_X6Y147_AQ;
  assign CLBLM_R_X3Y143_SLICE_X2Y143_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign LIOI3_X0Y61_ILOGIC_X0Y61_D = LIOB33_X0Y61_IOB_X0Y61_I;
  assign CLBLM_R_X3Y143_SLICE_X2Y143_D1 = 1'b1;
  assign CLBLM_R_X3Y143_SLICE_X2Y143_D2 = 1'b1;
  assign CLBLM_R_X3Y143_SLICE_X2Y143_D3 = 1'b1;
  assign CLBLM_R_X3Y143_SLICE_X2Y143_D4 = 1'b1;
  assign CLBLM_R_X3Y143_SLICE_X2Y143_D5 = 1'b1;
  assign CLBLM_R_X3Y143_SLICE_X2Y143_D6 = 1'b1;
  assign RIOI3_X105Y105_ILOGIC_X1Y106_D = RIOB33_X105Y105_IOB_X1Y106_I;
  assign RIOI3_X105Y105_ILOGIC_X1Y105_D = RIOB33_X105Y105_IOB_X1Y105_I;
  assign RIOI3_TBYTETERM_X105Y113_ILOGIC_X1Y113_D = RIOB33_X105Y113_IOB_X1Y113_I;
  assign RIOB33_X105Y173_IOB_X1Y174_O = CLBLM_R_X5Y152_SLICE_X7Y152_DO6;
  assign RIOB33_X105Y173_IOB_X1Y173_O = CLBLM_R_X5Y152_SLICE_X7Y152_DQ;
  assign CLBLM_R_X5Y154_SLICE_X7Y154_A1 = CLBLL_L_X4Y150_SLICE_X4Y150_A5Q;
  assign CLBLM_R_X5Y154_SLICE_X7Y154_A2 = CLBLM_R_X5Y150_SLICE_X7Y150_BO6;
  assign CLBLM_R_X5Y154_SLICE_X7Y154_A3 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X5Y154_SLICE_X7Y154_A4 = CLBLM_R_X5Y154_SLICE_X6Y154_BQ;
  assign CLBLM_R_X5Y154_SLICE_X7Y154_A5 = 1'b1;
  assign CLBLM_R_X5Y154_SLICE_X7Y154_A6 = CLBLM_R_X3Y149_SLICE_X2Y149_AQ;
  assign CLBLM_R_X5Y154_SLICE_X7Y154_B1 = 1'b1;
  assign CLBLM_R_X5Y154_SLICE_X7Y154_B2 = 1'b1;
  assign CLBLM_R_X5Y154_SLICE_X7Y154_B3 = 1'b1;
  assign CLBLM_R_X5Y154_SLICE_X7Y154_B4 = 1'b1;
  assign CLBLM_R_X5Y154_SLICE_X7Y154_B5 = 1'b1;
  assign CLBLM_R_X5Y154_SLICE_X7Y154_B6 = 1'b1;
  assign CLBLM_R_X5Y154_SLICE_X7Y154_C1 = 1'b1;
  assign CLBLM_R_X5Y154_SLICE_X7Y154_C2 = 1'b1;
  assign CLBLM_R_X5Y154_SLICE_X7Y154_C3 = 1'b1;
  assign CLBLM_R_X5Y154_SLICE_X7Y154_C4 = 1'b1;
  assign CLBLM_R_X5Y154_SLICE_X7Y154_C5 = 1'b1;
  assign CLBLM_R_X5Y154_SLICE_X7Y154_C6 = 1'b1;
  assign CLBLM_R_X3Y144_SLICE_X3Y144_A1 = CLBLM_R_X3Y144_SLICE_X3Y144_DO6;
  assign CLBLM_R_X3Y144_SLICE_X3Y144_A2 = CLBLL_L_X2Y144_SLICE_X1Y144_AO6;
  assign CLBLM_R_X5Y154_SLICE_X7Y154_CLK = CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O;
  assign CLBLM_R_X3Y144_SLICE_X3Y144_A3 = CLBLM_R_X3Y144_SLICE_X2Y144_AO6;
  assign CLBLM_R_X3Y144_SLICE_X3Y144_A4 = CLBLL_L_X4Y153_SLICE_X4Y153_BQ;
  assign CLBLM_R_X3Y144_SLICE_X3Y144_A5 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X3Y144_SLICE_X3Y144_A6 = CLBLM_R_X5Y147_SLICE_X6Y147_B5Q;
  assign CLBLM_R_X5Y154_SLICE_X7Y154_D1 = 1'b1;
  assign CLBLM_R_X5Y154_SLICE_X7Y154_D2 = 1'b1;
  assign CLBLM_R_X5Y154_SLICE_X7Y154_D3 = 1'b1;
  assign CLBLM_R_X5Y154_SLICE_X7Y154_D4 = 1'b1;
  assign CLBLM_R_X5Y154_SLICE_X7Y154_D5 = 1'b1;
  assign CLBLM_R_X5Y154_SLICE_X7Y154_D6 = 1'b1;
  assign CLBLM_R_X3Y144_SLICE_X3Y144_B3 = CLBLM_R_X3Y144_SLICE_X3Y144_AQ;
  assign CLBLM_R_X3Y144_SLICE_X3Y144_B4 = CLBLM_R_X3Y142_SLICE_X3Y142_BO6;
  assign CLBLM_R_X3Y144_SLICE_X3Y144_B6 = CLBLM_R_X3Y145_SLICE_X3Y145_CQ;
  assign CLBLM_R_X3Y144_SLICE_X3Y144_C1 = CLBLM_R_X3Y143_SLICE_X3Y143_CQ;
  assign CLBLM_R_X3Y144_SLICE_X3Y144_C2 = CLBLM_R_X3Y145_SLICE_X3Y145_CQ;
  assign CLBLM_R_X3Y144_SLICE_X3Y144_C3 = LIOB33_X0Y57_IOB_X0Y58_I;
  assign CLBLM_R_X3Y144_SLICE_X3Y144_C4 = CLBLM_R_X3Y143_SLICE_X2Y143_A5Q;
  assign CLBLM_R_X3Y144_SLICE_X3Y144_C5 = CLBLM_R_X3Y144_SLICE_X3Y144_AQ;
  assign CLBLM_R_X5Y154_SLICE_X6Y154_A4 = CLBLM_R_X5Y154_SLICE_X6Y154_AQ;
  assign CLBLM_R_X3Y144_SLICE_X3Y144_C6 = CLBLL_L_X2Y146_SLICE_X1Y146_B5Q;
  assign CLBLM_R_X5Y154_SLICE_X6Y154_A6 = CLBLM_L_X10Y153_SLICE_X12Y153_BQ;
  assign CLBLM_R_X3Y144_SLICE_X3Y144_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X5Y154_SLICE_X6Y154_A1 = CLBLL_L_X2Y150_SLICE_X1Y150_AQ;
  assign CLBLM_R_X5Y154_SLICE_X6Y154_A2 = CLBLM_R_X5Y154_SLICE_X6Y154_BQ;
  assign CLBLM_R_X5Y154_SLICE_X6Y154_B1 = CLBLL_L_X2Y150_SLICE_X1Y150_AQ;
  assign CLBLM_R_X5Y154_SLICE_X6Y154_B2 = CLBLM_R_X5Y154_SLICE_X6Y154_BQ;
  assign CLBLM_R_X5Y154_SLICE_X6Y154_B3 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X5Y154_SLICE_X6Y154_B4 = CLBLM_R_X5Y148_SLICE_X7Y148_CQ;
  assign CLBLM_R_X5Y154_SLICE_X6Y154_B5 = CLBLL_L_X4Y153_SLICE_X5Y153_BO5;
  assign CLBLM_R_X5Y154_SLICE_X6Y154_B6 = 1'b1;
  assign CLBLM_R_X3Y144_SLICE_X3Y144_D3 = CLBLM_R_X3Y144_SLICE_X2Y144_BO6;
  assign CLBLM_R_X3Y144_SLICE_X3Y144_D4 = CLBLM_R_X3Y145_SLICE_X3Y145_CQ;
  assign CLBLM_R_X3Y144_SLICE_X3Y144_D6 = CLBLM_R_X3Y142_SLICE_X3Y142_BO6;
  assign CLBLM_R_X5Y154_SLICE_X6Y154_C1 = 1'b1;
  assign CLBLM_R_X5Y154_SLICE_X6Y154_C2 = 1'b1;
  assign CLBLM_R_X5Y154_SLICE_X6Y154_C3 = 1'b1;
  assign CLBLM_R_X5Y154_SLICE_X6Y154_C4 = 1'b1;
  assign CLBLM_R_X5Y154_SLICE_X6Y154_C5 = 1'b1;
  assign CLBLM_R_X5Y154_SLICE_X6Y154_C6 = 1'b1;
  assign CLBLM_R_X3Y144_SLICE_X2Y144_A1 = CLBLM_R_X3Y145_SLICE_X3Y145_CQ;
  assign CLBLM_R_X3Y144_SLICE_X2Y144_AX = CLBLM_R_X3Y144_SLICE_X2Y144_BO5;
  assign CLBLM_R_X3Y144_SLICE_X2Y144_A2 = CLBLL_L_X2Y146_SLICE_X1Y146_B5Q;
  assign CLBLM_R_X3Y144_SLICE_X2Y144_B1 = CLBLM_R_X3Y143_SLICE_X2Y143_A5Q;
  assign CLBLM_R_X3Y144_SLICE_X2Y144_B2 = LIOB33_X0Y57_IOB_X0Y58_I;
  assign CLBLM_R_X3Y144_SLICE_X2Y144_B3 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X5Y154_SLICE_X6Y154_CLK = CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O;
  assign CLBLM_R_X3Y144_SLICE_X2Y144_B4 = CLBLM_R_X3Y150_SLICE_X2Y150_AQ;
  assign CLBLM_R_X3Y144_SLICE_X2Y144_B5 = CLBLM_R_X3Y143_SLICE_X3Y143_CQ;
  assign CLBLM_R_X5Y154_SLICE_X6Y154_D1 = 1'b1;
  assign CLBLM_R_X5Y154_SLICE_X6Y154_D2 = 1'b1;
  assign CLBLM_R_X5Y154_SLICE_X6Y154_D3 = 1'b1;
  assign CLBLM_R_X5Y154_SLICE_X6Y154_D4 = 1'b1;
  assign CLBLM_R_X5Y154_SLICE_X6Y154_D5 = 1'b1;
  assign CLBLM_R_X5Y154_SLICE_X6Y154_D6 = 1'b1;
  assign CLBLM_R_X3Y144_SLICE_X2Y144_C3 = CLBLM_R_X3Y144_SLICE_X3Y144_AQ;
  assign CLBLM_R_X3Y144_SLICE_X2Y144_C4 = CLBLM_R_X5Y143_SLICE_X6Y143_D5Q;
  assign CLBLM_R_X3Y144_SLICE_X2Y144_C1 = CLBLL_L_X2Y146_SLICE_X1Y146_B5Q;
  assign CLBLM_R_X3Y144_SLICE_X2Y144_C2 = CLBLM_R_X3Y145_SLICE_X3Y145_CQ;
  assign CLBLM_R_X3Y144_SLICE_X2Y144_C5 = CLBLM_R_X3Y144_SLICE_X2Y144_DO6;
  assign CLBLM_R_X3Y144_SLICE_X2Y144_C6 = CLBLM_R_X3Y144_SLICE_X2Y144_BO6;
  assign CLBLM_R_X3Y144_SLICE_X2Y144_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X3Y144_SLICE_X2Y144_D1 = CLBLM_R_X5Y153_SLICE_X6Y153_B5Q;
  assign CLBLM_R_X3Y144_SLICE_X2Y144_D2 = CLBLL_L_X2Y146_SLICE_X0Y146_DQ;
  assign CLBLM_R_X3Y144_SLICE_X2Y144_D3 = CLBLM_R_X3Y144_SLICE_X3Y144_AQ;
  assign CLBLM_R_X3Y144_SLICE_X2Y144_D4 = CLBLL_L_X2Y146_SLICE_X1Y146_B5Q;
  assign CLBLM_R_X3Y144_SLICE_X2Y144_D5 = CLBLM_R_X3Y145_SLICE_X3Y145_CQ;
  assign CLBLM_R_X3Y144_SLICE_X2Y144_D6 = 1'b1;
  assign RIOB33_X105Y175_IOB_X1Y176_O = CLBLL_L_X2Y148_SLICE_X1Y148_BO6;
  assign RIOB33_X105Y175_IOB_X1Y175_O = CLBLM_L_X10Y144_SLICE_X12Y144_BO6;
  assign CLBLM_R_X7Y145_SLICE_X8Y145_B2 = CLBLM_L_X8Y152_SLICE_X10Y152_A5Q;
  assign CLBLM_R_X7Y145_SLICE_X8Y145_B3 = CLBLM_R_X7Y149_SLICE_X8Y149_AQ;
  assign CLBLM_R_X7Y145_SLICE_X8Y145_B4 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X7Y145_SLICE_X8Y145_B5 = 1'b1;
  assign CLBLM_R_X7Y145_SLICE_X8Y145_B6 = 1'b1;
  assign CLBLM_R_X7Y145_SLICE_X8Y145_C1 = CLBLM_L_X8Y153_SLICE_X10Y153_D5Q;
  assign LIOI3_X0Y185_OLOGIC_X0Y186_D1 = RIOB33_X105Y119_IOB_X1Y120_I;
  assign LIOI3_X0Y185_OLOGIC_X0Y186_T1 = 1'b1;
  assign LIOI3_X0Y125_OLOGIC_X0Y126_D1 = CLBLL_L_X4Y147_SLICE_X5Y147_CQ;
  assign LIOI3_X0Y185_OLOGIC_X0Y185_D1 = RIOB33_X105Y133_IOB_X1Y133_I;
  assign LIOI3_X0Y125_OLOGIC_X0Y126_T1 = 1'b1;
  assign RIOI3_X105Y171_OLOGIC_X1Y172_D1 = CLBLL_L_X2Y148_SLICE_X0Y148_AQ;
  assign LIOI3_X0Y65_OLOGIC_X0Y66_D1 = CLBLL_L_X4Y151_SLICE_X4Y151_CQ;
  assign LIOI3_X0Y185_OLOGIC_X0Y185_T1 = 1'b1;
  assign LIOI3_X0Y125_OLOGIC_X0Y125_D1 = CLBLL_L_X4Y151_SLICE_X4Y151_BQ;
  assign RIOI3_X105Y171_OLOGIC_X1Y172_T1 = 1'b1;
  assign LIOI3_X0Y65_OLOGIC_X0Y66_T1 = 1'b1;
  assign CLBLM_R_X3Y145_SLICE_X3Y145_A1 = CLBLL_L_X4Y152_SLICE_X4Y152_DQ;
  assign CLBLM_R_X3Y145_SLICE_X3Y145_A2 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X3Y145_SLICE_X3Y145_A3 = CLBLL_L_X4Y145_SLICE_X4Y145_B5Q;
  assign CLBLM_R_X3Y145_SLICE_X3Y145_A4 = CLBLM_R_X3Y145_SLICE_X3Y145_AQ;
  assign CLBLM_R_X3Y145_SLICE_X3Y145_A5 = CLBLL_L_X4Y142_SLICE_X5Y142_DQ;
  assign CLBLM_R_X3Y145_SLICE_X3Y145_A6 = CLBLL_L_X4Y147_SLICE_X5Y147_CQ;
  assign LIOI3_X0Y65_OLOGIC_X0Y65_D1 = CLBLM_R_X7Y141_SLICE_X8Y141_BO6;
  assign LIOI3_X0Y125_OLOGIC_X0Y125_T1 = 1'b1;
  assign RIOI3_X105Y171_OLOGIC_X1Y171_D1 = CLBLM_L_X8Y153_SLICE_X11Y153_DO6;
  assign CLBLM_R_X3Y145_SLICE_X3Y145_B1 = CLBLL_L_X4Y145_SLICE_X4Y145_DO6;
  assign CLBLM_R_X3Y145_SLICE_X3Y145_B2 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X3Y145_SLICE_X3Y145_B3 = CLBLM_R_X3Y146_SLICE_X2Y146_C5Q;
  assign CLBLM_R_X3Y145_SLICE_X3Y145_B4 = 1'b1;
  assign CLBLM_R_X3Y145_SLICE_X3Y145_B5 = CLBLM_R_X3Y145_SLICE_X3Y145_BQ;
  assign CLBLM_R_X3Y145_SLICE_X3Y145_B6 = CLBLM_R_X3Y145_SLICE_X2Y145_CQ;
  assign LIOI3_TBYTESRC_X0Y119_OLOGIC_X0Y120_D1 = CLBLL_L_X4Y147_SLICE_X4Y147_AQ;
  assign LIOI3_X0Y65_OLOGIC_X0Y65_T1 = 1'b1;
  assign RIOI3_X105Y171_OLOGIC_X1Y171_T1 = 1'b1;
  assign CLBLM_R_X3Y145_SLICE_X3Y145_C1 = CLBLM_R_X3Y143_SLICE_X2Y143_A5Q;
  assign CLBLM_R_X3Y145_SLICE_X3Y145_C2 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X3Y145_SLICE_X3Y145_C3 = CLBLM_R_X3Y144_SLICE_X3Y144_BO6;
  assign CLBLM_R_X3Y145_SLICE_X3Y145_C4 = CLBLM_R_X3Y144_SLICE_X3Y144_CO6;
  assign CLBLM_R_X3Y145_SLICE_X3Y145_C5 = CLBLM_L_X10Y151_SLICE_X13Y151_A5Q;
  assign CLBLM_R_X3Y145_SLICE_X3Y145_C6 = 1'b1;
  assign LIOI3_TBYTESRC_X0Y119_OLOGIC_X0Y120_T1 = 1'b1;
  assign CLBLM_R_X3Y145_SLICE_X3Y145_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X3Y145_SLICE_X3Y145_D1 = CLBLL_L_X4Y151_SLICE_X4Y151_BQ;
  assign CLBLM_R_X3Y145_SLICE_X3Y145_D2 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X3Y145_SLICE_X3Y145_D3 = 1'b1;
  assign CLBLM_R_X3Y145_SLICE_X3Y145_D4 = CLBLM_R_X3Y146_SLICE_X2Y146_BQ;
  assign CLBLM_R_X3Y145_SLICE_X3Y145_D5 = CLBLM_R_X7Y146_SLICE_X8Y146_CQ;
  assign CLBLM_R_X3Y145_SLICE_X3Y145_D6 = 1'b1;
  assign LIOI3_TBYTESRC_X0Y119_OLOGIC_X0Y119_D1 = CLBLL_L_X2Y146_SLICE_X0Y146_CQ;
  assign CLBLM_R_X3Y145_SLICE_X2Y145_A1 = CLBLM_L_X10Y145_SLICE_X12Y145_AQ;
  assign CLBLM_R_X3Y145_SLICE_X2Y145_A2 = CLBLM_R_X3Y145_SLICE_X2Y145_BQ;
  assign CLBLM_R_X3Y145_SLICE_X2Y145_A3 = CLBLM_R_X3Y145_SLICE_X2Y145_AQ;
  assign CLBLM_R_X3Y145_SLICE_X2Y145_A4 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X3Y145_SLICE_X2Y145_A5 = CLBLM_R_X3Y143_SLICE_X2Y143_AQ;
  assign CLBLM_R_X3Y145_SLICE_X2Y145_A6 = CLBLM_R_X5Y142_SLICE_X7Y142_BQ;
  assign LIOI3_TBYTESRC_X0Y119_OLOGIC_X0Y119_T1 = 1'b1;
  assign CLBLM_R_X3Y145_SLICE_X2Y145_B1 = CLBLL_L_X4Y146_SLICE_X4Y146_C5Q;
  assign CLBLM_R_X3Y145_SLICE_X2Y145_B2 = CLBLM_R_X3Y145_SLICE_X2Y145_BQ;
  assign CLBLM_R_X3Y145_SLICE_X2Y145_B3 = CLBLL_L_X4Y145_SLICE_X4Y145_B5Q;
  assign CLBLM_R_X3Y145_SLICE_X2Y145_B4 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X3Y145_SLICE_X2Y145_B5 = CLBLM_R_X3Y151_SLICE_X3Y151_BQ;
  assign CLBLM_R_X3Y145_SLICE_X2Y145_B6 = 1'b1;
  assign CLBLM_R_X3Y145_SLICE_X2Y145_C1 = CLBLM_R_X5Y143_SLICE_X6Y143_C5Q;
  assign CLBLM_R_X3Y145_SLICE_X2Y145_C2 = CLBLL_L_X4Y147_SLICE_X5Y147_BQ;
  assign CLBLM_R_X3Y145_SLICE_X2Y145_C3 = CLBLL_L_X4Y147_SLICE_X5Y147_C5Q;
  assign CLBLM_R_X3Y145_SLICE_X2Y145_C4 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X3Y145_SLICE_X2Y145_C5 = CLBLM_R_X7Y144_SLICE_X9Y144_A5Q;
  assign CLBLM_R_X3Y145_SLICE_X2Y145_C6 = 1'b1;
  assign CLBLM_R_X3Y145_SLICE_X2Y145_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X3Y145_SLICE_X2Y145_D1 = CLBLM_R_X3Y148_SLICE_X2Y148_A5Q;
  assign CLBLM_R_X3Y145_SLICE_X2Y145_D2 = CLBLL_L_X4Y145_SLICE_X4Y145_C5Q;
  assign CLBLM_R_X3Y145_SLICE_X2Y145_D3 = CLBLM_R_X3Y147_SLICE_X2Y147_DQ;
  assign CLBLM_R_X3Y145_SLICE_X2Y145_D4 = CLBLM_L_X10Y153_SLICE_X13Y153_CQ;
  assign CLBLM_R_X3Y145_SLICE_X2Y145_D5 = CLBLM_R_X5Y145_SLICE_X6Y145_B5Q;
  assign CLBLM_R_X3Y145_SLICE_X2Y145_D6 = CLBLL_L_X4Y145_SLICE_X5Y145_CQ;
  assign RIOB33_X105Y177_IOB_X1Y178_O = CLBLM_R_X5Y147_SLICE_X6Y147_AQ;
  assign RIOB33_X105Y177_IOB_X1Y177_O = CLBLL_L_X2Y146_SLICE_X1Y146_B5Q;
  assign RIOI3_X105Y109_ILOGIC_X1Y110_D = RIOB33_X105Y109_IOB_X1Y110_I;
  assign RIOI3_X105Y109_ILOGIC_X1Y109_D = RIOB33_X105Y109_IOB_X1Y109_I;
  assign RIOI3_TBYTETERM_X105Y137_ILOGIC_X1Y138_D = RIOB33_X105Y137_IOB_X1Y138_I;
  assign RIOI3_TBYTETERM_X105Y137_ILOGIC_X1Y137_D = RIOB33_X105Y137_IOB_X1Y137_I;
  assign CLBLM_R_X3Y146_SLICE_X3Y146_A1 = 1'b1;
  assign CLBLM_R_X3Y146_SLICE_X3Y146_A2 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X3Y146_SLICE_X3Y146_A3 = CLBLM_R_X7Y146_SLICE_X8Y146_BQ;
  assign CLBLM_R_X3Y146_SLICE_X3Y146_A4 = CLBLM_R_X3Y146_SLICE_X2Y146_BQ;
  assign CLBLM_R_X3Y146_SLICE_X3Y146_A5 = CLBLM_R_X3Y145_SLICE_X3Y145_AQ;
  assign CLBLM_R_X3Y146_SLICE_X3Y146_A6 = CLBLM_R_X3Y146_SLICE_X3Y146_CO6;
  assign CLBLM_R_X3Y146_SLICE_X3Y146_B1 = CLBLM_R_X3Y146_SLICE_X2Y146_DQ;
  assign CLBLM_R_X3Y146_SLICE_X3Y146_B2 = CLBLM_R_X3Y146_SLICE_X3Y146_BQ;
  assign CLBLM_R_X3Y146_SLICE_X3Y146_B3 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X3Y146_SLICE_X3Y146_B4 = CLBLL_L_X4Y152_SLICE_X4Y152_DQ;
  assign CLBLM_R_X3Y146_SLICE_X3Y146_B5 = CLBLL_L_X4Y146_SLICE_X5Y146_AQ;
  assign CLBLM_R_X3Y146_SLICE_X3Y146_B6 = CLBLM_R_X3Y149_SLICE_X3Y149_CQ;
  assign CLBLM_R_X3Y146_SLICE_X3Y146_C1 = CLBLL_L_X4Y146_SLICE_X4Y146_DO5;
  assign CLBLM_R_X3Y146_SLICE_X3Y146_C2 = CLBLL_L_X2Y145_SLICE_X1Y145_CQ;
  assign CLBLM_R_X3Y146_SLICE_X3Y146_C3 = CLBLM_R_X3Y149_SLICE_X3Y149_DQ;
  assign CLBLM_R_X3Y146_SLICE_X3Y146_C4 = CLBLM_R_X5Y146_SLICE_X6Y146_CO6;
  assign CLBLM_R_X3Y146_SLICE_X3Y146_C5 = CLBLM_R_X3Y146_SLICE_X3Y146_DO6;
  assign CLBLM_R_X3Y146_SLICE_X3Y146_C6 = 1'b1;
  assign CLBLM_R_X3Y146_SLICE_X3Y146_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X3Y146_SLICE_X3Y146_D1 = CLBLL_L_X2Y145_SLICE_X1Y145_BQ;
  assign CLBLM_R_X3Y146_SLICE_X3Y146_D2 = CLBLM_R_X3Y148_SLICE_X3Y148_C5Q;
  assign CLBLM_R_X3Y146_SLICE_X3Y146_D3 = CLBLL_L_X4Y149_SLICE_X4Y149_AQ;
  assign CLBLM_R_X3Y146_SLICE_X3Y146_D4 = CLBLM_R_X5Y150_SLICE_X7Y150_A5Q;
  assign CLBLM_R_X3Y146_SLICE_X3Y146_D5 = 1'b1;
  assign CLBLM_R_X3Y146_SLICE_X3Y146_D6 = 1'b1;
  assign CLBLM_R_X3Y146_SLICE_X2Y146_A1 = CLBLM_R_X5Y142_SLICE_X7Y142_BQ;
  assign CLBLM_R_X3Y146_SLICE_X2Y146_A2 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X3Y146_SLICE_X2Y146_A3 = CLBLM_R_X3Y146_SLICE_X2Y146_AQ;
  assign CLBLM_R_X3Y146_SLICE_X2Y146_A4 = CLBLM_L_X10Y145_SLICE_X12Y145_AQ;
  assign CLBLM_R_X3Y146_SLICE_X2Y146_A5 = CLBLM_R_X3Y143_SLICE_X3Y143_C5Q;
  assign CLBLM_R_X3Y146_SLICE_X2Y146_A6 = CLBLM_R_X3Y145_SLICE_X2Y145_C5Q;
  assign LIOB33_X0Y139_IOB_X0Y139_O = CLBLM_R_X3Y147_SLICE_X2Y147_DQ;
  assign LIOB33_X0Y139_IOB_X0Y140_O = CLBLL_L_X4Y145_SLICE_X4Y145_C5Q;
  assign CLBLM_R_X3Y146_SLICE_X2Y146_B1 = CLBLM_R_X5Y149_SLICE_X6Y149_B5Q;
  assign CLBLM_R_X3Y146_SLICE_X2Y146_B2 = CLBLM_R_X3Y146_SLICE_X2Y146_BQ;
  assign CLBLM_R_X3Y146_SLICE_X2Y146_B3 = CLBLL_L_X4Y143_SLICE_X4Y143_D5Q;
  assign CLBLM_R_X3Y146_SLICE_X2Y146_B4 = 1'b1;
  assign CLBLM_R_X3Y146_SLICE_X2Y146_B5 = CLBLL_L_X2Y146_SLICE_X1Y146_DO6;
  assign CLBLM_R_X3Y146_SLICE_X2Y146_B6 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X3Y146_SLICE_X2Y146_C1 = CLBLM_R_X5Y150_SLICE_X6Y150_C5Q;
  assign CLBLM_R_X3Y146_SLICE_X2Y146_C2 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X3Y146_SLICE_X2Y146_C3 = CLBLM_R_X3Y147_SLICE_X2Y147_D5Q;
  assign CLBLM_R_X3Y146_SLICE_X2Y146_C4 = CLBLM_R_X7Y142_SLICE_X9Y142_CQ;
  assign CLBLM_R_X3Y146_SLICE_X2Y146_C5 = CLBLL_L_X4Y149_SLICE_X5Y149_CQ;
  assign CLBLM_R_X3Y146_SLICE_X2Y146_C6 = 1'b1;
  assign CLBLM_R_X3Y146_SLICE_X2Y146_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X3Y146_SLICE_X2Y146_D1 = CLBLL_L_X4Y147_SLICE_X4Y147_AQ;
  assign CLBLM_R_X3Y146_SLICE_X2Y146_D2 = CLBLM_R_X11Y148_SLICE_X14Y148_AO6;
  assign CLBLM_R_X3Y146_SLICE_X2Y146_D3 = CLBLL_L_X2Y145_SLICE_X1Y145_BQ;
  assign CLBLM_R_X3Y146_SLICE_X2Y146_D4 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X3Y146_SLICE_X2Y146_D5 = 1'b1;
  assign CLBLM_R_X3Y146_SLICE_X2Y146_D6 = 1'b1;
  assign RIOB33_X105Y179_IOB_X1Y180_O = CLBLM_L_X8Y145_SLICE_X11Y145_DQ;
  assign RIOB33_X105Y179_IOB_X1Y179_O = CLBLM_L_X8Y147_SLICE_X10Y147_BQ;
  assign CLBLL_L_X2Y166_SLICE_X0Y166_A1 = 1'b1;
  assign CLBLL_L_X2Y166_SLICE_X0Y166_A2 = 1'b1;
  assign CLBLL_L_X2Y166_SLICE_X0Y166_A3 = CLBLM_L_X12Y146_SLICE_X17Y146_AQ;
  assign CLBLL_L_X2Y166_SLICE_X0Y166_A4 = 1'b1;
  assign CLBLL_L_X2Y166_SLICE_X0Y166_A5 = 1'b1;
  assign CLBLL_L_X2Y166_SLICE_X0Y166_A6 = 1'b1;
  assign CLBLL_L_X2Y166_SLICE_X0Y166_B1 = 1'b1;
  assign CLBLL_L_X2Y166_SLICE_X0Y166_B2 = 1'b1;
  assign CLBLL_L_X2Y166_SLICE_X0Y166_B3 = 1'b1;
  assign CLBLL_L_X2Y166_SLICE_X0Y166_B4 = 1'b1;
  assign CLBLL_L_X2Y166_SLICE_X0Y166_B5 = 1'b1;
  assign CLBLL_L_X2Y166_SLICE_X0Y166_B6 = 1'b1;
  assign CLBLL_L_X2Y166_SLICE_X0Y166_C1 = 1'b1;
  assign CLBLL_L_X2Y166_SLICE_X0Y166_C2 = 1'b1;
  assign CLBLL_L_X2Y166_SLICE_X0Y166_C3 = 1'b1;
  assign CLBLL_L_X2Y166_SLICE_X0Y166_C4 = 1'b1;
  assign CLBLL_L_X2Y166_SLICE_X0Y166_C5 = 1'b1;
  assign CLBLL_L_X2Y166_SLICE_X0Y166_C6 = 1'b1;
  assign CLBLL_L_X2Y166_SLICE_X0Y166_D1 = 1'b1;
  assign CLBLL_L_X2Y166_SLICE_X0Y166_D2 = 1'b1;
  assign CLBLL_L_X2Y166_SLICE_X0Y166_D3 = 1'b1;
  assign CLBLL_L_X2Y166_SLICE_X0Y166_D4 = 1'b1;
  assign CLBLL_L_X2Y166_SLICE_X0Y166_D5 = 1'b1;
  assign CLBLL_L_X2Y166_SLICE_X0Y166_D6 = 1'b1;
  assign CLBLL_L_X2Y166_SLICE_X1Y166_A1 = 1'b1;
  assign CLBLL_L_X2Y166_SLICE_X1Y166_A2 = 1'b1;
  assign CLBLL_L_X2Y166_SLICE_X1Y166_A3 = 1'b1;
  assign CLBLL_L_X2Y166_SLICE_X1Y166_A4 = 1'b1;
  assign CLBLL_L_X2Y166_SLICE_X1Y166_A5 = 1'b1;
  assign CLBLL_L_X2Y166_SLICE_X1Y166_A6 = 1'b1;
  assign CLBLL_L_X2Y166_SLICE_X1Y166_B1 = 1'b1;
  assign CLBLL_L_X2Y166_SLICE_X1Y166_B2 = 1'b1;
  assign CLBLL_L_X2Y166_SLICE_X1Y166_B3 = 1'b1;
  assign CLBLL_L_X2Y166_SLICE_X1Y166_B4 = 1'b1;
  assign CLBLL_L_X2Y166_SLICE_X1Y166_B5 = 1'b1;
  assign CLBLL_L_X2Y166_SLICE_X1Y166_B6 = 1'b1;
  assign CLBLL_L_X2Y166_SLICE_X1Y166_C1 = 1'b1;
  assign CLBLL_L_X2Y166_SLICE_X1Y166_C2 = 1'b1;
  assign CLBLL_L_X2Y166_SLICE_X1Y166_C3 = 1'b1;
  assign CLBLL_L_X2Y166_SLICE_X1Y166_C4 = 1'b1;
  assign CLBLL_L_X2Y166_SLICE_X1Y166_C5 = 1'b1;
  assign CLBLL_L_X2Y166_SLICE_X1Y166_C6 = 1'b1;
  assign CLBLM_R_X3Y147_SLICE_X3Y147_A1 = CLBLM_R_X3Y147_SLICE_X3Y147_AQ;
  assign CLBLM_R_X3Y147_SLICE_X3Y147_A2 = CLBLM_R_X11Y148_SLICE_X15Y148_AO6;
  assign CLBLM_R_X3Y147_SLICE_X3Y147_A3 = CLBLM_R_X3Y143_SLICE_X3Y143_C5Q;
  assign CLBLM_R_X3Y147_SLICE_X3Y147_A4 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X3Y147_SLICE_X3Y147_A5 = CLBLM_R_X3Y145_SLICE_X3Y145_AQ;
  assign CLBLM_R_X3Y147_SLICE_X3Y147_A6 = 1'b1;
  assign CLBLL_L_X2Y166_SLICE_X1Y166_D1 = 1'b1;
  assign CLBLL_L_X2Y166_SLICE_X1Y166_D2 = 1'b1;
  assign CLBLL_L_X2Y166_SLICE_X1Y166_D3 = 1'b1;
  assign CLBLL_L_X2Y166_SLICE_X1Y166_D4 = 1'b1;
  assign CLBLL_L_X2Y166_SLICE_X1Y166_D5 = 1'b1;
  assign CLBLL_L_X2Y166_SLICE_X1Y166_D6 = 1'b1;
  assign CLBLM_R_X3Y147_SLICE_X3Y147_B4 = CLBLM_R_X3Y145_SLICE_X3Y145_BQ;
  assign CLBLM_R_X3Y147_SLICE_X3Y147_B5 = CLBLM_R_X5Y151_SLICE_X6Y151_C5Q;
  assign CLBLM_R_X3Y147_SLICE_X3Y147_B6 = 1'b1;
  assign CLBLM_R_X3Y147_SLICE_X3Y147_C1 = CLBLL_L_X4Y147_SLICE_X5Y147_C5Q;
  assign CLBLM_R_X3Y147_SLICE_X3Y147_C2 = CLBLM_R_X5Y147_SLICE_X6Y147_CQ;
  assign CLBLM_R_X3Y147_SLICE_X3Y147_C3 = 1'b1;
  assign CLBLM_R_X3Y147_SLICE_X3Y147_C4 = CLBLM_R_X7Y146_SLICE_X8Y146_DQ;
  assign CLBLM_R_X3Y147_SLICE_X3Y147_C5 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X3Y147_SLICE_X3Y147_C6 = 1'b1;
  assign CLBLM_R_X3Y147_SLICE_X3Y147_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X3Y147_SLICE_X3Y147_D1 = 1'b1;
  assign CLBLM_R_X3Y147_SLICE_X3Y147_D2 = CLBLM_R_X5Y146_SLICE_X7Y146_BQ;
  assign CLBLM_R_X3Y147_SLICE_X3Y147_D3 = CLBLL_L_X4Y150_SLICE_X4Y150_DO6;
  assign CLBLM_R_X3Y147_SLICE_X3Y147_D4 = 1'b1;
  assign CLBLM_R_X3Y147_SLICE_X3Y147_D5 = CLBLL_L_X2Y150_SLICE_X1Y150_AQ;
  assign CLBLM_R_X3Y147_SLICE_X3Y147_D6 = CLBLL_L_X4Y146_SLICE_X5Y146_BQ;
  assign CLBLM_L_X10Y148_SLICE_X13Y148_A2 = CLBLM_L_X10Y145_SLICE_X12Y145_AQ;
  assign CLBLM_R_X3Y147_SLICE_X2Y147_A1 = CLBLL_L_X2Y150_SLICE_X1Y150_AQ;
  assign CLBLM_R_X3Y147_SLICE_X2Y147_A2 = CLBLM_R_X3Y152_SLICE_X2Y152_AO6;
  assign CLBLM_R_X3Y147_SLICE_X2Y147_A3 = CLBLM_R_X3Y147_SLICE_X2Y147_AQ;
  assign CLBLM_R_X3Y147_SLICE_X2Y147_A4 = CLBLM_R_X3Y147_SLICE_X2Y147_D5Q;
  assign CLBLM_R_X3Y147_SLICE_X2Y147_A5 = 1'b1;
  assign CLBLM_R_X3Y147_SLICE_X2Y147_A6 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X3Y147_SLICE_X2Y147_B1 = CLBLM_R_X3Y148_SLICE_X2Y148_A5Q;
  assign CLBLM_R_X3Y147_SLICE_X2Y147_B2 = CLBLM_R_X3Y147_SLICE_X2Y147_BQ;
  assign CLBLM_R_X3Y147_SLICE_X2Y147_B3 = CLBLM_R_X3Y147_SLICE_X2Y147_AQ;
  assign CLBLM_R_X3Y147_SLICE_X2Y147_B4 = CLBLL_L_X2Y150_SLICE_X1Y150_AQ;
  assign CLBLM_R_X3Y147_SLICE_X2Y147_B5 = CLBLM_R_X3Y152_SLICE_X2Y152_AO6;
  assign CLBLM_R_X3Y147_SLICE_X2Y147_B6 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign LIOI3_X0Y189_OLOGIC_X0Y190_D1 = CLBLM_L_X10Y154_SLICE_X12Y154_CO5;
  assign CLBLM_R_X3Y147_SLICE_X2Y147_C1 = CLBLL_L_X2Y146_SLICE_X1Y146_AQ;
  assign CLBLM_R_X3Y147_SLICE_X2Y147_C2 = CLBLM_R_X3Y147_SLICE_X2Y147_CQ;
  assign CLBLM_R_X3Y147_SLICE_X2Y147_C3 = CLBLL_L_X4Y143_SLICE_X4Y143_D5Q;
  assign CLBLM_R_X3Y147_SLICE_X2Y147_C4 = CLBLL_L_X4Y149_SLICE_X5Y149_CQ;
  assign CLBLM_R_X3Y147_SLICE_X2Y147_C5 = CLBLM_R_X3Y149_SLICE_X3Y149_DQ;
  assign CLBLM_R_X3Y147_SLICE_X2Y147_C6 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign LIOI3_X0Y189_OLOGIC_X0Y190_T1 = 1'b1;
  assign CLBLM_R_X3Y147_SLICE_X2Y147_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign LIOI3_X0Y127_OLOGIC_X0Y128_D1 = CLBLM_L_X10Y145_SLICE_X12Y145_AQ;
  assign CLBLM_R_X3Y147_SLICE_X2Y147_D1 = CLBLM_R_X7Y152_SLICE_X8Y152_CQ;
  assign CLBLM_R_X3Y147_SLICE_X2Y147_D2 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X3Y147_SLICE_X2Y147_D3 = CLBLM_L_X10Y153_SLICE_X13Y153_CQ;
  assign CLBLM_R_X3Y147_SLICE_X2Y147_D4 = CLBLM_L_X8Y147_SLICE_X10Y147_BQ;
  assign CLBLM_R_X3Y147_SLICE_X2Y147_D5 = CLBLL_L_X4Y142_SLICE_X5Y142_D5Q;
  assign CLBLM_R_X3Y147_SLICE_X2Y147_D6 = 1'b1;
  assign LIOI3_X0Y127_OLOGIC_X0Y128_T1 = 1'b1;
  assign LIOI3_X0Y189_OLOGIC_X0Y189_D1 = CLBLM_L_X8Y147_SLICE_X10Y147_BQ;
  assign RIOI3_X105Y173_OLOGIC_X1Y174_D1 = CLBLM_R_X5Y152_SLICE_X7Y152_DO6;
  assign LIOI3_X0Y189_OLOGIC_X0Y189_T1 = 1'b1;
  assign LIOI3_X0Y127_OLOGIC_X0Y127_D1 = CLBLM_R_X7Y152_SLICE_X8Y152_D5Q;
  assign RIOB33_X105Y181_IOB_X1Y182_O = CLBLM_R_X11Y146_SLICE_X14Y146_BO5;
  assign RIOB33_X105Y181_IOB_X1Y181_O = CLBLM_L_X10Y154_SLICE_X12Y154_CO5;
  assign RIOI3_X105Y173_OLOGIC_X1Y174_T1 = 1'b1;
  assign LIOI3_X0Y127_OLOGIC_X0Y127_T1 = 1'b1;
  assign RIOI3_X105Y173_OLOGIC_X1Y173_D1 = CLBLM_R_X5Y152_SLICE_X7Y152_DQ;
  assign LIOI3_TBYTESRC_X0Y131_OLOGIC_X0Y132_D1 = CLBLM_R_X3Y143_SLICE_X2Y143_BO5;
  assign RIOI3_X105Y173_OLOGIC_X1Y173_T1 = 1'b1;
  assign LIOI3_TBYTESRC_X0Y131_OLOGIC_X0Y132_T1 = 1'b1;
  assign RIOI3_TBYTETERM_X105Y163_OLOGIC_X1Y164_D1 = CLBLM_L_X10Y153_SLICE_X12Y153_AQ;
  assign LIOI3_TBYTESRC_X0Y131_OLOGIC_X0Y131_D1 = CLBLL_L_X2Y75_SLICE_X0Y75_AO6;
  assign RIOI3_TBYTETERM_X105Y163_OLOGIC_X1Y164_T1 = 1'b1;
  assign LIOI3_TBYTESRC_X0Y131_OLOGIC_X0Y131_T1 = 1'b1;
  assign RIOI3_TBYTETERM_X105Y163_OLOGIC_X1Y163_D1 = CLBLM_R_X7Y151_SLICE_X9Y151_D5Q;
  assign RIOI3_TBYTETERM_X105Y163_OLOGIC_X1Y163_T1 = 1'b1;
  assign RIOI3_X105Y111_ILOGIC_X1Y112_D = RIOB33_X105Y111_IOB_X1Y112_I;
  assign CLBLM_R_X3Y148_SLICE_X3Y148_A1 = CLBLM_R_X5Y142_SLICE_X7Y142_BQ;
  assign CLBLM_R_X3Y148_SLICE_X3Y148_A2 = CLBLM_L_X10Y145_SLICE_X12Y145_AQ;
  assign CLBLM_R_X3Y148_SLICE_X3Y148_A3 = CLBLM_R_X3Y148_SLICE_X3Y148_AQ;
  assign CLBLM_R_X3Y148_SLICE_X3Y148_A4 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X3Y148_SLICE_X3Y148_A5 = CLBLM_R_X3Y150_SLICE_X3Y150_A5Q;
  assign CLBLM_R_X3Y148_SLICE_X3Y148_A6 = CLBLM_R_X3Y149_SLICE_X2Y149_CQ;
  assign RIOI3_X105Y111_ILOGIC_X1Y111_D = RIOB33_X105Y111_IOB_X1Y111_I;
  assign CLBLM_R_X3Y148_SLICE_X3Y148_B1 = CLBLL_L_X4Y148_SLICE_X5Y148_A5Q;
  assign CLBLM_R_X3Y148_SLICE_X3Y148_B2 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X3Y148_SLICE_X3Y148_B3 = CLBLL_L_X4Y146_SLICE_X4Y146_C5Q;
  assign CLBLM_R_X3Y148_SLICE_X3Y148_B4 = CLBLM_R_X5Y145_SLICE_X6Y145_C5Q;
  assign CLBLM_R_X3Y148_SLICE_X3Y148_B5 = CLBLM_R_X7Y148_SLICE_X9Y148_AQ;
  assign CLBLM_R_X3Y148_SLICE_X3Y148_B6 = 1'b1;
  assign CLBLM_R_X3Y148_SLICE_X3Y148_C1 = CLBLL_L_X4Y153_SLICE_X4Y153_AQ;
  assign CLBLM_R_X3Y148_SLICE_X3Y148_C2 = CLBLM_L_X12Y146_SLICE_X17Y146_AQ;
  assign CLBLM_R_X3Y148_SLICE_X3Y148_C3 = CLBLM_L_X10Y151_SLICE_X13Y151_A5Q;
  assign CLBLM_R_X3Y148_SLICE_X3Y148_C4 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X3Y148_SLICE_X3Y148_C5 = RIOB33_X105Y101_IOB_X1Y101_I;
  assign CLBLM_R_X3Y148_SLICE_X3Y148_C6 = 1'b1;
  assign CLBLM_R_X3Y148_SLICE_X3Y148_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X11Y153_SLICE_X15Y153_D5 = 1'b1;
  assign CLBLM_R_X3Y148_SLICE_X3Y148_D1 = 1'b1;
  assign CLBLM_R_X3Y148_SLICE_X3Y148_D2 = CLBLM_R_X3Y149_SLICE_X3Y149_CQ;
  assign CLBLM_R_X3Y148_SLICE_X3Y148_D3 = CLBLL_L_X4Y148_SLICE_X4Y148_C5Q;
  assign CLBLM_R_X3Y148_SLICE_X3Y148_D4 = CLBLM_R_X3Y149_SLICE_X2Y149_CQ;
  assign CLBLM_R_X3Y148_SLICE_X3Y148_D5 = CLBLL_L_X4Y152_SLICE_X4Y152_DQ;
  assign CLBLM_R_X3Y148_SLICE_X3Y148_D6 = 1'b1;
  assign CLBLM_R_X3Y148_SLICE_X2Y148_A1 = CLBLM_R_X3Y147_SLICE_X2Y147_DQ;
  assign CLBLM_R_X3Y148_SLICE_X2Y148_A2 = CLBLM_R_X7Y148_SLICE_X9Y148_AQ;
  assign CLBLM_R_X3Y148_SLICE_X2Y148_A3 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X3Y148_SLICE_X2Y148_A4 = CLBLM_R_X3Y151_SLICE_X3Y151_CQ;
  assign CLBLM_R_X3Y148_SLICE_X2Y148_A5 = CLBLM_R_X3Y145_SLICE_X2Y145_AQ;
  assign CLBLM_R_X3Y148_SLICE_X2Y148_A6 = 1'b1;
  assign CLBLM_R_X11Y153_SLICE_X15Y153_D6 = CLBLM_R_X11Y153_SLICE_X15Y153_AQ;
  assign CLBLM_R_X3Y148_SLICE_X2Y148_B1 = CLBLM_R_X3Y148_SLICE_X2Y148_BQ;
  assign CLBLM_R_X3Y148_SLICE_X2Y148_B2 = CLBLM_R_X3Y148_SLICE_X3Y148_B5Q;
  assign CLBLM_R_X3Y148_SLICE_X2Y148_B3 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X3Y148_SLICE_X2Y148_B4 = CLBLM_L_X10Y154_SLICE_X12Y154_B5Q;
  assign CLBLM_R_X3Y148_SLICE_X2Y148_B5 = CLBLM_R_X3Y148_SLICE_X2Y148_CO5;
  assign CLBLM_R_X3Y148_SLICE_X2Y148_B6 = 1'b1;
  assign CLBLM_R_X3Y148_SLICE_X2Y148_C1 = CLBLM_R_X3Y149_SLICE_X2Y149_DQ;
  assign CLBLM_R_X3Y148_SLICE_X2Y148_C2 = 1'b1;
  assign CLBLM_R_X3Y148_SLICE_X2Y148_C3 = CLBLL_L_X2Y146_SLICE_X1Y146_BQ;
  assign CLBLM_R_X3Y148_SLICE_X2Y148_C4 = CLBLL_L_X4Y149_SLICE_X4Y149_D5Q;
  assign CLBLM_R_X3Y148_SLICE_X2Y148_C5 = CLBLL_L_X4Y149_SLICE_X4Y149_DQ;
  assign CLBLM_R_X3Y148_SLICE_X2Y148_C6 = 1'b1;
  assign RIOB33_X105Y183_IOB_X1Y183_O = 1'b0;
  assign RIOB33_X105Y183_IOB_X1Y184_O = CLBLM_R_X3Y148_SLICE_X3Y148_DO5;
  assign CLBLM_R_X3Y148_SLICE_X2Y148_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X3Y148_SLICE_X2Y148_D1 = CLBLM_R_X5Y147_SLICE_X6Y147_CQ;
  assign CLBLM_R_X3Y148_SLICE_X2Y148_D2 = CLBLL_L_X4Y146_SLICE_X4Y146_B5Q;
  assign CLBLM_R_X3Y148_SLICE_X2Y148_D3 = CLBLM_R_X3Y150_SLICE_X3Y150_B5Q;
  assign CLBLM_R_X3Y148_SLICE_X2Y148_D4 = 1'b1;
  assign CLBLM_R_X3Y148_SLICE_X2Y148_D5 = 1'b1;
  assign CLBLM_R_X3Y148_SLICE_X2Y148_D6 = CLBLM_R_X3Y148_SLICE_X2Y148_AQ;
  assign CLBLM_R_X11Y144_SLICE_X14Y144_A6 = CLBLL_L_X4Y147_SLICE_X4Y147_CQ;
  assign CLBLM_R_X3Y149_SLICE_X3Y149_A1 = CLBLL_L_X2Y150_SLICE_X1Y150_AQ;
  assign CLBLM_R_X3Y149_SLICE_X3Y149_A2 = CLBLM_R_X3Y149_SLICE_X3Y149_BQ;
  assign CLBLM_R_X3Y149_SLICE_X3Y149_A3 = CLBLM_R_X3Y149_SLICE_X3Y149_AQ;
  assign CLBLM_R_X3Y149_SLICE_X3Y149_A4 = CLBLM_R_X7Y153_SLICE_X9Y153_AQ;
  assign CLBLM_R_X3Y149_SLICE_X3Y149_A5 = CLBLM_R_X3Y149_SLICE_X2Y149_AQ;
  assign CLBLM_R_X3Y149_SLICE_X3Y149_A6 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign RIOI3_X105Y189_OLOGIC_X1Y190_D1 = CLBLM_L_X12Y151_SLICE_X16Y151_AO5;
  assign CLBLM_R_X3Y149_SLICE_X3Y149_B1 = CLBLM_R_X3Y149_SLICE_X3Y149_CQ;
  assign CLBLM_R_X3Y149_SLICE_X3Y149_B2 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X3Y149_SLICE_X3Y149_B3 = CLBLL_L_X4Y142_SLICE_X5Y142_C5Q;
  assign CLBLM_R_X3Y149_SLICE_X3Y149_B4 = CLBLM_R_X7Y146_SLICE_X8Y146_CQ;
  assign CLBLM_R_X3Y149_SLICE_X3Y149_B5 = 1'b1;
  assign CLBLM_R_X3Y149_SLICE_X3Y149_B6 = CLBLM_R_X3Y147_SLICE_X3Y147_CQ;
  assign CLBLM_R_X3Y149_SLICE_X3Y149_C1 = CLBLM_R_X3Y149_SLICE_X3Y149_BQ;
  assign CLBLM_R_X3Y149_SLICE_X3Y149_C2 = CLBLM_R_X3Y149_SLICE_X3Y149_CQ;
  assign CLBLM_R_X3Y149_SLICE_X3Y149_C3 = CLBLM_R_X7Y146_SLICE_X8Y146_CQ;
  assign CLBLM_R_X3Y149_SLICE_X3Y149_C4 = CLBLM_R_X3Y147_SLICE_X3Y147_CQ;
  assign CLBLM_R_X3Y149_SLICE_X3Y149_C5 = CLBLM_R_X5Y153_SLICE_X6Y153_A5Q;
  assign CLBLM_R_X3Y149_SLICE_X3Y149_C6 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X3Y149_SLICE_X3Y149_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X3Y149_SLICE_X3Y149_D1 = CLBLM_R_X3Y146_SLICE_X2Y146_D5Q;
  assign CLBLM_R_X3Y149_SLICE_X3Y149_D2 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X3Y149_SLICE_X3Y149_D3 = CLBLM_R_X3Y150_SLICE_X3Y150_A5Q;
  assign CLBLM_R_X3Y149_SLICE_X3Y149_D4 = 1'b1;
  assign CLBLM_R_X3Y149_SLICE_X3Y149_D5 = CLBLM_R_X3Y150_SLICE_X2Y150_CQ;
  assign CLBLM_R_X3Y149_SLICE_X3Y149_D6 = 1'b1;
  assign CLBLM_R_X11Y144_SLICE_X14Y144_B3 = CLBLM_R_X5Y142_SLICE_X6Y142_D5Q;
  assign RIOB33_X105Y185_IOB_X1Y186_O = CLBLM_L_X10Y149_SLICE_X13Y149_BO6;
  assign CLBLM_R_X11Y144_SLICE_X14Y144_B4 = CLBLM_R_X7Y151_SLICE_X8Y151_D5Q;
  assign RIOB33_X105Y185_IOB_X1Y185_O = CLBLM_L_X10Y153_SLICE_X12Y153_DO6;
  assign CLBLM_R_X3Y149_SLICE_X2Y149_A1 = CLBLL_L_X2Y150_SLICE_X1Y150_AQ;
  assign CLBLM_R_X3Y149_SLICE_X2Y149_A2 = CLBLM_R_X3Y149_SLICE_X2Y149_DQ;
  assign CLBLM_R_X3Y149_SLICE_X2Y149_A3 = CLBLM_R_X3Y149_SLICE_X2Y149_AQ;
  assign CLBLM_R_X3Y149_SLICE_X2Y149_A4 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X3Y149_SLICE_X2Y149_A5 = CLBLM_R_X7Y153_SLICE_X9Y153_AQ;
  assign CLBLM_R_X3Y149_SLICE_X2Y149_A6 = 1'b1;
  assign CLBLM_R_X11Y144_SLICE_X14Y144_B5 = CLBLM_R_X7Y149_SLICE_X8Y149_AQ;
  assign CLBLM_R_X11Y144_SLICE_X14Y144_B6 = CLBLL_L_X4Y147_SLICE_X4Y147_CQ;
  assign CLBLM_R_X3Y149_SLICE_X2Y149_B1 = CLBLL_L_X4Y149_SLICE_X4Y149_AQ;
  assign CLBLM_R_X3Y149_SLICE_X2Y149_B2 = CLBLM_R_X3Y149_SLICE_X2Y149_BQ;
  assign CLBLM_R_X3Y149_SLICE_X2Y149_B3 = CLBLL_L_X4Y143_SLICE_X4Y143_D5Q;
  assign CLBLM_R_X3Y149_SLICE_X2Y149_B4 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X3Y149_SLICE_X2Y149_B5 = CLBLL_L_X4Y146_SLICE_X4Y146_DO6;
  assign CLBLM_R_X3Y149_SLICE_X2Y149_B6 = CLBLM_R_X3Y150_SLICE_X2Y150_DQ;
  assign RIOI3_X105Y189_OLOGIC_X1Y190_T1 = 1'b1;
  assign CLBLM_R_X3Y149_SLICE_X2Y149_C1 = CLBLM_R_X3Y148_SLICE_X2Y148_BQ;
  assign CLBLM_R_X3Y149_SLICE_X2Y149_C2 = CLBLM_R_X3Y150_SLICE_X2Y150_DQ;
  assign CLBLM_R_X3Y149_SLICE_X2Y149_C3 = CLBLM_R_X3Y148_SLICE_X3Y148_AQ;
  assign CLBLM_R_X3Y149_SLICE_X2Y149_C4 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X3Y149_SLICE_X2Y149_C5 = RIOB33_X105Y121_IOB_X1Y121_I;
  assign CLBLM_R_X3Y149_SLICE_X2Y149_C6 = 1'b1;
  assign CLBLM_R_X3Y149_SLICE_X2Y149_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X3Y149_SLICE_X2Y149_D1 = CLBLM_R_X3Y148_SLICE_X2Y148_BQ;
  assign CLBLM_R_X3Y149_SLICE_X2Y149_D2 = LIOB33_X0Y55_IOB_X0Y55_I;
  assign CLBLM_R_X3Y149_SLICE_X2Y149_D3 = CLBLM_R_X3Y149_SLICE_X2Y149_DQ;
  assign CLBLM_R_X3Y149_SLICE_X2Y149_D4 = CLBLM_R_X3Y148_SLICE_X2Y148_CO6;
  assign CLBLM_R_X3Y149_SLICE_X2Y149_D5 = CLBLM_R_X3Y150_SLICE_X3Y150_DQ;
  assign CLBLM_R_X3Y149_SLICE_X2Y149_D6 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X7Y146_SLICE_X8Y146_A6 = 1'b1;
  assign LIOI3_X0Y191_OLOGIC_X0Y192_D1 = CLBLL_L_X4Y153_SLICE_X4Y153_DO5;
  assign LIOI3_X0Y191_OLOGIC_X0Y192_T1 = 1'b1;
  assign LIOI3_X0Y129_OLOGIC_X0Y130_D1 = CLBLL_L_X2Y145_SLICE_X0Y145_BQ;
  assign LIOI3_X0Y191_OLOGIC_X0Y191_D1 = CLBLL_L_X2Y148_SLICE_X1Y148_CO6;
  assign LIOI3_X0Y129_OLOGIC_X0Y130_T1 = 1'b1;
  assign RIOI3_X105Y175_OLOGIC_X1Y176_D1 = CLBLL_L_X2Y148_SLICE_X1Y148_BO6;
  assign LIOI3_X0Y191_OLOGIC_X0Y191_T1 = 1'b1;
  assign CLBLM_R_X7Y146_SLICE_X8Y146_B3 = CLBLM_R_X5Y154_SLICE_X6Y154_AQ;
  assign LIOI3_X0Y129_OLOGIC_X0Y129_D1 = CLBLL_L_X2Y146_SLICE_X0Y146_CQ;
  assign CLBLM_R_X7Y146_SLICE_X8Y146_B4 = CLBLM_L_X10Y149_SLICE_X13Y149_AQ;
  assign RIOI3_X105Y175_OLOGIC_X1Y176_T1 = 1'b1;
  assign CLBLM_R_X7Y146_SLICE_X8Y146_B5 = 1'b1;
  assign CLBLM_R_X7Y146_SLICE_X8Y146_B6 = 1'b1;
  assign LIOI3_X0Y129_OLOGIC_X0Y129_T1 = 1'b1;
  assign RIOI3_X105Y175_OLOGIC_X1Y175_D1 = CLBLM_L_X10Y144_SLICE_X12Y144_BO6;
  assign LIOI3_TBYTESRC_X0Y143_OLOGIC_X0Y144_D1 = CLBLM_R_X5Y147_SLICE_X7Y147_DO6;
  assign RIOI3_X105Y175_OLOGIC_X1Y175_T1 = 1'b1;
  assign LIOI3_TBYTESRC_X0Y143_OLOGIC_X0Y144_T1 = 1'b1;
  assign CLBLM_R_X11Y151_SLICE_X15Y151_D5 = 1'b1;
  assign RIOI3_TBYTETERM_X105Y187_OLOGIC_X1Y188_D1 = CLBLM_R_X11Y146_SLICE_X14Y146_BO5;
  assign LIOI3_TBYTESRC_X0Y143_OLOGIC_X0Y143_D1 = CLBLM_R_X3Y151_SLICE_X2Y151_BO5;
  assign RIOI3_TBYTETERM_X105Y187_OLOGIC_X1Y188_T1 = 1'b1;
  assign LIOI3_TBYTESRC_X0Y143_OLOGIC_X0Y143_T1 = 1'b1;
  assign RIOI3_TBYTETERM_X105Y187_OLOGIC_X1Y187_D1 = CLBLM_R_X103Y178_SLICE_X163Y178_AO6;
  assign CLBLM_R_X11Y151_SLICE_X15Y151_D6 = 1'b1;
  assign LIOB33_X0Y101_IOB_X0Y102_O = CLBLM_R_X5Y141_SLICE_X6Y141_DQ;
  assign LIOB33_X0Y101_IOB_X0Y101_O = CLBLM_L_X8Y145_SLICE_X11Y145_C5Q;
  assign RIOI3_TBYTETERM_X105Y187_OLOGIC_X1Y187_T1 = 1'b1;
  assign CLBLM_R_X7Y146_SLICE_X8Y146_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X3Y150_SLICE_X3Y150_A1 = CLBLM_R_X3Y143_SLICE_X3Y143_BQ;
  assign CLBLM_R_X3Y150_SLICE_X3Y150_A2 = 1'b1;
  assign CLBLM_R_X3Y150_SLICE_X3Y150_A3 = CLBLM_L_X10Y149_SLICE_X12Y149_BQ;
  assign CLBLM_R_X3Y150_SLICE_X3Y150_A4 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X3Y150_SLICE_X3Y150_A5 = CLBLL_L_X4Y151_SLICE_X4Y151_AQ;
  assign CLBLM_R_X3Y150_SLICE_X3Y150_A6 = 1'b1;
  assign CLBLM_R_X3Y150_SLICE_X3Y150_B1 = CLBLL_L_X4Y151_SLICE_X5Y151_CQ;
  assign CLBLM_R_X3Y150_SLICE_X3Y150_B2 = CLBLM_R_X3Y149_SLICE_X3Y149_D5Q;
  assign CLBLM_R_X3Y150_SLICE_X3Y150_B3 = CLBLM_R_X3Y150_SLICE_X3Y150_CQ;
  assign CLBLM_R_X3Y150_SLICE_X3Y150_B4 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X3Y150_SLICE_X3Y150_B5 = CLBLM_R_X7Y151_SLICE_X9Y151_AQ;
  assign CLBLM_R_X3Y150_SLICE_X3Y150_B6 = 1'b1;
  assign RIOB33_X105Y187_IOB_X1Y187_O = CLBLM_R_X103Y178_SLICE_X163Y178_AO6;
  assign RIOB33_X105Y187_IOB_X1Y188_O = CLBLM_R_X11Y146_SLICE_X14Y146_BO5;
  assign CLBLM_R_X3Y150_SLICE_X3Y150_C1 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X3Y150_SLICE_X3Y150_C2 = CLBLM_R_X3Y150_SLICE_X3Y150_CQ;
  assign CLBLM_R_X3Y150_SLICE_X3Y150_C3 = CLBLM_R_X5Y153_SLICE_X6Y153_D5Q;
  assign CLBLM_R_X3Y150_SLICE_X3Y150_C4 = CLBLM_R_X3Y150_SLICE_X2Y150_CQ;
  assign CLBLM_R_X3Y150_SLICE_X3Y150_C5 = CLBLM_R_X3Y150_SLICE_X2Y150_BQ;
  assign CLBLM_R_X3Y150_SLICE_X3Y150_C6 = CLBLL_L_X4Y150_SLICE_X4Y150_CQ;
  assign CLBLM_R_X3Y150_SLICE_X3Y150_CLK = CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O;
  assign CLBLM_R_X3Y150_SLICE_X3Y150_D1 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X3Y150_SLICE_X3Y150_D2 = CLBLL_L_X4Y152_SLICE_X4Y152_AQ;
  assign CLBLM_R_X3Y150_SLICE_X3Y150_D3 = CLBLM_R_X3Y150_SLICE_X2Y150_D5Q;
  assign CLBLM_R_X3Y150_SLICE_X3Y150_D4 = CLBLM_R_X3Y151_SLICE_X3Y151_BQ;
  assign CLBLM_R_X3Y150_SLICE_X3Y150_D5 = CLBLM_R_X3Y150_SLICE_X3Y150_AQ;
  assign CLBLM_R_X3Y150_SLICE_X3Y150_D6 = 1'b1;
  assign CLBLM_R_X3Y150_SLICE_X2Y150_A1 = CLBLM_R_X5Y142_SLICE_X7Y142_BQ;
  assign CLBLM_R_X3Y150_SLICE_X2Y150_A2 = CLBLL_L_X4Y152_SLICE_X5Y152_AQ;
  assign CLBLM_R_X3Y150_SLICE_X2Y150_A3 = CLBLM_R_X3Y150_SLICE_X2Y150_AQ;
  assign CLBLM_R_X3Y150_SLICE_X2Y150_A4 = CLBLM_R_X3Y150_SLICE_X3Y150_BQ;
  assign CLBLM_R_X3Y150_SLICE_X2Y150_A5 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X3Y150_SLICE_X2Y150_A6 = CLBLM_L_X10Y145_SLICE_X12Y145_AQ;
  assign CLBLM_R_X3Y150_SLICE_X2Y150_B1 = CLBLM_R_X5Y153_SLICE_X6Y153_D5Q;
  assign CLBLM_R_X3Y150_SLICE_X2Y150_B2 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X3Y150_SLICE_X2Y150_B3 = CLBLM_R_X3Y148_SLICE_X2Y148_AQ;
  assign CLBLM_R_X3Y150_SLICE_X2Y150_B4 = CLBLM_R_X3Y150_SLICE_X2Y150_CQ;
  assign CLBLM_R_X3Y150_SLICE_X2Y150_B5 = CLBLM_R_X3Y150_SLICE_X3Y150_CQ;
  assign CLBLM_R_X3Y150_SLICE_X2Y150_B6 = CLBLM_R_X3Y150_SLICE_X2Y150_BQ;
  assign CLBLM_R_X3Y150_SLICE_X2Y150_C1 = CLBLM_R_X3Y150_SLICE_X2Y150_CQ;
  assign CLBLM_R_X3Y150_SLICE_X2Y150_C2 = CLBLL_L_X4Y144_SLICE_X5Y144_CQ;
  assign CLBLM_R_X3Y150_SLICE_X2Y150_C3 = CLBLM_R_X3Y150_SLICE_X2Y150_BQ;
  assign CLBLM_R_X3Y150_SLICE_X2Y150_C4 = CLBLM_R_X3Y150_SLICE_X3Y150_CQ;
  assign CLBLM_R_X3Y150_SLICE_X2Y150_C5 = CLBLM_R_X5Y153_SLICE_X6Y153_D5Q;
  assign CLBLM_R_X3Y150_SLICE_X2Y150_C6 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X3Y150_SLICE_X2Y150_CLK = CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O;
  assign CLBLM_R_X3Y150_SLICE_X2Y150_D1 = CLBLM_R_X3Y152_SLICE_X3Y152_AQ;
  assign CLBLM_R_X3Y150_SLICE_X2Y150_D2 = CLBLM_L_X10Y151_SLICE_X13Y151_AQ;
  assign CLBLM_R_X3Y150_SLICE_X2Y150_D3 = CLBLM_R_X3Y150_SLICE_X3Y150_B5Q;
  assign CLBLM_R_X3Y150_SLICE_X2Y150_D4 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X3Y150_SLICE_X2Y150_D5 = 1'b1;
  assign CLBLM_R_X3Y150_SLICE_X2Y150_D6 = 1'b1;
  assign CLBLM_L_X12Y145_SLICE_X17Y145_A1 = CLBLM_R_X7Y149_SLICE_X8Y149_AQ;
  assign CLBLM_L_X12Y145_SLICE_X17Y145_A2 = CLBLM_R_X7Y153_SLICE_X8Y153_A5Q;
  assign CLBLM_L_X12Y145_SLICE_X17Y145_A3 = CLBLM_R_X7Y144_SLICE_X9Y144_B5Q;
  assign CLBLM_L_X12Y145_SLICE_X17Y145_A4 = CLBLL_L_X4Y148_SLICE_X4Y148_CQ;
  assign CLBLM_L_X12Y145_SLICE_X17Y145_A5 = CLBLM_L_X12Y145_SLICE_X17Y145_DO6;
  assign CLBLM_L_X12Y145_SLICE_X17Y145_A6 = 1'b1;
  assign CLBLM_L_X12Y145_SLICE_X17Y145_B1 = RIOB33_X105Y141_IOB_X1Y142_I;
  assign CLBLM_L_X12Y145_SLICE_X17Y145_B2 = CLBLM_L_X12Y146_SLICE_X16Y146_CQ;
  assign CLBLM_L_X12Y145_SLICE_X17Y145_B3 = RIOB33_X105Y143_IOB_X1Y144_I;
  assign CLBLM_L_X12Y145_SLICE_X17Y145_B4 = RIOB33_X105Y143_IOB_X1Y143_I;
  assign CLBLM_L_X12Y145_SLICE_X17Y145_B5 = CLBLM_R_X5Y148_SLICE_X6Y148_CQ;
  assign CLBLM_L_X12Y145_SLICE_X17Y145_B6 = CLBLM_L_X12Y146_SLICE_X16Y146_AQ;
  assign CLBLM_L_X12Y145_SLICE_X17Y145_C1 = CLBLM_R_X5Y142_SLICE_X6Y142_D5Q;
  assign CLBLM_L_X12Y145_SLICE_X17Y145_C2 = CLBLL_L_X4Y147_SLICE_X4Y147_CQ;
  assign CLBLM_L_X12Y145_SLICE_X17Y145_C3 = CLBLM_R_X7Y149_SLICE_X8Y149_AQ;
  assign CLBLM_L_X12Y145_SLICE_X17Y145_C4 = CLBLM_R_X7Y151_SLICE_X8Y151_D5Q;
  assign CLBLM_L_X12Y145_SLICE_X17Y145_C5 = CLBLM_L_X10Y146_SLICE_X12Y146_DQ;
  assign CLBLM_L_X12Y145_SLICE_X17Y145_C6 = CLBLL_L_X4Y148_SLICE_X4Y148_CQ;
  assign RIOI3_X105Y115_ILOGIC_X1Y116_D = RIOB33_X105Y115_IOB_X1Y116_I;
  assign RIOI3_X105Y115_ILOGIC_X1Y115_D = RIOB33_X105Y115_IOB_X1Y115_I;
  assign CLBLM_L_X12Y145_SLICE_X17Y145_D1 = CLBLM_R_X5Y142_SLICE_X6Y142_D5Q;
  assign CLBLM_L_X12Y145_SLICE_X17Y145_D2 = CLBLL_L_X4Y147_SLICE_X4Y147_CQ;
  assign CLBLM_L_X12Y145_SLICE_X17Y145_D3 = CLBLM_L_X10Y146_SLICE_X12Y146_DQ;
  assign CLBLM_L_X12Y145_SLICE_X17Y145_D4 = CLBLM_R_X7Y151_SLICE_X8Y151_D5Q;
  assign CLBLM_L_X12Y145_SLICE_X17Y145_D5 = 1'b1;
  assign CLBLM_L_X12Y145_SLICE_X17Y145_D6 = 1'b1;
  assign CLBLM_L_X12Y145_SLICE_X16Y145_A1 = RIOB33_X105Y141_IOB_X1Y142_I;
  assign CLBLM_L_X12Y145_SLICE_X16Y145_A2 = CLBLM_R_X7Y144_SLICE_X9Y144_B5Q;
  assign CLBLM_L_X12Y145_SLICE_X16Y145_A3 = CLBLM_L_X12Y145_SLICE_X17Y145_CO6;
  assign CLBLM_L_X12Y145_SLICE_X16Y145_A4 = CLBLM_L_X12Y146_SLICE_X16Y146_CQ;
  assign CLBLM_L_X12Y145_SLICE_X16Y145_A5 = CLBLM_R_X7Y153_SLICE_X8Y153_A5Q;
  assign CLBLM_L_X12Y145_SLICE_X16Y145_A6 = 1'b1;
  assign CLBLM_L_X12Y145_SLICE_X16Y145_AX = CLBLM_R_X11Y145_SLICE_X15Y145_AQ;
  assign CLBLM_L_X12Y145_SLICE_X16Y145_B1 = CLBLM_R_X7Y149_SLICE_X8Y149_AQ;
  assign CLBLM_L_X12Y145_SLICE_X16Y145_B2 = CLBLL_L_X4Y148_SLICE_X4Y148_CQ;
  assign CLBLM_L_X12Y145_SLICE_X16Y145_B3 = CLBLM_L_X12Y145_SLICE_X17Y145_DO6;
  assign CLBLM_L_X12Y145_SLICE_X16Y145_B4 = CLBLM_R_X7Y146_SLICE_X9Y146_CO6;
  assign CLBLM_L_X12Y145_SLICE_X16Y145_B5 = CLBLM_R_X7Y144_SLICE_X9Y144_B5Q;
  assign CLBLM_L_X12Y145_SLICE_X16Y145_B6 = CLBLM_R_X7Y153_SLICE_X8Y153_A5Q;
  assign CLBLM_L_X12Y145_SLICE_X16Y145_C1 = CLBLM_L_X12Y145_SLICE_X16Y145_AO6;
  assign CLBLM_L_X12Y145_SLICE_X16Y145_C2 = CLBLM_L_X12Y145_SLICE_X17Y145_AO5;
  assign CLBLM_L_X12Y145_SLICE_X16Y145_C3 = CLBLM_L_X10Y143_SLICE_X13Y143_AQ;
  assign CLBLM_L_X12Y145_SLICE_X16Y145_C4 = RIOB33_X105Y133_IOB_X1Y134_I;
  assign CLBLM_L_X12Y145_SLICE_X16Y145_C5 = CLBLM_L_X12Y146_SLICE_X16Y146_CO6;
  assign CLBLM_L_X12Y145_SLICE_X16Y145_C6 = 1'b1;
  assign CLBLM_L_X12Y145_SLICE_X16Y145_CE = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_L_X12Y145_SLICE_X16Y145_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X12Y145_SLICE_X16Y145_D1 = CLBLM_R_X7Y147_SLICE_X8Y147_AQ;
  assign CLBLM_L_X12Y145_SLICE_X16Y145_D2 = CLBLM_L_X12Y145_SLICE_X16Y145_AQ;
  assign CLBLM_L_X12Y145_SLICE_X16Y145_D3 = RIOB33_X105Y135_IOB_X1Y136_I;
  assign CLBLM_L_X12Y145_SLICE_X16Y145_D4 = 1'b1;
  assign CLBLM_L_X12Y145_SLICE_X16Y145_D5 = 1'b1;
  assign CLBLM_L_X12Y145_SLICE_X16Y145_D6 = RIOB33_X105Y137_IOB_X1Y137_I;
  assign LIOB33_X0Y141_IOB_X0Y142_O = CLBLL_L_X2Y146_SLICE_X0Y146_CQ;
  assign LIOB33_X0Y141_IOB_X0Y141_O = CLBLL_L_X4Y145_SLICE_X5Y145_CQ;
  assign LIOB33_X0Y103_IOB_X0Y104_O = CLBLM_R_X3Y145_SLICE_X2Y145_C5Q;
  assign LIOB33_X0Y103_IOB_X0Y103_O = CLBLM_R_X5Y145_SLICE_X7Y145_BQ;
  assign RIOB33_X105Y189_IOB_X1Y190_O = CLBLM_L_X12Y151_SLICE_X16Y151_AO5;
  assign RIOB33_X105Y189_IOB_X1Y189_O = CLBLM_R_X103Y178_SLICE_X163Y178_AO6;
  assign CLBLM_R_X3Y151_SLICE_X3Y151_A1 = CLBLM_R_X3Y151_SLICE_X3Y151_CQ;
  assign CLBLM_R_X3Y151_SLICE_X3Y151_A2 = CLBLM_R_X3Y145_SLICE_X2Y145_CQ;
  assign CLBLM_R_X3Y151_SLICE_X3Y151_A3 = CLBLM_R_X3Y151_SLICE_X3Y151_AQ;
  assign CLBLM_R_X3Y151_SLICE_X3Y151_A4 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X3Y151_SLICE_X3Y151_A5 = CLBLL_L_X4Y147_SLICE_X5Y147_DO6;
  assign CLBLM_R_X3Y151_SLICE_X3Y151_A6 = CLBLM_L_X8Y154_SLICE_X10Y154_AQ;
  assign CLBLM_R_X3Y151_SLICE_X3Y151_AX = CLBLM_R_X3Y151_SLICE_X2Y151_BO6;
  assign CLBLM_R_X3Y151_SLICE_X3Y151_B1 = CLBLM_R_X3Y145_SLICE_X2Y145_CQ;
  assign CLBLM_R_X3Y151_SLICE_X3Y151_B2 = CLBLM_R_X3Y151_SLICE_X3Y151_BQ;
  assign CLBLM_R_X3Y151_SLICE_X3Y151_B3 = CLBLM_R_X5Y146_SLICE_X6Y146_BQ;
  assign CLBLM_R_X3Y151_SLICE_X3Y151_B4 = CLBLM_R_X3Y151_SLICE_X3Y151_DO5;
  assign CLBLM_R_X3Y151_SLICE_X3Y151_B5 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X3Y151_SLICE_X3Y151_B6 = CLBLL_L_X4Y147_SLICE_X4Y147_AQ;
  assign CLBLM_R_X3Y151_SLICE_X3Y151_C1 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X3Y151_SLICE_X3Y151_C2 = CLBLM_R_X3Y151_SLICE_X3Y151_CQ;
  assign CLBLM_R_X3Y151_SLICE_X3Y151_C3 = CLBLL_L_X4Y147_SLICE_X5Y147_DO6;
  assign CLBLM_R_X3Y151_SLICE_X3Y151_C4 = CLBLL_L_X4Y152_SLICE_X4Y152_CQ;
  assign CLBLM_R_X3Y151_SLICE_X3Y151_C5 = 1'b1;
  assign CLBLM_R_X3Y151_SLICE_X3Y151_C6 = CLBLM_R_X3Y145_SLICE_X2Y145_CQ;
  assign CLBLM_R_X3Y151_SLICE_X3Y151_CLK = CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O;
  assign CLBLM_R_X3Y151_SLICE_X3Y151_D1 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X3Y151_SLICE_X3Y151_D2 = CLBLM_R_X3Y151_SLICE_X3Y151_CQ;
  assign CLBLM_R_X3Y151_SLICE_X3Y151_D3 = CLBLM_R_X3Y151_SLICE_X3Y151_AQ;
  assign CLBLM_R_X3Y151_SLICE_X3Y151_D4 = CLBLL_L_X4Y147_SLICE_X5Y147_DO6;
  assign CLBLM_R_X3Y151_SLICE_X3Y151_D5 = CLBLM_L_X10Y150_SLICE_X12Y150_AQ;
  assign CLBLM_R_X3Y151_SLICE_X3Y151_D6 = 1'b1;
  assign CLBLM_R_X3Y151_SLICE_X2Y151_A1 = CLBLM_R_X3Y151_SLICE_X3Y151_A5Q;
  assign CLBLM_R_X3Y151_SLICE_X2Y151_A2 = CLBLL_L_X4Y144_SLICE_X4Y144_B5Q;
  assign CLBLM_R_X3Y151_SLICE_X2Y151_A3 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X3Y151_SLICE_X2Y151_A4 = CLBLM_R_X5Y148_SLICE_X6Y148_BQ;
  assign CLBLM_R_X3Y151_SLICE_X2Y151_A5 = 1'b1;
  assign CLBLM_R_X3Y151_SLICE_X2Y151_A6 = 1'b1;
  assign CLBLM_R_X3Y151_SLICE_X2Y151_AX = CLBLL_L_X4Y151_SLICE_X4Y151_DQ;
  assign CLBLM_R_X3Y151_SLICE_X2Y151_B1 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X3Y151_SLICE_X2Y151_B2 = CLBLL_L_X4Y142_SLICE_X4Y142_AQ;
  assign CLBLM_R_X3Y151_SLICE_X2Y151_B3 = CLBLL_L_X4Y151_SLICE_X4Y151_DQ;
  assign CLBLM_R_X3Y151_SLICE_X2Y151_B4 = CLBLM_R_X3Y143_SLICE_X3Y143_BQ;
  assign CLBLM_R_X3Y151_SLICE_X2Y151_B5 = CLBLM_R_X3Y149_SLICE_X2Y149_C5Q;
  assign CLBLM_R_X3Y151_SLICE_X2Y151_B6 = 1'b1;
  assign CLBLM_R_X3Y151_SLICE_X2Y151_C1 = CLBLM_R_X3Y151_SLICE_X3Y151_AQ;
  assign CLBLM_R_X3Y151_SLICE_X2Y151_C2 = CLBLL_L_X4Y147_SLICE_X5Y147_DO6;
  assign CLBLM_R_X3Y151_SLICE_X2Y151_C3 = CLBLM_R_X3Y151_SLICE_X3Y151_CQ;
  assign CLBLM_R_X3Y151_SLICE_X2Y151_C4 = CLBLL_L_X4Y150_SLICE_X4Y150_B5Q;
  assign CLBLM_R_X3Y151_SLICE_X2Y151_C5 = CLBLL_L_X4Y147_SLICE_X4Y147_AQ;
  assign CLBLM_R_X3Y151_SLICE_X2Y151_C6 = CLBLM_R_X3Y151_SLICE_X3Y151_BQ;
  assign CLBLM_R_X3Y151_SLICE_X2Y151_CE = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X3Y151_SLICE_X2Y151_CLK = CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O;
  assign CLBLM_R_X3Y151_SLICE_X2Y151_D1 = 1'b1;
  assign CLBLM_R_X3Y151_SLICE_X2Y151_D2 = 1'b1;
  assign CLBLM_R_X3Y151_SLICE_X2Y151_D3 = 1'b1;
  assign CLBLM_R_X3Y151_SLICE_X2Y151_D4 = 1'b1;
  assign CLBLM_R_X3Y151_SLICE_X2Y151_D5 = 1'b1;
  assign CLBLM_R_X3Y151_SLICE_X2Y151_D6 = 1'b1;
  assign CLBLM_L_X12Y146_SLICE_X17Y146_A1 = CLBLM_R_X11Y150_SLICE_X14Y150_AQ;
  assign CLBLM_L_X12Y146_SLICE_X17Y146_A2 = CLBLM_R_X13Y146_SLICE_X18Y146_CO6;
  assign CLBLM_L_X12Y146_SLICE_X17Y146_A3 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_L_X12Y146_SLICE_X17Y146_A4 = CLBLM_L_X12Y146_SLICE_X17Y146_BO6;
  assign CLBLM_L_X12Y146_SLICE_X17Y146_A5 = CLBLM_R_X7Y145_SLICE_X8Y145_DQ;
  assign CLBLM_L_X12Y146_SLICE_X17Y146_A6 = RIOB33_X105Y139_IOB_X1Y139_I;
  assign CLBLM_L_X12Y146_SLICE_X17Y146_B1 = CLBLM_L_X12Y146_SLICE_X16Y146_DQ;
  assign CLBLM_L_X12Y146_SLICE_X17Y146_B2 = CLBLM_L_X12Y145_SLICE_X16Y145_DO6;
  assign CLBLM_L_X12Y146_SLICE_X17Y146_B3 = CLBLM_L_X12Y145_SLICE_X17Y145_BO6;
  assign CLBLM_L_X12Y146_SLICE_X17Y146_B4 = CLBLM_R_X11Y146_SLICE_X15Y146_AO5;
  assign CLBLM_L_X12Y146_SLICE_X17Y146_B5 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_L_X12Y146_SLICE_X17Y146_B6 = CLBLM_L_X12Y147_SLICE_X17Y147_CO6;
  assign CLBLM_L_X12Y146_SLICE_X17Y146_C1 = CLBLM_R_X13Y146_SLICE_X18Y146_AO6;
  assign CLBLM_L_X12Y146_SLICE_X17Y146_C2 = CLBLM_L_X12Y147_SLICE_X17Y147_AO6;
  assign CLBLM_L_X12Y146_SLICE_X17Y146_C3 = CLBLM_R_X11Y146_SLICE_X14Y146_AQ;
  assign CLBLM_L_X12Y146_SLICE_X17Y146_C4 = CLBLM_L_X10Y147_SLICE_X12Y147_AQ;
  assign CLBLM_L_X12Y146_SLICE_X17Y146_C5 = RIOB33_X105Y139_IOB_X1Y140_I;
  assign CLBLM_L_X12Y146_SLICE_X17Y146_C6 = CLBLM_L_X12Y145_SLICE_X17Y145_AO6;
  assign CLBLM_L_X12Y146_SLICE_X17Y146_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X12Y146_SLICE_X17Y146_D1 = CLBLM_L_X10Y147_SLICE_X13Y147_AQ;
  assign CLBLM_L_X12Y146_SLICE_X17Y146_D2 = CLBLM_L_X12Y147_SLICE_X17Y147_AO6;
  assign CLBLM_L_X12Y146_SLICE_X17Y146_D3 = CLBLM_L_X12Y145_SLICE_X17Y145_AO6;
  assign CLBLM_L_X12Y146_SLICE_X17Y146_D4 = CLBLM_R_X11Y150_SLICE_X14Y150_AQ;
  assign CLBLM_L_X12Y146_SLICE_X17Y146_D5 = RIOB33_X105Y139_IOB_X1Y139_I;
  assign CLBLM_L_X12Y146_SLICE_X17Y146_D6 = CLBLM_R_X13Y146_SLICE_X18Y146_AO6;
  assign CLBLM_L_X12Y146_SLICE_X16Y146_A1 = CLBLM_R_X7Y153_SLICE_X8Y153_A5Q;
  assign CLBLM_L_X12Y146_SLICE_X16Y146_A2 = CLBLM_L_X10Y146_SLICE_X13Y146_DO6;
  assign CLBLM_L_X12Y146_SLICE_X16Y146_A3 = CLBLM_L_X12Y145_SLICE_X17Y145_CO6;
  assign CLBLM_L_X12Y146_SLICE_X16Y146_A4 = CLBLM_R_X7Y144_SLICE_X9Y144_B5Q;
  assign CLBLM_L_X12Y146_SLICE_X16Y146_A5 = RIOB33_X105Y141_IOB_X1Y141_I;
  assign CLBLM_L_X12Y146_SLICE_X16Y146_A6 = 1'b1;
  assign CLBLM_L_X12Y146_SLICE_X16Y146_AX = CLBLM_R_X5Y144_SLICE_X6Y144_CQ;
  assign CLBLM_L_X12Y146_SLICE_X16Y146_B1 = CLBLM_R_X11Y144_SLICE_X14Y144_DO6;
  assign CLBLM_L_X12Y146_SLICE_X16Y146_B2 = CLBLM_L_X12Y145_SLICE_X16Y145_CO6;
  assign CLBLM_L_X12Y146_SLICE_X16Y146_B3 = CLBLM_L_X12Y146_SLICE_X17Y146_CO6;
  assign CLBLM_L_X12Y146_SLICE_X16Y146_B4 = CLBLM_L_X12Y145_SLICE_X16Y145_BO6;
  assign CLBLM_L_X12Y146_SLICE_X16Y146_B5 = CLBLM_R_X13Y146_SLICE_X18Y146_BO6;
  assign CLBLM_L_X12Y146_SLICE_X16Y146_B6 = CLBLM_L_X10Y146_SLICE_X13Y146_CQ;
  assign CLBLM_L_X12Y146_SLICE_X16Y146_BX = CLBLM_L_X12Y146_SLICE_X16Y146_AQ;
  assign CLBLM_L_X12Y146_SLICE_X16Y146_C1 = CLBLM_R_X5Y142_SLICE_X6Y142_D5Q;
  assign CLBLM_L_X12Y146_SLICE_X16Y146_C2 = CLBLL_L_X4Y147_SLICE_X4Y147_CQ;
  assign CLBLM_L_X12Y146_SLICE_X16Y146_C3 = CLBLM_L_X10Y147_SLICE_X12Y147_BO6;
  assign CLBLM_L_X12Y146_SLICE_X16Y146_C4 = CLBLM_L_X10Y146_SLICE_X12Y146_DQ;
  assign CLBLM_L_X12Y146_SLICE_X16Y146_C5 = CLBLM_R_X7Y149_SLICE_X8Y149_AQ;
  assign CLBLM_L_X12Y146_SLICE_X16Y146_C6 = CLBLM_R_X7Y151_SLICE_X8Y151_D5Q;
  assign CLBLM_L_X12Y146_SLICE_X16Y146_CE = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_L_X12Y146_SLICE_X16Y146_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X12Y146_SLICE_X16Y146_CX = CLBLM_L_X8Y152_SLICE_X11Y152_D5Q;
  assign CLBLM_L_X12Y146_SLICE_X16Y146_D1 = CLBLM_L_X12Y145_SLICE_X17Y145_AO5;
  assign CLBLM_L_X12Y146_SLICE_X16Y146_D2 = RIOB33_X105Y147_IOB_X1Y147_I;
  assign CLBLM_L_X12Y146_SLICE_X16Y146_D3 = CLBLM_R_X11Y146_SLICE_X15Y146_CO6;
  assign CLBLM_L_X12Y146_SLICE_X16Y146_D4 = CLBLM_L_X12Y146_SLICE_X16Y146_AO5;
  assign CLBLM_L_X12Y146_SLICE_X16Y146_D5 = CLBLM_R_X11Y146_SLICE_X14Y146_DO6;
  assign CLBLM_L_X12Y146_SLICE_X16Y146_D6 = CLBLM_L_X12Y145_SLICE_X16Y145_BO6;
  assign CLBLM_L_X12Y146_SLICE_X16Y146_DX = CLBLM_L_X12Y146_SLICE_X16Y146_CQ;
  assign LIOB33_X0Y105_IOB_X0Y106_O = CLBLM_R_X3Y146_SLICE_X3Y146_BQ;
  assign LIOB33_X0Y105_IOB_X0Y105_O = CLBLL_L_X4Y150_SLICE_X4Y150_C5Q;
  assign CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_CE = 1'b1;
  assign RIOB33_X105Y191_IOB_X1Y192_O = CLBLM_L_X12Y153_SLICE_X16Y153_AO6;
  assign RIOB33_X105Y191_IOB_X1Y191_O = CLBLM_L_X12Y149_SLICE_X17Y149_AO5;
  assign LIOI3_X0Y195_OLOGIC_X0Y196_D1 = CLBLM_R_X3Y148_SLICE_X3Y148_DO5;
  assign LIOI3_X0Y195_OLOGIC_X0Y196_T1 = 1'b1;
  assign LIOI3_X0Y133_OLOGIC_X0Y134_D1 = CLBLL_L_X2Y145_SLICE_X0Y145_BQ;
  assign CLBLM_R_X3Y152_SLICE_X3Y152_A1 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X3Y152_SLICE_X3Y152_A2 = CLBLL_L_X4Y152_SLICE_X5Y152_A5Q;
  assign CLBLM_R_X3Y152_SLICE_X3Y152_A3 = CLBLM_R_X3Y152_SLICE_X3Y152_AQ;
  assign CLBLM_R_X3Y152_SLICE_X3Y152_A4 = CLBLL_L_X4Y151_SLICE_X5Y151_AQ;
  assign CLBLM_R_X3Y152_SLICE_X3Y152_A5 = CLBLL_L_X2Y150_SLICE_X1Y150_AQ;
  assign CLBLM_R_X3Y152_SLICE_X3Y152_A6 = CLBLL_L_X4Y152_SLICE_X5Y152_DO6;
  assign LIOI3_X0Y133_OLOGIC_X0Y134_T1 = 1'b1;
  assign LIOI3_X0Y195_OLOGIC_X0Y195_D1 = CLBLM_R_X3Y151_SLICE_X2Y151_AO5;
  assign RIOI3_X105Y177_OLOGIC_X1Y178_D1 = CLBLM_R_X5Y147_SLICE_X6Y147_AQ;
  assign CLBLM_R_X3Y152_SLICE_X3Y152_B1 = CLBLM_R_X3Y152_SLICE_X3Y152_DO6;
  assign CLBLM_R_X3Y152_SLICE_X3Y152_B2 = CLBLM_R_X3Y152_SLICE_X3Y152_BQ;
  assign CLBLM_R_X3Y152_SLICE_X3Y152_B3 = CLBLM_R_X3Y152_SLICE_X3Y152_CQ;
  assign CLBLM_R_X3Y152_SLICE_X3Y152_B4 = CLBLM_R_X5Y153_SLICE_X6Y153_D5Q;
  assign CLBLM_R_X3Y152_SLICE_X3Y152_B5 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X3Y152_SLICE_X3Y152_B6 = CLBLL_L_X4Y150_SLICE_X4Y150_AQ;
  assign LIOI3_X0Y133_OLOGIC_X0Y133_D1 = CLBLL_L_X4Y140_SLICE_X4Y140_BO5;
  assign LIOI3_X0Y195_OLOGIC_X0Y195_T1 = 1'b1;
  assign RIOI3_X105Y177_OLOGIC_X1Y178_T1 = 1'b1;
  assign CLBLM_R_X3Y152_SLICE_X3Y152_C1 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X3Y152_SLICE_X3Y152_C2 = CLBLM_R_X3Y152_SLICE_X3Y152_CQ;
  assign CLBLM_R_X3Y152_SLICE_X3Y152_C3 = CLBLM_R_X5Y153_SLICE_X6Y153_D5Q;
  assign CLBLM_R_X3Y152_SLICE_X3Y152_C4 = CLBLM_R_X3Y150_SLICE_X2Y150_CQ;
  assign CLBLM_R_X3Y152_SLICE_X3Y152_C5 = CLBLM_R_X5Y152_SLICE_X7Y152_CQ;
  assign CLBLM_R_X3Y152_SLICE_X3Y152_C6 = CLBLM_R_X3Y150_SLICE_X2Y150_BQ;
  assign CLBLM_R_X3Y152_SLICE_X3Y152_CLK = CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O;
  assign LIOI3_X0Y133_OLOGIC_X0Y133_T1 = 1'b1;
  assign RIOI3_X105Y177_OLOGIC_X1Y177_D1 = CLBLL_L_X2Y146_SLICE_X1Y146_B5Q;
  assign CLBLM_R_X3Y152_SLICE_X3Y152_D1 = CLBLM_R_X3Y150_SLICE_X2Y150_BQ;
  assign CLBLM_R_X3Y152_SLICE_X3Y152_D2 = CLBLM_R_X3Y150_SLICE_X2Y150_CQ;
  assign CLBLM_R_X3Y152_SLICE_X3Y152_D3 = 1'b1;
  assign CLBLM_R_X3Y152_SLICE_X3Y152_D4 = 1'b1;
  assign CLBLM_R_X3Y152_SLICE_X3Y152_D5 = 1'b1;
  assign CLBLM_R_X3Y152_SLICE_X3Y152_D6 = 1'b1;
  assign LIOI3_TBYTESRC_X0Y157_OLOGIC_X0Y158_D1 = RIOB33_X105Y133_IOB_X1Y134_I;
  assign RIOI3_X105Y177_OLOGIC_X1Y177_T1 = 1'b1;
  assign CLBLM_R_X3Y152_SLICE_X2Y152_A1 = CLBLL_L_X4Y152_SLICE_X5Y152_AQ;
  assign CLBLM_R_X3Y152_SLICE_X2Y152_A2 = 1'b1;
  assign CLBLM_R_X3Y152_SLICE_X2Y152_A3 = 1'b1;
  assign CLBLM_R_X3Y152_SLICE_X2Y152_A4 = CLBLL_L_X4Y152_SLICE_X5Y152_DO6;
  assign CLBLM_R_X3Y152_SLICE_X2Y152_A5 = CLBLM_R_X3Y152_SLICE_X3Y152_AQ;
  assign CLBLM_R_X3Y152_SLICE_X2Y152_A6 = CLBLL_L_X4Y152_SLICE_X5Y152_A5Q;
  assign LIOI3_TBYTESRC_X0Y157_OLOGIC_X0Y158_T1 = 1'b1;
  assign CLBLM_R_X3Y152_SLICE_X2Y152_B1 = 1'b1;
  assign CLBLM_R_X3Y152_SLICE_X2Y152_B2 = 1'b1;
  assign CLBLM_R_X3Y152_SLICE_X2Y152_B3 = 1'b1;
  assign CLBLM_R_X3Y152_SLICE_X2Y152_B4 = 1'b1;
  assign CLBLM_R_X3Y152_SLICE_X2Y152_B5 = 1'b1;
  assign CLBLM_R_X3Y152_SLICE_X2Y152_B6 = 1'b1;
  assign LIOI3_TBYTESRC_X0Y157_OLOGIC_X0Y157_D1 = CLBLM_R_X3Y152_SLICE_X3Y152_BQ;
  assign CLBLM_R_X3Y152_SLICE_X2Y152_C1 = 1'b1;
  assign CLBLM_R_X3Y152_SLICE_X2Y152_C2 = 1'b1;
  assign CLBLM_R_X3Y152_SLICE_X2Y152_C3 = 1'b1;
  assign CLBLM_R_X3Y152_SLICE_X2Y152_C4 = 1'b1;
  assign CLBLM_R_X3Y152_SLICE_X2Y152_C5 = 1'b1;
  assign CLBLM_R_X3Y152_SLICE_X2Y152_C6 = 1'b1;
  assign LIOI3_TBYTESRC_X0Y157_OLOGIC_X0Y157_T1 = 1'b1;
  assign CLBLM_R_X3Y152_SLICE_X2Y152_D1 = 1'b1;
  assign CLBLM_R_X3Y152_SLICE_X2Y152_D2 = 1'b1;
  assign CLBLM_R_X3Y152_SLICE_X2Y152_D3 = 1'b1;
  assign CLBLM_R_X3Y152_SLICE_X2Y152_D4 = 1'b1;
  assign CLBLM_R_X3Y152_SLICE_X2Y152_D5 = 1'b1;
  assign CLBLM_R_X3Y152_SLICE_X2Y152_D6 = 1'b1;
  assign CLBLM_L_X12Y147_SLICE_X17Y147_A1 = CLBLM_R_X7Y148_SLICE_X8Y148_AQ;
  assign CLBLM_L_X12Y147_SLICE_X17Y147_A2 = CLBLM_R_X7Y153_SLICE_X8Y153_A5Q;
  assign CLBLM_L_X12Y147_SLICE_X17Y147_A3 = CLBLM_R_X7Y144_SLICE_X9Y144_B5Q;
  assign CLBLM_L_X12Y147_SLICE_X17Y147_A4 = CLBLM_L_X12Y146_SLICE_X16Y146_BQ;
  assign CLBLM_L_X12Y147_SLICE_X17Y147_A5 = CLBLM_L_X12Y145_SLICE_X17Y145_CO6;
  assign CLBLM_L_X12Y147_SLICE_X17Y147_A6 = 1'b1;
  assign CLBLM_L_X12Y147_SLICE_X17Y147_B1 = CLBLM_R_X13Y146_SLICE_X18Y146_AO6;
  assign CLBLM_L_X12Y147_SLICE_X17Y147_B2 = CLBLM_L_X12Y147_SLICE_X16Y147_BO6;
  assign CLBLM_L_X12Y147_SLICE_X17Y147_B3 = CLBLM_L_X12Y145_SLICE_X17Y145_AO5;
  assign CLBLM_L_X12Y147_SLICE_X17Y147_B4 = RIOB33_SING_X105Y149_IOB_X1Y149_I;
  assign CLBLM_L_X12Y147_SLICE_X17Y147_B5 = RIOB33_X105Y137_IOB_X1Y138_I;
  assign CLBLM_L_X12Y147_SLICE_X17Y147_B6 = CLBLM_L_X12Y147_SLICE_X17Y147_AO5;
  assign CLBLM_L_X12Y147_SLICE_X17Y147_C1 = CLBLM_L_X8Y149_SLICE_X10Y149_AQ;
  assign CLBLM_L_X12Y147_SLICE_X17Y147_C2 = 1'b1;
  assign CLBLM_L_X12Y147_SLICE_X17Y147_C3 = CLBLM_R_X7Y148_SLICE_X8Y148_AQ;
  assign CLBLM_L_X12Y147_SLICE_X17Y147_C4 = 1'b1;
  assign CLBLM_L_X12Y147_SLICE_X17Y147_C5 = RIOB33_X105Y135_IOB_X1Y135_I;
  assign CLBLM_L_X12Y147_SLICE_X17Y147_C6 = RIOB33_X105Y137_IOB_X1Y138_I;
  assign CLBLM_L_X12Y147_SLICE_X17Y147_D1 = CLBLM_L_X12Y145_SLICE_X17Y145_AO5;
  assign CLBLM_L_X12Y147_SLICE_X17Y147_D2 = 1'b1;
  assign CLBLM_L_X12Y147_SLICE_X17Y147_D3 = CLBLM_R_X13Y146_SLICE_X18Y146_AO6;
  assign CLBLM_L_X12Y147_SLICE_X17Y147_D4 = 1'b1;
  assign CLBLM_L_X12Y147_SLICE_X17Y147_D5 = RIOB33_SING_X105Y149_IOB_X1Y149_I;
  assign CLBLM_L_X12Y147_SLICE_X17Y147_D6 = RIOB33_X105Y137_IOB_X1Y138_I;
  assign CLBLM_L_X12Y147_SLICE_X16Y147_A1 = CLBLM_R_X7Y153_SLICE_X8Y153_A5Q;
  assign CLBLM_L_X12Y147_SLICE_X16Y147_A2 = CLBLM_L_X8Y149_SLICE_X10Y149_AQ;
  assign CLBLM_L_X12Y147_SLICE_X16Y147_A3 = CLBLM_L_X12Y145_SLICE_X17Y145_CO6;
  assign CLBLM_L_X12Y147_SLICE_X16Y147_A4 = CLBLM_R_X7Y144_SLICE_X9Y144_B5Q;
  assign CLBLM_L_X12Y147_SLICE_X16Y147_A5 = RIOB33_X105Y135_IOB_X1Y135_I;
  assign CLBLM_L_X12Y147_SLICE_X16Y147_A6 = 1'b1;
  assign CLBLM_L_X12Y147_SLICE_X16Y147_B1 = RIOB33_X105Y145_IOB_X1Y145_I;
  assign CLBLM_L_X12Y147_SLICE_X16Y147_B2 = CLBLM_R_X11Y147_SLICE_X14Y147_AO5;
  assign CLBLM_L_X12Y147_SLICE_X16Y147_B3 = CLBLM_L_X8Y147_SLICE_X11Y147_AQ;
  assign CLBLM_L_X12Y147_SLICE_X16Y147_B4 = CLBLM_R_X7Y146_SLICE_X9Y146_CO6;
  assign CLBLM_L_X12Y147_SLICE_X16Y147_B5 = CLBLM_L_X12Y145_SLICE_X17Y145_CO6;
  assign CLBLM_L_X12Y147_SLICE_X16Y147_B6 = CLBLM_L_X12Y147_SLICE_X16Y147_AO5;
  assign CLBLM_L_X12Y147_SLICE_X16Y147_C1 = CLBLM_L_X8Y147_SLICE_X11Y147_AQ;
  assign CLBLM_L_X12Y147_SLICE_X16Y147_C2 = CLBLM_L_X12Y147_SLICE_X17Y147_AO5;
  assign CLBLM_L_X12Y147_SLICE_X16Y147_C3 = RIOB33_X105Y145_IOB_X1Y145_I;
  assign CLBLM_L_X12Y147_SLICE_X16Y147_C4 = CLBLM_L_X12Y146_SLICE_X16Y146_CO6;
  assign CLBLM_L_X12Y147_SLICE_X16Y147_C5 = 1'b1;
  assign CLBLM_L_X12Y147_SLICE_X16Y147_C6 = CLBLM_L_X12Y148_SLICE_X16Y148_AO6;
  assign CLBLM_L_X12Y147_SLICE_X16Y147_D1 = 1'b1;
  assign CLBLM_L_X12Y147_SLICE_X16Y147_D2 = CLBLM_R_X7Y151_SLICE_X8Y151_D5Q;
  assign CLBLM_L_X12Y147_SLICE_X16Y147_D3 = CLBLM_L_X10Y146_SLICE_X12Y146_DQ;
  assign CLBLM_L_X12Y147_SLICE_X16Y147_D4 = CLBLL_L_X4Y147_SLICE_X4Y147_CQ;
  assign CLBLM_L_X12Y147_SLICE_X16Y147_D5 = 1'b1;
  assign CLBLM_L_X12Y147_SLICE_X16Y147_D6 = CLBLM_R_X5Y142_SLICE_X6Y142_D5Q;
  assign LIOB33_X0Y107_IOB_X0Y108_O = CLBLL_L_X4Y143_SLICE_X4Y143_DQ;
  assign LIOB33_X0Y107_IOB_X0Y107_O = CLBLM_R_X7Y146_SLICE_X8Y146_DQ;
  assign RIOI3_X105Y117_ILOGIC_X1Y118_D = RIOB33_X105Y117_IOB_X1Y118_I;
  assign RIOI3_X105Y117_ILOGIC_X1Y117_D = RIOB33_X105Y117_IOB_X1Y117_I;
  assign RIOB33_X105Y193_IOB_X1Y194_O = CLBLM_L_X12Y151_SLICE_X16Y151_BO6;
  assign RIOB33_X105Y193_IOB_X1Y193_O = CLBLM_L_X12Y151_SLICE_X16Y151_BO5;
  assign CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_I = CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_O;
  assign CLBLM_R_X3Y153_SLICE_X3Y153_A1 = 1'b1;
  assign CLBLM_R_X3Y153_SLICE_X3Y153_A2 = 1'b1;
  assign CLBLM_R_X3Y153_SLICE_X3Y153_A3 = 1'b1;
  assign CLBLM_R_X3Y153_SLICE_X3Y153_A4 = 1'b1;
  assign CLBLM_R_X3Y153_SLICE_X3Y153_A5 = 1'b1;
  assign CLBLM_R_X3Y153_SLICE_X3Y153_A6 = 1'b1;
  assign CLBLM_R_X3Y153_SLICE_X3Y153_B1 = 1'b1;
  assign CLBLM_R_X3Y153_SLICE_X3Y153_B2 = 1'b1;
  assign CLBLM_R_X3Y153_SLICE_X3Y153_B3 = 1'b1;
  assign CLBLM_R_X3Y153_SLICE_X3Y153_B4 = 1'b1;
  assign CLBLM_R_X3Y153_SLICE_X3Y153_B5 = 1'b1;
  assign CLBLM_R_X3Y153_SLICE_X3Y153_B6 = 1'b1;
  assign CLBLM_R_X3Y153_SLICE_X3Y153_C1 = 1'b1;
  assign CLBLM_R_X3Y153_SLICE_X3Y153_C2 = 1'b1;
  assign CLBLM_R_X3Y153_SLICE_X3Y153_C3 = 1'b1;
  assign CLBLM_R_X3Y153_SLICE_X3Y153_C4 = 1'b1;
  assign CLBLM_R_X3Y153_SLICE_X3Y153_C5 = 1'b1;
  assign CLBLM_R_X3Y153_SLICE_X3Y153_C6 = 1'b1;
  assign CLBLM_R_X3Y153_SLICE_X3Y153_D1 = 1'b1;
  assign CLBLM_R_X3Y153_SLICE_X3Y153_D2 = 1'b1;
  assign CLBLM_R_X3Y153_SLICE_X3Y153_D3 = 1'b1;
  assign CLBLM_R_X3Y153_SLICE_X3Y153_D4 = 1'b1;
  assign CLBLM_R_X3Y153_SLICE_X3Y153_D5 = 1'b1;
  assign CLBLM_R_X3Y153_SLICE_X3Y153_D6 = 1'b1;
  assign LIOI3_X0Y155_OLOGIC_X0Y155_D1 = CLBLM_R_X5Y154_SLICE_X7Y154_AQ;
  assign CLBLM_R_X3Y153_SLICE_X2Y153_A1 = 1'b1;
  assign CLBLM_R_X3Y153_SLICE_X2Y153_A2 = 1'b1;
  assign CLBLM_R_X3Y153_SLICE_X2Y153_A3 = 1'b1;
  assign CLBLM_R_X3Y153_SLICE_X2Y153_A4 = 1'b1;
  assign CLBLM_R_X3Y153_SLICE_X2Y153_A5 = 1'b1;
  assign CLBLM_R_X3Y153_SLICE_X2Y153_A6 = 1'b1;
  assign CLBLM_R_X3Y153_SLICE_X2Y153_AX = CLBLM_R_X3Y151_SLICE_X2Y151_AO6;
  assign CLBLM_R_X3Y153_SLICE_X2Y153_B1 = 1'b1;
  assign CLBLM_R_X3Y153_SLICE_X2Y153_B2 = 1'b1;
  assign CLBLM_R_X3Y153_SLICE_X2Y153_B3 = 1'b1;
  assign CLBLM_R_X3Y153_SLICE_X2Y153_B4 = 1'b1;
  assign CLBLM_R_X3Y153_SLICE_X2Y153_B5 = 1'b1;
  assign CLBLM_R_X3Y153_SLICE_X2Y153_B6 = 1'b1;
  assign CLBLM_R_X3Y153_SLICE_X2Y153_C1 = 1'b1;
  assign CLBLM_R_X3Y153_SLICE_X2Y153_C2 = 1'b1;
  assign CLBLM_R_X3Y153_SLICE_X2Y153_C3 = 1'b1;
  assign CLBLM_R_X3Y153_SLICE_X2Y153_C4 = 1'b1;
  assign CLBLM_R_X3Y153_SLICE_X2Y153_C5 = 1'b1;
  assign CLBLM_R_X3Y153_SLICE_X2Y153_C6 = 1'b1;
  assign CLBLM_R_X3Y153_SLICE_X2Y153_CLK = CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O;
  assign CLBLM_R_X3Y153_SLICE_X2Y153_D1 = 1'b1;
  assign CLBLM_R_X3Y153_SLICE_X2Y153_D2 = 1'b1;
  assign CLBLM_R_X3Y153_SLICE_X2Y153_D3 = 1'b1;
  assign CLBLM_R_X3Y153_SLICE_X2Y153_D4 = 1'b1;
  assign CLBLM_R_X3Y153_SLICE_X2Y153_D5 = 1'b1;
  assign CLBLM_R_X3Y153_SLICE_X2Y153_D6 = 1'b1;
  assign CLBLM_L_X12Y148_SLICE_X17Y148_A1 = CLBLM_L_X12Y145_SLICE_X17Y145_AO5;
  assign CLBLM_L_X12Y148_SLICE_X17Y148_A2 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_L_X12Y148_SLICE_X17Y148_A3 = CLBLM_R_X7Y144_SLICE_X9Y144_B5Q;
  assign CLBLM_L_X12Y148_SLICE_X17Y148_A4 = RIOB33_X105Y147_IOB_X1Y148_I;
  assign CLBLM_L_X12Y148_SLICE_X17Y148_A5 = CLBLM_L_X12Y145_SLICE_X17Y145_CO6;
  assign CLBLM_L_X12Y148_SLICE_X17Y148_A6 = CLBLM_R_X7Y153_SLICE_X8Y153_A5Q;
  assign CLBLM_L_X12Y148_SLICE_X17Y148_B1 = 1'b1;
  assign CLBLM_L_X12Y148_SLICE_X17Y148_B2 = 1'b1;
  assign CLBLM_L_X12Y148_SLICE_X17Y148_B3 = 1'b1;
  assign CLBLM_L_X12Y148_SLICE_X17Y148_B4 = 1'b1;
  assign CLBLM_L_X12Y148_SLICE_X17Y148_B5 = 1'b1;
  assign CLBLM_L_X12Y148_SLICE_X17Y148_B6 = 1'b1;
  assign CLBLM_R_X7Y155_SLICE_X8Y155_C4 = 1'b1;
  assign CLBLM_L_X12Y148_SLICE_X17Y148_C1 = 1'b1;
  assign CLBLM_L_X12Y148_SLICE_X17Y148_C2 = 1'b1;
  assign CLBLM_L_X12Y148_SLICE_X17Y148_C3 = 1'b1;
  assign CLBLM_L_X12Y148_SLICE_X17Y148_C4 = 1'b1;
  assign CLBLM_L_X12Y148_SLICE_X17Y148_C5 = 1'b1;
  assign CLBLM_L_X12Y148_SLICE_X17Y148_C6 = 1'b1;
  assign CLBLM_L_X12Y148_SLICE_X17Y148_D1 = 1'b1;
  assign CLBLM_L_X12Y148_SLICE_X17Y148_D2 = 1'b1;
  assign CLBLM_L_X12Y148_SLICE_X17Y148_D3 = 1'b1;
  assign CLBLM_L_X12Y148_SLICE_X17Y148_D4 = 1'b1;
  assign CLBLM_L_X12Y148_SLICE_X17Y148_D5 = 1'b1;
  assign CLBLM_L_X12Y148_SLICE_X17Y148_D6 = 1'b1;
  assign CLBLM_R_X7Y155_SLICE_X8Y155_C5 = 1'b1;
  assign CLBLM_L_X12Y148_SLICE_X16Y148_A1 = CLBLM_L_X12Y146_SLICE_X16Y146_DQ;
  assign CLBLM_L_X12Y148_SLICE_X16Y148_A2 = CLBLM_R_X7Y153_SLICE_X8Y153_A5Q;
  assign CLBLM_L_X12Y148_SLICE_X16Y148_A3 = CLBLM_L_X12Y145_SLICE_X17Y145_CO6;
  assign CLBLM_L_X12Y148_SLICE_X16Y148_A4 = CLBLM_R_X7Y144_SLICE_X9Y144_B5Q;
  assign CLBLM_L_X12Y148_SLICE_X16Y148_A5 = CLBLM_R_X7Y147_SLICE_X8Y147_AQ;
  assign CLBLM_L_X12Y148_SLICE_X16Y148_A6 = 1'b1;
  assign CLBLM_L_X12Y148_SLICE_X16Y148_B1 = CLBLM_L_X12Y148_SLICE_X16Y148_CO6;
  assign CLBLM_L_X12Y148_SLICE_X16Y148_B2 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_L_X12Y148_SLICE_X16Y148_B3 = RIOB33_X105Y147_IOB_X1Y148_I;
  assign CLBLM_L_X12Y148_SLICE_X16Y148_B4 = CLBLM_L_X12Y145_SLICE_X17Y145_AO5;
  assign CLBLM_L_X12Y148_SLICE_X16Y148_B5 = CLBLM_L_X12Y148_SLICE_X16Y148_AO6;
  assign CLBLM_L_X12Y148_SLICE_X16Y148_B6 = CLBLM_L_X12Y148_SLICE_X16Y148_AO5;
  assign CLBLM_R_X7Y155_SLICE_X8Y155_C6 = 1'b1;
  assign CLBLM_L_X12Y148_SLICE_X16Y148_C1 = CLBLM_L_X12Y145_SLICE_X17Y145_CO6;
  assign CLBLM_L_X12Y148_SLICE_X16Y148_C2 = CLBLM_L_X10Y147_SLICE_X12Y147_BO6;
  assign CLBLM_L_X12Y148_SLICE_X16Y148_C3 = CLBLM_R_X7Y149_SLICE_X8Y149_AQ;
  assign CLBLM_L_X12Y148_SLICE_X16Y148_C4 = RIOB33_X105Y137_IOB_X1Y137_I;
  assign CLBLM_L_X12Y148_SLICE_X16Y148_C5 = CLBLM_R_X7Y146_SLICE_X9Y146_CO6;
  assign CLBLM_L_X12Y148_SLICE_X16Y148_C6 = CLBLM_R_X5Y144_SLICE_X7Y144_AQ;
  assign LIOB33_X0Y109_IOB_X0Y109_O = CLBLM_R_X5Y141_SLICE_X6Y141_BQ;
  assign LIOB33_X0Y109_IOB_X0Y110_O = CLBLM_R_X5Y145_SLICE_X7Y145_AQ;
  assign CLBLM_L_X12Y148_SLICE_X16Y148_D1 = CLBLM_R_X13Y146_SLICE_X18Y146_AO6;
  assign CLBLM_L_X12Y148_SLICE_X16Y148_D2 = CLBLM_L_X12Y146_SLICE_X16Y146_CO6;
  assign CLBLM_L_X12Y148_SLICE_X16Y148_D3 = 1'b1;
  assign CLBLM_L_X12Y148_SLICE_X16Y148_D4 = CLBLM_L_X12Y148_SLICE_X16Y148_AO5;
  assign CLBLM_L_X12Y148_SLICE_X16Y148_D5 = CLBLM_R_X5Y144_SLICE_X7Y144_AQ;
  assign CLBLM_L_X12Y148_SLICE_X16Y148_D6 = RIOB33_X105Y137_IOB_X1Y137_I;
  assign RIOB33_X105Y195_IOB_X1Y196_O = CLBLM_L_X12Y150_SLICE_X16Y150_AO6;
  assign RIOB33_X105Y195_IOB_X1Y195_O = CLBLM_L_X10Y149_SLICE_X13Y149_AO5;
  assign CLBLM_R_X11Y145_SLICE_X14Y145_A4 = RIOB33_X105Y143_IOB_X1Y144_I;
  assign CLBLM_R_X11Y145_SLICE_X14Y145_B1 = CLBLM_L_X12Y145_SLICE_X17Y145_CO6;
  assign CLBLM_R_X11Y145_SLICE_X14Y145_B2 = CLBLM_L_X12Y145_SLICE_X17Y145_DO6;
  assign CLBLM_R_X11Y145_SLICE_X14Y145_B3 = CLBLM_L_X10Y147_SLICE_X12Y147_BO6;
  assign CLBLM_R_X11Y145_SLICE_X14Y145_B6 = CLBLM_R_X11Y146_SLICE_X14Y146_CO5;
  assign LIOI3_X0Y197_OLOGIC_X0Y198_D1 = 1'b1;
  assign CLBLM_L_X12Y149_SLICE_X17Y149_A1 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_L_X12Y149_SLICE_X17Y149_A2 = CLBLM_R_X11Y149_SLICE_X15Y149_AO6;
  assign CLBLM_L_X12Y149_SLICE_X17Y149_A3 = CLBLM_L_X10Y148_SLICE_X12Y148_AQ;
  assign CLBLM_L_X12Y149_SLICE_X17Y149_A4 = 1'b1;
  assign CLBLM_L_X12Y149_SLICE_X17Y149_A5 = CLBLM_L_X10Y148_SLICE_X13Y148_BQ;
  assign CLBLM_L_X12Y149_SLICE_X17Y149_A6 = 1'b1;
  assign LIOI3_X0Y197_OLOGIC_X0Y198_T1 = 1'b1;
  assign CLBLM_L_X12Y149_SLICE_X17Y149_B1 = CLBLM_R_X7Y149_SLICE_X8Y149_AQ;
  assign CLBLM_L_X12Y149_SLICE_X17Y149_B2 = CLBLL_L_X4Y148_SLICE_X4Y148_CQ;
  assign CLBLM_L_X12Y149_SLICE_X17Y149_B3 = CLBLM_R_X7Y153_SLICE_X8Y153_A5Q;
  assign CLBLM_L_X12Y149_SLICE_X17Y149_B4 = CLBLM_L_X12Y147_SLICE_X16Y147_DO6;
  assign CLBLM_L_X12Y149_SLICE_X17Y149_B5 = CLBLM_R_X7Y144_SLICE_X9Y144_B5Q;
  assign CLBLM_L_X12Y149_SLICE_X17Y149_B6 = 1'b1;
  assign LIOI3_X0Y135_OLOGIC_X0Y136_D1 = CLBLM_L_X10Y153_SLICE_X13Y153_CQ;
  assign CLBLM_L_X12Y149_SLICE_X17Y149_C1 = CLBLM_L_X12Y147_SLICE_X16Y147_DO6;
  assign CLBLM_L_X12Y149_SLICE_X17Y149_C2 = CLBLL_L_X4Y148_SLICE_X4Y148_CQ;
  assign CLBLM_L_X12Y149_SLICE_X17Y149_C3 = CLBLM_R_X7Y149_SLICE_X8Y149_AQ;
  assign CLBLM_L_X12Y149_SLICE_X17Y149_C4 = CLBLM_R_X7Y153_SLICE_X8Y153_A5Q;
  assign CLBLM_L_X12Y149_SLICE_X17Y149_C5 = CLBLM_L_X10Y146_SLICE_X13Y146_DO6;
  assign CLBLM_L_X12Y149_SLICE_X17Y149_C6 = CLBLM_R_X7Y144_SLICE_X9Y144_B5Q;
  assign CLBLM_R_X11Y145_SLICE_X14Y145_C5 = CLBLM_L_X12Y145_SLICE_X17Y145_DO6;
  assign CLBLM_R_X11Y145_SLICE_X14Y145_C6 = CLBLM_R_X11Y146_SLICE_X14Y146_CO5;
  assign LIOI3_X0Y135_OLOGIC_X0Y136_T1 = 1'b1;
  assign LIOI3_X0Y197_OLOGIC_X0Y197_D1 = CLBLL_L_X4Y153_SLICE_X4Y153_CO5;
  assign RIOI3_X105Y179_OLOGIC_X1Y180_D1 = CLBLM_L_X8Y145_SLICE_X11Y145_DQ;
  assign LIOI3_X0Y197_OLOGIC_X0Y197_T1 = 1'b1;
  assign CLBLM_L_X12Y149_SLICE_X17Y149_D1 = CLBLM_L_X8Y152_SLICE_X11Y152_CQ;
  assign CLBLM_L_X12Y149_SLICE_X17Y149_D2 = 1'b1;
  assign CLBLM_L_X12Y149_SLICE_X17Y149_D3 = CLBLM_L_X10Y146_SLICE_X12Y146_AQ;
  assign CLBLM_L_X12Y149_SLICE_X17Y149_D4 = CLBLM_L_X10Y146_SLICE_X13Y146_DO6;
  assign CLBLM_L_X12Y149_SLICE_X17Y149_D5 = CLBLM_L_X12Y149_SLICE_X17Y149_BO5;
  assign CLBLM_L_X12Y149_SLICE_X17Y149_D6 = CLBLM_L_X12Y149_SLICE_X17Y149_BO6;
  assign LIOB33_X0Y111_IOB_X0Y111_O = CLBLM_R_X3Y145_SLICE_X2Y145_B5Q;
  assign LIOB33_X0Y111_IOB_X0Y112_O = CLBLL_L_X4Y146_SLICE_X4Y146_C5Q;
  assign LIOI3_X0Y135_OLOGIC_X0Y135_D1 = CLBLL_L_X2Y145_SLICE_X0Y145_BQ;
  assign RIOI3_X105Y179_OLOGIC_X1Y180_T1 = 1'b1;
  assign CLBLM_L_X12Y149_SLICE_X16Y149_A1 = CLBLM_L_X12Y147_SLICE_X16Y147_DO6;
  assign CLBLM_L_X12Y149_SLICE_X16Y149_A2 = CLBLM_R_X11Y150_SLICE_X14Y150_BO6;
  assign CLBLM_L_X12Y149_SLICE_X16Y149_A3 = CLBLM_L_X12Y146_SLICE_X16Y146_BO6;
  assign CLBLM_L_X12Y149_SLICE_X16Y149_A4 = CLBLM_L_X12Y149_SLICE_X16Y149_BO6;
  assign CLBLM_L_X12Y149_SLICE_X16Y149_A5 = CLBLM_L_X8Y145_SLICE_X10Y145_BO6;
  assign CLBLM_L_X12Y149_SLICE_X16Y149_A6 = CLBLM_R_X7Y148_SLICE_X8Y148_CO6;
  assign LIOI3_X0Y135_OLOGIC_X0Y135_T1 = 1'b1;
  assign RIOI3_X105Y179_OLOGIC_X1Y179_D1 = CLBLM_L_X8Y147_SLICE_X10Y147_BQ;
  assign CLBLM_L_X12Y149_SLICE_X16Y149_B1 = CLBLL_L_X4Y144_SLICE_X4Y144_D5Q;
  assign CLBLM_L_X12Y149_SLICE_X16Y149_B2 = CLBLM_R_X7Y144_SLICE_X9Y144_B5Q;
  assign CLBLM_L_X12Y149_SLICE_X16Y149_B3 = CLBLM_R_X7Y149_SLICE_X9Y149_BQ;
  assign CLBLM_L_X12Y149_SLICE_X16Y149_B4 = CLBLM_L_X8Y149_SLICE_X10Y149_AO6;
  assign CLBLM_L_X12Y149_SLICE_X16Y149_B5 = CLBLM_R_X7Y153_SLICE_X8Y153_A5Q;
  assign CLBLM_L_X12Y149_SLICE_X16Y149_B6 = CLBLM_R_X11Y144_SLICE_X14Y144_AO6;
  assign LIOI3_TBYTESRC_X0Y169_OLOGIC_X0Y170_D1 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign RIOI3_X105Y179_OLOGIC_X1Y179_T1 = 1'b1;
  assign CLBLM_L_X12Y149_SLICE_X16Y149_C1 = CLBLM_L_X12Y146_SLICE_X16Y146_BO6;
  assign CLBLM_L_X12Y149_SLICE_X16Y149_C2 = CLBLM_L_X12Y147_SLICE_X16Y147_DO6;
  assign CLBLM_L_X12Y149_SLICE_X16Y149_C3 = CLBLM_R_X11Y149_SLICE_X14Y149_DO6;
  assign CLBLM_L_X12Y149_SLICE_X16Y149_C4 = CLBLM_R_X11Y149_SLICE_X15Y149_DO6;
  assign CLBLM_L_X12Y149_SLICE_X16Y149_C5 = CLBLM_R_X11Y147_SLICE_X14Y147_DO6;
  assign CLBLM_L_X12Y149_SLICE_X16Y149_C6 = CLBLM_L_X8Y145_SLICE_X10Y145_BO6;
  assign LIOI3_TBYTESRC_X0Y169_OLOGIC_X0Y170_T1 = 1'b1;
  assign RIOB33_X105Y197_IOB_X1Y198_O = CLBLM_L_X12Y150_SLICE_X16Y150_AO5;
  assign RIOB33_X105Y197_IOB_X1Y197_O = CLBLM_L_X12Y152_SLICE_X16Y152_AO5;
  assign CLBLM_R_X7Y147_SLICE_X8Y147_A4 = CLBLM_L_X8Y153_SLICE_X10Y153_C5Q;
  assign LIOI3_TBYTESRC_X0Y169_OLOGIC_X0Y169_D1 = RIOB33_X105Y117_IOB_X1Y117_I;
  assign CLBLM_L_X12Y149_SLICE_X16Y149_D1 = CLBLM_R_X7Y149_SLICE_X9Y149_BQ;
  assign CLBLM_L_X12Y149_SLICE_X16Y149_D2 = 1'b1;
  assign CLBLM_L_X12Y149_SLICE_X16Y149_D3 = CLBLM_R_X11Y144_SLICE_X14Y144_AO6;
  assign CLBLM_L_X12Y149_SLICE_X16Y149_D4 = CLBLM_R_X7Y153_SLICE_X8Y153_A5Q;
  assign CLBLM_L_X12Y149_SLICE_X16Y149_D5 = CLBLL_L_X4Y144_SLICE_X4Y144_D5Q;
  assign CLBLM_L_X12Y149_SLICE_X16Y149_D6 = CLBLM_R_X7Y144_SLICE_X9Y144_B5Q;
  assign LIOI3_TBYTESRC_X0Y169_OLOGIC_X0Y169_T1 = 1'b1;
  assign CLBLM_R_X7Y147_SLICE_X8Y147_AX = CLBLL_L_X2Y150_SLICE_X1Y150_AQ;
  assign CLBLM_R_X7Y147_SLICE_X8Y147_B1 = CLBLL_L_X4Y144_SLICE_X4Y144_AQ;
  assign CLBLM_R_X7Y147_SLICE_X8Y147_B2 = CLBLM_L_X10Y146_SLICE_X13Y146_DO6;
  assign CLBLM_R_X7Y147_SLICE_X8Y147_B3 = CLBLM_R_X5Y144_SLICE_X6Y144_BQ;
  assign CLBLM_R_X7Y147_SLICE_X8Y147_B6 = CLBLM_R_X11Y144_SLICE_X14Y144_CO6;
  assign CLBLM_R_X7Y147_SLICE_X8Y147_C5 = CLBLM_R_X11Y144_SLICE_X14Y144_AO6;
  assign CLBLM_R_X7Y147_SLICE_X8Y147_C6 = CLBLM_R_X5Y144_SLICE_X7Y144_BQ;
  assign CLBLM_R_X7Y147_SLICE_X8Y147_CE = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X7Y147_SLICE_X8Y147_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X7Y153_SLICE_X8Y153_C4 = CLBLL_L_X4Y147_SLICE_X5Y147_CQ;
  assign RIOI3_X105Y121_ILOGIC_X1Y122_D = RIOB33_X105Y121_IOB_X1Y122_I;
  assign RIOI3_X105Y121_ILOGIC_X1Y121_D = RIOB33_X105Y121_IOB_X1Y121_I;
  assign CLBLM_R_X7Y153_SLICE_X8Y153_C5 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X7Y153_SLICE_X8Y153_C6 = CLBLM_R_X7Y153_SLICE_X8Y153_AQ;
  assign CLBLM_L_X12Y150_SLICE_X17Y150_A1 = 1'b1;
  assign CLBLM_L_X12Y150_SLICE_X17Y150_A2 = 1'b1;
  assign CLBLM_L_X12Y150_SLICE_X17Y150_A3 = 1'b1;
  assign CLBLM_L_X12Y150_SLICE_X17Y150_A4 = 1'b1;
  assign CLBLM_L_X12Y150_SLICE_X17Y150_A5 = 1'b1;
  assign CLBLM_L_X12Y150_SLICE_X17Y150_A6 = 1'b1;
  assign LIOB33_X0Y113_IOB_X0Y113_O = CLBLM_R_X3Y147_SLICE_X3Y147_C5Q;
  assign CLBLM_L_X12Y150_SLICE_X17Y150_B1 = 1'b1;
  assign CLBLM_L_X12Y150_SLICE_X17Y150_B2 = 1'b1;
  assign CLBLM_L_X12Y150_SLICE_X17Y150_B3 = 1'b1;
  assign CLBLM_L_X12Y150_SLICE_X17Y150_B4 = 1'b1;
  assign CLBLM_L_X12Y150_SLICE_X17Y150_B5 = 1'b1;
  assign CLBLM_L_X12Y150_SLICE_X17Y150_B6 = 1'b1;
  assign LIOB33_X0Y113_IOB_X0Y114_O = CLBLM_L_X8Y142_SLICE_X10Y142_A5Q;
  assign CLBLM_L_X12Y150_SLICE_X17Y150_C1 = 1'b1;
  assign CLBLM_L_X12Y150_SLICE_X17Y150_C2 = 1'b1;
  assign CLBLM_L_X12Y150_SLICE_X17Y150_C3 = 1'b1;
  assign CLBLM_L_X12Y150_SLICE_X17Y150_C4 = 1'b1;
  assign CLBLM_L_X12Y150_SLICE_X17Y150_C5 = 1'b1;
  assign CLBLM_L_X12Y150_SLICE_X17Y150_C6 = 1'b1;
  assign CLBLM_L_X12Y150_SLICE_X17Y150_D1 = 1'b1;
  assign CLBLM_L_X12Y150_SLICE_X17Y150_D2 = 1'b1;
  assign CLBLM_L_X12Y150_SLICE_X17Y150_D3 = 1'b1;
  assign CLBLM_L_X12Y150_SLICE_X17Y150_D4 = 1'b1;
  assign CLBLM_L_X12Y150_SLICE_X17Y150_D5 = 1'b1;
  assign CLBLM_L_X12Y150_SLICE_X17Y150_D6 = 1'b1;
  assign CLBLM_L_X12Y150_SLICE_X16Y150_A1 = 1'b1;
  assign CLBLM_L_X12Y150_SLICE_X16Y150_A2 = 1'b1;
  assign CLBLM_L_X12Y150_SLICE_X16Y150_A3 = CLBLM_L_X8Y149_SLICE_X11Y149_BO6;
  assign CLBLM_L_X12Y150_SLICE_X16Y150_A4 = CLBLM_L_X10Y148_SLICE_X12Y148_AQ;
  assign CLBLM_L_X12Y150_SLICE_X16Y150_A5 = CLBLM_R_X11Y149_SLICE_X15Y149_CO6;
  assign CLBLM_L_X12Y150_SLICE_X16Y150_A6 = 1'b1;
  assign CLBLM_L_X12Y150_SLICE_X16Y150_B1 = CLBLM_L_X8Y152_SLICE_X10Y152_DQ;
  assign CLBLM_L_X12Y150_SLICE_X16Y150_B2 = CLBLM_L_X12Y147_SLICE_X16Y147_AO5;
  assign CLBLM_L_X12Y150_SLICE_X16Y150_B3 = CLBLM_R_X11Y144_SLICE_X14Y144_CO6;
  assign CLBLM_L_X12Y150_SLICE_X16Y150_B4 = CLBLL_L_X4Y150_SLICE_X4Y150_CQ;
  assign CLBLM_L_X12Y150_SLICE_X16Y150_B5 = CLBLM_L_X10Y146_SLICE_X13Y146_DO6;
  assign CLBLM_L_X12Y150_SLICE_X16Y150_B6 = CLBLM_R_X7Y148_SLICE_X8Y148_AO5;
  assign CLBLM_L_X12Y150_SLICE_X16Y150_C1 = CLBLM_R_X7Y149_SLICE_X8Y149_AQ;
  assign CLBLM_L_X12Y150_SLICE_X16Y150_C2 = CLBLM_L_X10Y146_SLICE_X12Y146_AQ;
  assign CLBLM_L_X12Y150_SLICE_X16Y150_C3 = CLBLL_L_X4Y148_SLICE_X4Y148_CQ;
  assign CLBLM_L_X12Y150_SLICE_X16Y150_C4 = CLBLM_R_X7Y144_SLICE_X9Y144_B5Q;
  assign CLBLM_L_X12Y150_SLICE_X16Y150_C5 = CLBLM_R_X7Y153_SLICE_X8Y153_A5Q;
  assign CLBLM_L_X12Y150_SLICE_X16Y150_C6 = CLBLM_L_X12Y147_SLICE_X16Y147_DO6;
  assign CLBLM_L_X12Y150_SLICE_X16Y150_D1 = 1'b1;
  assign CLBLM_L_X12Y150_SLICE_X16Y150_D2 = 1'b1;
  assign CLBLM_L_X12Y150_SLICE_X16Y150_D3 = 1'b1;
  assign CLBLM_L_X12Y150_SLICE_X16Y150_D4 = 1'b1;
  assign CLBLM_L_X12Y150_SLICE_X16Y150_D5 = 1'b1;
  assign CLBLM_L_X12Y150_SLICE_X16Y150_D6 = 1'b1;
  assign LIOB33_SING_X0Y100_IOB_X0Y100_O = CLBLM_R_X3Y148_SLICE_X2Y148_B5Q;
  assign LIOI3_X0Y103_OLOGIC_X0Y104_T1 = 1'b1;
  assign LIOI3_X0Y77_ILOGIC_X0Y78_D = LIOB33_X0Y77_IOB_X0Y78_I;
  assign LIOI3_X0Y103_OLOGIC_X0Y103_D1 = CLBLM_R_X5Y145_SLICE_X7Y145_BQ;
  assign LIOB33_X0Y115_IOB_X0Y116_O = CLBLM_R_X7Y143_SLICE_X9Y143_B5Q;
  assign LIOB33_X0Y115_IOB_X0Y115_O = CLBLM_R_X5Y147_SLICE_X6Y147_C5Q;
  assign CLBLM_L_X12Y151_SLICE_X17Y151_A1 = 1'b1;
  assign CLBLM_L_X12Y151_SLICE_X17Y151_A2 = 1'b1;
  assign CLBLM_L_X12Y151_SLICE_X17Y151_A3 = 1'b1;
  assign CLBLM_L_X12Y151_SLICE_X17Y151_A4 = 1'b1;
  assign CLBLM_L_X12Y151_SLICE_X17Y151_A5 = 1'b1;
  assign CLBLM_L_X12Y151_SLICE_X17Y151_A6 = 1'b1;
  assign CLBLM_L_X12Y151_SLICE_X17Y151_B1 = 1'b1;
  assign CLBLM_L_X12Y151_SLICE_X17Y151_B2 = 1'b1;
  assign CLBLM_L_X12Y151_SLICE_X17Y151_B3 = 1'b1;
  assign CLBLM_L_X12Y151_SLICE_X17Y151_B4 = 1'b1;
  assign CLBLM_L_X12Y151_SLICE_X17Y151_B5 = 1'b1;
  assign CLBLM_L_X12Y151_SLICE_X17Y151_B6 = 1'b1;
  assign CLBLM_L_X12Y151_SLICE_X17Y151_C1 = 1'b1;
  assign CLBLM_L_X12Y151_SLICE_X17Y151_C2 = 1'b1;
  assign CLBLM_L_X12Y151_SLICE_X17Y151_C3 = 1'b1;
  assign CLBLM_L_X12Y151_SLICE_X17Y151_C4 = 1'b1;
  assign CLBLM_L_X12Y151_SLICE_X17Y151_C5 = 1'b1;
  assign CLBLM_L_X12Y151_SLICE_X17Y151_C6 = 1'b1;
  assign LIOB33_SING_X0Y149_IOB_X0Y149_O = RIOB33_X105Y115_IOB_X1Y115_I;
  assign LIOI3_X0Y103_OLOGIC_X0Y103_T1 = 1'b1;
  assign CLBLM_L_X12Y151_SLICE_X17Y151_D1 = 1'b1;
  assign CLBLM_L_X12Y151_SLICE_X17Y151_D2 = 1'b1;
  assign CLBLM_L_X12Y151_SLICE_X17Y151_D3 = 1'b1;
  assign CLBLM_L_X12Y151_SLICE_X17Y151_D4 = 1'b1;
  assign CLBLM_L_X12Y151_SLICE_X17Y151_D5 = 1'b1;
  assign CLBLM_L_X12Y151_SLICE_X17Y151_D6 = 1'b1;
  assign CLBLM_L_X12Y151_SLICE_X16Y151_A1 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_L_X12Y151_SLICE_X16Y151_A2 = 1'b1;
  assign CLBLM_L_X12Y151_SLICE_X16Y151_A3 = CLBLM_L_X12Y149_SLICE_X16Y149_AO6;
  assign CLBLM_L_X12Y151_SLICE_X16Y151_A4 = CLBLM_R_X11Y151_SLICE_X15Y151_A5Q;
  assign CLBLM_L_X12Y151_SLICE_X16Y151_A5 = CLBLM_L_X10Y148_SLICE_X12Y148_AQ;
  assign CLBLM_L_X12Y151_SLICE_X16Y151_A6 = 1'b1;
  assign CLBLM_L_X12Y151_SLICE_X16Y151_B1 = 1'b1;
  assign CLBLM_L_X12Y151_SLICE_X16Y151_B2 = 1'b1;
  assign CLBLM_L_X12Y151_SLICE_X16Y151_B3 = CLBLM_L_X10Y149_SLICE_X12Y149_CO6;
  assign CLBLM_L_X12Y151_SLICE_X16Y151_B4 = CLBLM_R_X11Y148_SLICE_X14Y148_AO6;
  assign CLBLM_L_X12Y151_SLICE_X16Y151_B5 = CLBLM_L_X10Y148_SLICE_X12Y148_AQ;
  assign CLBLM_L_X12Y151_SLICE_X16Y151_B6 = 1'b1;
  assign CLBLM_L_X12Y151_SLICE_X16Y151_C1 = 1'b1;
  assign CLBLM_L_X12Y151_SLICE_X16Y151_C2 = 1'b1;
  assign CLBLM_L_X12Y151_SLICE_X16Y151_C3 = 1'b1;
  assign CLBLM_L_X12Y151_SLICE_X16Y151_C4 = 1'b1;
  assign CLBLM_L_X12Y151_SLICE_X16Y151_C5 = 1'b1;
  assign CLBLM_L_X12Y151_SLICE_X16Y151_C6 = 1'b1;
  assign CLBLM_L_X12Y151_SLICE_X16Y151_CLK = CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O;
  assign CLBLM_L_X12Y151_SLICE_X16Y151_D1 = 1'b1;
  assign CLBLM_L_X12Y151_SLICE_X16Y151_D2 = 1'b1;
  assign CLBLM_L_X12Y151_SLICE_X16Y151_D3 = 1'b1;
  assign CLBLM_L_X12Y151_SLICE_X16Y151_D4 = 1'b1;
  assign CLBLM_L_X12Y151_SLICE_X16Y151_D5 = 1'b1;
  assign CLBLM_L_X12Y151_SLICE_X16Y151_D6 = 1'b1;
  assign LIOI3_X0Y139_OLOGIC_X0Y140_D1 = CLBLL_L_X4Y145_SLICE_X4Y145_C5Q;
  assign LIOI3_X0Y139_OLOGIC_X0Y140_T1 = 1'b1;
  assign RIOI3_X105Y183_OLOGIC_X1Y184_D1 = CLBLM_R_X3Y148_SLICE_X3Y148_DO5;
  assign LIOI3_X0Y139_OLOGIC_X0Y139_D1 = CLBLM_R_X3Y147_SLICE_X2Y147_DQ;
  assign RIOI3_X105Y183_OLOGIC_X1Y184_T1 = 1'b1;
  assign LIOI3_X0Y139_OLOGIC_X0Y139_T1 = 1'b1;
  assign RIOI3_X105Y183_OLOGIC_X1Y183_D1 = 1'b0;
  assign LIOB33_SING_X0Y150_IOB_X0Y150_O = CLBLM_R_X3Y144_SLICE_X2Y144_AO5;
  assign LIOI3_TBYTESRC_X0Y181_OLOGIC_X0Y182_D1 = RIOB33_X105Y129_IOB_X1Y129_I;
  assign RIOI3_X105Y183_OLOGIC_X1Y183_T1 = 1'b1;
  assign LIOI3_TBYTESRC_X0Y181_OLOGIC_X0Y182_T1 = 1'b1;
  assign LIOI3_TBYTESRC_X0Y181_OLOGIC_X0Y181_D1 = RIOB33_X105Y127_IOB_X1Y128_I;
  assign LIOI3_TBYTESRC_X0Y181_OLOGIC_X0Y181_T1 = 1'b1;
  assign LIOB33_X0Y117_IOB_X0Y118_O = CLBLM_R_X7Y142_SLICE_X9Y142_BQ;
  assign LIOB33_X0Y117_IOB_X0Y117_O = CLBLM_L_X10Y143_SLICE_X13Y143_C5Q;
  assign LIOB33_SING_X0Y199_IOB_X0Y199_O = 1'b1;
  assign CLBLM_L_X12Y152_SLICE_X17Y152_A1 = 1'b1;
  assign CLBLM_L_X12Y152_SLICE_X17Y152_A2 = 1'b1;
  assign CLBLM_L_X12Y152_SLICE_X17Y152_A3 = 1'b1;
  assign CLBLM_L_X12Y152_SLICE_X17Y152_A4 = 1'b1;
  assign CLBLM_L_X12Y152_SLICE_X17Y152_A5 = 1'b1;
  assign CLBLM_L_X12Y152_SLICE_X17Y152_A6 = 1'b1;
  assign CLBLM_L_X12Y152_SLICE_X17Y152_B1 = 1'b1;
  assign CLBLM_L_X12Y152_SLICE_X17Y152_B2 = 1'b1;
  assign CLBLM_L_X12Y152_SLICE_X17Y152_B3 = 1'b1;
  assign CLBLM_L_X12Y152_SLICE_X17Y152_B4 = 1'b1;
  assign CLBLM_L_X12Y152_SLICE_X17Y152_B5 = 1'b1;
  assign CLBLM_L_X12Y152_SLICE_X17Y152_B6 = 1'b1;
  assign CLBLM_L_X10Y142_SLICE_X13Y142_A1 = CLBLM_R_X11Y146_SLICE_X14Y146_AQ;
  assign CLBLM_L_X12Y152_SLICE_X17Y152_C2 = 1'b1;
  assign CLBLM_L_X12Y152_SLICE_X17Y152_C3 = 1'b1;
  assign CLBLM_L_X12Y152_SLICE_X17Y152_C4 = 1'b1;
  assign CLBLM_L_X12Y152_SLICE_X17Y152_C5 = 1'b1;
  assign CLBLM_L_X12Y152_SLICE_X17Y152_C6 = 1'b1;
  assign CLBLM_L_X10Y142_SLICE_X13Y142_A2 = CLBLM_L_X8Y142_SLICE_X10Y142_BQ;
  assign CLBLM_L_X10Y142_SLICE_X13Y142_A3 = CLBLM_L_X10Y142_SLICE_X13Y142_AQ;
  assign CLBLM_L_X10Y142_SLICE_X13Y142_A4 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_L_X10Y142_SLICE_X13Y142_A5 = CLBLM_L_X8Y144_SLICE_X10Y144_AO6;
  assign CLBLM_L_X10Y142_SLICE_X13Y142_A6 = CLBLM_L_X10Y144_SLICE_X12Y144_AO6;
  assign CLBLM_L_X10Y142_SLICE_X13Y142_B1 = CLBLM_L_X10Y144_SLICE_X13Y144_CQ;
  assign CLBLM_L_X10Y142_SLICE_X13Y142_B2 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X10Y142_SLICE_X13Y142_B3 = CLBLM_R_X7Y142_SLICE_X9Y142_BQ;
  assign CLBLM_L_X10Y142_SLICE_X13Y142_B4 = CLBLM_L_X10Y147_SLICE_X12Y147_AO5;
  assign CLBLM_L_X10Y142_SLICE_X13Y142_B5 = CLBLM_L_X8Y147_SLICE_X10Y147_C5Q;
  assign CLBLM_L_X10Y142_SLICE_X13Y142_B6 = CLBLM_L_X10Y142_SLICE_X13Y142_CO6;
  assign CLBLM_L_X12Y152_SLICE_X17Y152_D1 = 1'b1;
  assign CLBLM_L_X12Y152_SLICE_X17Y152_D2 = 1'b1;
  assign CLBLM_L_X10Y142_SLICE_X13Y142_C1 = CLBLM_L_X10Y145_SLICE_X12Y145_AQ;
  assign CLBLM_L_X10Y142_SLICE_X13Y142_C2 = CLBLM_R_X5Y142_SLICE_X7Y142_BQ;
  assign CLBLM_L_X10Y142_SLICE_X13Y142_C3 = 1'b1;
  assign CLBLM_L_X10Y142_SLICE_X13Y142_C4 = 1'b1;
  assign CLBLM_L_X10Y142_SLICE_X13Y142_C5 = 1'b1;
  assign CLBLM_L_X10Y142_SLICE_X13Y142_C6 = 1'b1;
  assign CLBLM_L_X10Y142_SLICE_X13Y142_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X12Y152_SLICE_X16Y152_A1 = RIOB33_X105Y133_IOB_X1Y133_I;
  assign CLBLM_L_X12Y152_SLICE_X16Y152_A2 = 1'b1;
  assign CLBLM_L_X12Y152_SLICE_X16Y152_A3 = CLBLM_L_X10Y148_SLICE_X12Y148_AQ;
  assign CLBLM_L_X12Y152_SLICE_X16Y152_A6 = 1'b1;
  assign CLBLM_L_X10Y142_SLICE_X13Y142_D1 = 1'b1;
  assign CLBLM_L_X10Y142_SLICE_X13Y142_D2 = 1'b1;
  assign CLBLM_L_X10Y142_SLICE_X13Y142_D3 = 1'b1;
  assign CLBLM_L_X10Y142_SLICE_X13Y142_D4 = 1'b1;
  assign CLBLM_L_X10Y142_SLICE_X13Y142_D5 = 1'b1;
  assign CLBLM_L_X12Y152_SLICE_X16Y152_B2 = 1'b1;
  assign CLBLM_L_X12Y152_SLICE_X16Y152_B3 = 1'b1;
  assign CLBLM_L_X12Y152_SLICE_X16Y152_B4 = 1'b1;
  assign CLBLM_L_X12Y152_SLICE_X16Y152_B5 = 1'b1;
  assign CLBLM_L_X12Y152_SLICE_X16Y152_B6 = 1'b1;
  assign CLBLM_L_X10Y142_SLICE_X13Y142_D6 = 1'b1;
  assign CLBLM_L_X12Y152_SLICE_X16Y152_B1 = 1'b1;
  assign CLBLM_L_X10Y142_SLICE_X12Y142_A1 = CLBLM_L_X8Y148_SLICE_X11Y148_B5Q;
  assign CLBLM_L_X10Y142_SLICE_X12Y142_A2 = CLBLM_L_X8Y147_SLICE_X10Y147_C5Q;
  assign CLBLM_L_X10Y142_SLICE_X12Y142_A3 = RIOB33_X105Y101_IOB_X1Y102_I;
  assign CLBLM_L_X12Y152_SLICE_X16Y152_C2 = 1'b1;
  assign CLBLM_L_X12Y152_SLICE_X16Y152_C3 = 1'b1;
  assign CLBLM_L_X12Y152_SLICE_X16Y152_C4 = 1'b1;
  assign CLBLM_L_X12Y152_SLICE_X16Y152_C5 = 1'b1;
  assign CLBLM_L_X12Y152_SLICE_X16Y152_C6 = 1'b1;
  assign CLBLM_L_X10Y142_SLICE_X12Y142_A4 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_L_X10Y142_SLICE_X12Y142_A5 = RIOB33_SING_X105Y100_IOB_X1Y100_I;
  assign CLBLM_L_X10Y142_SLICE_X12Y142_A6 = CLBLM_L_X10Y147_SLICE_X12Y147_CO6;
  assign CLBLM_L_X10Y142_SLICE_X12Y142_B1 = CLBLM_R_X7Y142_SLICE_X9Y142_CQ;
  assign CLBLM_L_X10Y142_SLICE_X12Y142_B2 = RIOB33_X105Y101_IOB_X1Y101_I;
  assign CLBLM_L_X10Y142_SLICE_X12Y142_B3 = RIOB33_SING_X105Y100_IOB_X1Y100_I;
  assign CLBLM_L_X10Y142_SLICE_X12Y142_B4 = RIOB33_X105Y103_IOB_X1Y104_I;
  assign CLBLM_L_X10Y142_SLICE_X12Y142_B5 = RIOB33_X105Y103_IOB_X1Y103_I;
  assign CLBLM_L_X10Y142_SLICE_X12Y142_B6 = RIOB33_X105Y131_IOB_X1Y131_I;
  assign CLBLM_L_X12Y152_SLICE_X16Y152_D1 = 1'b1;
  assign CLBLM_L_X12Y152_SLICE_X16Y152_D2 = 1'b1;
  assign CLBLM_L_X12Y152_SLICE_X16Y152_D3 = 1'b1;
  assign CLBLM_L_X10Y142_SLICE_X12Y142_C1 = CLBLL_L_X4Y151_SLICE_X4Y151_CQ;
  assign CLBLM_L_X10Y142_SLICE_X12Y142_C2 = 1'b1;
  assign CLBLM_L_X10Y142_SLICE_X12Y142_C3 = 1'b1;
  assign CLBLM_L_X10Y142_SLICE_X12Y142_C4 = RIOB33_X105Y131_IOB_X1Y131_I;
  assign CLBLM_L_X10Y142_SLICE_X12Y142_C5 = 1'b1;
  assign CLBLM_L_X10Y142_SLICE_X12Y142_C6 = CLBLM_L_X8Y142_SLICE_X11Y142_BQ;
  assign CLBLM_L_X12Y152_SLICE_X16Y152_D4 = 1'b1;
  assign CLBLM_L_X12Y152_SLICE_X16Y152_D5 = 1'b1;
  assign CLBLM_L_X12Y152_SLICE_X16Y152_D6 = 1'b1;
  assign CLBLM_L_X10Y142_SLICE_X12Y142_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign RIOI3_TBYTESRC_X105Y107_ILOGIC_X1Y108_D = RIOB33_X105Y107_IOB_X1Y108_I;
  assign RIOI3_TBYTESRC_X105Y107_ILOGIC_X1Y107_D = RIOB33_X105Y107_IOB_X1Y107_I;
  assign CLBLM_L_X10Y142_SLICE_X12Y142_D1 = 1'b1;
  assign CLBLM_L_X10Y142_SLICE_X12Y142_D2 = 1'b1;
  assign CLBLM_L_X10Y142_SLICE_X12Y142_D3 = 1'b1;
  assign CLBLM_L_X10Y142_SLICE_X12Y142_D4 = 1'b1;
  assign CLBLM_L_X10Y142_SLICE_X12Y142_D5 = 1'b1;
  assign CLBLM_L_X10Y142_SLICE_X12Y142_D6 = 1'b1;
  assign CLBLM_R_X13Y146_SLICE_X19Y146_A1 = 1'b1;
  assign CLBLM_R_X13Y146_SLICE_X19Y146_A2 = 1'b1;
  assign CLBLM_R_X13Y146_SLICE_X19Y146_A3 = 1'b1;
  assign CLBLM_R_X13Y146_SLICE_X19Y146_A4 = 1'b1;
  assign CLBLM_R_X13Y146_SLICE_X19Y146_A5 = 1'b1;
  assign CLBLM_R_X13Y146_SLICE_X19Y146_A6 = 1'b1;
  assign LIOI3_X0Y165_OLOGIC_X0Y165_T1 = 1'b1;
  assign CLBLM_R_X13Y146_SLICE_X19Y146_B1 = 1'b1;
  assign CLBLM_R_X13Y146_SLICE_X19Y146_B2 = 1'b1;
  assign CLBLM_R_X13Y146_SLICE_X19Y146_B3 = 1'b1;
  assign CLBLM_R_X13Y146_SLICE_X19Y146_B4 = 1'b1;
  assign CLBLM_R_X13Y146_SLICE_X19Y146_B5 = 1'b1;
  assign CLBLM_R_X13Y146_SLICE_X19Y146_B6 = 1'b1;
  assign CLBLM_R_X13Y146_SLICE_X19Y146_C1 = 1'b1;
  assign CLBLM_R_X13Y146_SLICE_X19Y146_C2 = 1'b1;
  assign CLBLM_R_X13Y146_SLICE_X19Y146_C3 = 1'b1;
  assign CLBLM_R_X13Y146_SLICE_X19Y146_C4 = 1'b1;
  assign CLBLM_R_X13Y146_SLICE_X19Y146_C5 = 1'b1;
  assign CLBLM_R_X13Y146_SLICE_X19Y146_C6 = 1'b1;
  assign CLBLM_R_X13Y146_SLICE_X19Y146_D1 = 1'b1;
  assign CLBLM_R_X13Y146_SLICE_X19Y146_D2 = 1'b1;
  assign CLBLM_R_X13Y146_SLICE_X19Y146_D3 = 1'b1;
  assign CLBLM_R_X13Y146_SLICE_X19Y146_D4 = 1'b1;
  assign CLBLM_R_X13Y146_SLICE_X19Y146_D5 = 1'b1;
  assign CLBLM_R_X13Y146_SLICE_X19Y146_D6 = 1'b1;
  assign CLBLM_R_X13Y146_SLICE_X18Y146_A1 = CLBLM_R_X7Y153_SLICE_X8Y153_A5Q;
  assign CLBLM_R_X13Y146_SLICE_X18Y146_A2 = CLBLM_R_X7Y144_SLICE_X9Y144_B5Q;
  assign CLBLM_R_X13Y146_SLICE_X18Y146_A3 = RIOB33_X105Y143_IOB_X1Y143_I;
  assign CLBLM_R_X13Y146_SLICE_X18Y146_A4 = CLBLM_L_X12Y146_SLICE_X16Y146_AQ;
  assign CLBLM_R_X13Y146_SLICE_X18Y146_A5 = CLBLM_L_X12Y145_SLICE_X17Y145_CO6;
  assign CLBLM_R_X13Y146_SLICE_X18Y146_A6 = 1'b1;
  assign CLBLM_R_X13Y146_SLICE_X18Y146_B1 = CLBLM_R_X7Y153_SLICE_X8Y153_A5Q;
  assign CLBLM_R_X13Y146_SLICE_X18Y146_B2 = CLBLM_R_X7Y144_SLICE_X9Y144_B5Q;
  assign CLBLM_R_X13Y146_SLICE_X18Y146_B3 = CLBLM_R_X7Y149_SLICE_X8Y149_AQ;
  assign CLBLM_R_X13Y146_SLICE_X18Y146_B4 = CLBLL_L_X4Y148_SLICE_X4Y148_CQ;
  assign CLBLM_R_X13Y146_SLICE_X18Y146_B5 = CLBLM_R_X7Y146_SLICE_X9Y146_CO6;
  assign CLBLM_R_X13Y146_SLICE_X18Y146_B6 = CLBLM_L_X10Y146_SLICE_X13Y146_DO6;
  assign CLBLM_R_X13Y146_SLICE_X18Y146_C1 = RIOB33_X105Y141_IOB_X1Y141_I;
  assign CLBLM_R_X13Y146_SLICE_X18Y146_C2 = 1'b1;
  assign CLBLM_R_X13Y146_SLICE_X18Y146_C3 = CLBLM_L_X10Y147_SLICE_X12Y147_AQ;
  assign CLBLM_R_X13Y146_SLICE_X18Y146_C4 = CLBLM_L_X10Y147_SLICE_X12Y147_CQ;
  assign CLBLM_R_X13Y146_SLICE_X18Y146_C5 = 1'b1;
  assign CLBLM_R_X13Y146_SLICE_X18Y146_C6 = RIOB33_X105Y139_IOB_X1Y140_I;
  assign LIOB33_X0Y119_IOB_X0Y119_O = CLBLL_L_X2Y146_SLICE_X0Y146_CQ;
  assign CLBLM_R_X13Y146_SLICE_X18Y146_D1 = 1'b1;
  assign CLBLM_R_X13Y146_SLICE_X18Y146_D2 = 1'b1;
  assign CLBLM_R_X13Y146_SLICE_X18Y146_D3 = 1'b1;
  assign CLBLM_R_X13Y146_SLICE_X18Y146_D4 = 1'b1;
  assign CLBLM_R_X13Y146_SLICE_X18Y146_D5 = 1'b1;
  assign CLBLM_R_X13Y146_SLICE_X18Y146_D6 = 1'b1;
  assign LIOB33_X0Y119_IOB_X0Y120_O = CLBLL_L_X4Y147_SLICE_X4Y147_AQ;
  assign CLBLM_L_X12Y153_SLICE_X17Y153_A1 = 1'b1;
  assign CLBLM_L_X12Y153_SLICE_X17Y153_A2 = 1'b1;
  assign CLBLM_L_X12Y153_SLICE_X17Y153_A3 = 1'b1;
  assign CLBLM_L_X12Y153_SLICE_X17Y153_A4 = 1'b1;
  assign CLBLM_L_X12Y153_SLICE_X17Y153_A5 = 1'b1;
  assign CLBLM_L_X12Y153_SLICE_X17Y153_A6 = 1'b1;
  assign RIOI3_X105Y141_ILOGIC_X1Y142_D = RIOB33_X105Y141_IOB_X1Y142_I;
  assign CLBLM_L_X12Y153_SLICE_X17Y153_B1 = 1'b1;
  assign CLBLM_L_X12Y153_SLICE_X17Y153_B2 = 1'b1;
  assign CLBLM_L_X12Y153_SLICE_X17Y153_B3 = 1'b1;
  assign CLBLM_L_X12Y153_SLICE_X17Y153_B4 = 1'b1;
  assign CLBLM_L_X12Y153_SLICE_X17Y153_B5 = 1'b1;
  assign CLBLM_L_X12Y153_SLICE_X17Y153_B6 = 1'b1;
  assign CLBLM_L_X10Y143_SLICE_X13Y143_A1 = CLBLM_L_X8Y146_SLICE_X11Y146_B5Q;
  assign CLBLM_L_X10Y143_SLICE_X13Y143_A2 = 1'b1;
  assign CLBLM_L_X10Y143_SLICE_X13Y143_A3 = CLBLM_L_X10Y143_SLICE_X13Y143_AQ;
  assign CLBLM_L_X12Y153_SLICE_X17Y153_C4 = 1'b1;
  assign CLBLM_L_X12Y153_SLICE_X17Y153_C5 = 1'b1;
  assign CLBLM_L_X12Y153_SLICE_X17Y153_C6 = 1'b1;
  assign CLBLM_L_X10Y143_SLICE_X13Y143_A4 = CLBLM_R_X11Y146_SLICE_X14Y146_DO6;
  assign CLBLM_L_X10Y143_SLICE_X13Y143_A5 = CLBLM_L_X8Y142_SLICE_X10Y142_AQ;
  assign CLBLM_L_X10Y143_SLICE_X13Y143_A6 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_L_X12Y153_SLICE_X17Y153_C1 = 1'b1;
  assign CLBLM_L_X12Y153_SLICE_X17Y153_C2 = 1'b1;
  assign CLBLM_L_X10Y143_SLICE_X13Y143_B1 = CLBLM_L_X10Y144_SLICE_X12Y144_AO6;
  assign CLBLM_L_X10Y143_SLICE_X13Y143_B2 = CLBLM_L_X10Y143_SLICE_X13Y143_BQ;
  assign CLBLM_L_X10Y143_SLICE_X13Y143_B3 = 1'b1;
  assign CLBLM_L_X10Y143_SLICE_X13Y143_B4 = CLBLM_L_X8Y143_SLICE_X11Y143_BQ;
  assign CLBLM_L_X12Y153_SLICE_X17Y153_D2 = 1'b1;
  assign CLBLM_L_X12Y153_SLICE_X17Y153_D3 = 1'b1;
  assign CLBLM_L_X12Y153_SLICE_X17Y153_D4 = 1'b1;
  assign CLBLM_L_X10Y143_SLICE_X13Y143_B5 = CLBLM_L_X10Y143_SLICE_X12Y143_DO6;
  assign CLBLM_L_X10Y143_SLICE_X13Y143_B6 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_L_X12Y153_SLICE_X17Y153_D1 = 1'b1;
  assign CLBLM_L_X12Y153_SLICE_X17Y153_D5 = 1'b1;
  assign CLBLM_L_X10Y143_SLICE_X13Y143_C1 = CLBLM_L_X10Y143_SLICE_X12Y143_AQ;
  assign CLBLM_L_X10Y143_SLICE_X13Y143_C2 = CLBLM_L_X10Y143_SLICE_X13Y143_CQ;
  assign CLBLM_L_X10Y143_SLICE_X13Y143_C3 = RIOB33_X105Y127_IOB_X1Y128_I;
  assign CLBLM_L_X10Y143_SLICE_X13Y143_C4 = CLBLM_L_X10Y146_SLICE_X12Y146_D5Q;
  assign CLBLM_L_X10Y143_SLICE_X13Y143_C5 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_L_X10Y143_SLICE_X13Y143_C6 = 1'b1;
  assign CLBLM_L_X10Y143_SLICE_X13Y143_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X12Y153_SLICE_X16Y153_A1 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_L_X12Y153_SLICE_X16Y153_A2 = CLBLM_R_X11Y149_SLICE_X14Y149_AO6;
  assign CLBLM_L_X12Y153_SLICE_X16Y153_A3 = CLBLM_R_X7Y153_SLICE_X9Y153_D5Q;
  assign CLBLM_L_X12Y153_SLICE_X16Y153_A4 = 1'b1;
  assign CLBLM_L_X12Y153_SLICE_X16Y153_A5 = CLBLM_L_X10Y148_SLICE_X12Y148_AQ;
  assign CLBLM_L_X10Y143_SLICE_X13Y143_D1 = CLBLM_L_X8Y144_SLICE_X10Y144_AO6;
  assign CLBLM_L_X10Y143_SLICE_X13Y143_D2 = CLBLM_L_X10Y142_SLICE_X13Y142_AQ;
  assign CLBLM_L_X10Y143_SLICE_X13Y143_D3 = CLBLM_L_X8Y144_SLICE_X11Y144_AQ;
  assign CLBLM_L_X10Y143_SLICE_X13Y143_D4 = CLBLM_L_X10Y143_SLICE_X13Y143_BQ;
  assign CLBLM_L_X12Y153_SLICE_X16Y153_B5 = 1'b1;
  assign CLBLM_L_X12Y153_SLICE_X16Y153_B6 = 1'b1;
  assign CLBLM_L_X10Y143_SLICE_X13Y143_D5 = CLBLM_L_X8Y142_SLICE_X10Y142_BQ;
  assign CLBLM_L_X10Y143_SLICE_X13Y143_D6 = 1'b1;
  assign CLBLM_L_X12Y153_SLICE_X16Y153_B1 = 1'b1;
  assign CLBLM_L_X12Y153_SLICE_X16Y153_B2 = 1'b1;
  assign CLBLM_L_X12Y153_SLICE_X16Y153_B3 = 1'b1;
  assign CLBLM_L_X12Y153_SLICE_X16Y153_B4 = 1'b1;
  assign CLBLM_L_X10Y143_SLICE_X12Y143_A1 = RIOB33_X105Y109_IOB_X1Y110_I;
  assign CLBLM_L_X12Y153_SLICE_X16Y153_C4 = 1'b1;
  assign CLBLM_L_X10Y143_SLICE_X12Y143_A2 = CLBLM_R_X7Y151_SLICE_X9Y151_A5Q;
  assign CLBLM_L_X12Y153_SLICE_X16Y153_C6 = 1'b1;
  assign CLBLM_L_X10Y143_SLICE_X12Y143_A3 = CLBLM_L_X10Y143_SLICE_X12Y143_AQ;
  assign CLBLM_L_X10Y143_SLICE_X12Y143_A4 = CLBLM_L_X10Y145_SLICE_X12Y145_A5Q;
  assign CLBLM_L_X10Y143_SLICE_X12Y143_A5 = CLBLM_L_X10Y144_SLICE_X12Y144_AQ;
  assign CLBLM_L_X10Y143_SLICE_X12Y143_A6 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_L_X12Y153_SLICE_X16Y153_C2 = 1'b1;
  assign CLBLM_L_X10Y143_SLICE_X12Y143_B1 = CLBLM_L_X8Y146_SLICE_X11Y146_B5Q;
  assign CLBLM_L_X10Y143_SLICE_X12Y143_B2 = CLBLM_L_X10Y143_SLICE_X12Y143_BQ;
  assign CLBLM_L_X10Y143_SLICE_X12Y143_B3 = CLBLM_R_X7Y153_SLICE_X9Y153_C5Q;
  assign CLBLM_L_X10Y143_SLICE_X12Y143_B4 = CLBLM_L_X8Y149_SLICE_X11Y149_AQ;
  assign CLBLM_L_X10Y143_SLICE_X12Y143_B5 = CLBLM_L_X10Y143_SLICE_X12Y143_CO5;
  assign CLBLM_L_X10Y143_SLICE_X12Y143_B6 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_L_X12Y153_SLICE_X16Y153_D1 = 1'b1;
  assign CLBLM_L_X12Y153_SLICE_X16Y153_D2 = 1'b1;
  assign CLBLM_L_X12Y153_SLICE_X16Y153_D3 = 1'b1;
  assign CLBLM_L_X10Y143_SLICE_X12Y143_C1 = CLBLM_L_X10Y143_SLICE_X12Y143_BQ;
  assign CLBLM_L_X10Y143_SLICE_X12Y143_C2 = 1'b1;
  assign CLBLM_L_X10Y143_SLICE_X12Y143_C3 = CLBLM_L_X10Y144_SLICE_X13Y144_DQ;
  assign CLBLM_L_X10Y143_SLICE_X12Y143_C4 = CLBLM_R_X7Y143_SLICE_X9Y143_AQ;
  assign CLBLM_L_X10Y143_SLICE_X12Y143_C5 = 1'b1;
  assign CLBLM_L_X10Y143_SLICE_X12Y143_C6 = 1'b1;
  assign CLBLM_L_X12Y153_SLICE_X16Y153_D5 = 1'b1;
  assign CLBLM_L_X12Y153_SLICE_X16Y153_D6 = 1'b1;
  assign CLBLM_L_X10Y143_SLICE_X12Y143_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X10Y143_SLICE_X12Y143_D1 = CLBLM_L_X8Y143_SLICE_X10Y143_AQ;
  assign CLBLM_L_X10Y143_SLICE_X12Y143_D2 = CLBLM_R_X3Y142_SLICE_X2Y142_BO5;
  assign CLBLM_L_X10Y143_SLICE_X12Y143_D3 = CLBLM_R_X5Y145_SLICE_X7Y145_B5Q;
  assign CLBLM_L_X10Y143_SLICE_X12Y143_D4 = CLBLM_L_X10Y142_SLICE_X13Y142_AQ;
  assign CLBLM_L_X10Y143_SLICE_X12Y143_D5 = CLBLM_L_X10Y144_SLICE_X13Y144_A5Q;
  assign CLBLM_L_X10Y143_SLICE_X12Y143_D6 = CLBLM_L_X8Y142_SLICE_X10Y142_BQ;
  assign RIOI3_X105Y197_OLOGIC_X1Y197_D1 = CLBLM_L_X12Y152_SLICE_X16Y152_AO5;
  assign LIOB33_X0Y121_IOB_X0Y122_O = CLBLL_L_X4Y144_SLICE_X5Y144_CQ;
  assign LIOB33_X0Y121_IOB_X0Y121_O = CLBLM_L_X8Y147_SLICE_X10Y147_C5Q;
  assign CLBLM_R_X11Y146_SLICE_X14Y146_A5 = CLBLM_L_X10Y146_SLICE_X13Y146_DO5;
  assign CLBLM_R_X11Y146_SLICE_X14Y146_A6 = CLBLM_L_X10Y144_SLICE_X13Y144_AQ;
  assign LIOI3_X0Y141_OLOGIC_X0Y142_D1 = CLBLL_L_X2Y146_SLICE_X0Y146_CQ;
  assign CLBLL_L_X4Y140_SLICE_X4Y140_A1 = 1'b1;
  assign CLBLL_L_X4Y140_SLICE_X4Y140_A2 = CLBLL_L_X4Y148_SLICE_X4Y148_AQ;
  assign CLBLL_L_X4Y140_SLICE_X4Y140_A3 = CLBLL_L_X4Y140_SLICE_X4Y140_AQ;
  assign CLBLL_L_X4Y140_SLICE_X4Y140_A4 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLL_L_X4Y140_SLICE_X4Y140_A5 = 1'b1;
  assign CLBLL_L_X4Y140_SLICE_X4Y140_A6 = CLBLL_L_X4Y140_SLICE_X4Y140_CO6;
  assign LIOI3_X0Y141_OLOGIC_X0Y142_T1 = 1'b1;
  assign RIOI3_X105Y185_OLOGIC_X1Y186_D1 = CLBLM_L_X10Y149_SLICE_X13Y149_BO6;
  assign CLBLL_L_X4Y140_SLICE_X4Y140_AX = CLBLL_L_X4Y140_SLICE_X4Y140_BO6;
  assign CLBLL_L_X4Y140_SLICE_X4Y140_B1 = LIOB33_X0Y59_IOB_X0Y60_I;
  assign CLBLL_L_X4Y140_SLICE_X4Y140_B2 = CLBLL_L_X4Y142_SLICE_X4Y142_CQ;
  assign CLBLL_L_X4Y140_SLICE_X4Y140_B3 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLL_L_X4Y140_SLICE_X4Y140_B4 = CLBLM_R_X3Y149_SLICE_X3Y149_D5Q;
  assign CLBLL_L_X4Y140_SLICE_X4Y140_B5 = CLBLL_L_X4Y140_SLICE_X4Y140_A5Q;
  assign CLBLL_L_X4Y140_SLICE_X4Y140_B6 = 1'b1;
  assign LIOI3_X0Y141_OLOGIC_X0Y141_D1 = CLBLL_L_X4Y145_SLICE_X5Y145_CQ;
  assign RIOI3_X105Y185_OLOGIC_X1Y186_T1 = 1'b1;
  assign CLBLL_L_X4Y140_SLICE_X4Y140_C1 = 1'b1;
  assign CLBLL_L_X4Y140_SLICE_X4Y140_C2 = 1'b1;
  assign CLBLL_L_X4Y140_SLICE_X4Y140_C3 = CLBLL_L_X4Y140_SLICE_X5Y140_DO6;
  assign CLBLL_L_X4Y140_SLICE_X4Y140_C4 = 1'b1;
  assign CLBLL_L_X4Y140_SLICE_X4Y140_C5 = LIOB33_X0Y53_IOB_X0Y54_I;
  assign CLBLL_L_X4Y140_SLICE_X4Y140_C6 = 1'b1;
  assign LIOI3_X0Y141_OLOGIC_X0Y141_T1 = 1'b1;
  assign CLBLL_L_X4Y140_SLICE_X4Y140_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign RIOI3_X105Y185_OLOGIC_X1Y185_D1 = CLBLM_L_X10Y153_SLICE_X12Y153_DO6;
  assign CLBLL_L_X4Y140_SLICE_X4Y140_D1 = 1'b1;
  assign CLBLL_L_X4Y140_SLICE_X4Y140_D2 = 1'b1;
  assign CLBLL_L_X4Y140_SLICE_X4Y140_D3 = 1'b1;
  assign CLBLL_L_X4Y140_SLICE_X4Y140_D4 = 1'b1;
  assign CLBLL_L_X4Y140_SLICE_X4Y140_D5 = 1'b1;
  assign CLBLL_L_X4Y140_SLICE_X4Y140_D6 = 1'b1;
  assign LIOI3_TBYTESRC_X0Y193_OLOGIC_X0Y194_D1 = RIOB33_X105Y103_IOB_X1Y103_I;
  assign RIOI3_X105Y185_OLOGIC_X1Y185_T1 = 1'b1;
  assign CLBLM_R_X11Y146_SLICE_X14Y146_B6 = 1'b1;
  assign LIOI3_TBYTESRC_X0Y193_OLOGIC_X0Y194_T1 = 1'b1;
  assign LIOI3_TBYTESRC_X0Y193_OLOGIC_X0Y193_D1 = CLBLL_L_X2Y166_SLICE_X0Y166_AO6;
  assign CLBLL_L_X4Y140_SLICE_X5Y140_A1 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLL_L_X4Y140_SLICE_X5Y140_A2 = CLBLM_R_X5Y152_SLICE_X6Y152_AQ;
  assign CLBLL_L_X4Y140_SLICE_X5Y140_A3 = CLBLL_L_X4Y140_SLICE_X5Y140_AQ;
  assign CLBLL_L_X4Y140_SLICE_X5Y140_A4 = 1'b1;
  assign CLBLL_L_X4Y140_SLICE_X5Y140_A5 = CLBLL_L_X4Y140_SLICE_X5Y140_CO5;
  assign CLBLL_L_X4Y140_SLICE_X5Y140_A6 = LIOB33_X0Y53_IOB_X0Y54_I;
  assign CLBLM_R_X11Y146_SLICE_X14Y146_C1 = CLBLM_R_X7Y149_SLICE_X8Y149_AQ;
  assign LIOI3_TBYTESRC_X0Y193_OLOGIC_X0Y193_T1 = 1'b1;
  assign CLBLL_L_X4Y140_SLICE_X5Y140_B1 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLL_L_X4Y140_SLICE_X5Y140_B2 = LIOB33_X0Y53_IOB_X0Y54_I;
  assign CLBLL_L_X4Y140_SLICE_X5Y140_B3 = 1'b1;
  assign CLBLL_L_X4Y140_SLICE_X5Y140_B4 = CLBLL_L_X4Y140_SLICE_X5Y140_BQ;
  assign CLBLL_L_X4Y140_SLICE_X5Y140_B5 = CLBLL_L_X4Y140_SLICE_X4Y140_AQ;
  assign CLBLL_L_X4Y140_SLICE_X5Y140_B6 = CLBLL_L_X4Y140_SLICE_X5Y140_CO6;
  assign CLBLM_L_X10Y144_SLICE_X13Y144_A1 = CLBLM_L_X10Y149_SLICE_X13Y149_AQ;
  assign CLBLM_L_X10Y144_SLICE_X13Y144_A4 = RIOB33_X105Y133_IOB_X1Y133_I;
  assign CLBLM_L_X10Y144_SLICE_X13Y144_A2 = CLBLM_R_X7Y144_SLICE_X8Y144_C5Q;
  assign CLBLM_L_X10Y144_SLICE_X13Y144_A6 = CLBLM_L_X10Y145_SLICE_X13Y145_CO6;
  assign CLBLM_L_X10Y144_SLICE_X13Y144_A3 = RIOB33_X105Y131_IOB_X1Y132_I;
  assign CLBLL_L_X4Y140_SLICE_X5Y140_C1 = CLBLL_L_X4Y140_SLICE_X4Y140_AQ;
  assign CLBLL_L_X4Y140_SLICE_X5Y140_C2 = CLBLM_R_X5Y140_SLICE_X6Y140_BQ;
  assign CLBLL_L_X4Y140_SLICE_X5Y140_C3 = CLBLM_R_X5Y140_SLICE_X6Y140_CQ;
  assign CLBLL_L_X4Y140_SLICE_X5Y140_C4 = CLBLL_L_X4Y140_SLICE_X5Y140_BQ;
  assign CLBLL_L_X4Y140_SLICE_X5Y140_C5 = CLBLM_R_X5Y140_SLICE_X6Y140_AQ;
  assign CLBLM_L_X10Y144_SLICE_X13Y144_B4 = CLBLM_L_X10Y145_SLICE_X12Y145_CO6;
  assign CLBLL_L_X4Y140_SLICE_X5Y140_C6 = 1'b1;
  assign CLBLM_L_X10Y144_SLICE_X13Y144_B5 = CLBLM_L_X10Y143_SLICE_X13Y143_C5Q;
  assign CLBLM_L_X10Y144_SLICE_X13Y144_B6 = CLBLM_R_X5Y148_SLICE_X7Y148_BQ;
  assign CLBLL_L_X4Y140_SLICE_X5Y140_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X10Y144_SLICE_X13Y144_B1 = CLBLM_L_X10Y144_SLICE_X12Y144_AO5;
  assign CLBLM_L_X10Y144_SLICE_X13Y144_C1 = CLBLM_L_X10Y143_SLICE_X13Y143_AQ;
  assign CLBLM_L_X10Y144_SLICE_X13Y144_B3 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLL_L_X4Y140_SLICE_X5Y140_D1 = CLBLL_L_X4Y140_SLICE_X4Y140_AQ;
  assign CLBLL_L_X4Y140_SLICE_X5Y140_D2 = CLBLM_R_X5Y140_SLICE_X6Y140_BQ;
  assign CLBLL_L_X4Y140_SLICE_X5Y140_D3 = CLBLL_L_X4Y140_SLICE_X5Y140_BQ;
  assign CLBLL_L_X4Y140_SLICE_X5Y140_D4 = CLBLM_R_X5Y140_SLICE_X6Y140_CQ;
  assign CLBLL_L_X4Y140_SLICE_X5Y140_D5 = CLBLL_L_X4Y140_SLICE_X5Y140_AQ;
  assign CLBLL_L_X4Y140_SLICE_X5Y140_D6 = CLBLM_R_X5Y140_SLICE_X6Y140_AQ;
  assign CLBLM_L_X10Y144_SLICE_X13Y144_C2 = CLBLM_L_X10Y143_SLICE_X13Y143_C5Q;
  assign CLBLM_L_X10Y144_SLICE_X13Y144_C3 = CLBLM_L_X8Y147_SLICE_X10Y147_C5Q;
  assign CLBLM_L_X10Y144_SLICE_X13Y144_C4 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_L_X10Y144_SLICE_X13Y144_C5 = 1'b1;
  assign CLBLM_L_X10Y144_SLICE_X13Y144_C6 = 1'b1;
  assign CLBLM_L_X10Y144_SLICE_X13Y144_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X10Y144_SLICE_X13Y144_D1 = CLBLM_R_X7Y143_SLICE_X9Y143_AQ;
  assign CLBLM_L_X10Y144_SLICE_X13Y144_D2 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_L_X10Y144_SLICE_X13Y144_D3 = CLBLM_L_X10Y144_SLICE_X13Y144_DQ;
  assign CLBLM_L_X10Y144_SLICE_X13Y144_D4 = CLBLM_L_X8Y151_SLICE_X10Y151_BQ;
  assign CLBLM_L_X10Y144_SLICE_X13Y144_D5 = CLBLM_L_X10Y144_SLICE_X13Y144_AQ;
  assign CLBLM_L_X10Y144_SLICE_X13Y144_D6 = CLBLM_L_X8Y149_SLICE_X11Y149_AQ;
  assign CLBLM_L_X10Y144_SLICE_X12Y144_A1 = CLBLM_L_X8Y145_SLICE_X11Y145_DQ;
  assign CLBLM_L_X10Y144_SLICE_X12Y144_A2 = CLBLM_L_X10Y147_SLICE_X12Y147_BQ;
  assign CLBLM_L_X10Y144_SLICE_X12Y144_A3 = CLBLM_L_X10Y144_SLICE_X13Y144_C5Q;
  assign CLBLM_L_X10Y144_SLICE_X12Y144_A4 = CLBLM_L_X10Y145_SLICE_X12Y145_CO6;
  assign CLBLM_L_X10Y144_SLICE_X12Y144_A5 = CLBLM_L_X10Y143_SLICE_X13Y143_C5Q;
  assign CLBLM_L_X10Y144_SLICE_X12Y144_A6 = 1'b1;
  assign CLBLM_L_X10Y144_SLICE_X12Y144_AX = CLBLM_R_X3Y145_SLICE_X3Y145_C5Q;
  assign CLBLM_L_X10Y144_SLICE_X12Y144_B1 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_L_X10Y144_SLICE_X12Y144_B2 = CLBLM_R_X3Y142_SLICE_X2Y142_BO5;
  assign CLBLM_L_X10Y144_SLICE_X12Y144_B3 = CLBLM_L_X10Y144_SLICE_X13Y144_A5Q;
  assign CLBLM_L_X10Y144_SLICE_X12Y144_B4 = CLBLM_L_X10Y144_SLICE_X13Y144_BQ;
  assign CLBLM_L_X10Y144_SLICE_X12Y144_B5 = CLBLM_L_X10Y144_SLICE_X12Y144_AO6;
  assign CLBLM_L_X10Y144_SLICE_X12Y144_B6 = 1'b1;
  assign CLBLM_L_X10Y144_SLICE_X12Y144_C1 = CLBLM_L_X10Y142_SLICE_X12Y142_AQ;
  assign CLBLM_L_X10Y144_SLICE_X12Y144_C2 = RIOB33_X105Y101_IOB_X1Y102_I;
  assign CLBLM_L_X10Y144_SLICE_X12Y144_C3 = RIOB33_SING_X105Y100_IOB_X1Y100_I;
  assign CLBLM_L_X10Y144_SLICE_X12Y144_C4 = CLBLM_L_X8Y148_SLICE_X11Y148_B5Q;
  assign CLBLM_L_X10Y144_SLICE_X12Y144_C5 = CLBLM_L_X10Y142_SLICE_X12Y142_BO6;
  assign CLBLM_L_X10Y144_SLICE_X12Y144_C6 = CLBLM_L_X8Y154_SLICE_X10Y154_BO5;
  assign CLBLM_L_X10Y144_SLICE_X12Y144_CE = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X7Y148_SLICE_X8Y148_A5 = CLBLM_R_X7Y149_SLICE_X8Y149_AQ;
  assign CLBLM_L_X10Y144_SLICE_X12Y144_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X7Y148_SLICE_X8Y148_A6 = 1'b1;
  assign CLBLM_L_X10Y144_SLICE_X12Y144_D1 = 1'b1;
  assign CLBLM_L_X10Y144_SLICE_X12Y144_D2 = 1'b1;
  assign CLBLM_L_X10Y144_SLICE_X12Y144_D3 = 1'b1;
  assign CLBLM_L_X10Y144_SLICE_X12Y144_D4 = 1'b1;
  assign CLBLM_L_X10Y144_SLICE_X12Y144_D5 = 1'b1;
  assign CLBLM_L_X10Y144_SLICE_X12Y144_D6 = 1'b1;
  assign CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_I = CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_O;
  assign RIOI3_X105Y125_ILOGIC_X1Y126_D = RIOB33_X105Y125_IOB_X1Y126_I;
  assign RIOI3_X105Y125_ILOGIC_X1Y125_D = RIOB33_X105Y125_IOB_X1Y125_I;
  assign LIOB33_X0Y123_IOB_X0Y124_O = CLBLL_L_X4Y151_SLICE_X4Y151_CQ;
  assign LIOB33_X0Y123_IOB_X0Y123_O = CLBLL_L_X2Y146_SLICE_X0Y146_CQ;
  assign CLBLM_R_X7Y148_SLICE_X8Y148_C1 = CLBLM_R_X7Y148_SLICE_X8Y148_AO6;
  assign CLBLM_R_X7Y148_SLICE_X8Y148_C2 = CLBLM_R_X7Y144_SLICE_X9Y144_A5Q;
  assign CLBLM_R_X7Y148_SLICE_X8Y148_C5 = CLBLM_R_X5Y142_SLICE_X6Y142_BQ;
  assign RIOI3_TBYTESRC_X105Y119_ILOGIC_X1Y120_D = RIOB33_X105Y119_IOB_X1Y120_I;
  assign RIOI3_TBYTESRC_X105Y119_ILOGIC_X1Y119_D = RIOB33_X105Y119_IOB_X1Y119_I;
  assign CLBLM_L_X10Y145_SLICE_X13Y145_A1 = CLBLM_L_X10Y143_SLICE_X13Y143_DO6;
  assign CLBLM_L_X10Y145_SLICE_X13Y145_A2 = CLBLM_L_X8Y144_SLICE_X11Y144_AQ;
  assign CLBLM_L_X10Y145_SLICE_X13Y145_A3 = CLBLM_L_X10Y145_SLICE_X13Y145_AQ;
  assign CLBLM_L_X10Y145_SLICE_X13Y145_A4 = CLBLM_R_X5Y145_SLICE_X6Y145_DQ;
  assign CLBLM_L_X10Y145_SLICE_X13Y145_A5 = CLBLM_L_X10Y144_SLICE_X12Y144_AO6;
  assign CLBLM_L_X10Y145_SLICE_X13Y145_A6 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_L_X10Y145_SLICE_X13Y145_B1 = CLBLM_L_X8Y144_SLICE_X10Y144_BO6;
  assign CLBLM_L_X10Y145_SLICE_X13Y145_B2 = CLBLM_L_X10Y149_SLICE_X13Y149_AQ;
  assign CLBLM_L_X10Y145_SLICE_X13Y145_B3 = CLBLM_L_X10Y151_SLICE_X13Y151_A5Q;
  assign CLBLM_L_X10Y145_SLICE_X13Y145_B4 = CLBLM_R_X7Y144_SLICE_X8Y144_C5Q;
  assign CLBLM_L_X10Y145_SLICE_X13Y145_B5 = CLBLM_L_X10Y153_SLICE_X13Y153_A5Q;
  assign CLBLM_L_X10Y145_SLICE_X13Y145_B6 = CLBLL_L_X4Y149_SLICE_X5Y149_C5Q;
  assign CLBLM_L_X10Y145_SLICE_X13Y145_C1 = CLBLM_L_X10Y153_SLICE_X13Y153_A5Q;
  assign CLBLM_L_X10Y145_SLICE_X13Y145_C2 = CLBLM_L_X10Y149_SLICE_X13Y149_AQ;
  assign CLBLM_L_X10Y145_SLICE_X13Y145_C3 = CLBLM_L_X8Y144_SLICE_X10Y144_BO6;
  assign CLBLM_L_X10Y145_SLICE_X13Y145_C4 = CLBLL_L_X4Y149_SLICE_X5Y149_C5Q;
  assign CLBLM_L_X10Y145_SLICE_X13Y145_C5 = 1'b1;
  assign CLBLM_L_X10Y145_SLICE_X13Y145_C6 = CLBLM_L_X10Y151_SLICE_X13Y151_A5Q;
  assign CLBLM_L_X10Y145_SLICE_X13Y145_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X10Y145_SLICE_X13Y145_D1 = 1'b1;
  assign CLBLM_L_X10Y145_SLICE_X13Y145_D2 = CLBLM_L_X10Y144_SLICE_X13Y144_A5Q;
  assign CLBLM_L_X10Y145_SLICE_X13Y145_D3 = CLBLM_L_X8Y146_SLICE_X10Y146_AQ;
  assign CLBLM_L_X10Y145_SLICE_X13Y145_D4 = 1'b1;
  assign CLBLM_L_X10Y145_SLICE_X13Y145_D5 = CLBLM_L_X10Y145_SLICE_X13Y145_AQ;
  assign CLBLM_L_X10Y145_SLICE_X13Y145_D6 = CLBLM_L_X10Y143_SLICE_X13Y143_DO5;
  assign CLBLM_L_X10Y145_SLICE_X12Y145_A1 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_L_X10Y145_SLICE_X12Y145_A2 = CLBLM_L_X8Y147_SLICE_X11Y147_AQ;
  assign CLBLM_L_X10Y145_SLICE_X12Y145_A3 = RIOB33_X105Y109_IOB_X1Y110_I;
  assign CLBLM_L_X10Y145_SLICE_X12Y145_A4 = CLBLM_L_X8Y153_SLICE_X10Y153_CQ;
  assign CLBLM_L_X10Y145_SLICE_X12Y145_A5 = 1'b1;
  assign CLBLM_L_X10Y145_SLICE_X12Y145_A6 = 1'b1;
  assign CLBLM_L_X10Y145_SLICE_X12Y145_B1 = CLBLM_L_X10Y142_SLICE_X12Y142_CO6;
  assign CLBLM_L_X10Y145_SLICE_X12Y145_B2 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_L_X10Y145_SLICE_X12Y145_B3 = CLBLM_L_X10Y144_SLICE_X12Y144_AQ;
  assign CLBLM_L_X10Y145_SLICE_X12Y145_B4 = CLBLM_L_X8Y145_SLICE_X11Y145_DQ;
  assign CLBLM_L_X10Y145_SLICE_X12Y145_B5 = 1'b1;
  assign CLBLM_L_X10Y145_SLICE_X12Y145_B6 = CLBLM_R_X3Y145_SLICE_X3Y145_DQ;
  assign CLBLM_L_X10Y145_SLICE_X12Y145_C1 = CLBLM_R_X3Y142_SLICE_X2Y142_BO5;
  assign CLBLM_L_X10Y145_SLICE_X12Y145_C2 = CLBLM_L_X8Y145_SLICE_X11Y145_DQ;
  assign CLBLM_L_X10Y145_SLICE_X12Y145_C3 = CLBLM_L_X10Y145_SLICE_X13Y145_DO6;
  assign CLBLM_L_X10Y145_SLICE_X12Y145_C4 = CLBLM_R_X5Y145_SLICE_X7Y145_B5Q;
  assign CLBLM_L_X10Y145_SLICE_X12Y145_C5 = CLBLM_L_X8Y146_SLICE_X10Y146_AQ;
  assign CLBLM_L_X10Y145_SLICE_X12Y145_C6 = CLBLM_L_X10Y147_SLICE_X12Y147_BQ;
  assign CLBLM_L_X10Y145_SLICE_X12Y145_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X10Y145_SLICE_X12Y145_D1 = CLBLM_L_X10Y151_SLICE_X13Y151_A5Q;
  assign CLBLM_L_X10Y145_SLICE_X12Y145_D2 = CLBLM_L_X10Y148_SLICE_X12Y148_AO5;
  assign CLBLM_L_X10Y145_SLICE_X12Y145_D3 = CLBLM_R_X7Y145_SLICE_X9Y145_DO6;
  assign CLBLM_L_X10Y145_SLICE_X12Y145_D4 = CLBLL_L_X4Y148_SLICE_X4Y148_CQ;
  assign CLBLM_L_X10Y145_SLICE_X12Y145_D5 = CLBLM_L_X12Y146_SLICE_X16Y146_CO6;
  assign CLBLM_L_X10Y145_SLICE_X12Y145_D6 = CLBLM_R_X3Y145_SLICE_X3Y145_C5Q;
  assign LIOB33_X0Y125_IOB_X0Y126_O = CLBLL_L_X4Y147_SLICE_X5Y147_CQ;
  assign LIOB33_X0Y125_IOB_X0Y125_O = CLBLL_L_X4Y151_SLICE_X4Y151_BQ;
  assign CLBLM_R_X13Y149_SLICE_X19Y149_A1 = 1'b1;
  assign CLBLM_R_X13Y149_SLICE_X19Y149_A2 = 1'b1;
  assign CLBLM_R_X13Y149_SLICE_X19Y149_A3 = 1'b1;
  assign CLBLM_R_X13Y149_SLICE_X19Y149_A4 = 1'b1;
  assign CLBLM_R_X13Y149_SLICE_X19Y149_A5 = 1'b1;
  assign CLBLM_R_X13Y149_SLICE_X19Y149_A6 = 1'b1;
  assign CLBLM_R_X13Y149_SLICE_X19Y149_B1 = 1'b1;
  assign CLBLM_R_X13Y149_SLICE_X19Y149_B2 = 1'b1;
  assign CLBLM_R_X13Y149_SLICE_X19Y149_B3 = 1'b1;
  assign CLBLM_R_X13Y149_SLICE_X19Y149_B4 = 1'b1;
  assign CLBLM_R_X13Y149_SLICE_X19Y149_B5 = 1'b1;
  assign CLBLM_R_X13Y149_SLICE_X19Y149_B6 = 1'b1;
  assign CLBLM_R_X13Y149_SLICE_X19Y149_C1 = 1'b1;
  assign CLBLM_R_X13Y149_SLICE_X19Y149_C2 = 1'b1;
  assign CLBLM_R_X13Y149_SLICE_X19Y149_C3 = 1'b1;
  assign CLBLM_R_X13Y149_SLICE_X19Y149_C4 = 1'b1;
  assign CLBLM_R_X13Y149_SLICE_X19Y149_C5 = 1'b1;
  assign CLBLM_R_X13Y149_SLICE_X19Y149_C6 = 1'b1;
  assign CLBLM_R_X13Y149_SLICE_X19Y149_D1 = 1'b1;
  assign CLBLM_R_X13Y149_SLICE_X19Y149_D2 = 1'b1;
  assign CLBLM_R_X13Y149_SLICE_X19Y149_D3 = 1'b1;
  assign CLBLM_R_X13Y149_SLICE_X19Y149_D4 = 1'b1;
  assign CLBLM_R_X13Y149_SLICE_X19Y149_D5 = 1'b1;
  assign CLBLM_R_X13Y149_SLICE_X19Y149_D6 = 1'b1;
  assign CLBLM_R_X13Y149_SLICE_X18Y149_A1 = CLBLM_R_X7Y144_SLICE_X9Y144_B5Q;
  assign CLBLM_R_X13Y149_SLICE_X18Y149_A2 = CLBLM_R_X7Y153_SLICE_X8Y153_A5Q;
  assign CLBLM_R_X13Y149_SLICE_X18Y149_A3 = CLBLM_R_X7Y149_SLICE_X8Y149_AQ;
  assign CLBLM_R_X13Y149_SLICE_X18Y149_A4 = CLBLL_L_X4Y148_SLICE_X4Y148_CQ;
  assign CLBLM_R_X13Y149_SLICE_X18Y149_A5 = CLBLM_L_X12Y147_SLICE_X16Y147_DO6;
  assign CLBLM_R_X13Y149_SLICE_X18Y149_A6 = CLBLM_L_X10Y146_SLICE_X13Y146_DO6;
  assign CLBLM_R_X13Y149_SLICE_X18Y149_B1 = 1'b1;
  assign CLBLM_R_X13Y149_SLICE_X18Y149_B2 = 1'b1;
  assign CLBLM_R_X13Y149_SLICE_X18Y149_B3 = 1'b1;
  assign CLBLM_R_X13Y149_SLICE_X18Y149_B4 = 1'b1;
  assign CLBLM_R_X13Y149_SLICE_X18Y149_B5 = 1'b1;
  assign CLBLM_R_X13Y149_SLICE_X18Y149_B6 = 1'b1;
  assign CLBLM_R_X13Y149_SLICE_X18Y149_C1 = 1'b1;
  assign CLBLM_R_X13Y149_SLICE_X18Y149_C2 = 1'b1;
  assign CLBLM_R_X13Y149_SLICE_X18Y149_C3 = 1'b1;
  assign CLBLM_R_X13Y149_SLICE_X18Y149_C4 = 1'b1;
  assign CLBLM_R_X13Y149_SLICE_X18Y149_C5 = 1'b1;
  assign CLBLM_R_X13Y149_SLICE_X18Y149_C6 = 1'b1;
  assign CLBLM_R_X13Y149_SLICE_X18Y149_D1 = 1'b1;
  assign CLBLM_R_X13Y149_SLICE_X18Y149_D2 = 1'b1;
  assign CLBLM_R_X13Y149_SLICE_X18Y149_D3 = 1'b1;
  assign CLBLM_R_X13Y149_SLICE_X18Y149_D4 = 1'b1;
  assign CLBLM_R_X13Y149_SLICE_X18Y149_D5 = 1'b1;
  assign CLBLM_R_X13Y149_SLICE_X18Y149_D6 = 1'b1;
  assign CLBLL_L_X4Y142_SLICE_X4Y142_A1 = LIOB33_X0Y59_IOB_X0Y60_I;
  assign CLBLL_L_X4Y142_SLICE_X4Y142_A2 = CLBLM_R_X3Y151_SLICE_X2Y151_BO5;
  assign CLBLL_L_X4Y142_SLICE_X4Y142_A3 = CLBLL_L_X4Y142_SLICE_X4Y142_CQ;
  assign CLBLL_L_X4Y142_SLICE_X4Y142_A4 = CLBLL_L_X4Y144_SLICE_X5Y144_BQ;
  assign CLBLL_L_X4Y142_SLICE_X4Y142_A5 = CLBLL_L_X4Y140_SLICE_X4Y140_A5Q;
  assign CLBLL_L_X4Y142_SLICE_X4Y142_A6 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLL_L_X4Y142_SLICE_X4Y142_AX = CLBLL_L_X4Y143_SLICE_X5Y143_CO6;
  assign CLBLL_L_X4Y142_SLICE_X4Y142_B1 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLL_L_X4Y142_SLICE_X4Y142_B2 = CLBLL_L_X4Y142_SLICE_X4Y142_BQ;
  assign CLBLL_L_X4Y142_SLICE_X4Y142_B3 = CLBLM_L_X10Y144_SLICE_X12Y144_AO6;
  assign CLBLL_L_X4Y142_SLICE_X4Y142_B4 = CLBLL_L_X4Y143_SLICE_X4Y143_C5Q;
  assign CLBLL_L_X4Y142_SLICE_X4Y142_B5 = CLBLM_R_X5Y147_SLICE_X6Y147_AQ;
  assign CLBLL_L_X4Y142_SLICE_X4Y142_B6 = CLBLM_R_X3Y142_SLICE_X3Y142_AQ;
  assign CLBLL_L_X4Y142_SLICE_X4Y142_C1 = 1'b1;
  assign CLBLL_L_X4Y142_SLICE_X4Y142_C2 = CLBLL_L_X4Y142_SLICE_X4Y142_CQ;
  assign CLBLL_L_X4Y142_SLICE_X4Y142_C3 = LIOB33_X0Y59_IOB_X0Y60_I;
  assign CLBLL_L_X4Y142_SLICE_X4Y142_C4 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLL_L_X4Y142_SLICE_X4Y142_C5 = CLBLM_R_X7Y142_SLICE_X8Y142_DQ;
  assign CLBLL_L_X4Y142_SLICE_X4Y142_C6 = 1'b1;
  assign CLBLL_L_X4Y142_SLICE_X4Y142_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLL_L_X2Y75_SLICE_X0Y75_A1 = 1'b1;
  assign CLBLL_L_X2Y75_SLICE_X0Y75_A2 = 1'b1;
  assign CLBLL_L_X2Y75_SLICE_X0Y75_A3 = LIOB33_X0Y55_IOB_X0Y56_I;
  assign CLBLL_L_X2Y75_SLICE_X0Y75_A4 = 1'b1;
  assign CLBLL_L_X4Y142_SLICE_X4Y142_D4 = 1'b1;
  assign CLBLL_L_X4Y142_SLICE_X4Y142_D5 = 1'b1;
  assign CLBLL_L_X4Y142_SLICE_X4Y142_D6 = 1'b1;
  assign CLBLL_L_X2Y75_SLICE_X0Y75_A5 = 1'b1;
  assign CLBLL_L_X2Y75_SLICE_X0Y75_A6 = 1'b1;
  assign CLBLL_L_X4Y142_SLICE_X4Y142_D1 = 1'b1;
  assign CLBLL_L_X4Y142_SLICE_X4Y142_D2 = 1'b1;
  assign CLBLL_L_X4Y142_SLICE_X4Y142_D3 = 1'b1;
  assign CLBLL_L_X2Y75_SLICE_X0Y75_B1 = 1'b1;
  assign CLBLL_L_X2Y75_SLICE_X0Y75_B2 = 1'b1;
  assign CLBLL_L_X2Y75_SLICE_X0Y75_B3 = 1'b1;
  assign CLBLL_L_X2Y75_SLICE_X0Y75_B4 = 1'b1;
  assign CLBLL_L_X2Y75_SLICE_X0Y75_B5 = 1'b1;
  assign CLBLL_L_X2Y75_SLICE_X0Y75_B6 = 1'b1;
  assign CLBLL_L_X2Y75_SLICE_X0Y75_C1 = 1'b1;
  assign CLBLL_L_X2Y75_SLICE_X0Y75_C2 = 1'b1;
  assign CLBLL_L_X2Y75_SLICE_X0Y75_C3 = 1'b1;
  assign CLBLL_L_X2Y75_SLICE_X0Y75_C4 = 1'b1;
  assign CLBLL_L_X2Y75_SLICE_X0Y75_C5 = 1'b1;
  assign CLBLL_L_X2Y75_SLICE_X0Y75_C6 = 1'b1;
  assign CLBLL_L_X2Y75_SLICE_X0Y75_D1 = 1'b1;
  assign CLBLL_L_X2Y75_SLICE_X0Y75_D2 = 1'b1;
  assign CLBLL_L_X2Y75_SLICE_X0Y75_D3 = 1'b1;
  assign CLBLL_L_X2Y75_SLICE_X0Y75_D4 = 1'b1;
  assign CLBLL_L_X2Y75_SLICE_X0Y75_D5 = 1'b1;
  assign CLBLL_L_X2Y75_SLICE_X0Y75_D6 = 1'b1;
  assign CLBLL_L_X4Y142_SLICE_X5Y142_A1 = CLBLL_L_X4Y142_SLICE_X5Y142_AQ;
  assign CLBLL_L_X4Y142_SLICE_X5Y142_A2 = CLBLL_L_X4Y143_SLICE_X4Y143_CQ;
  assign CLBLL_L_X4Y142_SLICE_X5Y142_A3 = CLBLM_L_X8Y147_SLICE_X10Y147_C5Q;
  assign CLBLL_L_X4Y142_SLICE_X5Y142_A4 = CLBLL_L_X4Y140_SLICE_X5Y140_BQ;
  assign CLBLL_L_X4Y142_SLICE_X5Y142_A5 = CLBLM_L_X10Y144_SLICE_X13Y144_CQ;
  assign CLBLL_L_X4Y142_SLICE_X5Y142_A6 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLL_L_X4Y142_SLICE_X5Y142_B1 = CLBLL_L_X4Y147_SLICE_X4Y147_BQ;
  assign CLBLL_L_X4Y142_SLICE_X5Y142_B2 = CLBLL_L_X4Y142_SLICE_X5Y142_BQ;
  assign CLBLL_L_X4Y142_SLICE_X5Y142_B3 = CLBLM_L_X8Y147_SLICE_X10Y147_C5Q;
  assign CLBLL_L_X4Y142_SLICE_X5Y142_B4 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLL_L_X4Y142_SLICE_X5Y142_B5 = CLBLM_L_X10Y144_SLICE_X13Y144_CQ;
  assign CLBLL_L_X4Y142_SLICE_X5Y142_B6 = CLBLM_L_X12Y145_SLICE_X16Y145_AQ;
  assign CLBLL_L_X4Y142_SLICE_X5Y142_C1 = 1'b1;
  assign CLBLL_L_X4Y142_SLICE_X5Y142_C2 = CLBLM_R_X5Y140_SLICE_X6Y140_BQ;
  assign CLBLL_L_X4Y142_SLICE_X5Y142_C3 = CLBLL_L_X4Y143_SLICE_X4Y143_DQ;
  assign CLBLL_L_X4Y142_SLICE_X5Y142_C4 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLL_L_X4Y142_SLICE_X5Y142_C5 = CLBLL_L_X4Y142_SLICE_X4Y142_BQ;
  assign CLBLL_L_X4Y142_SLICE_X5Y142_C6 = 1'b1;
  assign CLBLM_L_X10Y146_SLICE_X13Y146_A1 = CLBLM_R_X11Y146_SLICE_X14Y146_DO6;
  assign CLBLM_L_X10Y146_SLICE_X13Y146_A2 = 1'b1;
  assign CLBLL_L_X4Y142_SLICE_X5Y142_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X10Y146_SLICE_X13Y146_A3 = CLBLM_L_X10Y146_SLICE_X13Y146_AQ;
  assign CLBLM_L_X10Y146_SLICE_X13Y146_A4 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_L_X10Y146_SLICE_X13Y146_A5 = CLBLL_L_X4Y146_SLICE_X4Y146_AQ;
  assign CLBLM_L_X10Y146_SLICE_X13Y146_A6 = CLBLL_L_X4Y150_SLICE_X5Y150_A5Q;
  assign CLBLL_L_X2Y75_SLICE_X1Y75_A1 = 1'b1;
  assign CLBLL_L_X2Y75_SLICE_X1Y75_A2 = 1'b1;
  assign CLBLL_L_X2Y75_SLICE_X1Y75_A3 = 1'b1;
  assign CLBLL_L_X4Y142_SLICE_X5Y142_D3 = CLBLL_L_X4Y142_SLICE_X5Y142_BQ;
  assign CLBLL_L_X4Y142_SLICE_X5Y142_D4 = CLBLL_L_X4Y147_SLICE_X5Y147_CQ;
  assign CLBLL_L_X4Y142_SLICE_X5Y142_D5 = CLBLL_L_X4Y148_SLICE_X4Y148_CQ;
  assign CLBLL_L_X4Y142_SLICE_X5Y142_D6 = 1'b1;
  assign CLBLL_L_X2Y75_SLICE_X1Y75_A4 = 1'b1;
  assign CLBLL_L_X2Y75_SLICE_X1Y75_A5 = 1'b1;
  assign CLBLL_L_X2Y75_SLICE_X1Y75_A6 = 1'b1;
  assign CLBLL_L_X4Y142_SLICE_X5Y142_D1 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLL_L_X4Y142_SLICE_X5Y142_D2 = CLBLM_R_X7Y142_SLICE_X9Y142_BQ;
  assign CLBLL_L_X2Y75_SLICE_X1Y75_B1 = 1'b1;
  assign CLBLL_L_X2Y75_SLICE_X1Y75_B2 = 1'b1;
  assign CLBLL_L_X2Y75_SLICE_X1Y75_B3 = 1'b1;
  assign CLBLL_L_X2Y75_SLICE_X1Y75_B4 = 1'b1;
  assign CLBLL_L_X2Y75_SLICE_X1Y75_B5 = 1'b1;
  assign CLBLL_L_X2Y75_SLICE_X1Y75_B6 = 1'b1;
  assign CLBLL_L_X2Y75_SLICE_X1Y75_C1 = 1'b1;
  assign CLBLL_L_X2Y75_SLICE_X1Y75_C2 = 1'b1;
  assign CLBLL_L_X2Y75_SLICE_X1Y75_C3 = 1'b1;
  assign CLBLL_L_X2Y75_SLICE_X1Y75_C4 = 1'b1;
  assign CLBLL_L_X2Y75_SLICE_X1Y75_C5 = 1'b1;
  assign CLBLL_L_X2Y75_SLICE_X1Y75_C6 = 1'b1;
  assign CLBLM_L_X10Y146_SLICE_X13Y146_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X10Y146_SLICE_X13Y146_D1 = RIOB33_X105Y133_IOB_X1Y133_I;
  assign CLBLM_L_X10Y146_SLICE_X13Y146_D2 = RIOB33_X105Y129_IOB_X1Y130_I;
  assign CLBLM_L_X10Y146_SLICE_X13Y146_D3 = RIOB33_X105Y129_IOB_X1Y129_I;
  assign CLBLM_L_X10Y146_SLICE_X13Y146_D4 = RIOB33_X105Y131_IOB_X1Y132_I;
  assign CLBLM_L_X10Y146_SLICE_X13Y146_D5 = CLBLM_L_X10Y144_SLICE_X13Y144_AQ;
  assign CLBLM_L_X10Y146_SLICE_X13Y146_D6 = 1'b1;
  assign CLBLL_L_X2Y75_SLICE_X1Y75_D1 = 1'b1;
  assign CLBLL_L_X2Y75_SLICE_X1Y75_D2 = 1'b1;
  assign CLBLL_L_X2Y75_SLICE_X1Y75_D3 = 1'b1;
  assign CLBLL_L_X2Y75_SLICE_X1Y75_D4 = 1'b1;
  assign CLBLL_L_X2Y75_SLICE_X1Y75_D5 = 1'b1;
  assign CLBLL_L_X2Y75_SLICE_X1Y75_D6 = 1'b1;
  assign CLBLM_L_X10Y146_SLICE_X12Y146_A1 = CLBLM_R_X5Y145_SLICE_X6Y145_DQ;
  assign CLBLM_L_X10Y146_SLICE_X12Y146_A2 = CLBLL_L_X4Y142_SLICE_X5Y142_DQ;
  assign CLBLM_L_X10Y146_SLICE_X12Y146_A3 = CLBLM_L_X10Y146_SLICE_X12Y146_AQ;
  assign CLBLM_L_X10Y146_SLICE_X12Y146_A4 = CLBLM_L_X8Y142_SLICE_X11Y142_AQ;
  assign CLBLM_L_X10Y146_SLICE_X12Y146_A5 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_L_X10Y146_SLICE_X12Y146_B1 = CLBLL_L_X4Y142_SLICE_X5Y142_DQ;
  assign CLBLM_L_X10Y146_SLICE_X12Y146_B2 = CLBLM_L_X10Y146_SLICE_X12Y146_BQ;
  assign CLBLM_L_X10Y146_SLICE_X12Y146_B3 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_L_X10Y146_SLICE_X12Y146_B4 = CLBLM_R_X7Y146_SLICE_X8Y146_AQ;
  assign CLBLM_L_X10Y146_SLICE_X12Y146_B5 = CLBLM_L_X10Y149_SLICE_X12Y149_AQ;
  assign CLBLM_L_X10Y146_SLICE_X12Y146_B6 = CLBLL_L_X4Y147_SLICE_X5Y147_CQ;
  assign RIOI3_X105Y189_OLOGIC_X1Y189_D1 = CLBLM_R_X103Y178_SLICE_X163Y178_AO6;
  assign CLBLM_L_X10Y146_SLICE_X12Y146_C1 = CLBLM_L_X8Y147_SLICE_X10Y147_C5Q;
  assign CLBLM_L_X10Y146_SLICE_X12Y146_C2 = CLBLM_L_X10Y146_SLICE_X12Y146_CQ;
  assign CLBLM_L_X10Y146_SLICE_X12Y146_C3 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_L_X10Y146_SLICE_X12Y146_C4 = CLBLM_L_X10Y145_SLICE_X12Y145_A5Q;
  assign CLBLM_L_X10Y146_SLICE_X12Y146_C5 = CLBLM_L_X10Y144_SLICE_X13Y144_CQ;
  assign CLBLM_L_X10Y146_SLICE_X12Y146_C6 = CLBLM_R_X7Y146_SLICE_X8Y146_AQ;
  assign RIOI3_X105Y189_OLOGIC_X1Y189_T1 = 1'b1;
  assign CLBLM_L_X10Y146_SLICE_X12Y146_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X10Y146_SLICE_X12Y146_D1 = CLBLM_L_X8Y145_SLICE_X11Y145_CQ;
  assign CLBLM_L_X10Y146_SLICE_X12Y146_D2 = CLBLM_L_X10Y146_SLICE_X12Y146_AQ;
  assign CLBLM_L_X10Y146_SLICE_X12Y146_D3 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_L_X10Y146_SLICE_X12Y146_D4 = CLBLL_L_X4Y149_SLICE_X5Y149_C5Q;
  assign CLBLM_L_X10Y146_SLICE_X12Y146_D5 = CLBLM_L_X8Y148_SLICE_X10Y148_B5Q;
  assign CLBLM_L_X10Y146_SLICE_X12Y146_D6 = 1'b1;
  assign LIOB33_X0Y127_IOB_X0Y127_O = CLBLM_R_X7Y152_SLICE_X8Y152_D5Q;
  assign LIOB33_X0Y127_IOB_X0Y128_O = CLBLM_L_X10Y145_SLICE_X12Y145_AQ;
  assign LIOI3_X0Y153_OLOGIC_X0Y154_D1 = CLBLM_R_X7Y153_SLICE_X9Y153_DQ;
  assign CLBLM_R_X11Y148_SLICE_X14Y148_A2 = CLBLM_R_X11Y150_SLICE_X15Y150_AO6;
  assign LIOI3_X0Y153_OLOGIC_X0Y154_T1 = 1'b1;
  assign CLBLL_L_X4Y143_SLICE_X4Y143_A1 = CLBLL_L_X4Y143_SLICE_X4Y143_BO5;
  assign CLBLL_L_X4Y143_SLICE_X4Y143_A2 = CLBLM_R_X5Y148_SLICE_X6Y148_BQ;
  assign CLBLL_L_X4Y143_SLICE_X4Y143_A3 = CLBLL_L_X4Y143_SLICE_X4Y143_AQ;
  assign CLBLL_L_X4Y143_SLICE_X4Y143_A4 = CLBLM_R_X3Y145_SLICE_X2Y145_CQ;
  assign CLBLL_L_X4Y143_SLICE_X4Y143_A5 = CLBLL_L_X4Y147_SLICE_X4Y147_AQ;
  assign CLBLL_L_X4Y143_SLICE_X4Y143_A6 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign LIOI3_X0Y153_OLOGIC_X0Y153_D1 = CLBLM_L_X8Y153_SLICE_X10Y153_A5Q;
  assign CLBLL_L_X4Y143_SLICE_X4Y143_AX = CLBLM_R_X3Y143_SLICE_X2Y143_CO6;
  assign CLBLL_L_X4Y143_SLICE_X4Y143_B1 = CLBLM_R_X5Y143_SLICE_X6Y143_CQ;
  assign CLBLL_L_X4Y143_SLICE_X4Y143_B2 = CLBLL_L_X4Y143_SLICE_X4Y143_BQ;
  assign CLBLL_L_X4Y143_SLICE_X4Y143_B3 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLL_L_X4Y143_SLICE_X4Y143_B4 = CLBLM_R_X3Y145_SLICE_X2Y145_CQ;
  assign CLBLL_L_X4Y143_SLICE_X4Y143_B5 = CLBLM_R_X5Y145_SLICE_X6Y145_D5Q;
  assign CLBLL_L_X4Y143_SLICE_X4Y143_B6 = 1'b1;
  assign CLBLL_L_X4Y143_SLICE_X4Y143_C1 = RIOB33_X105Y121_IOB_X1Y122_I;
  assign CLBLL_L_X4Y143_SLICE_X4Y143_C2 = CLBLL_L_X4Y143_SLICE_X4Y143_CQ;
  assign CLBLL_L_X4Y143_SLICE_X4Y143_C3 = CLBLL_L_X2Y145_SLICE_X1Y145_AQ;
  assign CLBLL_L_X4Y143_SLICE_X4Y143_C4 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLL_L_X4Y143_SLICE_X4Y143_C5 = CLBLL_L_X4Y146_SLICE_X4Y146_CQ;
  assign CLBLL_L_X4Y143_SLICE_X4Y143_C6 = 1'b1;
  assign CLBLL_L_X4Y143_SLICE_X4Y143_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLL_L_X4Y143_SLICE_X4Y143_D1 = CLBLM_R_X7Y149_SLICE_X9Y149_AQ;
  assign CLBLL_L_X4Y143_SLICE_X4Y143_D2 = CLBLM_R_X5Y146_SLICE_X7Y146_C5Q;
  assign CLBLL_L_X4Y143_SLICE_X4Y143_D3 = CLBLL_L_X4Y143_SLICE_X4Y143_DQ;
  assign CLBLL_L_X4Y143_SLICE_X4Y143_D4 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLL_L_X4Y143_SLICE_X4Y143_D5 = CLBLM_R_X5Y141_SLICE_X6Y141_BQ;
  assign CLBLL_L_X4Y143_SLICE_X4Y143_D6 = 1'b1;
  assign RIOI3_X105Y127_ILOGIC_X1Y128_D = RIOB33_X105Y127_IOB_X1Y128_I;
  assign RIOI3_X105Y127_ILOGIC_X1Y127_D = RIOB33_X105Y127_IOB_X1Y127_I;
  assign LIOI3_X0Y153_OLOGIC_X0Y153_T1 = 1'b1;
  assign CLBLL_L_X4Y143_SLICE_X5Y143_A1 = CLBLL_L_X4Y144_SLICE_X5Y144_DQ;
  assign CLBLL_L_X4Y143_SLICE_X5Y143_A2 = CLBLL_L_X4Y151_SLICE_X4Y151_BQ;
  assign CLBLL_L_X4Y143_SLICE_X5Y143_A3 = CLBLL_L_X4Y143_SLICE_X5Y143_AQ;
  assign CLBLL_L_X4Y143_SLICE_X5Y143_A4 = CLBLM_R_X3Y145_SLICE_X3Y145_D5Q;
  assign CLBLL_L_X4Y143_SLICE_X5Y143_A5 = CLBLL_L_X4Y143_SLICE_X5Y143_B5Q;
  assign CLBLL_L_X4Y143_SLICE_X5Y143_A6 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLL_L_X4Y143_SLICE_X5Y143_B1 = LIOB33_X0Y59_IOB_X0Y59_I;
  assign CLBLL_L_X4Y143_SLICE_X5Y143_B2 = CLBLM_R_X5Y144_SLICE_X7Y144_BQ;
  assign CLBLL_L_X4Y143_SLICE_X5Y143_B3 = CLBLM_R_X7Y151_SLICE_X8Y151_C5Q;
  assign CLBLL_L_X4Y143_SLICE_X5Y143_B4 = CLBLM_R_X5Y143_SLICE_X7Y143_BQ;
  assign CLBLL_L_X4Y143_SLICE_X5Y143_B5 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLL_L_X4Y143_SLICE_X5Y143_B6 = 1'b1;
  assign RIOI3_TBYTESRC_X105Y131_ILOGIC_X1Y132_D = RIOB33_X105Y131_IOB_X1Y132_I;
  assign CLBLL_L_X4Y143_SLICE_X5Y143_C1 = CLBLL_L_X4Y143_SLICE_X4Y143_AQ;
  assign CLBLL_L_X4Y143_SLICE_X5Y143_C2 = CLBLM_R_X5Y145_SLICE_X6Y145_D5Q;
  assign CLBLL_L_X4Y143_SLICE_X5Y143_C3 = CLBLL_L_X4Y148_SLICE_X5Y148_DQ;
  assign CLBLL_L_X4Y143_SLICE_X5Y143_C4 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLL_L_X4Y143_SLICE_X5Y143_C5 = CLBLL_L_X4Y143_SLICE_X4Y143_BQ;
  assign CLBLL_L_X4Y143_SLICE_X5Y143_C6 = 1'b1;
  assign RIOI3_TBYTESRC_X105Y131_ILOGIC_X1Y131_D = RIOB33_X105Y131_IOB_X1Y131_I;
  assign CLBLL_L_X4Y143_SLICE_X5Y143_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X10Y147_SLICE_X13Y147_A1 = CLBLM_L_X10Y146_SLICE_X13Y146_DO5;
  assign CLBLM_L_X10Y147_SLICE_X13Y147_A2 = CLBLM_L_X10Y145_SLICE_X13Y145_BO6;
  assign CLBLM_L_X10Y147_SLICE_X13Y147_A3 = CLBLM_L_X10Y147_SLICE_X13Y147_AQ;
  assign CLBLM_L_X10Y147_SLICE_X13Y147_A4 = CLBLM_R_X7Y147_SLICE_X9Y147_A5Q;
  assign CLBLM_L_X10Y147_SLICE_X13Y147_A5 = RIOB33_X105Y131_IOB_X1Y132_I;
  assign CLBLL_L_X4Y143_SLICE_X5Y143_D1 = 1'b1;
  assign CLBLL_L_X4Y143_SLICE_X5Y143_D2 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLL_L_X4Y143_SLICE_X5Y143_D3 = LIOB33_X0Y63_IOB_X0Y63_I;
  assign CLBLL_L_X4Y143_SLICE_X5Y143_D4 = CLBLL_L_X4Y151_SLICE_X4Y151_AQ;
  assign CLBLL_L_X4Y143_SLICE_X5Y143_D5 = CLBLL_L_X4Y144_SLICE_X5Y144_DQ;
  assign CLBLL_L_X4Y143_SLICE_X5Y143_D6 = 1'b1;
  assign CLBLM_L_X10Y147_SLICE_X13Y147_A6 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_L_X10Y147_SLICE_X13Y147_B1 = CLBLM_L_X10Y146_SLICE_X12Y146_DQ;
  assign CLBLM_L_X10Y147_SLICE_X13Y147_B2 = CLBLM_R_X5Y142_SLICE_X6Y142_D5Q;
  assign CLBLM_L_X10Y147_SLICE_X13Y147_B5 = CLBLL_L_X4Y148_SLICE_X4Y148_CQ;
  assign CLBLM_L_X10Y147_SLICE_X13Y147_B6 = CLBLM_R_X7Y149_SLICE_X8Y149_AQ;
  assign CLBLM_L_X10Y147_SLICE_X13Y147_C1 = CLBLM_L_X8Y148_SLICE_X11Y148_CO6;
  assign CLBLM_L_X10Y147_SLICE_X13Y147_C2 = CLBLM_L_X8Y145_SLICE_X10Y145_CO6;
  assign CLBLM_L_X10Y147_SLICE_X13Y147_C3 = CLBLM_R_X11Y145_SLICE_X14Y145_DO6;
  assign CLBLM_L_X10Y147_SLICE_X13Y147_C4 = CLBLM_L_X10Y150_SLICE_X13Y150_DO6;
  assign CLBLM_L_X10Y147_SLICE_X13Y147_C5 = CLBLM_L_X8Y147_SLICE_X10Y147_DO6;
  assign CLBLM_L_X10Y147_SLICE_X13Y147_C6 = CLBLM_L_X12Y147_SLICE_X16Y147_DO6;
  assign CLBLM_L_X10Y147_SLICE_X13Y147_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign RIOI3_X105Y155_OLOGIC_X1Y156_D1 = 1'b1;
  assign CLBLM_L_X10Y147_SLICE_X13Y147_D1 = CLBLM_L_X8Y147_SLICE_X11Y147_C5Q;
  assign CLBLM_L_X10Y147_SLICE_X13Y147_D2 = CLBLM_L_X10Y143_SLICE_X13Y143_CQ;
  assign CLBLM_L_X10Y147_SLICE_X13Y147_D3 = CLBLM_R_X7Y144_SLICE_X9Y144_B5Q;
  assign CLBLM_L_X10Y147_SLICE_X13Y147_D4 = 1'b1;
  assign CLBLM_L_X10Y147_SLICE_X13Y147_D5 = CLBLM_R_X7Y153_SLICE_X8Y153_A5Q;
  assign CLBLM_L_X10Y147_SLICE_X13Y147_D6 = CLBLM_R_X11Y147_SLICE_X15Y147_BO6;
  assign CLBLM_L_X10Y147_SLICE_X12Y147_A1 = CLBLL_L_X4Y142_SLICE_X5Y142_DQ;
  assign CLBLM_L_X10Y147_SLICE_X12Y147_A2 = CLBLL_L_X4Y147_SLICE_X5Y147_CQ;
  assign CLBLM_L_X10Y147_SLICE_X12Y147_A3 = 1'b1;
  assign CLBLM_L_X10Y147_SLICE_X12Y147_A4 = CLBLM_L_X10Y146_SLICE_X13Y146_DO6;
  assign CLBLM_L_X10Y147_SLICE_X12Y147_A5 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_L_X10Y147_SLICE_X12Y147_A6 = 1'b1;
  assign CLBLM_R_X3Y142_SLICE_X2Y142_B1 = CLBLL_L_X4Y142_SLICE_X4Y142_BQ;
  assign LIOB33_X0Y129_IOB_X0Y130_O = CLBLL_L_X2Y145_SLICE_X0Y145_BQ;
  assign CLBLM_R_X3Y142_SLICE_X2Y142_B2 = CLBLM_R_X3Y142_SLICE_X3Y142_AQ;
  assign CLBLM_L_X10Y147_SLICE_X12Y147_AX = CLBLM_L_X8Y146_SLICE_X10Y146_AQ;
  assign LIOB33_X0Y129_IOB_X0Y129_O = CLBLL_L_X2Y146_SLICE_X0Y146_CQ;
  assign CLBLM_L_X10Y147_SLICE_X12Y147_B1 = CLBLM_R_X7Y153_SLICE_X8Y153_A5Q;
  assign CLBLM_L_X10Y147_SLICE_X12Y147_B2 = CLBLM_R_X7Y153_SLICE_X9Y153_A5Q;
  assign CLBLM_L_X10Y147_SLICE_X12Y147_B3 = CLBLM_R_X11Y147_SLICE_X15Y147_BO6;
  assign CLBLM_L_X10Y147_SLICE_X12Y147_B4 = CLBLM_R_X7Y144_SLICE_X9Y144_B5Q;
  assign CLBLM_L_X10Y147_SLICE_X12Y147_B5 = CLBLM_L_X10Y144_SLICE_X12Y144_AQ;
  assign CLBLM_L_X10Y147_SLICE_X12Y147_B6 = 1'b1;
  assign CLBLM_R_X3Y142_SLICE_X2Y142_B4 = CLBLM_R_X3Y143_SLICE_X2Y143_AQ;
  assign CLBLM_L_X10Y147_SLICE_X12Y147_BX = CLBLM_R_X7Y143_SLICE_X9Y143_BQ;
  assign CLBLM_L_X10Y147_SLICE_X12Y147_C1 = RIOB33_X105Y131_IOB_X1Y131_I;
  assign CLBLM_L_X10Y147_SLICE_X12Y147_C2 = CLBLL_L_X4Y153_SLICE_X5Y153_A5Q;
  assign CLBLM_L_X10Y147_SLICE_X12Y147_C3 = CLBLL_L_X4Y150_SLICE_X5Y150_A5Q;
  assign CLBLM_L_X10Y147_SLICE_X12Y147_C4 = CLBLM_R_X5Y142_SLICE_X7Y142_CO6;
  assign CLBLM_L_X10Y147_SLICE_X12Y147_C5 = CLBLM_L_X8Y145_SLICE_X11Y145_DQ;
  assign CLBLM_L_X10Y147_SLICE_X12Y147_C6 = CLBLM_L_X10Y149_SLICE_X12Y149_BO6;
  assign CLBLM_L_X10Y147_SLICE_X12Y147_CE = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_L_X10Y147_SLICE_X12Y147_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X10Y147_SLICE_X12Y147_CX = CLBLL_L_X4Y143_SLICE_X5Y143_AQ;
  assign CLBLM_L_X10Y147_SLICE_X12Y147_D1 = CLBLL_L_X4Y148_SLICE_X4Y148_CQ;
  assign CLBLM_L_X10Y147_SLICE_X12Y147_D2 = CLBLM_L_X10Y151_SLICE_X13Y151_AQ;
  assign CLBLM_L_X10Y147_SLICE_X12Y147_D3 = CLBLM_L_X12Y146_SLICE_X16Y146_CO6;
  assign CLBLM_L_X10Y147_SLICE_X12Y147_D4 = CLBLM_L_X10Y148_SLICE_X12Y148_AO5;
  assign CLBLM_L_X10Y147_SLICE_X12Y147_D5 = CLBLM_R_X7Y145_SLICE_X9Y145_AO6;
  assign CLBLM_L_X10Y147_SLICE_X12Y147_D6 = CLBLM_L_X8Y152_SLICE_X11Y152_D5Q;
  assign RIOI3_X105Y155_OLOGIC_X1Y156_T1 = 1'b1;
  assign CLBLL_L_X4Y144_SLICE_X4Y144_A1 = CLBLL_L_X2Y145_SLICE_X0Y145_BQ;
  assign CLBLL_L_X4Y144_SLICE_X4Y144_A2 = CLBLL_L_X4Y144_SLICE_X4Y144_BQ;
  assign CLBLL_L_X4Y144_SLICE_X4Y144_A3 = CLBLL_L_X4Y144_SLICE_X4Y144_AQ;
  assign CLBLL_L_X4Y144_SLICE_X4Y144_A4 = CLBLM_R_X7Y152_SLICE_X8Y152_D5Q;
  assign CLBLL_L_X4Y144_SLICE_X4Y144_A5 = CLBLM_R_X7Y142_SLICE_X8Y142_C5Q;
  assign CLBLL_L_X4Y144_SLICE_X4Y144_A6 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLL_L_X4Y144_SLICE_X4Y144_B1 = CLBLM_R_X5Y145_SLICE_X6Y145_B5Q;
  assign CLBLL_L_X4Y144_SLICE_X4Y144_B2 = CLBLL_L_X4Y150_SLICE_X4Y150_B5Q;
  assign CLBLL_L_X4Y144_SLICE_X4Y144_B3 = CLBLL_L_X4Y144_SLICE_X4Y144_CQ;
  assign CLBLL_L_X4Y144_SLICE_X4Y144_B4 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLL_L_X4Y144_SLICE_X4Y144_B5 = CLBLM_R_X5Y144_SLICE_X7Y144_BQ;
  assign CLBLL_L_X4Y144_SLICE_X4Y144_B6 = 1'b1;
  assign CLBLL_L_X4Y144_SLICE_X4Y144_C1 = CLBLM_L_X8Y145_SLICE_X11Y145_C5Q;
  assign CLBLL_L_X4Y144_SLICE_X4Y144_C2 = CLBLL_L_X4Y144_SLICE_X5Y144_BQ;
  assign CLBLL_L_X4Y144_SLICE_X4Y144_C3 = CLBLL_L_X4Y147_SLICE_X4Y147_BQ;
  assign CLBLL_L_X4Y144_SLICE_X4Y144_C4 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLL_L_X4Y144_SLICE_X4Y144_C5 = CLBLL_L_X4Y147_SLICE_X5Y147_B5Q;
  assign CLBLL_L_X4Y144_SLICE_X4Y144_C6 = 1'b1;
  assign CLBLL_L_X4Y144_SLICE_X4Y144_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLL_L_X4Y144_SLICE_X4Y144_D1 = CLBLL_L_X4Y140_SLICE_X5Y140_AQ;
  assign CLBLL_L_X4Y144_SLICE_X4Y144_D2 = 1'b1;
  assign CLBLL_L_X4Y144_SLICE_X4Y144_D3 = CLBLM_R_X3Y146_SLICE_X2Y146_CQ;
  assign CLBLL_L_X4Y144_SLICE_X4Y144_D4 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLL_L_X4Y144_SLICE_X4Y144_D5 = CLBLM_L_X12Y151_SLICE_X16Y151_AQ;
  assign CLBLL_L_X4Y144_SLICE_X4Y144_D6 = 1'b1;
  assign CLBLL_L_X4Y144_SLICE_X5Y144_A1 = CLBLL_L_X4Y142_SLICE_X5Y142_DQ;
  assign CLBLL_L_X4Y144_SLICE_X5Y144_A2 = CLBLL_L_X4Y148_SLICE_X5Y148_DQ;
  assign CLBLL_L_X4Y144_SLICE_X5Y144_A3 = CLBLL_L_X4Y144_SLICE_X5Y144_AQ;
  assign CLBLL_L_X4Y144_SLICE_X5Y144_A4 = CLBLL_L_X4Y142_SLICE_X5Y142_D5Q;
  assign CLBLL_L_X4Y144_SLICE_X5Y144_A5 = CLBLL_L_X4Y147_SLICE_X5Y147_CQ;
  assign CLBLL_L_X4Y144_SLICE_X5Y144_A6 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLL_L_X4Y144_SLICE_X5Y144_B1 = CLBLM_R_X11Y146_SLICE_X15Y146_AO6;
  assign CLBLL_L_X4Y144_SLICE_X5Y144_B2 = CLBLL_L_X4Y152_SLICE_X4Y152_B5Q;
  assign CLBLL_L_X4Y144_SLICE_X5Y144_B3 = CLBLL_L_X4Y147_SLICE_X5Y147_BQ;
  assign CLBLL_L_X4Y144_SLICE_X5Y144_B4 = CLBLL_L_X4Y144_SLICE_X5Y144_CQ;
  assign CLBLL_L_X4Y144_SLICE_X5Y144_B5 = CLBLM_L_X8Y148_SLICE_X11Y148_AQ;
  assign CLBLL_L_X4Y144_SLICE_X5Y144_B6 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLL_L_X4Y144_SLICE_X5Y144_C1 = CLBLL_L_X4Y147_SLICE_X5Y147_BQ;
  assign CLBLL_L_X4Y144_SLICE_X5Y144_C2 = CLBLL_L_X4Y144_SLICE_X5Y144_CQ;
  assign CLBLL_L_X4Y144_SLICE_X5Y144_C3 = CLBLM_R_X5Y145_SLICE_X6Y145_B5Q;
  assign CLBLL_L_X4Y144_SLICE_X5Y144_C4 = CLBLM_R_X11Y146_SLICE_X15Y146_AO6;
  assign CLBLL_L_X4Y144_SLICE_X5Y144_C5 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLL_L_X4Y144_SLICE_X5Y144_C6 = CLBLM_R_X3Y145_SLICE_X3Y145_D5Q;
  assign CLBLL_L_X4Y144_SLICE_X5Y144_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X10Y148_SLICE_X13Y148_A1 = CLBLM_L_X10Y148_SLICE_X13Y148_CQ;
  assign CLBLL_L_X4Y144_SLICE_X5Y144_D1 = CLBLM_L_X10Y145_SLICE_X12Y145_AQ;
  assign CLBLM_L_X10Y148_SLICE_X13Y148_A3 = CLBLM_L_X10Y148_SLICE_X13Y148_AQ;
  assign CLBLM_L_X10Y148_SLICE_X13Y148_A4 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLL_L_X4Y144_SLICE_X5Y144_D2 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_L_X10Y148_SLICE_X13Y148_A6 = CLBLM_R_X5Y142_SLICE_X7Y142_BQ;
  assign CLBLL_L_X4Y144_SLICE_X5Y144_D3 = 1'b1;
  assign CLBLL_L_X4Y144_SLICE_X5Y144_D4 = CLBLL_L_X4Y145_SLICE_X5Y145_BQ;
  assign CLBLL_L_X4Y144_SLICE_X5Y144_D5 = CLBLL_L_X4Y144_SLICE_X5Y144_AQ;
  assign CLBLL_L_X4Y144_SLICE_X5Y144_D6 = 1'b1;
  assign CLBLM_L_X10Y148_SLICE_X13Y148_A5 = CLBLM_L_X10Y148_SLICE_X12Y148_AQ;
  assign CLBLM_L_X10Y148_SLICE_X13Y148_B3 = CLBLM_L_X8Y147_SLICE_X11Y147_BQ;
  assign CLBLM_L_X10Y148_SLICE_X13Y148_B4 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_L_X10Y148_SLICE_X13Y148_B5 = CLBLM_R_X13Y149_SLICE_X18Y149_AO6;
  assign CLBLM_L_X10Y148_SLICE_X13Y148_B6 = CLBLM_R_X7Y151_SLICE_X8Y151_BQ;
  assign CLBLM_L_X10Y148_SLICE_X13Y148_B1 = 1'b1;
  assign CLBLM_L_X10Y148_SLICE_X13Y148_B2 = CLBLM_L_X10Y148_SLICE_X13Y148_BQ;
  assign CLBLM_L_X10Y148_SLICE_X13Y148_C1 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_L_X10Y148_SLICE_X13Y148_C2 = CLBLM_R_X3Y151_SLICE_X3Y151_CQ;
  assign CLBLM_L_X10Y148_SLICE_X13Y148_C3 = 1'b1;
  assign CLBLM_L_X10Y148_SLICE_X13Y148_C4 = CLBLM_L_X8Y143_SLICE_X11Y143_D5Q;
  assign CLBLM_L_X10Y148_SLICE_X13Y148_C5 = CLBLM_L_X12Y146_SLICE_X16Y146_DQ;
  assign CLBLM_L_X10Y148_SLICE_X13Y148_C6 = 1'b1;
  assign LIOB33_X0Y131_IOB_X0Y131_O = CLBLL_L_X2Y75_SLICE_X0Y75_AO6;
  assign LIOB33_X0Y131_IOB_X0Y132_O = CLBLM_R_X3Y143_SLICE_X2Y143_BO5;
  assign CLBLM_L_X10Y148_SLICE_X13Y148_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X10Y148_SLICE_X13Y148_D1 = CLBLM_L_X10Y142_SLICE_X13Y142_BO6;
  assign CLBLM_L_X10Y148_SLICE_X13Y148_D2 = CLBLM_L_X12Y145_SLICE_X17Y145_BO6;
  assign CLBLM_L_X10Y148_SLICE_X13Y148_D3 = CLBLM_R_X5Y148_SLICE_X6Y148_DO6;
  assign CLBLM_L_X10Y148_SLICE_X13Y148_D4 = CLBLM_R_X3Y142_SLICE_X2Y142_BO5;
  assign CLBLM_L_X10Y148_SLICE_X13Y148_D5 = CLBLM_L_X10Y144_SLICE_X13Y144_A5Q;
  assign CLBLM_L_X10Y148_SLICE_X13Y148_D6 = CLBLM_R_X11Y152_SLICE_X14Y152_AO6;
  assign CLBLM_L_X10Y148_SLICE_X12Y148_A1 = CLBLM_R_X7Y153_SLICE_X8Y153_A5Q;
  assign CLBLM_L_X10Y148_SLICE_X12Y148_A2 = CLBLM_R_X7Y149_SLICE_X8Y149_AQ;
  assign CLBLM_L_X10Y148_SLICE_X12Y148_A3 = CLBLL_L_X4Y148_SLICE_X4Y148_CQ;
  assign CLBLM_L_X10Y148_SLICE_X12Y148_A4 = CLBLM_R_X7Y146_SLICE_X9Y146_CO6;
  assign CLBLM_L_X10Y148_SLICE_X12Y148_A5 = CLBLM_R_X7Y144_SLICE_X9Y144_B5Q;
  assign CLBLM_L_X10Y148_SLICE_X12Y148_A6 = 1'b1;
  assign CLBLM_L_X10Y148_SLICE_X12Y148_AX = CLBLM_L_X10Y147_SLICE_X12Y147_AO6;
  assign CLBLM_L_X10Y148_SLICE_X12Y148_B1 = CLBLM_R_X7Y149_SLICE_X8Y149_AQ;
  assign CLBLM_L_X10Y148_SLICE_X12Y148_B2 = CLBLM_L_X12Y147_SLICE_X16Y147_DO6;
  assign CLBLM_L_X10Y148_SLICE_X12Y148_B3 = CLBLM_R_X5Y146_SLICE_X6Y146_B5Q;
  assign CLBLM_L_X10Y148_SLICE_X12Y148_B4 = CLBLM_L_X10Y148_SLICE_X13Y148_BQ;
  assign CLBLM_L_X10Y148_SLICE_X12Y148_B5 = CLBLM_L_X10Y147_SLICE_X12Y147_BO6;
  assign CLBLM_L_X10Y148_SLICE_X12Y148_B6 = CLBLL_L_X4Y148_SLICE_X4Y148_CQ;
  assign CLBLM_L_X10Y148_SLICE_X12Y148_C1 = CLBLM_R_X7Y148_SLICE_X9Y148_BQ;
  assign CLBLM_L_X10Y148_SLICE_X12Y148_C2 = CLBLM_L_X10Y149_SLICE_X13Y149_CO6;
  assign CLBLM_L_X10Y148_SLICE_X12Y148_C3 = CLBLM_L_X10Y151_SLICE_X13Y151_BO6;
  assign CLBLM_L_X10Y148_SLICE_X12Y148_C4 = CLBLM_L_X10Y147_SLICE_X12Y147_BO5;
  assign CLBLM_L_X10Y148_SLICE_X12Y148_C5 = CLBLM_L_X12Y149_SLICE_X17Y149_BO5;
  assign CLBLM_L_X10Y148_SLICE_X12Y148_C6 = CLBLM_R_X5Y146_SLICE_X6Y146_AQ;
  assign CLBLM_L_X10Y148_SLICE_X12Y148_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X10Y148_SLICE_X12Y148_D1 = CLBLM_L_X8Y147_SLICE_X11Y147_CQ;
  assign CLBLM_L_X10Y148_SLICE_X12Y148_D2 = CLBLL_L_X4Y148_SLICE_X4Y148_CQ;
  assign CLBLM_L_X10Y148_SLICE_X12Y148_D3 = CLBLM_L_X10Y153_SLICE_X13Y153_A5Q;
  assign CLBLM_L_X10Y148_SLICE_X12Y148_D4 = CLBLM_L_X10Y148_SLICE_X12Y148_AO5;
  assign CLBLM_L_X10Y148_SLICE_X12Y148_D5 = 1'b1;
  assign CLBLM_L_X10Y148_SLICE_X12Y148_D6 = CLBLM_L_X12Y146_SLICE_X16Y146_CO6;
  assign LIOI3_X0Y147_OLOGIC_X0Y148_D1 = CLBLL_L_X2Y147_SLICE_X1Y147_AO6;
  assign LIOI3_X0Y147_OLOGIC_X0Y148_T1 = 1'b1;
  assign RIOI3_X105Y191_OLOGIC_X1Y192_D1 = CLBLM_L_X12Y153_SLICE_X16Y153_AO6;
  assign CLBLM_R_X11Y147_SLICE_X15Y147_D4 = 1'b1;
  assign LIOI3_X0Y147_OLOGIC_X0Y147_D1 = CLBLM_R_X5Y141_SLICE_X6Y141_CO5;
  assign CLBLM_R_X11Y147_SLICE_X15Y147_D5 = CLBLM_R_X11Y144_SLICE_X14Y144_DO6;
  assign RIOI3_X105Y191_OLOGIC_X1Y192_T1 = 1'b1;
  assign CLBLM_R_X11Y147_SLICE_X15Y147_D6 = CLBLM_R_X11Y145_SLICE_X14Y145_CO6;
  assign LIOI3_X0Y147_OLOGIC_X0Y147_T1 = 1'b1;
  assign RIOI3_X105Y191_OLOGIC_X1Y191_D1 = CLBLM_L_X12Y149_SLICE_X17Y149_AO5;
  assign RIOI3_X105Y191_OLOGIC_X1Y191_T1 = 1'b1;
  assign CLBLM_R_X11Y147_SLICE_X14Y147_A1 = CLBLM_R_X7Y153_SLICE_X8Y153_A5Q;
  assign CLBLL_L_X4Y145_SLICE_X4Y145_A1 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLL_L_X4Y145_SLICE_X4Y145_A2 = CLBLL_L_X4Y145_SLICE_X4Y145_BQ;
  assign CLBLL_L_X4Y145_SLICE_X4Y145_A3 = CLBLL_L_X4Y145_SLICE_X4Y145_AQ;
  assign CLBLL_L_X4Y145_SLICE_X4Y145_A4 = CLBLM_R_X7Y142_SLICE_X8Y142_C5Q;
  assign CLBLL_L_X4Y145_SLICE_X4Y145_A5 = CLBLM_L_X8Y149_SLICE_X11Y149_AQ;
  assign CLBLL_L_X4Y145_SLICE_X4Y145_A6 = CLBLM_R_X7Y152_SLICE_X8Y152_D5Q;
  assign CLBLM_R_X11Y147_SLICE_X14Y147_A2 = CLBLM_L_X12Y147_SLICE_X16Y147_DO6;
  assign CLBLM_R_X11Y147_SLICE_X14Y147_A3 = CLBLM_R_X7Y149_SLICE_X8Y149_AQ;
  assign CLBLL_L_X4Y145_SLICE_X4Y145_B1 = CLBLL_L_X4Y151_SLICE_X5Y151_CQ;
  assign CLBLL_L_X4Y145_SLICE_X4Y145_B2 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLL_L_X4Y145_SLICE_X4Y145_B3 = CLBLL_L_X4Y146_SLICE_X4Y146_AQ;
  assign CLBLL_L_X4Y145_SLICE_X4Y145_B4 = CLBLM_R_X5Y141_SLICE_X6Y141_B5Q;
  assign CLBLL_L_X4Y145_SLICE_X4Y145_B5 = 1'b1;
  assign CLBLL_L_X4Y145_SLICE_X4Y145_B6 = 1'b1;
  assign CLBLL_L_X4Y145_SLICE_X4Y145_C1 = CLBLM_R_X3Y148_SLICE_X2Y148_A5Q;
  assign CLBLL_L_X4Y145_SLICE_X4Y145_C2 = CLBLL_L_X4Y145_SLICE_X4Y145_CQ;
  assign CLBLL_L_X4Y145_SLICE_X4Y145_C3 = CLBLM_R_X5Y148_SLICE_X6Y148_CQ;
  assign CLBLL_L_X4Y145_SLICE_X4Y145_C4 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLL_L_X4Y145_SLICE_X4Y145_C5 = CLBLM_L_X10Y153_SLICE_X13Y153_A5Q;
  assign CLBLL_L_X4Y145_SLICE_X4Y145_C6 = 1'b1;
  assign CLBLL_L_X4Y145_SLICE_X4Y145_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLL_L_X4Y145_SLICE_X4Y145_D1 = CLBLL_L_X4Y143_SLICE_X4Y143_AQ;
  assign CLBLL_L_X4Y145_SLICE_X4Y145_D2 = CLBLL_L_X4Y151_SLICE_X4Y151_AQ;
  assign CLBLL_L_X4Y145_SLICE_X4Y145_D3 = CLBLL_L_X4Y151_SLICE_X5Y151_CQ;
  assign CLBLL_L_X4Y145_SLICE_X4Y145_D4 = CLBLM_R_X5Y145_SLICE_X6Y145_D5Q;
  assign CLBLL_L_X4Y145_SLICE_X4Y145_D5 = CLBLL_L_X4Y143_SLICE_X4Y143_BQ;
  assign CLBLL_L_X4Y145_SLICE_X4Y145_D6 = 1'b1;
  assign CLBLL_L_X4Y145_SLICE_X5Y145_A1 = CLBLM_R_X3Y146_SLICE_X2Y146_DQ;
  assign CLBLL_L_X4Y145_SLICE_X5Y145_A2 = CLBLM_L_X10Y144_SLICE_X13Y144_CQ;
  assign CLBLL_L_X4Y145_SLICE_X5Y145_A3 = CLBLL_L_X4Y145_SLICE_X5Y145_AQ;
  assign CLBLL_L_X4Y145_SLICE_X5Y145_A4 = CLBLM_R_X7Y145_SLICE_X8Y145_C5Q;
  assign CLBLL_L_X4Y145_SLICE_X5Y145_A5 = CLBLM_L_X8Y147_SLICE_X10Y147_C5Q;
  assign CLBLL_L_X4Y145_SLICE_X5Y145_A6 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLL_L_X4Y145_SLICE_X5Y145_B1 = CLBLL_L_X4Y145_SLICE_X5Y145_DO6;
  assign CLBLL_L_X4Y145_SLICE_X5Y145_B2 = CLBLL_L_X4Y145_SLICE_X5Y145_BQ;
  assign CLBLL_L_X4Y145_SLICE_X5Y145_B3 = CLBLL_L_X4Y147_SLICE_X5Y147_DO6;
  assign CLBLL_L_X4Y145_SLICE_X5Y145_B4 = CLBLM_R_X5Y145_SLICE_X7Y145_AQ;
  assign CLBLL_L_X4Y145_SLICE_X5Y145_B5 = CLBLM_R_X3Y145_SLICE_X2Y145_CQ;
  assign CLBLL_L_X4Y145_SLICE_X5Y145_B6 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLL_L_X4Y145_SLICE_X5Y145_C1 = CLBLM_R_X5Y147_SLICE_X6Y147_C5Q;
  assign CLBLL_L_X4Y145_SLICE_X5Y145_C2 = CLBLL_L_X4Y145_SLICE_X4Y145_C5Q;
  assign CLBLL_L_X4Y145_SLICE_X5Y145_C3 = CLBLM_R_X5Y146_SLICE_X7Y146_DQ;
  assign CLBLL_L_X4Y145_SLICE_X5Y145_C4 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLL_L_X4Y145_SLICE_X5Y145_C5 = CLBLM_R_X7Y153_SLICE_X9Y153_CQ;
  assign CLBLL_L_X4Y145_SLICE_X5Y145_C6 = 1'b1;
  assign LIOB33_X0Y147_IOB_X0Y147_O = CLBLM_R_X5Y141_SLICE_X6Y141_CO5;
  assign LIOB33_X0Y147_IOB_X0Y148_O = CLBLL_L_X2Y147_SLICE_X1Y147_AO6;
  assign CLBLL_L_X4Y145_SLICE_X5Y145_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign LIOB33_X0Y133_IOB_X0Y134_O = CLBLL_L_X2Y145_SLICE_X0Y145_BQ;
  assign LIOB33_X0Y133_IOB_X0Y133_O = CLBLL_L_X4Y140_SLICE_X4Y140_BO5;
  assign CLBLL_L_X4Y145_SLICE_X5Y145_D1 = CLBLM_R_X3Y145_SLICE_X3Y145_BQ;
  assign CLBLL_L_X4Y145_SLICE_X5Y145_D2 = CLBLM_R_X5Y152_SLICE_X6Y152_DQ;
  assign CLBLL_L_X4Y145_SLICE_X5Y145_D3 = CLBLL_L_X4Y151_SLICE_X5Y151_CQ;
  assign CLBLL_L_X4Y145_SLICE_X5Y145_D4 = CLBLL_L_X4Y143_SLICE_X5Y143_CO5;
  assign CLBLL_L_X4Y145_SLICE_X5Y145_D5 = CLBLM_R_X5Y152_SLICE_X6Y152_CQ;
  assign CLBLL_L_X4Y145_SLICE_X5Y145_D6 = CLBLL_L_X4Y151_SLICE_X4Y151_AQ;
  assign CLBLM_L_X10Y149_SLICE_X13Y149_A1 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_L_X10Y149_SLICE_X13Y149_A2 = CLBLM_L_X10Y147_SLICE_X13Y147_CO6;
  assign CLBLM_L_X10Y149_SLICE_X13Y149_A3 = CLBLM_L_X10Y148_SLICE_X12Y148_AQ;
  assign CLBLM_L_X10Y149_SLICE_X13Y149_A4 = CLBLM_R_X7Y145_SLICE_X8Y145_AQ;
  assign CLBLM_L_X10Y149_SLICE_X13Y149_A5 = 1'b1;
  assign CLBLM_L_X10Y149_SLICE_X13Y149_A6 = 1'b1;
  assign CLBLM_L_X10Y149_SLICE_X13Y149_B1 = CLBLL_L_X4Y151_SLICE_X4Y151_CQ;
  assign CLBLM_L_X10Y149_SLICE_X13Y149_B2 = RIOB33_X105Y101_IOB_X1Y101_I;
  assign CLBLM_L_X10Y149_SLICE_X13Y149_B3 = CLBLM_L_X8Y142_SLICE_X11Y142_BQ;
  assign CLBLM_L_X10Y149_SLICE_X13Y149_B4 = CLBLM_L_X10Y149_SLICE_X12Y149_BO5;
  assign CLBLM_L_X10Y149_SLICE_X13Y149_B5 = RIOB33_SING_X105Y100_IOB_X1Y100_I;
  assign CLBLM_L_X10Y149_SLICE_X13Y149_B6 = RIOB33_X105Y131_IOB_X1Y131_I;
  assign CLBLM_R_X7Y149_SLICE_X9Y149_D4 = CLBLM_R_X7Y144_SLICE_X9Y144_B5Q;
  assign CLBLM_L_X10Y149_SLICE_X13Y149_C1 = CLBLM_R_X11Y144_SLICE_X14Y144_CO6;
  assign CLBLM_L_X10Y149_SLICE_X13Y149_C2 = CLBLM_L_X10Y150_SLICE_X13Y150_AQ;
  assign CLBLM_L_X10Y149_SLICE_X13Y149_C3 = CLBLM_R_X7Y151_SLICE_X8Y151_DQ;
  assign CLBLM_L_X10Y149_SLICE_X13Y149_C4 = CLBLM_R_X11Y144_SLICE_X14Y144_BO6;
  assign CLBLM_L_X10Y149_SLICE_X13Y149_C5 = CLBLM_L_X10Y146_SLICE_X13Y146_DO6;
  assign CLBLM_L_X10Y149_SLICE_X13Y149_C6 = CLBLM_L_X10Y147_SLICE_X12Y147_BO6;
  assign CLBLM_R_X7Y149_SLICE_X9Y149_D5 = 1'b1;
  assign CLBLM_R_X7Y149_SLICE_X9Y149_D6 = CLBLM_R_X7Y153_SLICE_X8Y153_A5Q;
  assign CLBLM_L_X10Y149_SLICE_X13Y149_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X10Y149_SLICE_X13Y149_D1 = CLBLM_R_X5Y149_SLICE_X7Y149_CQ;
  assign CLBLM_L_X10Y149_SLICE_X13Y149_D2 = CLBLM_R_X7Y151_SLICE_X8Y151_BQ;
  assign CLBLM_L_X10Y149_SLICE_X13Y149_D3 = CLBLM_L_X10Y148_SLICE_X12Y148_AO6;
  assign CLBLM_L_X10Y149_SLICE_X13Y149_D4 = CLBLM_L_X10Y147_SLICE_X13Y147_DO6;
  assign CLBLM_L_X10Y149_SLICE_X13Y149_D5 = 1'b1;
  assign CLBLM_L_X10Y149_SLICE_X13Y149_D6 = CLBLM_L_X12Y149_SLICE_X17Y149_CO6;
  assign CLBLM_L_X10Y149_SLICE_X12Y149_A1 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_L_X10Y149_SLICE_X12Y149_A2 = CLBLL_L_X4Y150_SLICE_X4Y150_B5Q;
  assign CLBLM_L_X10Y149_SLICE_X12Y149_A3 = CLBLM_R_X3Y145_SLICE_X3Y145_BQ;
  assign CLBLM_L_X10Y149_SLICE_X12Y149_A4 = CLBLM_L_X10Y152_SLICE_X12Y152_AQ;
  assign CLBLM_L_X10Y149_SLICE_X12Y149_A5 = CLBLM_L_X10Y146_SLICE_X13Y146_AQ;
  assign CLBLM_L_X10Y149_SLICE_X12Y149_A6 = 1'b1;
  assign RIOI3_X105Y129_ILOGIC_X1Y130_D = RIOB33_X105Y129_IOB_X1Y130_I;
  assign RIOI3_X105Y129_ILOGIC_X1Y129_D = RIOB33_X105Y129_IOB_X1Y129_I;
  assign CLBLM_L_X10Y149_SLICE_X12Y149_B1 = CLBLM_L_X10Y145_SLICE_X12Y145_BQ;
  assign CLBLM_L_X10Y149_SLICE_X12Y149_B2 = CLBLM_L_X8Y154_SLICE_X10Y154_BO5;
  assign CLBLM_L_X10Y149_SLICE_X12Y149_B3 = CLBLL_L_X4Y153_SLICE_X5Y153_A5Q;
  assign CLBLM_L_X10Y149_SLICE_X12Y149_B4 = CLBLM_R_X7Y145_SLICE_X8Y145_A5Q;
  assign CLBLM_L_X10Y149_SLICE_X12Y149_B5 = RIOB33_X105Y131_IOB_X1Y131_I;
  assign CLBLM_L_X10Y149_SLICE_X12Y149_B6 = 1'b1;
  assign CLBLM_L_X10Y149_SLICE_X12Y149_BX = CLBLM_L_X12Y149_SLICE_X17Y149_AO6;
  assign CLBLM_L_X10Y149_SLICE_X12Y149_C1 = CLBLM_L_X12Y147_SLICE_X16Y147_DO6;
  assign CLBLM_L_X10Y149_SLICE_X12Y149_C2 = CLBLM_R_X11Y148_SLICE_X15Y148_BO6;
  assign CLBLM_L_X10Y149_SLICE_X12Y149_C3 = CLBLM_L_X10Y147_SLICE_X12Y147_DO6;
  assign CLBLM_L_X10Y149_SLICE_X12Y149_C4 = CLBLM_R_X7Y149_SLICE_X8Y149_DO6;
  assign CLBLM_L_X10Y149_SLICE_X12Y149_C5 = CLBLM_L_X10Y150_SLICE_X12Y150_CO6;
  assign CLBLM_L_X10Y149_SLICE_X12Y149_C6 = CLBLM_R_X7Y150_SLICE_X9Y150_BO6;
  assign CLBLM_L_X10Y149_SLICE_X12Y149_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X7Y149_SLICE_X8Y149_A4 = CLBLM_L_X10Y151_SLICE_X13Y151_AQ;
  assign CLBLM_R_X7Y149_SLICE_X8Y149_A5 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_L_X10Y149_SLICE_X12Y149_D1 = 1'b1;
  assign CLBLM_L_X10Y149_SLICE_X12Y149_D2 = CLBLM_L_X10Y150_SLICE_X12Y150_AO5;
  assign CLBLM_L_X10Y149_SLICE_X12Y149_D3 = 1'b1;
  assign CLBLM_L_X10Y149_SLICE_X12Y149_D4 = CLBLM_R_X7Y149_SLICE_X8Y149_DO6;
  assign CLBLM_L_X10Y149_SLICE_X12Y149_D5 = CLBLM_L_X8Y149_SLICE_X11Y149_DO6;
  assign CLBLM_L_X10Y149_SLICE_X12Y149_D6 = CLBLM_R_X7Y150_SLICE_X9Y150_BO6;
  assign LIOI3_SING_X0Y150_OLOGIC_X0Y150_D1 = CLBLM_R_X3Y144_SLICE_X2Y144_AO5;
  assign CLBLM_R_X103Y178_SLICE_X163Y178_A1 = 1'b1;
  assign CLBLM_R_X103Y178_SLICE_X163Y178_A2 = RIOB33_X105Y125_IOB_X1Y125_I;
  assign CLBLM_R_X103Y178_SLICE_X163Y178_A3 = 1'b1;
  assign CLBLM_R_X103Y178_SLICE_X163Y178_A4 = RIOB33_X105Y125_IOB_X1Y126_I;
  assign CLBLM_R_X103Y178_SLICE_X163Y178_A5 = 1'b1;
  assign CLBLM_R_X103Y178_SLICE_X163Y178_A6 = RIOB33_X105Y127_IOB_X1Y127_I;
  assign RIOI3_TBYTESRC_X105Y143_ILOGIC_X1Y144_D = RIOB33_X105Y143_IOB_X1Y144_I;
  assign CLBLM_R_X103Y178_SLICE_X163Y178_B1 = 1'b1;
  assign CLBLM_R_X103Y178_SLICE_X163Y178_B2 = 1'b1;
  assign CLBLM_R_X103Y178_SLICE_X163Y178_B3 = 1'b1;
  assign CLBLM_R_X103Y178_SLICE_X163Y178_B4 = 1'b1;
  assign CLBLM_R_X103Y178_SLICE_X163Y178_B5 = 1'b1;
  assign CLBLM_R_X103Y178_SLICE_X163Y178_B6 = 1'b1;
  assign RIOI3_TBYTESRC_X105Y143_ILOGIC_X1Y143_D = RIOB33_X105Y143_IOB_X1Y143_I;
  assign CLBLM_R_X103Y178_SLICE_X163Y178_C1 = 1'b1;
  assign CLBLM_R_X103Y178_SLICE_X163Y178_C2 = 1'b1;
  assign CLBLM_R_X103Y178_SLICE_X163Y178_C3 = 1'b1;
  assign CLBLM_R_X103Y178_SLICE_X163Y178_C4 = 1'b1;
  assign CLBLM_R_X103Y178_SLICE_X163Y178_C5 = 1'b1;
  assign CLBLM_R_X103Y178_SLICE_X163Y178_C6 = 1'b1;
  assign CLBLM_R_X103Y178_SLICE_X163Y178_D1 = 1'b1;
  assign CLBLM_R_X103Y178_SLICE_X163Y178_D2 = 1'b1;
  assign CLBLM_R_X103Y178_SLICE_X163Y178_D3 = 1'b1;
  assign CLBLM_R_X103Y178_SLICE_X163Y178_D4 = 1'b1;
  assign CLBLM_R_X103Y178_SLICE_X163Y178_D5 = 1'b1;
  assign CLBLM_R_X103Y178_SLICE_X163Y178_D6 = 1'b1;
  assign CLBLM_R_X7Y149_SLICE_X8Y149_B5 = CLBLM_R_X7Y153_SLICE_X8Y153_A5Q;
  assign CLBLM_R_X103Y178_SLICE_X162Y178_A1 = 1'b1;
  assign CLBLM_R_X103Y178_SLICE_X162Y178_A2 = 1'b1;
  assign CLBLM_R_X103Y178_SLICE_X162Y178_A3 = 1'b1;
  assign CLBLM_R_X103Y178_SLICE_X162Y178_A4 = 1'b1;
  assign CLBLM_R_X7Y149_SLICE_X8Y149_B6 = CLBLM_R_X7Y149_SLICE_X9Y149_CQ;
  assign CLBLM_R_X103Y178_SLICE_X162Y178_A5 = 1'b1;
  assign CLBLM_R_X103Y178_SLICE_X162Y178_A6 = 1'b1;
  assign CLBLM_R_X103Y178_SLICE_X162Y178_B1 = 1'b1;
  assign CLBLM_R_X103Y178_SLICE_X162Y178_B2 = 1'b1;
  assign CLBLM_R_X103Y178_SLICE_X162Y178_B3 = 1'b1;
  assign CLBLM_R_X103Y178_SLICE_X162Y178_B4 = 1'b1;
  assign CLBLM_R_X103Y178_SLICE_X162Y178_B5 = 1'b1;
  assign CLBLM_R_X103Y178_SLICE_X162Y178_B6 = 1'b1;
  assign LIOI3_SING_X0Y150_OLOGIC_X0Y150_T1 = 1'b1;
  assign CLBLM_R_X103Y178_SLICE_X162Y178_C1 = 1'b1;
  assign CLBLM_R_X103Y178_SLICE_X162Y178_C2 = 1'b1;
  assign CLBLM_R_X103Y178_SLICE_X162Y178_C3 = 1'b1;
  assign CLBLM_R_X103Y178_SLICE_X162Y178_C4 = 1'b1;
  assign CLBLM_R_X103Y178_SLICE_X162Y178_C5 = 1'b1;
  assign CLBLM_R_X103Y178_SLICE_X162Y178_C6 = 1'b1;
  assign CLBLM_R_X103Y178_SLICE_X162Y178_D1 = 1'b1;
  assign CLBLM_R_X103Y178_SLICE_X162Y178_D2 = 1'b1;
  assign CLBLM_R_X103Y178_SLICE_X162Y178_D3 = 1'b1;
  assign CLBLM_R_X103Y178_SLICE_X162Y178_D4 = 1'b1;
  assign CLBLM_R_X103Y178_SLICE_X162Y178_D5 = 1'b1;
  assign CLBLM_R_X103Y178_SLICE_X162Y178_D6 = 1'b1;
  assign CLBLL_L_X4Y146_SLICE_X4Y146_A1 = CLBLL_L_X4Y144_SLICE_X4Y144_DQ;
  assign CLBLL_L_X4Y146_SLICE_X4Y146_A2 = CLBLM_L_X10Y145_SLICE_X12Y145_AQ;
  assign CLBLL_L_X4Y146_SLICE_X4Y146_A3 = CLBLL_L_X4Y146_SLICE_X4Y146_AQ;
  assign CLBLL_L_X4Y146_SLICE_X4Y146_A4 = CLBLM_R_X5Y142_SLICE_X7Y142_BQ;
  assign CLBLL_L_X4Y146_SLICE_X4Y146_A5 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLL_L_X4Y146_SLICE_X4Y146_A6 = CLBLL_L_X4Y149_SLICE_X4Y149_BQ;
  assign CLBLL_L_X4Y146_SLICE_X4Y146_B1 = CLBLM_R_X3Y151_SLICE_X3Y151_AQ;
  assign CLBLL_L_X4Y146_SLICE_X4Y146_B2 = CLBLL_L_X4Y145_SLICE_X4Y145_CQ;
  assign CLBLL_L_X4Y146_SLICE_X4Y146_B3 = CLBLM_R_X3Y147_SLICE_X2Y147_AQ;
  assign CLBLL_L_X4Y146_SLICE_X4Y146_B4 = CLBLL_L_X4Y144_SLICE_X4Y144_D5Q;
  assign CLBLL_L_X4Y146_SLICE_X4Y146_B5 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLL_L_X4Y146_SLICE_X4Y146_B6 = 1'b1;
  assign CLBLL_L_X4Y146_SLICE_X4Y146_C1 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLL_L_X4Y146_SLICE_X4Y146_C2 = 1'b1;
  assign CLBLL_L_X4Y146_SLICE_X4Y146_C3 = CLBLM_R_X3Y147_SLICE_X3Y147_C5Q;
  assign CLBLL_L_X4Y146_SLICE_X4Y146_C4 = CLBLM_L_X12Y151_SLICE_X16Y151_AQ;
  assign CLBLL_L_X4Y146_SLICE_X4Y146_C5 = CLBLM_R_X3Y149_SLICE_X3Y149_CQ;
  assign CLBLL_L_X4Y146_SLICE_X4Y146_C6 = 1'b1;
  assign CLBLL_L_X4Y146_SLICE_X4Y146_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLL_L_X4Y146_SLICE_X4Y146_D1 = CLBLL_L_X2Y146_SLICE_X1Y146_AQ;
  assign CLBLL_L_X4Y146_SLICE_X4Y146_D2 = CLBLL_L_X4Y149_SLICE_X5Y149_CQ;
  assign CLBLL_L_X4Y146_SLICE_X4Y146_D3 = CLBLM_R_X7Y144_SLICE_X8Y144_DQ;
  assign CLBLL_L_X4Y146_SLICE_X4Y146_D4 = CLBLM_R_X3Y147_SLICE_X2Y147_CQ;
  assign CLBLL_L_X4Y146_SLICE_X4Y146_D5 = CLBLM_R_X5Y146_SLICE_X7Y146_C5Q;
  assign CLBLL_L_X4Y146_SLICE_X4Y146_D6 = 1'b1;
  assign CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_CE = 1'b1;
  assign CLBLL_L_X4Y146_SLICE_X5Y146_A1 = CLBLL_L_X4Y153_SLICE_X4Y153_AQ;
  assign CLBLL_L_X4Y146_SLICE_X5Y146_A2 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLL_L_X4Y146_SLICE_X5Y146_A3 = CLBLL_L_X4Y146_SLICE_X5Y146_AQ;
  assign CLBLL_L_X4Y146_SLICE_X5Y146_A4 = CLBLL_L_X4Y146_SLICE_X5Y146_CQ;
  assign CLBLL_L_X4Y146_SLICE_X5Y146_A5 = CLBLM_L_X8Y146_SLICE_X11Y146_C5Q;
  assign CLBLL_L_X4Y146_SLICE_X5Y146_A6 = 1'b1;
  assign LIOB33_X0Y135_IOB_X0Y136_O = CLBLM_L_X10Y153_SLICE_X13Y153_CQ;
  assign LIOB33_X0Y135_IOB_X0Y135_O = CLBLL_L_X2Y145_SLICE_X0Y145_BQ;
  assign CLBLL_L_X4Y146_SLICE_X5Y146_B1 = 1'b1;
  assign CLBLL_L_X4Y146_SLICE_X5Y146_B2 = CLBLL_L_X4Y145_SLICE_X4Y145_DO5;
  assign CLBLL_L_X4Y146_SLICE_X5Y146_B3 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLL_L_X4Y146_SLICE_X5Y146_B4 = CLBLM_R_X5Y145_SLICE_X6Y145_D5Q;
  assign CLBLL_L_X4Y146_SLICE_X5Y146_B5 = CLBLL_L_X4Y143_SLICE_X4Y143_BQ;
  assign CLBLL_L_X4Y146_SLICE_X5Y146_B6 = CLBLL_L_X4Y146_SLICE_X5Y146_DQ;
  assign CLBLL_L_X4Y146_SLICE_X5Y146_C1 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLL_L_X4Y146_SLICE_X5Y146_C2 = CLBLM_L_X8Y142_SLICE_X10Y142_CQ;
  assign CLBLL_L_X4Y146_SLICE_X5Y146_C3 = CLBLL_L_X4Y153_SLICE_X4Y153_AQ;
  assign CLBLL_L_X4Y146_SLICE_X5Y146_C4 = 1'b1;
  assign CLBLL_L_X4Y146_SLICE_X5Y146_C5 = CLBLL_L_X4Y146_SLICE_X5Y146_AQ;
  assign CLBLL_L_X4Y146_SLICE_X5Y146_C6 = CLBLL_L_X4Y146_SLICE_X5Y146_CQ;
  assign CLBLL_L_X4Y146_SLICE_X5Y146_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLL_L_X4Y146_SLICE_X5Y146_D1 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLL_L_X4Y146_SLICE_X5Y146_D2 = CLBLL_L_X4Y142_SLICE_X4Y142_AQ;
  assign CLBLL_L_X4Y146_SLICE_X5Y146_D3 = CLBLM_L_X10Y151_SLICE_X13Y151_AQ;
  assign CLBLL_L_X4Y146_SLICE_X5Y146_D4 = CLBLL_L_X4Y148_SLICE_X4Y148_AQ;
  assign CLBLL_L_X4Y146_SLICE_X5Y146_D5 = CLBLM_R_X3Y143_SLICE_X3Y143_BQ;
  assign CLBLL_L_X4Y146_SLICE_X5Y146_D6 = CLBLL_L_X4Y146_SLICE_X5Y146_CQ;
  assign CLBLM_L_X10Y150_SLICE_X13Y150_A1 = CLBLM_R_X7Y151_SLICE_X8Y151_DQ;
  assign CLBLM_L_X10Y150_SLICE_X13Y150_A2 = 1'b1;
  assign CLBLM_L_X10Y150_SLICE_X13Y150_A3 = CLBLM_L_X10Y150_SLICE_X13Y150_AQ;
  assign CLBLM_L_X10Y150_SLICE_X13Y150_A4 = CLBLL_L_X4Y150_SLICE_X5Y150_BQ;
  assign CLBLM_L_X10Y150_SLICE_X13Y150_A5 = CLBLM_R_X13Y149_SLICE_X18Y149_AO6;
  assign CLBLM_L_X10Y150_SLICE_X13Y150_A6 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_L_X10Y150_SLICE_X13Y150_B1 = CLBLM_R_X11Y150_SLICE_X14Y150_DO6;
  assign CLBLM_L_X10Y150_SLICE_X13Y150_B2 = CLBLM_L_X10Y151_SLICE_X13Y151_BO6;
  assign CLBLM_L_X10Y150_SLICE_X13Y150_B3 = CLBLM_R_X5Y148_SLICE_X7Y148_BQ;
  assign CLBLM_L_X10Y150_SLICE_X13Y150_B4 = CLBLM_L_X10Y151_SLICE_X13Y151_BO5;
  assign CLBLM_L_X10Y150_SLICE_X13Y150_B5 = CLBLM_L_X10Y150_SLICE_X12Y150_AQ;
  assign CLBLM_L_X10Y150_SLICE_X13Y150_B6 = 1'b1;
  assign CLBLM_L_X10Y150_SLICE_X13Y150_C1 = CLBLM_R_X7Y149_SLICE_X8Y149_AQ;
  assign CLBLM_L_X10Y150_SLICE_X13Y150_C2 = CLBLM_L_X12Y147_SLICE_X16Y147_DO6;
  assign CLBLM_L_X10Y150_SLICE_X13Y150_C3 = CLBLM_R_X7Y153_SLICE_X8Y153_A5Q;
  assign CLBLM_L_X10Y150_SLICE_X13Y150_C4 = CLBLL_L_X4Y148_SLICE_X4Y148_CQ;
  assign CLBLM_L_X10Y150_SLICE_X13Y150_C5 = CLBLM_R_X7Y144_SLICE_X9Y144_B5Q;
  assign CLBLM_L_X10Y150_SLICE_X13Y150_C6 = CLBLM_L_X8Y149_SLICE_X11Y149_A5Q;
  assign CLBLM_L_X10Y150_SLICE_X13Y150_CLK = CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O;
  assign CLBLM_L_X10Y150_SLICE_X13Y150_D1 = CLBLM_L_X8Y145_SLICE_X11Y145_CQ;
  assign CLBLM_L_X10Y150_SLICE_X13Y150_D2 = CLBLM_L_X10Y146_SLICE_X13Y146_DO6;
  assign CLBLM_L_X10Y150_SLICE_X13Y150_D3 = CLBLM_L_X10Y150_SLICE_X12Y150_BO5;
  assign CLBLM_L_X10Y150_SLICE_X13Y150_D4 = CLBLM_L_X10Y150_SLICE_X13Y150_CO6;
  assign CLBLM_L_X10Y150_SLICE_X13Y150_D5 = CLBLM_L_X10Y147_SLICE_X12Y147_BQ;
  assign CLBLM_L_X10Y150_SLICE_X13Y150_D6 = CLBLM_L_X10Y151_SLICE_X13Y151_BO5;
  assign CLBLM_L_X10Y150_SLICE_X12Y150_A1 = CLBLM_L_X10Y150_SLICE_X12Y150_DO6;
  assign CLBLM_L_X10Y150_SLICE_X12Y150_A2 = CLBLM_L_X10Y151_SLICE_X13Y151_BO5;
  assign CLBLM_L_X10Y150_SLICE_X12Y150_A3 = CLBLM_L_X12Y149_SLICE_X17Y149_CO6;
  assign CLBLM_L_X10Y150_SLICE_X12Y150_A4 = CLBLM_L_X8Y151_SLICE_X10Y151_AQ;
  assign CLBLM_L_X10Y150_SLICE_X12Y150_A5 = CLBLM_L_X8Y150_SLICE_X11Y150_AQ;
  assign CLBLM_L_X10Y150_SLICE_X12Y150_A6 = 1'b1;
  assign CLBLM_L_X10Y150_SLICE_X12Y150_AX = CLBLM_L_X10Y151_SLICE_X12Y151_BQ;
  assign CLBLM_L_X10Y150_SLICE_X12Y150_B1 = CLBLM_R_X7Y153_SLICE_X8Y153_A5Q;
  assign CLBLM_L_X10Y150_SLICE_X12Y150_B2 = CLBLM_L_X12Y147_SLICE_X16Y147_DO6;
  assign CLBLM_L_X10Y150_SLICE_X12Y150_B3 = CLBLM_R_X7Y149_SLICE_X8Y149_AQ;
  assign CLBLM_L_X10Y150_SLICE_X12Y150_B4 = CLBLL_L_X4Y148_SLICE_X4Y148_CQ;
  assign CLBLM_L_X10Y150_SLICE_X12Y150_B5 = CLBLM_R_X7Y144_SLICE_X9Y144_B5Q;
  assign CLBLM_L_X10Y150_SLICE_X12Y150_B6 = 1'b1;
  assign CLBLM_L_X10Y150_SLICE_X12Y150_C1 = CLBLM_L_X10Y150_SLICE_X12Y150_AO6;
  assign CLBLM_L_X10Y150_SLICE_X12Y150_C2 = CLBLM_L_X8Y151_SLICE_X10Y151_C5Q;
  assign CLBLM_L_X10Y150_SLICE_X12Y150_C3 = CLBLM_L_X10Y148_SLICE_X12Y148_AO6;
  assign CLBLM_L_X10Y150_SLICE_X12Y150_C4 = CLBLM_L_X8Y149_SLICE_X11Y149_DO6;
  assign CLBLM_L_X10Y150_SLICE_X12Y150_C5 = CLBLM_R_X7Y147_SLICE_X9Y147_D5Q;
  assign CLBLM_L_X10Y150_SLICE_X12Y150_C6 = CLBLM_L_X10Y150_SLICE_X12Y150_BO6;
  assign CLBLM_L_X10Y150_SLICE_X12Y150_CE = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_L_X10Y150_SLICE_X12Y150_CLK = CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O;
  assign CLBLM_L_X10Y150_SLICE_X12Y150_D1 = CLBLM_R_X11Y144_SLICE_X14Y144_BO6;
  assign CLBLM_L_X10Y150_SLICE_X12Y150_D2 = CLBLM_R_X7Y144_SLICE_X9Y144_B5Q;
  assign CLBLM_L_X10Y150_SLICE_X12Y150_D3 = CLBLM_R_X11Y147_SLICE_X15Y147_BO6;
  assign CLBLM_L_X10Y150_SLICE_X12Y150_D4 = CLBLM_R_X7Y147_SLICE_X9Y147_D5Q;
  assign CLBLM_L_X10Y150_SLICE_X12Y150_D5 = CLBLM_R_X7Y153_SLICE_X8Y153_A5Q;
  assign CLBLM_L_X10Y150_SLICE_X12Y150_D6 = CLBLM_L_X8Y151_SLICE_X10Y151_C5Q;
  assign CLBLM_R_X11Y144_SLICE_X15Y144_A1 = 1'b1;
  assign CLBLM_R_X11Y144_SLICE_X15Y144_A2 = 1'b1;
  assign CLBLM_R_X11Y144_SLICE_X15Y144_A3 = 1'b1;
  assign CLBLM_R_X11Y144_SLICE_X15Y144_A4 = 1'b1;
  assign CLBLM_R_X11Y144_SLICE_X15Y144_A5 = 1'b1;
  assign CLBLM_R_X11Y144_SLICE_X15Y144_A6 = 1'b1;
  assign CLBLM_R_X11Y144_SLICE_X15Y144_B1 = 1'b1;
  assign CLBLM_R_X11Y144_SLICE_X15Y144_B2 = 1'b1;
  assign CLBLM_R_X11Y144_SLICE_X15Y144_B3 = 1'b1;
  assign CLBLM_R_X11Y144_SLICE_X15Y144_B4 = 1'b1;
  assign CLBLM_R_X11Y144_SLICE_X15Y144_B5 = 1'b1;
  assign CLBLM_R_X11Y144_SLICE_X15Y144_B6 = 1'b1;
  assign CLBLM_R_X11Y144_SLICE_X15Y144_C1 = 1'b1;
  assign CLBLM_R_X11Y144_SLICE_X15Y144_C2 = 1'b1;
  assign CLBLM_R_X11Y144_SLICE_X15Y144_C3 = 1'b1;
  assign CLBLM_R_X11Y144_SLICE_X15Y144_C4 = 1'b1;
  assign CLBLM_R_X11Y144_SLICE_X15Y144_C5 = 1'b1;
  assign CLBLM_R_X11Y144_SLICE_X15Y144_C6 = 1'b1;
  assign CLBLM_R_X11Y144_SLICE_X15Y144_D1 = 1'b1;
  assign CLBLM_R_X11Y144_SLICE_X15Y144_D2 = 1'b1;
  assign CLBLM_R_X11Y144_SLICE_X15Y144_D3 = 1'b1;
  assign CLBLM_R_X11Y144_SLICE_X15Y144_D4 = 1'b1;
  assign CLBLM_R_X11Y144_SLICE_X15Y144_D5 = 1'b1;
  assign CLBLM_R_X11Y144_SLICE_X15Y144_D6 = 1'b1;
  assign CLBLM_R_X11Y144_SLICE_X14Y144_A1 = CLBLM_L_X10Y146_SLICE_X12Y146_DQ;
  assign CLBLM_R_X11Y144_SLICE_X14Y144_A2 = CLBLM_R_X7Y149_SLICE_X8Y149_AQ;
  assign CLBLL_L_X4Y147_SLICE_X4Y147_A1 = CLBLL_L_X4Y150_SLICE_X4Y150_DO6;
  assign CLBLL_L_X4Y147_SLICE_X4Y147_A2 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLL_L_X4Y147_SLICE_X4Y147_A3 = CLBLM_R_X5Y146_SLICE_X7Y146_BQ;
  assign CLBLL_L_X4Y147_SLICE_X4Y147_A4 = CLBLL_L_X4Y143_SLICE_X5Y143_BQ;
  assign CLBLL_L_X4Y147_SLICE_X4Y147_A5 = 1'b1;
  assign CLBLL_L_X4Y147_SLICE_X4Y147_A6 = 1'b1;
  assign CLBLM_R_X11Y144_SLICE_X14Y144_A3 = CLBLM_R_X5Y142_SLICE_X6Y142_D5Q;
  assign CLBLM_R_X11Y144_SLICE_X14Y144_A4 = CLBLM_R_X7Y151_SLICE_X8Y151_D5Q;
  assign CLBLM_R_X11Y144_SLICE_X14Y144_A5 = CLBLL_L_X4Y148_SLICE_X4Y148_CQ;
  assign CLBLL_L_X4Y147_SLICE_X4Y147_B1 = CLBLM_R_X5Y150_SLICE_X6Y150_B5Q;
  assign CLBLL_L_X4Y147_SLICE_X4Y147_B2 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLL_L_X4Y147_SLICE_X4Y147_B3 = CLBLL_L_X2Y146_SLICE_X1Y146_AQ;
  assign CLBLL_L_X4Y147_SLICE_X4Y147_B4 = CLBLM_R_X7Y143_SLICE_X9Y143_B5Q;
  assign CLBLL_L_X4Y147_SLICE_X4Y147_B5 = 1'b1;
  assign CLBLL_L_X4Y147_SLICE_X4Y147_B6 = 1'b1;
  assign CLBLM_R_X11Y144_SLICE_X14Y144_B1 = CLBLM_L_X10Y146_SLICE_X12Y146_DQ;
  assign CLBLM_R_X11Y144_SLICE_X14Y144_B2 = CLBLL_L_X4Y148_SLICE_X4Y148_CQ;
  assign CLBLL_L_X4Y147_SLICE_X4Y147_C1 = CLBLM_L_X10Y149_SLICE_X13Y149_AQ;
  assign CLBLL_L_X4Y147_SLICE_X4Y147_C2 = 1'b1;
  assign CLBLL_L_X4Y147_SLICE_X4Y147_C3 = CLBLL_L_X4Y147_SLICE_X4Y147_DQ;
  assign CLBLL_L_X4Y147_SLICE_X4Y147_C4 = CLBLM_R_X7Y149_SLICE_X9Y149_A5Q;
  assign CLBLL_L_X4Y147_SLICE_X4Y147_C5 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLL_L_X4Y147_SLICE_X4Y147_C6 = 1'b1;
  assign CLBLM_R_X11Y144_SLICE_X14Y144_C1 = CLBLM_R_X5Y142_SLICE_X6Y142_D5Q;
  assign CLBLL_L_X4Y147_SLICE_X4Y147_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X11Y144_SLICE_X14Y144_C2 = CLBLL_L_X4Y147_SLICE_X4Y147_CQ;
  assign CLBLM_R_X11Y144_SLICE_X14Y144_C3 = CLBLM_R_X7Y149_SLICE_X8Y149_AQ;
  assign CLBLM_R_X11Y144_SLICE_X14Y144_C4 = CLBLM_R_X7Y151_SLICE_X8Y151_D5Q;
  assign CLBLM_R_X11Y144_SLICE_X14Y144_C5 = CLBLM_L_X10Y146_SLICE_X12Y146_DQ;
  assign CLBLM_R_X11Y144_SLICE_X14Y144_C6 = CLBLL_L_X4Y148_SLICE_X4Y148_CQ;
  assign CLBLL_L_X4Y147_SLICE_X4Y147_D1 = CLBLM_R_X3Y146_SLICE_X3Y146_AQ;
  assign CLBLL_L_X4Y147_SLICE_X4Y147_D2 = CLBLM_R_X7Y153_SLICE_X9Y153_DQ;
  assign CLBLL_L_X4Y147_SLICE_X4Y147_D3 = CLBLL_L_X4Y144_SLICE_X4Y144_AQ;
  assign CLBLL_L_X4Y147_SLICE_X4Y147_D4 = CLBLM_R_X3Y147_SLICE_X3Y147_B5Q;
  assign CLBLL_L_X4Y147_SLICE_X4Y147_D5 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLL_L_X4Y147_SLICE_X4Y147_D6 = 1'b1;
  assign CLBLM_R_X11Y144_SLICE_X14Y144_D1 = CLBLM_R_X5Y142_SLICE_X6Y142_D5Q;
  assign CLBLM_R_X11Y144_SLICE_X14Y144_D2 = CLBLL_L_X4Y147_SLICE_X4Y147_CQ;
  assign CLBLM_R_X11Y144_SLICE_X14Y144_D3 = CLBLM_R_X7Y149_SLICE_X8Y149_AQ;
  assign CLBLM_R_X11Y144_SLICE_X14Y144_D4 = CLBLM_R_X7Y151_SLICE_X8Y151_D5Q;
  assign CLBLM_R_X11Y144_SLICE_X14Y144_D5 = CLBLM_L_X10Y146_SLICE_X12Y146_DQ;
  assign CLBLM_R_X11Y144_SLICE_X14Y144_D6 = CLBLL_L_X4Y148_SLICE_X4Y148_CQ;
  assign LIOB33_X0Y137_IOB_X0Y138_O = CLBLM_R_X3Y148_SLICE_X2Y148_A5Q;
  assign LIOB33_X0Y137_IOB_X0Y137_O = CLBLM_R_X5Y153_SLICE_X6Y153_B5Q;
  assign LIOI3_X0Y151_OLOGIC_X0Y152_D1 = CLBLL_L_X4Y147_SLICE_X5Y147_C5Q;
  assign LIOI3_SING_X0Y50_ILOGIC_X0Y50_D = LIOB33_SING_X0Y50_IOB_X0Y50_I;
  assign LIOI3_X0Y151_OLOGIC_X0Y152_T1 = 1'b1;
  assign RIOI3_X105Y195_OLOGIC_X1Y196_D1 = CLBLM_L_X12Y150_SLICE_X16Y150_AO6;
  assign CLBLL_L_X4Y147_SLICE_X5Y147_A1 = CLBLM_L_X8Y149_SLICE_X11Y149_AQ;
  assign CLBLL_L_X4Y147_SLICE_X5Y147_A2 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLL_L_X4Y147_SLICE_X5Y147_A3 = CLBLL_L_X4Y147_SLICE_X5Y147_AQ;
  assign CLBLL_L_X4Y147_SLICE_X5Y147_A4 = CLBLL_L_X4Y143_SLICE_X5Y143_BQ;
  assign CLBLL_L_X4Y147_SLICE_X5Y147_A5 = CLBLM_R_X5Y148_SLICE_X6Y148_AO6;
  assign CLBLL_L_X4Y147_SLICE_X5Y147_A6 = CLBLM_R_X5Y147_SLICE_X7Y147_BQ;
  assign CLBLM_R_X5Y141_SLICE_X7Y141_B1 = 1'b1;
  assign LIOI3_X0Y151_OLOGIC_X0Y151_D1 = CLBLL_L_X2Y146_SLICE_X0Y146_CQ;
  assign CLBLM_R_X5Y141_SLICE_X7Y141_B2 = 1'b1;
  assign CLBLL_L_X4Y147_SLICE_X5Y147_B1 = CLBLM_R_X3Y148_SLICE_X2Y148_B5Q;
  assign CLBLL_L_X4Y147_SLICE_X5Y147_B2 = CLBLL_L_X4Y148_SLICE_X5Y148_D5Q;
  assign CLBLL_L_X4Y147_SLICE_X5Y147_B3 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLL_L_X4Y147_SLICE_X5Y147_B4 = CLBLM_R_X7Y153_SLICE_X9Y153_DQ;
  assign CLBLL_L_X4Y147_SLICE_X5Y147_B5 = CLBLM_L_X8Y153_SLICE_X11Y153_CO6;
  assign CLBLL_L_X4Y147_SLICE_X5Y147_B6 = 1'b1;
  assign CLBLM_R_X5Y141_SLICE_X7Y141_B3 = 1'b1;
  assign RIOI3_X105Y195_OLOGIC_X1Y196_T1 = 1'b1;
  assign LIOI3_X0Y151_OLOGIC_X0Y151_T1 = 1'b1;
  assign CLBLL_L_X4Y147_SLICE_X5Y147_C1 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLL_L_X4Y147_SLICE_X5Y147_C2 = CLBLM_R_X7Y143_SLICE_X9Y143_B5Q;
  assign CLBLL_L_X4Y147_SLICE_X5Y147_C3 = CLBLL_L_X4Y148_SLICE_X5Y148_CQ;
  assign CLBLL_L_X4Y147_SLICE_X5Y147_C4 = CLBLM_R_X5Y147_SLICE_X6Y147_B5Q;
  assign CLBLL_L_X4Y147_SLICE_X5Y147_C5 = RIOB33_X105Y109_IOB_X1Y109_I;
  assign CLBLL_L_X4Y147_SLICE_X5Y147_C6 = 1'b1;
  assign RIOI3_X105Y195_OLOGIC_X1Y195_D1 = CLBLM_L_X10Y149_SLICE_X13Y149_AO5;
  assign CLBLL_L_X4Y147_SLICE_X5Y147_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign RIOI3_X105Y195_OLOGIC_X1Y195_T1 = 1'b1;
  assign CLBLL_L_X4Y147_SLICE_X5Y147_D1 = CLBLM_R_X5Y145_SLICE_X6Y145_D5Q;
  assign CLBLL_L_X4Y147_SLICE_X5Y147_D2 = CLBLL_L_X4Y150_SLICE_X5Y150_CO5;
  assign CLBLL_L_X4Y147_SLICE_X5Y147_D3 = CLBLL_L_X4Y143_SLICE_X4Y143_BQ;
  assign CLBLL_L_X4Y147_SLICE_X5Y147_D4 = CLBLL_L_X4Y145_SLICE_X5Y145_BQ;
  assign CLBLL_L_X4Y147_SLICE_X5Y147_D5 = 1'b1;
  assign CLBLL_L_X4Y147_SLICE_X5Y147_D6 = CLBLL_L_X4Y145_SLICE_X4Y145_DO5;
  assign CLBLM_L_X10Y151_SLICE_X13Y151_A1 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_L_X10Y151_SLICE_X13Y151_A2 = CLBLM_R_X11Y148_SLICE_X14Y148_BO6;
  assign CLBLM_L_X10Y151_SLICE_X13Y151_A3 = CLBLM_L_X10Y149_SLICE_X12Y149_CO6;
  assign CLBLM_L_X10Y151_SLICE_X13Y151_A4 = CLBLM_R_X7Y151_SLICE_X8Y151_CQ;
  assign CLBLM_L_X10Y151_SLICE_X13Y151_A5 = CLBLM_L_X10Y145_SLICE_X13Y145_AQ;
  assign CLBLM_L_X10Y151_SLICE_X13Y151_A6 = 1'b1;
  assign CLBLM_R_X5Y141_SLICE_X7Y141_C1 = 1'b1;
  assign CLBLM_L_X10Y151_SLICE_X13Y151_B1 = CLBLM_R_X7Y149_SLICE_X8Y149_AQ;
  assign CLBLM_L_X10Y151_SLICE_X13Y151_B2 = CLBLM_L_X12Y147_SLICE_X16Y147_DO6;
  assign CLBLM_L_X10Y151_SLICE_X13Y151_B3 = CLBLM_R_X7Y153_SLICE_X8Y153_A5Q;
  assign CLBLM_L_X10Y151_SLICE_X13Y151_B4 = CLBLL_L_X4Y148_SLICE_X4Y148_CQ;
  assign CLBLM_L_X10Y151_SLICE_X13Y151_B5 = CLBLM_R_X7Y144_SLICE_X9Y144_B5Q;
  assign CLBLM_L_X10Y151_SLICE_X13Y151_B6 = 1'b1;
  assign CLBLM_R_X5Y141_SLICE_X7Y141_C2 = 1'b1;
  assign CLBLM_R_X5Y141_SLICE_X7Y141_C3 = 1'b1;
  assign RIOI3_TBYTESRC_X105Y157_OLOGIC_X1Y158_D1 = 1'b1;
  assign CLBLM_L_X10Y151_SLICE_X13Y151_C1 = CLBLM_R_X3Y150_SLICE_X2Y150_AQ;
  assign CLBLM_L_X10Y151_SLICE_X13Y151_C2 = CLBLM_L_X12Y149_SLICE_X17Y149_CO6;
  assign CLBLM_L_X10Y151_SLICE_X13Y151_C3 = CLBLM_R_X5Y153_SLICE_X7Y153_DO6;
  assign CLBLM_L_X10Y151_SLICE_X13Y151_C4 = CLBLM_L_X10Y148_SLICE_X13Y148_DO6;
  assign CLBLM_L_X10Y151_SLICE_X13Y151_C5 = CLBLM_L_X10Y151_SLICE_X12Y151_DQ;
  assign CLBLM_L_X10Y151_SLICE_X13Y151_C6 = CLBLM_R_X13Y146_SLICE_X18Y146_BO6;
  assign RIOI3_TBYTESRC_X105Y157_OLOGIC_X1Y158_T1 = 1'b1;
  assign CLBLM_L_X10Y151_SLICE_X13Y151_CLK = CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O;
  assign CLBLM_L_X10Y151_SLICE_X13Y151_D1 = CLBLM_L_X8Y151_SLICE_X11Y151_AQ;
  assign CLBLM_L_X10Y151_SLICE_X13Y151_D2 = CLBLM_R_X7Y153_SLICE_X8Y153_A5Q;
  assign CLBLM_L_X10Y151_SLICE_X13Y151_D3 = CLBLM_L_X10Y147_SLICE_X13Y147_BO6;
  assign CLBLM_L_X10Y151_SLICE_X13Y151_D4 = CLBLM_L_X10Y146_SLICE_X13Y146_DO6;
  assign CLBLM_L_X10Y151_SLICE_X13Y151_D5 = CLBLM_L_X10Y151_SLICE_X12Y151_DQ;
  assign CLBLM_L_X10Y151_SLICE_X13Y151_D6 = CLBLM_R_X7Y144_SLICE_X9Y144_B5Q;
  assign RIOI3_TBYTESRC_X105Y157_OLOGIC_X1Y157_D1 = 1'b1;
  assign CLBLM_L_X10Y151_SLICE_X12Y151_A1 = CLBLM_L_X10Y152_SLICE_X13Y152_CQ;
  assign CLBLM_L_X10Y151_SLICE_X12Y151_A2 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_L_X10Y151_SLICE_X12Y151_A3 = CLBLM_L_X10Y151_SLICE_X12Y151_AQ;
  assign CLBLM_L_X10Y151_SLICE_X12Y151_A4 = CLBLM_L_X10Y149_SLICE_X12Y149_A5Q;
  assign CLBLM_L_X10Y151_SLICE_X12Y151_A5 = CLBLM_L_X10Y145_SLICE_X12Y145_AQ;
  assign CLBLM_L_X10Y151_SLICE_X12Y151_A6 = CLBLM_R_X5Y142_SLICE_X7Y142_BQ;
  assign RIOI3_TBYTESRC_X105Y157_OLOGIC_X1Y157_T1 = 1'b1;
  assign CLBLM_L_X10Y151_SLICE_X12Y151_B1 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_L_X10Y151_SLICE_X12Y151_B2 = CLBLM_L_X8Y143_SLICE_X11Y143_D5Q;
  assign CLBLM_L_X10Y151_SLICE_X12Y151_B3 = CLBLL_L_X4Y147_SLICE_X5Y147_CQ;
  assign CLBLM_L_X10Y151_SLICE_X12Y151_B4 = CLBLL_L_X4Y142_SLICE_X5Y142_DQ;
  assign CLBLM_L_X10Y151_SLICE_X12Y151_B5 = CLBLM_L_X8Y146_SLICE_X11Y146_D5Q;
  assign CLBLM_L_X10Y151_SLICE_X12Y151_B6 = CLBLM_L_X10Y151_SLICE_X12Y151_BQ;
  assign CLBLM_L_X10Y151_SLICE_X12Y151_C1 = CLBLM_L_X8Y152_SLICE_X11Y152_AQ;
  assign CLBLM_L_X10Y151_SLICE_X12Y151_C2 = CLBLM_L_X10Y151_SLICE_X12Y151_CQ;
  assign CLBLM_L_X10Y151_SLICE_X12Y151_C3 = CLBLM_L_X10Y151_SLICE_X12Y151_BQ;
  assign CLBLM_L_X10Y151_SLICE_X12Y151_C4 = CLBLM_R_X11Y148_SLICE_X15Y148_AO6;
  assign CLBLM_L_X10Y151_SLICE_X12Y151_C5 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_L_X10Y151_SLICE_X12Y151_C6 = 1'b1;
  assign CLBLM_L_X10Y151_SLICE_X12Y151_CLK = CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O;
  assign CLBLM_L_X10Y151_SLICE_X12Y151_D1 = CLBLM_L_X8Y151_SLICE_X11Y151_AQ;
  assign CLBLM_L_X10Y151_SLICE_X12Y151_D2 = 1'b1;
  assign CLBLM_L_X10Y151_SLICE_X12Y151_D3 = CLBLM_L_X10Y151_SLICE_X12Y151_DQ;
  assign CLBLM_L_X10Y151_SLICE_X12Y151_D4 = CLBLM_L_X12Y149_SLICE_X17Y149_CO6;
  assign CLBLM_L_X10Y151_SLICE_X12Y151_D5 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_L_X10Y151_SLICE_X12Y151_D6 = CLBLM_L_X8Y142_SLICE_X11Y142_AQ;
  assign CLBLM_R_X3Y143_SLICE_X3Y143_B1 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X3Y143_SLICE_X3Y143_B2 = CLBLM_R_X3Y143_SLICE_X3Y143_BQ;
  assign CLBLM_R_X11Y145_SLICE_X15Y145_A1 = CLBLM_L_X10Y144_SLICE_X13Y144_DQ;
  assign CLBLM_R_X11Y145_SLICE_X15Y145_A2 = CLBLM_L_X10Y146_SLICE_X13Y146_BQ;
  assign CLBLM_R_X11Y145_SLICE_X15Y145_A3 = CLBLM_R_X11Y145_SLICE_X15Y145_AQ;
  assign CLBLM_R_X3Y143_SLICE_X3Y143_B5 = CLBLL_L_X4Y142_SLICE_X4Y142_AQ;
  assign CLBLM_R_X11Y145_SLICE_X15Y145_A4 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X11Y145_SLICE_X15Y145_A5 = CLBLM_R_X11Y146_SLICE_X14Y146_DO6;
  assign CLBLM_R_X11Y145_SLICE_X15Y145_A6 = 1'b1;
  assign CLBLM_R_X11Y145_SLICE_X15Y145_B1 = CLBLM_R_X7Y146_SLICE_X9Y146_CO6;
  assign CLBLM_R_X11Y145_SLICE_X15Y145_B2 = CLBLM_R_X11Y146_SLICE_X15Y146_BO6;
  assign CLBLM_R_X11Y145_SLICE_X15Y145_B3 = CLBLM_L_X12Y145_SLICE_X16Y145_AQ;
  assign CLBLM_R_X11Y145_SLICE_X15Y145_B4 = CLBLM_R_X11Y145_SLICE_X15Y145_AQ;
  assign CLBLM_R_X11Y145_SLICE_X15Y145_B5 = CLBLM_L_X12Y145_SLICE_X17Y145_CO6;
  assign CLBLM_R_X11Y145_SLICE_X15Y145_B6 = CLBLM_R_X11Y147_SLICE_X14Y147_AO5;
  assign CLBLM_R_X11Y145_SLICE_X15Y145_C1 = CLBLM_R_X5Y141_SLICE_X6Y141_AQ;
  assign CLBLM_R_X11Y145_SLICE_X15Y145_C2 = CLBLM_R_X5Y148_SLICE_X6Y148_CQ;
  assign CLBLM_R_X11Y145_SLICE_X15Y145_C3 = CLBLM_R_X11Y146_SLICE_X15Y146_BO5;
  assign CLBLM_R_X11Y145_SLICE_X15Y145_C4 = CLBLM_L_X12Y146_SLICE_X16Y146_CO6;
  assign CLBLM_R_X11Y145_SLICE_X15Y145_C5 = CLBLM_L_X12Y145_SLICE_X16Y145_AO5;
  assign CLBLM_R_X11Y145_SLICE_X15Y145_C6 = 1'b1;
  assign RIOI3_X105Y133_ILOGIC_X1Y134_D = RIOB33_X105Y133_IOB_X1Y134_I;
  assign RIOI3_X105Y133_ILOGIC_X1Y133_D = RIOB33_X105Y133_IOB_X1Y133_I;
  assign CLBLM_R_X11Y145_SLICE_X15Y145_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X11Y145_SLICE_X15Y145_D1 = 1'b1;
  assign CLBLM_R_X11Y145_SLICE_X15Y145_D2 = 1'b1;
  assign CLBLM_R_X11Y145_SLICE_X15Y145_D3 = 1'b1;
  assign CLBLM_R_X11Y145_SLICE_X15Y145_D4 = 1'b1;
  assign CLBLM_R_X11Y145_SLICE_X15Y145_D5 = 1'b1;
  assign CLBLM_R_X11Y145_SLICE_X15Y145_D6 = 1'b1;
  assign CLBLL_L_X4Y148_SLICE_X4Y148_A1 = CLBLM_R_X3Y146_SLICE_X2Y146_D5Q;
  assign CLBLL_L_X4Y148_SLICE_X4Y148_A2 = CLBLL_L_X4Y148_SLICE_X4Y148_BQ;
  assign CLBLL_L_X4Y148_SLICE_X4Y148_A3 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLL_L_X4Y148_SLICE_X4Y148_A4 = CLBLM_R_X3Y143_SLICE_X3Y143_BQ;
  assign CLBLL_L_X4Y148_SLICE_X4Y148_A5 = CLBLL_L_X4Y142_SLICE_X4Y142_AQ;
  assign CLBLL_L_X4Y148_SLICE_X4Y148_A6 = CLBLM_R_X3Y152_SLICE_X3Y152_CQ;
  assign CLBLM_R_X11Y145_SLICE_X14Y145_A1 = CLBLM_R_X7Y153_SLICE_X8Y153_A5Q;
  assign CLBLM_R_X11Y145_SLICE_X14Y145_A2 = CLBLM_L_X12Y145_SLICE_X17Y145_CO6;
  assign CLBLM_R_X11Y145_SLICE_X14Y145_A3 = LIOB33_X0Y51_IOB_X0Y52_I;
  assign CLBLL_L_X4Y148_SLICE_X4Y148_B1 = CLBLL_L_X4Y149_SLICE_X5Y149_BQ;
  assign CLBLL_L_X4Y148_SLICE_X4Y148_B2 = CLBLM_R_X3Y143_SLICE_X3Y143_BQ;
  assign CLBLL_L_X4Y148_SLICE_X4Y148_B3 = CLBLL_L_X4Y147_SLICE_X4Y147_C5Q;
  assign CLBLL_L_X4Y148_SLICE_X4Y148_B4 = CLBLM_L_X10Y149_SLICE_X13Y149_AQ;
  assign CLBLL_L_X4Y148_SLICE_X4Y148_B5 = CLBLL_L_X4Y142_SLICE_X4Y142_AQ;
  assign CLBLL_L_X4Y148_SLICE_X4Y148_B6 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X11Y145_SLICE_X14Y145_A5 = CLBLM_R_X7Y144_SLICE_X9Y144_B5Q;
  assign CLBLM_R_X11Y145_SLICE_X14Y145_A6 = CLBLM_L_X12Y145_SLICE_X17Y145_AO5;
  assign CLBLL_L_X4Y148_SLICE_X4Y148_C1 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLL_L_X4Y148_SLICE_X4Y148_C2 = CLBLL_L_X4Y148_SLICE_X5Y148_A5Q;
  assign CLBLL_L_X4Y148_SLICE_X4Y148_C3 = CLBLL_L_X4Y143_SLICE_X4Y143_A5Q;
  assign CLBLL_L_X4Y148_SLICE_X4Y148_C4 = 1'b1;
  assign CLBLL_L_X4Y148_SLICE_X4Y148_C5 = CLBLM_L_X10Y153_SLICE_X13Y153_A5Q;
  assign CLBLL_L_X4Y148_SLICE_X4Y148_C6 = 1'b1;
  assign CLBLM_R_X11Y145_SLICE_X14Y145_B4 = RIOB33_X105Y135_IOB_X1Y136_I;
  assign CLBLM_R_X11Y145_SLICE_X14Y145_B5 = LIOB33_SING_X0Y50_IOB_X0Y50_I;
  assign CLBLL_L_X4Y148_SLICE_X4Y148_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X11Y145_SLICE_X14Y145_C1 = CLBLM_R_X5Y144_SLICE_X6Y144_AQ;
  assign CLBLM_R_X11Y145_SLICE_X14Y145_C2 = CLBLM_R_X11Y147_SLICE_X14Y147_AO5;
  assign CLBLM_R_X11Y145_SLICE_X14Y145_C3 = CLBLM_R_X7Y146_SLICE_X9Y146_CO6;
  assign CLBLM_R_X11Y145_SLICE_X14Y145_C4 = LIOB33_X0Y51_IOB_X0Y51_I;
  assign CLBLL_L_X4Y148_SLICE_X4Y148_D1 = CLBLL_L_X4Y151_SLICE_X4Y151_AQ;
  assign CLBLL_L_X4Y148_SLICE_X4Y148_D2 = CLBLM_R_X5Y145_SLICE_X6Y145_D5Q;
  assign CLBLL_L_X4Y148_SLICE_X4Y148_D3 = CLBLL_L_X4Y143_SLICE_X4Y143_AQ;
  assign CLBLL_L_X4Y148_SLICE_X4Y148_D4 = CLBLL_L_X4Y143_SLICE_X4Y143_BQ;
  assign CLBLL_L_X4Y148_SLICE_X4Y148_D5 = CLBLL_L_X4Y151_SLICE_X5Y151_CQ;
  assign CLBLL_L_X4Y148_SLICE_X4Y148_D6 = CLBLM_R_X3Y145_SLICE_X3Y145_BQ;
  assign CLBLM_R_X11Y145_SLICE_X14Y145_D1 = CLBLM_R_X11Y146_SLICE_X14Y146_DO6;
  assign CLBLM_R_X11Y145_SLICE_X14Y145_D2 = 1'b1;
  assign CLBLM_R_X11Y145_SLICE_X14Y145_D3 = CLBLM_R_X11Y145_SLICE_X15Y145_BO6;
  assign CLBLM_R_X11Y145_SLICE_X14Y145_D4 = CLBLM_L_X12Y145_SLICE_X16Y145_BO6;
  assign CLBLM_R_X11Y145_SLICE_X14Y145_D5 = CLBLM_R_X11Y144_SLICE_X14Y144_DO6;
  assign CLBLM_R_X11Y145_SLICE_X14Y145_D6 = CLBLM_R_X11Y145_SLICE_X14Y145_BO6;
  assign CLBLL_L_X4Y148_SLICE_X5Y148_A1 = CLBLL_L_X4Y148_SLICE_X5Y148_CQ;
  assign CLBLL_L_X4Y148_SLICE_X5Y148_A2 = CLBLL_L_X4Y153_SLICE_X5Y153_AQ;
  assign CLBLL_L_X4Y148_SLICE_X5Y148_A3 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLL_L_X4Y148_SLICE_X5Y148_A4 = RIOB33_X105Y117_IOB_X1Y117_I;
  assign CLBLL_L_X4Y148_SLICE_X5Y148_A5 = CLBLM_R_X5Y145_SLICE_X7Y145_B5Q;
  assign CLBLL_L_X4Y148_SLICE_X5Y148_A6 = 1'b1;
  assign CLBLL_L_X4Y148_SLICE_X5Y148_B1 = CLBLL_L_X4Y140_SLICE_X5Y140_DO6;
  assign CLBLL_L_X4Y148_SLICE_X5Y148_B2 = CLBLL_L_X4Y148_SLICE_X5Y148_BQ;
  assign CLBLL_L_X4Y148_SLICE_X5Y148_B3 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLL_L_X4Y148_SLICE_X5Y148_B4 = CLBLL_L_X4Y153_SLICE_X5Y153_A5Q;
  assign CLBLL_L_X4Y148_SLICE_X5Y148_B5 = CLBLM_R_X5Y152_SLICE_X7Y152_BQ;
  assign CLBLL_L_X4Y148_SLICE_X5Y148_B6 = 1'b1;
  assign CLBLL_L_X4Y148_SLICE_X5Y148_C1 = CLBLM_R_X7Y153_SLICE_X9Y153_AQ;
  assign CLBLL_L_X4Y148_SLICE_X5Y148_C2 = CLBLM_R_X5Y148_SLICE_X6Y148_BO6;
  assign CLBLL_L_X4Y148_SLICE_X5Y148_C3 = 1'b1;
  assign CLBLL_L_X4Y148_SLICE_X5Y148_C4 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLL_L_X4Y148_SLICE_X5Y148_C5 = CLBLL_L_X4Y148_SLICE_X5Y148_B5Q;
  assign CLBLL_L_X4Y148_SLICE_X5Y148_C6 = 1'b1;
  assign CLBLL_L_X4Y148_SLICE_X5Y148_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLL_L_X4Y148_SLICE_X5Y148_D1 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLL_L_X4Y148_SLICE_X5Y148_D2 = CLBLM_R_X5Y152_SLICE_X6Y152_DQ;
  assign CLBLL_L_X4Y148_SLICE_X5Y148_D3 = CLBLM_R_X3Y148_SLICE_X3Y148_C5Q;
  assign CLBLL_L_X4Y148_SLICE_X5Y148_D4 = CLBLM_R_X5Y149_SLICE_X6Y149_CQ;
  assign CLBLL_L_X4Y148_SLICE_X5Y148_D5 = 1'b1;
  assign CLBLL_L_X4Y148_SLICE_X5Y148_D6 = 1'b1;
  assign CLBLM_L_X10Y152_SLICE_X13Y152_A1 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_L_X10Y152_SLICE_X13Y152_A2 = CLBLM_L_X8Y151_SLICE_X10Y151_C5Q;
  assign CLBLM_L_X10Y152_SLICE_X13Y152_A3 = CLBLM_L_X10Y152_SLICE_X13Y152_AQ;
  assign CLBLM_L_X10Y152_SLICE_X13Y152_A4 = CLBLM_L_X10Y152_SLICE_X13Y152_DO6;
  assign CLBLM_L_X10Y152_SLICE_X13Y152_A5 = 1'b1;
  assign CLBLM_L_X10Y152_SLICE_X13Y152_A6 = CLBLM_L_X10Y153_SLICE_X13Y153_DO6;
  assign CLBLM_L_X10Y152_SLICE_X13Y152_B1 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_L_X10Y152_SLICE_X13Y152_B2 = CLBLM_L_X10Y152_SLICE_X13Y152_BQ;
  assign CLBLM_L_X10Y152_SLICE_X13Y152_B3 = CLBLM_L_X10Y152_SLICE_X13Y152_AQ;
  assign CLBLM_L_X10Y152_SLICE_X13Y152_B4 = CLBLM_L_X10Y152_SLICE_X13Y152_DO6;
  assign CLBLM_L_X10Y152_SLICE_X13Y152_B5 = CLBLM_L_X8Y149_SLICE_X11Y149_A5Q;
  assign CLBLM_L_X10Y152_SLICE_X13Y152_B6 = CLBLM_L_X10Y153_SLICE_X13Y153_DO6;
  assign CLBLM_L_X8Y142_SLICE_X11Y142_A1 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_L_X8Y142_SLICE_X11Y142_A2 = CLBLM_R_X3Y145_SLICE_X3Y145_D5Q;
  assign CLBLM_L_X8Y142_SLICE_X11Y142_A3 = CLBLM_L_X8Y142_SLICE_X11Y142_AQ;
  assign CLBLM_L_X10Y152_SLICE_X13Y152_C4 = CLBLM_R_X11Y148_SLICE_X15Y148_AO6;
  assign CLBLM_L_X10Y152_SLICE_X13Y152_C5 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_L_X8Y142_SLICE_X11Y142_A4 = CLBLL_L_X4Y151_SLICE_X4Y151_BQ;
  assign CLBLM_L_X8Y142_SLICE_X11Y142_A5 = CLBLL_L_X4Y142_SLICE_X4Y142_A5Q;
  assign CLBLM_L_X8Y142_SLICE_X11Y142_A6 = CLBLM_L_X8Y144_SLICE_X11Y144_CQ;
  assign CLBLM_L_X10Y152_SLICE_X13Y152_C1 = 1'b1;
  assign CLBLM_L_X10Y152_SLICE_X13Y152_C2 = CLBLM_L_X10Y152_SLICE_X13Y152_CQ;
  assign CLBLM_L_X10Y152_SLICE_X13Y152_C3 = CLBLM_R_X5Y146_SLICE_X7Y146_AQ;
  assign CLBLM_L_X8Y142_SLICE_X11Y142_B1 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_L_X8Y142_SLICE_X11Y142_B2 = CLBLM_L_X10Y144_SLICE_X12Y144_CO6;
  assign CLBLM_L_X8Y142_SLICE_X11Y142_B3 = 1'b1;
  assign CLBLM_L_X8Y142_SLICE_X11Y142_B4 = CLBLM_L_X8Y142_SLICE_X11Y142_DO6;
  assign CLBLM_L_X8Y142_SLICE_X11Y142_B5 = CLBLM_L_X8Y142_SLICE_X11Y142_CO5;
  assign CLBLM_L_X8Y142_SLICE_X11Y142_B6 = CLBLL_L_X4Y150_SLICE_X4Y150_B5Q;
  assign CLBLM_L_X10Y152_SLICE_X13Y152_D1 = CLBLM_L_X10Y152_SLICE_X12Y152_AQ;
  assign CLBLM_L_X8Y142_SLICE_X11Y142_C1 = CLBLM_L_X10Y142_SLICE_X13Y142_AQ;
  assign CLBLM_L_X8Y142_SLICE_X11Y142_C2 = RIOB33_X105Y131_IOB_X1Y131_I;
  assign CLBLM_L_X8Y142_SLICE_X11Y142_C3 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_L_X8Y142_SLICE_X11Y142_C4 = CLBLL_L_X4Y150_SLICE_X5Y150_A5Q;
  assign CLBLM_L_X8Y142_SLICE_X11Y142_C5 = CLBLM_R_X5Y142_SLICE_X7Y142_CO6;
  assign CLBLM_L_X8Y142_SLICE_X11Y142_C6 = 1'b1;
  assign CLBLM_L_X10Y152_SLICE_X13Y152_D4 = CLBLM_L_X8Y152_SLICE_X10Y152_CQ;
  assign CLBLM_L_X8Y142_SLICE_X11Y142_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X10Y152_SLICE_X12Y152_A1 = CLBLM_R_X5Y147_SLICE_X6Y147_AQ;
  assign CLBLM_L_X10Y152_SLICE_X12Y152_A2 = CLBLM_L_X10Y149_SLICE_X12Y149_AQ;
  assign CLBLM_L_X10Y152_SLICE_X12Y152_A3 = CLBLM_L_X10Y152_SLICE_X12Y152_AQ;
  assign CLBLM_L_X10Y152_SLICE_X12Y152_A4 = CLBLM_R_X7Y146_SLICE_X8Y146_A5Q;
  assign CLBLM_L_X10Y152_SLICE_X12Y152_A5 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_L_X8Y142_SLICE_X11Y142_D1 = CLBLM_L_X8Y142_SLICE_X11Y142_BQ;
  assign CLBLM_L_X8Y142_SLICE_X11Y142_D2 = CLBLL_L_X4Y151_SLICE_X4Y151_CQ;
  assign CLBLM_L_X8Y142_SLICE_X11Y142_D3 = RIOB33_X105Y131_IOB_X1Y131_I;
  assign CLBLM_L_X8Y142_SLICE_X11Y142_D4 = CLBLM_L_X8Y142_SLICE_X10Y142_CQ;
  assign CLBLM_L_X8Y142_SLICE_X11Y142_D5 = CLBLM_R_X7Y141_SLICE_X9Y141_AQ;
  assign CLBLM_L_X8Y142_SLICE_X11Y142_D6 = CLBLM_R_X7Y143_SLICE_X9Y143_CQ;
  assign CLBLM_L_X10Y152_SLICE_X12Y152_A6 = CLBLM_L_X10Y153_SLICE_X13Y153_CQ;
  assign CLBLM_L_X10Y152_SLICE_X12Y152_B1 = CLBLL_L_X4Y142_SLICE_X5Y142_DQ;
  assign CLBLM_L_X10Y152_SLICE_X12Y152_B2 = CLBLM_L_X10Y152_SLICE_X12Y152_BQ;
  assign CLBLM_L_X10Y152_SLICE_X12Y152_B3 = CLBLM_L_X8Y146_SLICE_X11Y146_D5Q;
  assign CLBLM_L_X10Y152_SLICE_X12Y152_B4 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_L_X8Y142_SLICE_X10Y142_A1 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_L_X8Y142_SLICE_X10Y142_A2 = CLBLM_L_X10Y145_SLICE_X12Y145_AQ;
  assign CLBLM_L_X8Y142_SLICE_X10Y142_A3 = CLBLM_L_X8Y142_SLICE_X10Y142_AQ;
  assign CLBLM_L_X8Y142_SLICE_X10Y142_A4 = CLBLM_R_X7Y142_SLICE_X8Y142_CQ;
  assign CLBLM_L_X8Y142_SLICE_X10Y142_A5 = CLBLM_L_X8Y143_SLICE_X11Y143_CQ;
  assign CLBLM_L_X8Y142_SLICE_X10Y142_A6 = CLBLM_R_X5Y142_SLICE_X7Y142_BQ;
  assign CLBLM_L_X10Y152_SLICE_X12Y152_C1 = CLBLM_L_X8Y152_SLICE_X11Y152_AQ;
  assign CLBLM_L_X10Y152_SLICE_X12Y152_C2 = CLBLM_L_X10Y152_SLICE_X12Y152_CQ;
  assign CLBLM_L_X8Y142_SLICE_X10Y142_AX = CLBLM_L_X8Y142_SLICE_X11Y142_CO6;
  assign CLBLM_L_X10Y152_SLICE_X12Y152_C3 = CLBLM_L_X10Y153_SLICE_X13Y153_AQ;
  assign CLBLM_L_X8Y142_SLICE_X10Y142_B1 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_L_X8Y142_SLICE_X10Y142_B2 = CLBLM_L_X8Y142_SLICE_X10Y142_BQ;
  assign CLBLM_L_X8Y142_SLICE_X10Y142_B3 = 1'b1;
  assign CLBLM_L_X8Y142_SLICE_X10Y142_B4 = CLBLM_R_X5Y143_SLICE_X6Y143_BQ;
  assign CLBLM_L_X8Y142_SLICE_X10Y142_B5 = CLBLM_L_X8Y144_SLICE_X10Y144_AO6;
  assign CLBLM_L_X8Y142_SLICE_X10Y142_B6 = CLBLM_L_X10Y144_SLICE_X12Y144_AO6;
  assign CLBLM_L_X10Y152_SLICE_X12Y152_CLK = CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O;
  assign CLBLM_L_X10Y152_SLICE_X12Y152_D1 = CLBLM_R_X7Y146_SLICE_X8Y146_A5Q;
  assign CLBLM_L_X10Y152_SLICE_X12Y152_D2 = CLBLM_L_X10Y152_SLICE_X12Y152_AQ;
  assign CLBLM_L_X8Y142_SLICE_X10Y142_C1 = CLBLM_R_X7Y141_SLICE_X9Y141_AQ;
  assign CLBLM_L_X8Y142_SLICE_X10Y142_C2 = CLBLM_L_X8Y142_SLICE_X10Y142_CQ;
  assign CLBLM_L_X8Y142_SLICE_X10Y142_C3 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_L_X8Y142_SLICE_X10Y142_C4 = CLBLM_R_X5Y142_SLICE_X7Y142_BQ;
  assign CLBLM_L_X8Y142_SLICE_X10Y142_C5 = CLBLM_L_X8Y142_SLICE_X10Y142_DO6;
  assign CLBLM_L_X8Y142_SLICE_X10Y142_C6 = CLBLL_L_X4Y151_SLICE_X4Y151_CQ;
  assign CLBLM_L_X10Y152_SLICE_X12Y152_D3 = CLBLM_R_X5Y147_SLICE_X6Y147_AQ;
  assign CLBLM_L_X10Y152_SLICE_X12Y152_D4 = CLBLM_L_X8Y152_SLICE_X10Y152_CQ;
  assign CLBLM_L_X10Y152_SLICE_X12Y152_D5 = CLBLM_L_X10Y153_SLICE_X13Y153_CQ;
  assign CLBLM_L_X8Y142_SLICE_X10Y142_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X10Y152_SLICE_X12Y152_D6 = 1'b1;
  assign CLBLM_L_X10Y152_SLICE_X13Y152_C6 = CLBLM_L_X10Y152_SLICE_X12Y152_BQ;
  assign CLBLM_L_X8Y142_SLICE_X10Y142_D1 = CLBLM_R_X7Y141_SLICE_X9Y141_AQ;
  assign CLBLM_L_X8Y142_SLICE_X10Y142_D2 = CLBLM_L_X8Y142_SLICE_X10Y142_CQ;
  assign CLBLM_L_X8Y142_SLICE_X10Y142_D3 = CLBLM_L_X10Y142_SLICE_X12Y142_CO6;
  assign CLBLM_L_X10Y152_SLICE_X13Y152_CLK = CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O;
  assign CLBLM_L_X8Y142_SLICE_X10Y142_D4 = CLBLM_R_X7Y143_SLICE_X9Y143_CQ;
  assign CLBLM_L_X8Y142_SLICE_X10Y142_D5 = CLBLM_L_X8Y145_SLICE_X11Y145_DQ;
  assign CLBLM_L_X8Y142_SLICE_X10Y142_D6 = RIOB33_X105Y131_IOB_X1Y131_I;
  assign RIOI3_X105Y141_ILOGIC_X1Y141_D = RIOB33_X105Y141_IOB_X1Y141_I;
  assign CLBLM_R_X11Y146_SLICE_X15Y146_A1 = CLBLM_R_X7Y146_SLICE_X8Y146_A5Q;
  assign CLBLM_R_X11Y146_SLICE_X15Y146_A2 = CLBLM_L_X12Y146_SLICE_X16Y146_BQ;
  assign CLBLM_R_X11Y146_SLICE_X15Y146_A3 = CLBLM_L_X8Y146_SLICE_X10Y146_BQ;
  assign CLBLM_R_X11Y146_SLICE_X15Y146_A4 = CLBLM_R_X5Y152_SLICE_X7Y152_C5Q;
  assign CLBLM_L_X10Y152_SLICE_X13Y152_D2 = CLBLM_L_X10Y153_SLICE_X13Y153_CQ;
  assign CLBLM_R_X11Y146_SLICE_X15Y146_A5 = RIOB33_X105Y145_IOB_X1Y145_I;
  assign CLBLM_R_X11Y146_SLICE_X15Y146_A6 = 1'b1;
  assign CLBLM_L_X10Y152_SLICE_X13Y152_D3 = CLBLM_R_X11Y153_SLICE_X14Y153_AQ;
  assign CLBLM_R_X11Y146_SLICE_X15Y146_B1 = CLBLM_R_X7Y153_SLICE_X8Y153_A5Q;
  assign CLBLM_R_X11Y146_SLICE_X15Y146_B2 = CLBLM_L_X12Y145_SLICE_X17Y145_CO6;
  assign CLBLM_R_X11Y146_SLICE_X15Y146_B3 = CLBLM_L_X8Y146_SLICE_X10Y146_BQ;
  assign CLBLM_R_X11Y146_SLICE_X15Y146_B4 = CLBLM_R_X7Y144_SLICE_X9Y144_B5Q;
  assign CLBLM_R_X11Y146_SLICE_X15Y146_B5 = CLBLM_R_X5Y152_SLICE_X7Y152_C5Q;
  assign CLBLM_R_X11Y146_SLICE_X15Y146_B6 = 1'b1;
  assign CLBLM_L_X10Y152_SLICE_X13Y152_D5 = CLBLM_R_X5Y147_SLICE_X6Y147_AQ;
  assign CLBLM_R_X11Y146_SLICE_X15Y146_C1 = CLBLM_L_X12Y145_SLICE_X17Y145_CO6;
  assign CLBLM_R_X11Y146_SLICE_X15Y146_C2 = CLBLM_L_X10Y146_SLICE_X13Y146_AQ;
  assign CLBLM_R_X11Y146_SLICE_X15Y146_C3 = CLBLM_R_X11Y147_SLICE_X14Y147_AO5;
  assign CLBLM_R_X11Y146_SLICE_X15Y146_C4 = CLBLM_L_X10Y147_SLICE_X12Y147_CQ;
  assign CLBLM_L_X10Y152_SLICE_X13Y152_D6 = CLBLM_R_X7Y146_SLICE_X8Y146_A5Q;
  assign CLBLM_R_X11Y146_SLICE_X15Y146_C5 = CLBLM_R_X7Y146_SLICE_X9Y146_CO6;
  assign CLBLM_R_X11Y146_SLICE_X15Y146_C6 = CLBLM_R_X11Y146_SLICE_X15Y146_BO6;
  assign CLBLM_R_X11Y146_SLICE_X15Y146_D1 = CLBLM_L_X12Y145_SLICE_X17Y145_AO5;
  assign CLBLM_R_X11Y146_SLICE_X15Y146_D2 = CLBLM_L_X12Y146_SLICE_X16Y146_CO6;
  assign CLBLM_R_X11Y146_SLICE_X15Y146_D3 = 1'b1;
  assign CLBLM_R_X11Y146_SLICE_X15Y146_D4 = CLBLM_R_X13Y146_SLICE_X18Y146_AO5;
  assign CLBLL_L_X4Y149_SLICE_X4Y149_A1 = CLBLL_L_X4Y146_SLICE_X4Y146_DO6;
  assign CLBLL_L_X4Y149_SLICE_X4Y149_A2 = 1'b1;
  assign CLBLL_L_X4Y149_SLICE_X4Y149_A3 = CLBLL_L_X4Y149_SLICE_X4Y149_AQ;
  assign CLBLL_L_X4Y149_SLICE_X4Y149_A4 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLL_L_X4Y149_SLICE_X4Y149_A5 = CLBLL_L_X4Y143_SLICE_X4Y143_D5Q;
  assign CLBLL_L_X4Y149_SLICE_X4Y149_A6 = CLBLM_R_X5Y149_SLICE_X6Y149_AQ;
  assign CLBLM_R_X11Y146_SLICE_X15Y146_D5 = LIOB33_X0Y53_IOB_X0Y53_I;
  assign CLBLM_R_X11Y146_SLICE_X15Y146_D6 = CLBLM_L_X8Y146_SLICE_X11Y146_AQ;
  assign CLBLM_R_X11Y146_SLICE_X14Y146_A1 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLL_L_X4Y149_SLICE_X4Y149_B1 = CLBLM_R_X3Y149_SLICE_X2Y149_AQ;
  assign CLBLL_L_X4Y149_SLICE_X4Y149_B2 = CLBLL_L_X4Y149_SLICE_X4Y149_BQ;
  assign CLBLL_L_X4Y149_SLICE_X4Y149_B3 = CLBLM_R_X5Y152_SLICE_X6Y152_DQ;
  assign CLBLL_L_X4Y149_SLICE_X4Y149_B4 = CLBLM_L_X8Y147_SLICE_X10Y147_BQ;
  assign CLBLL_L_X4Y149_SLICE_X4Y149_B5 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLL_L_X4Y149_SLICE_X4Y149_B6 = 1'b1;
  assign CLBLM_R_X11Y146_SLICE_X14Y146_A2 = CLBLM_L_X10Y147_SLICE_X12Y147_CQ;
  assign CLBLM_R_X11Y146_SLICE_X14Y146_A3 = CLBLM_R_X11Y146_SLICE_X14Y146_AQ;
  assign CLBLM_R_X11Y146_SLICE_X14Y146_A4 = 1'b1;
  assign CLBLL_L_X4Y149_SLICE_X4Y149_C1 = CLBLL_L_X4Y147_SLICE_X5Y147_C5Q;
  assign CLBLL_L_X4Y149_SLICE_X4Y149_C2 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLL_L_X4Y149_SLICE_X4Y149_C3 = CLBLL_L_X4Y149_SLICE_X4Y149_DQ;
  assign CLBLL_L_X4Y149_SLICE_X4Y149_C4 = CLBLM_L_X8Y145_SLICE_X11Y145_DQ;
  assign CLBLL_L_X4Y149_SLICE_X4Y149_C5 = 1'b1;
  assign CLBLL_L_X4Y149_SLICE_X4Y149_C6 = CLBLM_L_X8Y151_SLICE_X10Y151_AQ;
  assign CLBLM_R_X11Y146_SLICE_X14Y146_B1 = CLBLM_L_X8Y142_SLICE_X11Y142_BQ;
  assign CLBLL_L_X4Y149_SLICE_X4Y149_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X11Y146_SLICE_X14Y146_B2 = RIOB33_X105Y131_IOB_X1Y131_I;
  assign CLBLM_R_X11Y146_SLICE_X14Y146_B3 = CLBLM_L_X8Y145_SLICE_X11Y145_DQ;
  assign CLBLM_R_X11Y146_SLICE_X14Y146_B4 = CLBLL_L_X4Y151_SLICE_X4Y151_CQ;
  assign CLBLM_R_X11Y146_SLICE_X14Y146_B5 = 1'b1;
  assign CLBLL_L_X4Y149_SLICE_X4Y149_D1 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLL_L_X4Y149_SLICE_X4Y149_D2 = CLBLM_L_X10Y151_SLICE_X12Y151_DQ;
  assign CLBLL_L_X4Y149_SLICE_X4Y149_D3 = CLBLL_L_X4Y149_SLICE_X4Y149_DQ;
  assign CLBLL_L_X4Y149_SLICE_X4Y149_D4 = CLBLM_L_X10Y148_SLICE_X13Y148_AQ;
  assign CLBLL_L_X4Y149_SLICE_X4Y149_D5 = CLBLL_L_X4Y149_SLICE_X4Y149_D5Q;
  assign CLBLL_L_X4Y149_SLICE_X4Y149_D6 = 1'b1;
  assign CLBLM_R_X11Y146_SLICE_X14Y146_C3 = CLBLL_L_X4Y148_SLICE_X4Y148_CQ;
  assign CLBLM_R_X11Y146_SLICE_X14Y146_C4 = CLBLM_R_X7Y153_SLICE_X8Y153_A5Q;
  assign CLBLM_R_X11Y146_SLICE_X14Y146_C6 = 1'b1;
  assign CLBLM_R_X11Y146_SLICE_X14Y146_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X11Y146_SLICE_X14Y146_D1 = CLBLM_L_X10Y146_SLICE_X13Y146_DO6;
  assign CLBLM_R_X11Y146_SLICE_X14Y146_D2 = CLBLM_R_X7Y153_SLICE_X8Y153_A5Q;
  assign CLBLM_R_X11Y146_SLICE_X14Y146_D3 = CLBLL_L_X4Y148_SLICE_X4Y148_CQ;
  assign CLBLM_R_X11Y146_SLICE_X14Y146_D4 = CLBLM_R_X7Y149_SLICE_X8Y149_AQ;
  assign CLBLM_R_X11Y146_SLICE_X14Y146_D5 = CLBLM_R_X7Y146_SLICE_X9Y146_CO6;
  assign CLBLM_R_X11Y146_SLICE_X14Y146_D6 = CLBLM_R_X7Y144_SLICE_X9Y144_B5Q;
  assign LIOI3_SING_X0Y100_OLOGIC_X0Y100_D1 = CLBLM_R_X3Y148_SLICE_X2Y148_B5Q;
  assign LIOI3_SING_X0Y100_OLOGIC_X0Y100_T1 = 1'b1;
  assign CLBLL_L_X4Y149_SLICE_X5Y149_A1 = 1'b1;
  assign CLBLL_L_X4Y149_SLICE_X5Y149_A2 = CLBLM_R_X3Y143_SLICE_X3Y143_BQ;
  assign CLBLL_L_X4Y149_SLICE_X5Y149_A3 = CLBLL_L_X4Y142_SLICE_X4Y142_AQ;
  assign CLBLL_L_X4Y149_SLICE_X5Y149_A4 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLL_L_X4Y149_SLICE_X5Y149_A5 = CLBLM_L_X10Y151_SLICE_X13Y151_A5Q;
  assign CLBLL_L_X4Y149_SLICE_X5Y149_A6 = CLBLM_R_X7Y142_SLICE_X8Y142_C5Q;
  assign CLBLL_L_X4Y149_SLICE_X5Y149_B1 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLL_L_X4Y149_SLICE_X5Y149_B2 = CLBLM_R_X7Y148_SLICE_X9Y148_BQ;
  assign CLBLL_L_X4Y149_SLICE_X5Y149_B3 = CLBLL_L_X4Y149_SLICE_X5Y149_AQ;
  assign CLBLL_L_X4Y149_SLICE_X5Y149_B4 = CLBLM_R_X3Y143_SLICE_X3Y143_BQ;
  assign CLBLL_L_X4Y149_SLICE_X5Y149_B5 = CLBLL_L_X4Y149_SLICE_X5Y149_C5Q;
  assign CLBLL_L_X4Y149_SLICE_X5Y149_B6 = CLBLL_L_X4Y142_SLICE_X4Y142_AQ;
  assign CLBLL_L_X4Y149_SLICE_X5Y149_C1 = 1'b1;
  assign CLBLL_L_X4Y149_SLICE_X5Y149_C2 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLL_L_X4Y149_SLICE_X5Y149_C3 = CLBLM_R_X5Y150_SLICE_X6Y150_C5Q;
  assign CLBLL_L_X4Y149_SLICE_X5Y149_C4 = CLBLM_R_X5Y149_SLICE_X6Y149_C5Q;
  assign CLBLL_L_X4Y149_SLICE_X5Y149_C5 = CLBLM_L_X8Y149_SLICE_X11Y149_BO6;
  assign CLBLL_L_X4Y149_SLICE_X5Y149_C6 = 1'b1;
  assign CLBLL_L_X4Y149_SLICE_X5Y149_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X10Y152_SLICE_X12Y152_B5 = CLBLM_R_X7Y146_SLICE_X8Y146_A5Q;
  assign CLBLL_L_X4Y149_SLICE_X5Y149_D1 = CLBLL_L_X4Y151_SLICE_X4Y151_AQ;
  assign CLBLL_L_X4Y149_SLICE_X5Y149_D2 = CLBLL_L_X4Y143_SLICE_X4Y143_AQ;
  assign CLBLL_L_X4Y149_SLICE_X5Y149_D3 = CLBLL_L_X4Y143_SLICE_X4Y143_BQ;
  assign CLBLL_L_X4Y149_SLICE_X5Y149_D4 = CLBLL_L_X4Y151_SLICE_X5Y151_CQ;
  assign CLBLL_L_X4Y149_SLICE_X5Y149_D5 = CLBLL_L_X2Y145_SLICE_X0Y145_AQ;
  assign CLBLL_L_X4Y149_SLICE_X5Y149_D6 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_L_X10Y152_SLICE_X12Y152_B6 = CLBLL_L_X4Y147_SLICE_X5Y147_CQ;
  assign CLBLM_L_X10Y153_SLICE_X13Y153_A1 = CLBLM_L_X10Y154_SLICE_X13Y154_BO5;
  assign CLBLM_L_X10Y153_SLICE_X13Y153_A2 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_L_X10Y153_SLICE_X13Y153_A3 = CLBLM_L_X10Y153_SLICE_X13Y153_AQ;
  assign CLBLM_L_X10Y153_SLICE_X13Y153_A4 = CLBLM_L_X10Y155_SLICE_X12Y155_BO5;
  assign CLBLM_L_X10Y153_SLICE_X13Y153_A5 = CLBLM_R_X7Y151_SLICE_X9Y151_BQ;
  assign CLBLM_L_X10Y153_SLICE_X13Y153_A6 = CLBLM_L_X10Y154_SLICE_X13Y154_CO6;
  assign CLBLM_L_X10Y153_SLICE_X13Y153_AX = CLBLM_L_X12Y153_SLICE_X16Y153_AO5;
  assign CLBLM_L_X10Y153_SLICE_X13Y153_B1 = CLBLM_R_X11Y153_SLICE_X15Y153_CO6;
  assign CLBLM_L_X10Y153_SLICE_X13Y153_B2 = CLBLM_L_X10Y153_SLICE_X13Y153_BQ;
  assign CLBLM_L_X10Y153_SLICE_X13Y153_B3 = CLBLM_R_X11Y153_SLICE_X15Y153_DO6;
  assign CLBLM_L_X10Y153_SLICE_X13Y153_B4 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_L_X10Y153_SLICE_X13Y153_B5 = CLBLL_L_X4Y151_SLICE_X5Y151_BQ;
  assign CLBLM_L_X10Y153_SLICE_X13Y153_B6 = CLBLM_R_X11Y153_SLICE_X15Y153_BO5;
  assign CLBLM_L_X8Y143_SLICE_X11Y143_A1 = CLBLM_R_X7Y152_SLICE_X8Y152_D5Q;
  assign CLBLM_L_X10Y153_SLICE_X13Y153_C2 = CLBLM_R_X7Y146_SLICE_X8Y146_A5Q;
  assign CLBLM_L_X10Y153_SLICE_X13Y153_C3 = CLBLM_L_X10Y153_SLICE_X13Y153_CQ;
  assign CLBLM_L_X10Y153_SLICE_X13Y153_C4 = CLBLM_L_X10Y154_SLICE_X13Y154_CO6;
  assign CLBLM_L_X10Y153_SLICE_X13Y153_C5 = CLBLM_L_X10Y153_SLICE_X13Y153_AQ;
  assign CLBLM_L_X10Y153_SLICE_X13Y153_C6 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_L_X8Y143_SLICE_X11Y143_A2 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_L_X8Y143_SLICE_X11Y143_A3 = CLBLM_L_X8Y143_SLICE_X11Y143_AQ;
  assign CLBLM_L_X8Y143_SLICE_X11Y143_A4 = CLBLM_L_X10Y143_SLICE_X12Y143_AQ;
  assign CLBLM_L_X8Y143_SLICE_X11Y143_A5 = CLBLM_R_X7Y142_SLICE_X8Y142_C5Q;
  assign CLBLM_L_X8Y143_SLICE_X11Y143_A6 = CLBLM_R_X7Y145_SLICE_X8Y145_D5Q;
  assign CLBLM_L_X10Y152_SLICE_X12Y152_C5 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_L_X8Y143_SLICE_X11Y143_B1 = CLBLM_R_X13Y149_SLICE_X18Y149_AO6;
  assign CLBLM_L_X8Y143_SLICE_X11Y143_B2 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_L_X10Y153_SLICE_X13Y153_D1 = CLBLM_L_X10Y155_SLICE_X12Y155_BO5;
  assign CLBLM_L_X10Y153_SLICE_X13Y153_D2 = CLBLM_L_X10Y155_SLICE_X13Y155_AO5;
  assign CLBLM_L_X8Y143_SLICE_X11Y143_B3 = 1'b1;
  assign CLBLM_L_X8Y143_SLICE_X11Y143_B4 = CLBLM_L_X8Y145_SLICE_X11Y145_BQ;
  assign CLBLM_L_X10Y153_SLICE_X13Y153_D5 = CLBLM_L_X10Y152_SLICE_X12Y152_AQ;
  assign CLBLM_L_X10Y153_SLICE_X13Y153_D6 = CLBLM_R_X11Y153_SLICE_X14Y153_AQ;
  assign CLBLM_L_X8Y143_SLICE_X11Y143_B5 = CLBLM_R_X7Y141_SLICE_X9Y141_AQ;
  assign CLBLM_L_X8Y143_SLICE_X11Y143_B6 = CLBLM_L_X8Y143_SLICE_X11Y143_BQ;
  assign CLBLM_L_X8Y143_SLICE_X11Y143_C1 = CLBLL_L_X4Y149_SLICE_X5Y149_C5Q;
  assign CLBLM_L_X8Y143_SLICE_X11Y143_C2 = CLBLM_L_X8Y143_SLICE_X11Y143_CQ;
  assign CLBLM_L_X8Y143_SLICE_X11Y143_C3 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_L_X8Y143_SLICE_X11Y143_C4 = CLBLM_L_X12Y149_SLICE_X17Y149_CO6;
  assign CLBLM_L_X8Y143_SLICE_X11Y143_C5 = CLBLM_L_X8Y143_SLICE_X10Y143_DQ;
  assign CLBLM_L_X8Y143_SLICE_X11Y143_C6 = 1'b1;
  assign CLBLM_L_X8Y143_SLICE_X11Y143_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X10Y153_SLICE_X12Y153_A1 = CLBLM_R_X7Y154_SLICE_X8Y154_DO6;
  assign CLBLM_L_X10Y153_SLICE_X12Y153_A2 = CLBLM_L_X10Y153_SLICE_X12Y153_BQ;
  assign CLBLM_L_X10Y153_SLICE_X12Y153_A3 = 1'b1;
  assign CLBLM_L_X10Y153_SLICE_X12Y153_A4 = CLBLM_L_X10Y153_SLICE_X13Y153_BQ;
  assign CLBLM_L_X10Y153_SLICE_X12Y153_A5 = 1'b1;
  assign CLBLM_L_X8Y143_SLICE_X11Y143_D1 = CLBLL_L_X4Y143_SLICE_X4Y143_AQ;
  assign CLBLM_L_X8Y143_SLICE_X11Y143_D2 = CLBLM_L_X10Y143_SLICE_X13Y143_BQ;
  assign CLBLM_L_X8Y143_SLICE_X11Y143_D3 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_L_X8Y143_SLICE_X11Y143_D4 = 1'b1;
  assign CLBLM_L_X8Y143_SLICE_X11Y143_D5 = CLBLM_L_X8Y143_SLICE_X10Y143_DQ;
  assign CLBLM_L_X10Y153_SLICE_X12Y153_B5 = CLBLM_L_X12Y146_SLICE_X16Y146_BQ;
  assign CLBLM_L_X10Y153_SLICE_X12Y153_B6 = CLBLM_R_X5Y150_SLICE_X6Y150_B5Q;
  assign CLBLM_L_X8Y143_SLICE_X11Y143_D6 = 1'b1;
  assign CLBLM_L_X10Y153_SLICE_X12Y153_AX = CLBLM_L_X10Y153_SLICE_X12Y153_CO6;
  assign CLBLM_L_X10Y153_SLICE_X12Y153_B2 = CLBLM_L_X10Y153_SLICE_X12Y153_BQ;
  assign CLBLM_L_X10Y153_SLICE_X12Y153_B3 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_L_X10Y153_SLICE_X12Y153_B4 = CLBLM_R_X5Y152_SLICE_X6Y152_BQ;
  assign CLBLM_L_X8Y143_SLICE_X10Y143_A1 = CLBLM_L_X10Y144_SLICE_X13Y144_A5Q;
  assign CLBLM_L_X8Y143_SLICE_X10Y143_A2 = CLBLM_L_X8Y151_SLICE_X10Y151_BQ;
  assign CLBLM_L_X10Y153_SLICE_X12Y153_C5 = CLBLM_R_X5Y152_SLICE_X6Y152_BQ;
  assign CLBLM_L_X10Y153_SLICE_X12Y153_C6 = 1'b1;
  assign CLBLM_L_X8Y143_SLICE_X10Y143_A3 = CLBLM_L_X8Y143_SLICE_X10Y143_AQ;
  assign CLBLM_L_X8Y143_SLICE_X10Y143_A4 = CLBLM_L_X10Y144_SLICE_X12Y144_AO6;
  assign CLBLM_L_X8Y143_SLICE_X10Y143_A5 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_L_X8Y143_SLICE_X10Y143_A6 = CLBLM_R_X3Y142_SLICE_X2Y142_BO5;
  assign CLBLM_L_X10Y153_SLICE_X12Y153_C2 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_L_X10Y153_SLICE_X12Y153_C3 = CLBLM_L_X10Y153_SLICE_X12Y153_A5Q;
  assign CLBLM_L_X8Y143_SLICE_X10Y143_B1 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_L_X8Y143_SLICE_X10Y143_B2 = CLBLM_L_X8Y143_SLICE_X10Y143_BQ;
  assign CLBLM_L_X8Y143_SLICE_X10Y143_B3 = CLBLM_L_X10Y144_SLICE_X13Y144_CQ;
  assign CLBLM_L_X8Y143_SLICE_X10Y143_B4 = CLBLM_L_X10Y143_SLICE_X12Y143_CO6;
  assign CLBLM_L_X8Y143_SLICE_X10Y143_B5 = CLBLM_L_X8Y149_SLICE_X11Y149_AQ;
  assign CLBLM_L_X8Y143_SLICE_X10Y143_B6 = CLBLM_L_X8Y151_SLICE_X10Y151_CQ;
  assign CLBLM_L_X10Y153_SLICE_X12Y153_D1 = CLBLM_L_X10Y145_SLICE_X12Y145_BQ;
  assign CLBLM_L_X10Y153_SLICE_X12Y153_D2 = CLBLM_L_X8Y154_SLICE_X10Y154_BO5;
  assign CLBLM_L_X8Y143_SLICE_X10Y143_C1 = CLBLM_L_X8Y142_SLICE_X10Y142_AQ;
  assign CLBLM_L_X8Y143_SLICE_X10Y143_C2 = CLBLM_L_X8Y143_SLICE_X10Y143_CQ;
  assign CLBLM_L_X8Y143_SLICE_X10Y143_C3 = CLBLL_L_X4Y142_SLICE_X5Y142_DQ;
  assign CLBLM_L_X8Y143_SLICE_X10Y143_C4 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_L_X8Y143_SLICE_X10Y143_C5 = CLBLM_R_X5Y143_SLICE_X7Y143_CQ;
  assign CLBLM_L_X8Y143_SLICE_X10Y143_C6 = CLBLL_L_X4Y147_SLICE_X5Y147_CQ;
  assign CLBLM_L_X10Y153_SLICE_X12Y153_D5 = RIOB33_SING_X105Y100_IOB_X1Y100_I;
  assign CLBLM_L_X8Y143_SLICE_X10Y143_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign RIOI3_X105Y197_OLOGIC_X1Y197_T1 = 1'b1;
  assign CLBLM_L_X8Y143_SLICE_X10Y143_D1 = CLBLL_L_X4Y151_SLICE_X4Y151_BQ;
  assign CLBLM_L_X8Y143_SLICE_X10Y143_D2 = CLBLM_R_X3Y145_SLICE_X3Y145_D5Q;
  assign CLBLM_L_X8Y143_SLICE_X10Y143_D3 = CLBLM_L_X8Y143_SLICE_X10Y143_DQ;
  assign CLBLM_L_X8Y143_SLICE_X10Y143_D4 = CLBLM_R_X5Y146_SLICE_X7Y146_DQ;
  assign CLBLM_L_X8Y143_SLICE_X10Y143_D5 = CLBLM_R_X7Y148_SLICE_X9Y148_C5Q;
  assign CLBLM_L_X8Y143_SLICE_X10Y143_D6 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign RIOI3_TBYTESRC_X105Y169_OLOGIC_X1Y170_D1 = CLBLM_R_X3Y152_SLICE_X3Y152_BQ;
  assign RIOI3_TBYTESRC_X105Y169_OLOGIC_X1Y170_T1 = 1'b1;
  assign CLBLM_R_X11Y147_SLICE_X15Y147_A1 = CLBLM_L_X10Y148_SLICE_X13Y148_AQ;
  assign CLBLM_R_X11Y147_SLICE_X15Y147_A2 = CLBLM_R_X11Y146_SLICE_X15Y146_DO6;
  assign CLBLM_R_X11Y147_SLICE_X15Y147_A3 = CLBLM_R_X11Y144_SLICE_X14Y144_DO6;
  assign CLBLM_R_X11Y147_SLICE_X15Y147_A4 = CLBLM_L_X12Y146_SLICE_X17Y146_DO6;
  assign CLBLM_R_X11Y147_SLICE_X15Y147_A5 = CLBLM_R_X13Y146_SLICE_X18Y146_BO6;
  assign CLBLM_R_X11Y147_SLICE_X15Y147_A6 = CLBLM_L_X12Y145_SLICE_X16Y145_BO6;
  assign RIOI3_TBYTESRC_X105Y169_OLOGIC_X1Y169_D1 = CLBLM_R_X3Y152_SLICE_X3Y152_CQ;
  assign CLBLM_R_X11Y148_SLICE_X15Y148_D2 = CLBLM_L_X12Y147_SLICE_X16Y147_DO6;
  assign CLBLM_R_X11Y147_SLICE_X15Y147_B1 = CLBLL_L_X4Y147_SLICE_X4Y147_CQ;
  assign CLBLM_R_X11Y147_SLICE_X15Y147_B2 = CLBLM_R_X7Y151_SLICE_X8Y151_D5Q;
  assign CLBLM_R_X11Y147_SLICE_X15Y147_B3 = CLBLM_R_X5Y142_SLICE_X6Y142_D5Q;
  assign CLBLM_R_X11Y147_SLICE_X15Y147_B4 = CLBLL_L_X4Y148_SLICE_X4Y148_CQ;
  assign CLBLM_R_X11Y147_SLICE_X15Y147_B5 = CLBLM_R_X7Y149_SLICE_X8Y149_AQ;
  assign CLBLM_R_X11Y147_SLICE_X15Y147_B6 = CLBLM_L_X10Y146_SLICE_X12Y146_DQ;
  assign CLBLM_R_X11Y148_SLICE_X15Y148_D3 = CLBLM_R_X11Y148_SLICE_X14Y148_DO6;
  assign LIOB33_X0Y143_IOB_X0Y143_O = CLBLM_R_X3Y151_SLICE_X2Y151_BO5;
  assign RIOI3_TBYTESRC_X105Y169_OLOGIC_X1Y169_T1 = 1'b1;
  assign CLBLM_R_X11Y147_SLICE_X15Y147_C1 = CLBLM_R_X11Y147_SLICE_X14Y147_BO6;
  assign CLBLM_R_X11Y147_SLICE_X15Y147_C2 = CLBLM_R_X11Y146_SLICE_X15Y146_DO6;
  assign CLBLM_R_X11Y147_SLICE_X15Y147_C3 = CLBLM_L_X8Y146_SLICE_X10Y146_BO5;
  assign CLBLM_R_X11Y147_SLICE_X15Y147_C4 = CLBLM_L_X12Y146_SLICE_X17Y146_DO6;
  assign CLBLM_R_X11Y147_SLICE_X15Y147_C5 = CLBLM_R_X11Y144_SLICE_X14Y144_DO6;
  assign CLBLM_R_X11Y147_SLICE_X15Y147_C6 = CLBLM_L_X8Y146_SLICE_X10Y146_CO6;
  assign CLBLM_R_X11Y148_SLICE_X15Y148_D5 = CLBLM_R_X7Y147_SLICE_X8Y147_DO6;
  assign CLBLM_R_X11Y148_SLICE_X15Y148_D6 = CLBLM_R_X11Y150_SLICE_X15Y150_BO6;
  assign CLBLL_L_X4Y150_SLICE_X4Y150_A1 = CLBLL_L_X4Y153_SLICE_X4Y153_B5Q;
  assign CLBLL_L_X4Y150_SLICE_X4Y150_A2 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLL_L_X4Y150_SLICE_X4Y150_A3 = CLBLM_L_X10Y149_SLICE_X12Y149_BQ;
  assign CLBLL_L_X4Y150_SLICE_X4Y150_A4 = CLBLL_L_X4Y145_SLICE_X4Y145_BQ;
  assign CLBLL_L_X4Y150_SLICE_X4Y150_A5 = 1'b1;
  assign CLBLL_L_X4Y150_SLICE_X4Y150_A6 = 1'b1;
  assign CLBLM_R_X11Y147_SLICE_X15Y147_D1 = CLBLM_L_X12Y147_SLICE_X16Y147_AO6;
  assign CLBLM_R_X11Y147_SLICE_X15Y147_D2 = CLBLM_L_X12Y145_SLICE_X16Y145_BO6;
  assign CLBLM_R_X11Y147_SLICE_X15Y147_D3 = CLBLM_R_X11Y146_SLICE_X14Y146_DO6;
  assign CLBLL_L_X4Y150_SLICE_X4Y150_B1 = CLBLM_R_X3Y151_SLICE_X2Y151_CO6;
  assign CLBLL_L_X4Y150_SLICE_X4Y150_B2 = CLBLM_R_X3Y145_SLICE_X2Y145_CQ;
  assign CLBLL_L_X4Y150_SLICE_X4Y150_B3 = CLBLL_L_X4Y149_SLICE_X5Y149_BQ;
  assign CLBLL_L_X4Y150_SLICE_X4Y150_B4 = CLBLM_R_X5Y143_SLICE_X7Y143_AQ;
  assign CLBLL_L_X4Y150_SLICE_X4Y150_B5 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLL_L_X4Y150_SLICE_X4Y150_B6 = 1'b1;
  assign CLBLM_R_X11Y147_SLICE_X14Y147_A4 = CLBLL_L_X4Y148_SLICE_X4Y148_CQ;
  assign CLBLM_R_X11Y147_SLICE_X14Y147_A5 = CLBLM_R_X7Y144_SLICE_X9Y144_B5Q;
  assign CLBLM_R_X11Y147_SLICE_X14Y147_A6 = 1'b1;
  assign CLBLL_L_X4Y150_SLICE_X4Y150_C1 = CLBLM_L_X10Y149_SLICE_X12Y149_BQ;
  assign CLBLL_L_X4Y150_SLICE_X4Y150_C2 = CLBLL_L_X4Y150_SLICE_X5Y150_BQ;
  assign CLBLL_L_X4Y150_SLICE_X4Y150_C3 = CLBLL_L_X4Y150_SLICE_X4Y150_BQ;
  assign CLBLL_L_X4Y150_SLICE_X4Y150_C4 = 1'b1;
  assign CLBLL_L_X4Y150_SLICE_X4Y150_C5 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLL_L_X4Y150_SLICE_X4Y150_C6 = 1'b1;
  assign CLBLM_R_X11Y147_SLICE_X14Y147_B1 = CLBLM_L_X10Y148_SLICE_X13Y148_AQ;
  assign CLBLL_L_X4Y150_SLICE_X4Y150_CLK = CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O;
  assign CLBLM_R_X11Y147_SLICE_X14Y147_B2 = CLBLM_R_X3Y146_SLICE_X2Y146_AQ;
  assign CLBLM_R_X11Y147_SLICE_X14Y147_B3 = CLBLM_R_X13Y146_SLICE_X18Y146_BO6;
  assign CLBLM_R_X11Y147_SLICE_X14Y147_B4 = CLBLM_L_X12Y145_SLICE_X16Y145_BO6;
  assign CLBLM_R_X11Y147_SLICE_X14Y147_B5 = 1'b1;
  assign CLBLM_R_X11Y147_SLICE_X14Y147_B6 = 1'b1;
  assign CLBLL_L_X4Y150_SLICE_X4Y150_D1 = CLBLM_R_X3Y151_SLICE_X3Y151_AQ;
  assign CLBLL_L_X4Y150_SLICE_X4Y150_D2 = CLBLL_L_X4Y145_SLICE_X5Y145_BQ;
  assign CLBLL_L_X4Y150_SLICE_X4Y150_D3 = CLBLL_L_X4Y150_SLICE_X5Y150_CO5;
  assign CLBLL_L_X4Y150_SLICE_X4Y150_D4 = CLBLM_R_X3Y151_SLICE_X3Y151_CQ;
  assign CLBLL_L_X4Y150_SLICE_X4Y150_D5 = CLBLL_L_X4Y150_SLICE_X4Y150_B5Q;
  assign CLBLL_L_X4Y150_SLICE_X4Y150_D6 = CLBLM_R_X3Y151_SLICE_X3Y151_BQ;
  assign CLBLM_R_X11Y147_SLICE_X14Y147_C1 = CLBLM_R_X11Y145_SLICE_X14Y145_AO6;
  assign CLBLM_R_X11Y147_SLICE_X14Y147_C2 = CLBLM_R_X11Y144_SLICE_X14Y144_DO6;
  assign CLBLM_R_X11Y147_SLICE_X14Y147_C3 = CLBLM_R_X13Y146_SLICE_X18Y146_BO6;
  assign CLBLM_R_X11Y147_SLICE_X14Y147_C4 = CLBLM_R_X11Y145_SLICE_X15Y145_CO6;
  assign CLBLM_R_X11Y147_SLICE_X14Y147_C5 = CLBLM_R_X3Y146_SLICE_X2Y146_AQ;
  assign CLBLM_R_X11Y147_SLICE_X14Y147_C6 = CLBLM_L_X12Y145_SLICE_X16Y145_BO6;
  assign CLBLM_R_X11Y148_SLICE_X14Y148_A3 = CLBLM_R_X11Y148_SLICE_X15Y148_CO6;
  assign CLBLM_R_X11Y147_SLICE_X14Y147_D1 = CLBLM_R_X11Y145_SLICE_X14Y145_AO6;
  assign CLBLM_R_X11Y147_SLICE_X14Y147_D2 = CLBLM_R_X11Y144_SLICE_X14Y144_DO6;
  assign CLBLM_R_X11Y147_SLICE_X14Y147_D3 = CLBLM_L_X10Y148_SLICE_X12Y148_DO6;
  assign CLBLM_R_X11Y147_SLICE_X14Y147_D4 = CLBLM_L_X8Y146_SLICE_X10Y146_DO6;
  assign CLBLM_R_X11Y147_SLICE_X14Y147_D5 = CLBLM_R_X11Y147_SLICE_X14Y147_BO5;
  assign CLBLM_R_X11Y147_SLICE_X14Y147_D6 = CLBLM_R_X11Y145_SLICE_X15Y145_CO6;
  assign CLBLM_R_X11Y148_SLICE_X14Y148_A4 = CLBLM_L_X8Y148_SLICE_X10Y148_CO6;
  assign CLBLL_L_X4Y150_SLICE_X5Y150_A1 = CLBLL_L_X4Y150_SLICE_X5Y150_DO6;
  assign CLBLL_L_X4Y150_SLICE_X5Y150_A2 = CLBLM_R_X5Y145_SLICE_X6Y145_CQ;
  assign CLBLL_L_X4Y150_SLICE_X5Y150_A3 = 1'b1;
  assign CLBLL_L_X4Y150_SLICE_X5Y150_A4 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLL_L_X4Y150_SLICE_X5Y150_A5 = 1'b1;
  assign CLBLL_L_X4Y150_SLICE_X5Y150_A6 = CLBLL_L_X4Y150_SLICE_X5Y150_CO6;
  assign CLBLL_L_X4Y150_SLICE_X5Y150_AX = CLBLL_L_X4Y153_SLICE_X4Y153_CO6;
  assign CLBLL_L_X4Y150_SLICE_X5Y150_B1 = CLBLM_R_X7Y152_SLICE_X8Y152_D5Q;
  assign CLBLL_L_X4Y150_SLICE_X5Y150_B2 = CLBLL_L_X4Y150_SLICE_X5Y150_BQ;
  assign CLBLL_L_X4Y150_SLICE_X5Y150_B3 = CLBLM_R_X7Y142_SLICE_X8Y142_C5Q;
  assign CLBLL_L_X4Y150_SLICE_X5Y150_B4 = CLBLL_L_X4Y148_SLICE_X5Y148_D5Q;
  assign CLBLL_L_X4Y150_SLICE_X5Y150_B5 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLL_L_X4Y150_SLICE_X5Y150_B6 = CLBLM_R_X5Y151_SLICE_X6Y151_BQ;
  assign CLBLM_R_X7Y150_SLICE_X9Y150_C4 = CLBLM_L_X12Y147_SLICE_X16Y147_DO6;
  assign CLBLM_R_X7Y150_SLICE_X9Y150_C5 = CLBLM_R_X3Y147_SLICE_X3Y147_AQ;
  assign CLBLL_L_X4Y150_SLICE_X5Y150_C1 = CLBLM_R_X3Y151_SLICE_X3Y151_AQ;
  assign CLBLL_L_X4Y150_SLICE_X5Y150_C2 = CLBLM_R_X3Y145_SLICE_X3Y145_BQ;
  assign CLBLL_L_X4Y150_SLICE_X5Y150_C3 = CLBLL_L_X4Y150_SLICE_X4Y150_B5Q;
  assign CLBLL_L_X4Y150_SLICE_X5Y150_C4 = CLBLM_R_X5Y152_SLICE_X6Y152_CQ;
  assign CLBLL_L_X4Y150_SLICE_X5Y150_C5 = CLBLM_R_X5Y152_SLICE_X6Y152_DQ;
  assign CLBLL_L_X4Y150_SLICE_X5Y150_C6 = 1'b1;
  assign CLBLM_R_X7Y150_SLICE_X9Y150_C6 = CLBLM_R_X7Y149_SLICE_X8Y149_AQ;
  assign CLBLM_R_X11Y148_SLICE_X14Y148_B1 = CLBLM_L_X10Y148_SLICE_X12Y148_CO6;
  assign CLBLL_L_X4Y150_SLICE_X5Y150_CLK = CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O;
  assign CLBLM_R_X11Y148_SLICE_X14Y148_B2 = CLBLM_L_X8Y148_SLICE_X10Y148_DO6;
  assign CLBLM_R_X11Y148_SLICE_X14Y148_B3 = CLBLM_L_X10Y145_SLICE_X12Y145_DO6;
  assign LIOI3_SING_X0Y149_OLOGIC_X0Y149_D1 = RIOB33_X105Y115_IOB_X1Y115_I;
  assign RIOI3_X105Y135_ILOGIC_X1Y136_D = RIOB33_X105Y135_IOB_X1Y136_I;
  assign CLBLL_L_X4Y150_SLICE_X5Y150_D1 = CLBLL_L_X4Y145_SLICE_X5Y145_BQ;
  assign CLBLL_L_X4Y150_SLICE_X5Y150_D2 = CLBLM_R_X3Y151_SLICE_X3Y151_CQ;
  assign CLBLL_L_X4Y150_SLICE_X5Y150_D3 = 1'b1;
  assign CLBLL_L_X4Y150_SLICE_X5Y150_D4 = CLBLM_R_X5Y152_SLICE_X6Y152_CQ;
  assign CLBLL_L_X4Y150_SLICE_X5Y150_D5 = 1'b1;
  assign CLBLL_L_X4Y150_SLICE_X5Y150_D6 = CLBLM_R_X3Y151_SLICE_X3Y151_BQ;
  assign CLBLM_R_X11Y148_SLICE_X14Y148_B4 = CLBLM_L_X12Y147_SLICE_X16Y147_DO6;
  assign LIOI3_SING_X0Y149_OLOGIC_X0Y149_T1 = 1'b1;
  assign RIOI3_X105Y135_ILOGIC_X1Y135_D = RIOB33_X105Y135_IOB_X1Y135_I;
  assign CLBLM_R_X11Y148_SLICE_X14Y148_B6 = CLBLM_R_X11Y144_SLICE_X14Y144_DO6;
  assign CLBLM_L_X10Y154_SLICE_X13Y154_A1 = CLBLM_L_X10Y154_SLICE_X13Y154_DO6;
  assign CLBLM_L_X10Y154_SLICE_X13Y154_A2 = 1'b1;
  assign CLBLM_L_X10Y154_SLICE_X13Y154_A3 = CLBLM_L_X10Y154_SLICE_X13Y154_AQ;
  assign CLBLM_L_X10Y154_SLICE_X13Y154_A4 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_L_X10Y154_SLICE_X13Y154_A5 = CLBLM_L_X10Y154_SLICE_X13Y154_CO5;
  assign CLBLM_L_X10Y154_SLICE_X13Y154_A6 = CLBLM_L_X8Y145_SLICE_X11Y145_CQ;
  assign CLBLM_L_X10Y154_SLICE_X13Y154_B1 = CLBLM_L_X10Y154_SLICE_X13Y154_AQ;
  assign CLBLM_L_X10Y154_SLICE_X13Y154_B2 = CLBLM_L_X10Y155_SLICE_X13Y155_AO6;
  assign CLBLM_L_X10Y154_SLICE_X13Y154_B3 = CLBLM_L_X10Y154_SLICE_X12Y154_A5Q;
  assign CLBLM_L_X10Y154_SLICE_X13Y154_B4 = CLBLM_L_X10Y154_SLICE_X12Y154_BQ;
  assign CLBLM_L_X10Y154_SLICE_X13Y154_B5 = CLBLM_L_X10Y154_SLICE_X12Y154_AQ;
  assign CLBLM_L_X10Y154_SLICE_X13Y154_B6 = 1'b1;
  assign CLBLM_L_X8Y144_SLICE_X11Y144_A1 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_L_X8Y144_SLICE_X11Y144_A2 = CLBLM_R_X7Y146_SLICE_X9Y146_AQ;
  assign CLBLM_L_X8Y144_SLICE_X11Y144_A3 = CLBLM_L_X8Y144_SLICE_X11Y144_AQ;
  assign CLBLM_L_X10Y154_SLICE_X13Y154_C4 = CLBLM_L_X10Y155_SLICE_X13Y155_CO6;
  assign CLBLM_L_X10Y154_SLICE_X13Y154_C5 = CLBLM_L_X10Y154_SLICE_X13Y154_AQ;
  assign CLBLM_L_X10Y154_SLICE_X13Y154_C6 = 1'b1;
  assign CLBLM_L_X8Y144_SLICE_X11Y144_A4 = CLBLM_L_X10Y143_SLICE_X13Y143_DO6;
  assign CLBLM_L_X8Y144_SLICE_X11Y144_A5 = CLBLM_L_X10Y144_SLICE_X12Y144_AO6;
  assign CLBLM_L_X8Y144_SLICE_X11Y144_A6 = 1'b1;
  assign CLBLM_L_X10Y154_SLICE_X13Y154_C1 = CLBLM_L_X10Y154_SLICE_X12Y154_AQ;
  assign CLBLM_L_X10Y154_SLICE_X13Y154_C2 = CLBLM_L_X10Y154_SLICE_X12Y154_A5Q;
  assign CLBLM_L_X8Y144_SLICE_X11Y144_B1 = CLBLM_L_X10Y142_SLICE_X12Y142_AQ;
  assign CLBLM_L_X8Y144_SLICE_X11Y144_B2 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_L_X8Y144_SLICE_X11Y144_B3 = CLBLM_R_X7Y143_SLICE_X9Y143_AQ;
  assign CLBLM_L_X8Y144_SLICE_X11Y144_B4 = 1'b1;
  assign CLBLM_L_X10Y154_SLICE_X13Y154_D2 = CLBLM_L_X10Y154_SLICE_X12Y154_A5Q;
  assign CLBLM_L_X8Y144_SLICE_X11Y144_B5 = CLBLM_L_X10Y149_SLICE_X13Y149_AQ;
  assign CLBLM_L_X8Y144_SLICE_X11Y144_B6 = 1'b1;
  assign CLBLM_L_X10Y154_SLICE_X13Y154_D5 = CLBLM_L_X10Y153_SLICE_X13Y153_CQ;
  assign CLBLM_L_X10Y154_SLICE_X13Y154_D6 = CLBLM_L_X10Y154_SLICE_X12Y154_BQ;
  assign CLBLM_L_X10Y154_SLICE_X13Y154_D1 = CLBLM_L_X10Y154_SLICE_X12Y154_AQ;
  assign CLBLM_L_X8Y144_SLICE_X11Y144_C1 = CLBLL_L_X4Y142_SLICE_X5Y142_AQ;
  assign CLBLM_L_X8Y144_SLICE_X11Y144_C2 = CLBLM_L_X8Y144_SLICE_X11Y144_CQ;
  assign CLBLM_L_X8Y144_SLICE_X11Y144_C3 = CLBLM_R_X13Y149_SLICE_X18Y149_AO6;
  assign CLBLM_L_X8Y144_SLICE_X11Y144_C4 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_L_X8Y144_SLICE_X11Y144_C5 = CLBLM_L_X10Y146_SLICE_X12Y146_DQ;
  assign CLBLM_L_X8Y144_SLICE_X11Y144_C6 = 1'b1;
  assign CLBLM_L_X8Y144_SLICE_X11Y144_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X10Y154_SLICE_X12Y154_A1 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_L_X10Y154_SLICE_X12Y154_A2 = CLBLM_L_X10Y154_SLICE_X13Y154_BO6;
  assign CLBLM_L_X10Y154_SLICE_X12Y154_A3 = CLBLM_L_X10Y154_SLICE_X12Y154_AQ;
  assign CLBLM_L_X10Y154_SLICE_X12Y154_A4 = CLBLM_L_X10Y155_SLICE_X13Y155_CO6;
  assign CLBLM_L_X10Y154_SLICE_X12Y154_A5 = CLBLM_R_X7Y154_SLICE_X9Y154_BQ;
  assign CLBLM_L_X8Y144_SLICE_X11Y144_D1 = CLBLM_L_X8Y142_SLICE_X11Y142_BQ;
  assign CLBLM_L_X8Y144_SLICE_X11Y144_D2 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_L_X8Y144_SLICE_X11Y144_D3 = CLBLM_L_X8Y144_SLICE_X11Y144_DQ;
  assign CLBLM_L_X8Y144_SLICE_X11Y144_D4 = CLBLM_R_X7Y142_SLICE_X9Y142_AQ;
  assign CLBLM_L_X8Y144_SLICE_X11Y144_D5 = 1'b1;
  assign CLBLM_L_X10Y154_SLICE_X12Y154_B5 = CLBLM_L_X10Y154_SLICE_X12Y154_A5Q;
  assign CLBLM_L_X10Y154_SLICE_X12Y154_B6 = CLBLM_L_X10Y155_SLICE_X13Y155_CO6;
  assign CLBLM_L_X8Y144_SLICE_X11Y144_D6 = CLBLM_L_X12Y149_SLICE_X17Y149_CO6;
  assign CLBLM_L_X10Y154_SLICE_X12Y154_AX = CLBLM_L_X10Y154_SLICE_X12Y154_CO6;
  assign CLBLM_L_X10Y154_SLICE_X12Y154_B1 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_L_X10Y154_SLICE_X12Y154_B2 = CLBLM_L_X10Y154_SLICE_X12Y154_BQ;
  assign CLBLM_L_X10Y154_SLICE_X12Y154_B3 = CLBLM_R_X7Y152_SLICE_X8Y152_B5Q;
  assign CLBLM_L_X10Y154_SLICE_X12Y154_B4 = CLBLM_L_X10Y155_SLICE_X13Y155_BO6;
  assign CLBLM_L_X8Y144_SLICE_X10Y144_A1 = CLBLM_R_X5Y145_SLICE_X7Y145_B5Q;
  assign CLBLM_L_X10Y154_SLICE_X12Y154_C4 = CLBLM_L_X10Y154_SLICE_X12Y154_A5Q;
  assign CLBLM_L_X10Y154_SLICE_X12Y154_C5 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_L_X10Y154_SLICE_X12Y154_C6 = 1'b1;
  assign CLBLM_L_X8Y144_SLICE_X10Y144_A2 = 1'b1;
  assign CLBLM_L_X8Y144_SLICE_X10Y144_A3 = CLBLM_R_X3Y142_SLICE_X2Y142_BO5;
  assign CLBLM_L_X8Y144_SLICE_X10Y144_A4 = CLBLM_L_X8Y143_SLICE_X10Y143_AQ;
  assign CLBLM_L_X8Y144_SLICE_X10Y144_A5 = CLBLM_L_X10Y144_SLICE_X13Y144_A5Q;
  assign CLBLM_L_X8Y144_SLICE_X10Y144_A6 = 1'b1;
  assign CLBLM_L_X8Y144_SLICE_X10Y144_AX = CLBLM_R_X7Y144_SLICE_X8Y144_DQ;
  assign CLBLM_L_X8Y144_SLICE_X10Y144_B1 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_L_X8Y144_SLICE_X10Y144_B2 = CLBLM_L_X12Y151_SLICE_X16Y151_AQ;
  assign CLBLM_L_X8Y144_SLICE_X10Y144_B3 = CLBLM_L_X10Y149_SLICE_X12Y149_BQ;
  assign CLBLM_L_X8Y144_SLICE_X10Y144_B4 = CLBLM_L_X10Y151_SLICE_X13Y151_AQ;
  assign CLBLM_L_X8Y144_SLICE_X10Y144_B5 = CLBLM_R_X3Y146_SLICE_X2Y146_D5Q;
  assign CLBLM_L_X8Y144_SLICE_X10Y144_B6 = 1'b1;
  assign CLBLM_L_X10Y154_SLICE_X12Y154_CLK = CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O;
  assign CLBLM_L_X10Y154_SLICE_X12Y154_D5 = CLBLM_L_X10Y154_SLICE_X12Y154_BQ;
  assign CLBLM_L_X10Y154_SLICE_X12Y154_D1 = RIOB33_X105Y131_IOB_X1Y131_I;
  assign CLBLM_L_X8Y144_SLICE_X10Y144_BX = CLBLM_R_X7Y142_SLICE_X9Y142_AQ;
  assign CLBLM_L_X10Y154_SLICE_X12Y154_D2 = CLBLM_R_X5Y142_SLICE_X7Y142_CO6;
  assign CLBLM_L_X8Y144_SLICE_X10Y144_C1 = CLBLM_R_X7Y144_SLICE_X8Y144_CQ;
  assign CLBLM_L_X8Y144_SLICE_X10Y144_C2 = CLBLM_R_X7Y146_SLICE_X9Y146_DO6;
  assign CLBLM_L_X8Y144_SLICE_X10Y144_C3 = CLBLM_R_X11Y144_SLICE_X14Y144_BO6;
  assign CLBLM_L_X8Y144_SLICE_X10Y144_C4 = CLBLM_R_X7Y153_SLICE_X8Y153_A5Q;
  assign CLBLM_L_X8Y144_SLICE_X10Y144_C5 = CLBLL_L_X4Y144_SLICE_X4Y144_DQ;
  assign CLBLM_L_X8Y144_SLICE_X10Y144_C6 = CLBLM_R_X7Y144_SLICE_X9Y144_B5Q;
  assign CLBLM_L_X8Y144_SLICE_X10Y144_CE = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_L_X8Y144_SLICE_X10Y144_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X8Y144_SLICE_X10Y144_D1 = CLBLM_L_X8Y143_SLICE_X11Y143_BQ;
  assign CLBLM_L_X8Y144_SLICE_X10Y144_D2 = CLBLM_R_X7Y153_SLICE_X8Y153_A5Q;
  assign CLBLM_L_X8Y144_SLICE_X10Y144_D3 = CLBLM_L_X8Y144_SLICE_X11Y144_B5Q;
  assign CLBLM_L_X8Y144_SLICE_X10Y144_D4 = CLBLM_R_X11Y144_SLICE_X14Y144_AO6;
  assign CLBLM_L_X8Y144_SLICE_X10Y144_D5 = CLBLM_R_X11Y144_SLICE_X14Y144_CO6;
  assign CLBLM_L_X8Y144_SLICE_X10Y144_D6 = CLBLM_R_X7Y144_SLICE_X9Y144_B5Q;
  assign LIOB33_X0Y145_IOB_X0Y146_O = CLBLM_R_X3Y143_SLICE_X3Y143_DO6;
  assign LIOB33_X0Y145_IOB_X0Y145_O = CLBLM_R_X3Y148_SLICE_X3Y148_DO6;
  assign CLBLM_R_X5Y152_SLICE_X7Y152_C4 = CLBLM_R_X5Y152_SLICE_X7Y152_A5Q;
  assign CLBLM_R_X5Y152_SLICE_X7Y152_C5 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X5Y152_SLICE_X7Y152_C6 = 1'b1;
  assign CLBLM_R_X11Y148_SLICE_X15Y148_A1 = CLBLM_R_X7Y153_SLICE_X8Y153_A5Q;
  assign CLBLM_R_X11Y148_SLICE_X15Y148_A2 = CLBLM_R_X7Y149_SLICE_X8Y149_AQ;
  assign CLBLM_R_X11Y148_SLICE_X15Y148_A3 = CLBLM_R_X7Y144_SLICE_X9Y144_B5Q;
  assign CLBLM_R_X11Y148_SLICE_X15Y148_A4 = CLBLL_L_X4Y148_SLICE_X4Y148_CQ;
  assign CLBLM_R_X11Y148_SLICE_X15Y148_A5 = CLBLM_L_X12Y147_SLICE_X16Y147_DO6;
  assign CLBLM_R_X11Y148_SLICE_X15Y148_A6 = CLBLM_L_X10Y146_SLICE_X13Y146_DO6;
  assign CLBLM_L_X10Y152_SLICE_X12Y152_C4 = CLBLM_R_X13Y149_SLICE_X18Y149_AO6;
  assign CLBLM_R_X7Y150_SLICE_X8Y150_B6 = 1'b1;
  assign CLBLM_R_X11Y148_SLICE_X15Y148_B1 = CLBLM_L_X12Y147_SLICE_X17Y147_DO6;
  assign CLBLM_R_X11Y148_SLICE_X15Y148_B2 = CLBLM_R_X11Y144_SLICE_X14Y144_DO6;
  assign CLBLM_R_X11Y148_SLICE_X15Y148_B3 = CLBLM_L_X12Y147_SLICE_X16Y147_CO6;
  assign CLBLM_R_X11Y148_SLICE_X15Y148_B4 = CLBLM_R_X13Y146_SLICE_X18Y146_BO6;
  assign CLBLM_R_X11Y148_SLICE_X15Y148_B5 = CLBLM_R_X3Y145_SLICE_X2Y145_AQ;
  assign CLBLM_R_X11Y148_SLICE_X15Y148_B6 = CLBLM_L_X12Y145_SLICE_X16Y145_BO6;
  assign CLBLM_R_X11Y148_SLICE_X15Y148_C1 = CLBLM_L_X12Y148_SLICE_X17Y148_AO6;
  assign CLBLM_R_X11Y148_SLICE_X15Y148_C2 = CLBLM_R_X11Y144_SLICE_X14Y144_DO6;
  assign CLBLM_R_X11Y148_SLICE_X15Y148_C3 = CLBLM_L_X10Y151_SLICE_X12Y151_AQ;
  assign CLBLM_R_X11Y148_SLICE_X15Y148_C4 = CLBLM_L_X12Y148_SLICE_X16Y148_DO6;
  assign CLBLM_R_X11Y148_SLICE_X15Y148_C5 = CLBLM_L_X12Y145_SLICE_X16Y145_BO6;
  assign CLBLM_R_X11Y148_SLICE_X15Y148_C6 = CLBLM_R_X13Y146_SLICE_X18Y146_BO6;
  assign CLBLL_L_X4Y151_SLICE_X4Y151_A1 = 1'b1;
  assign CLBLL_L_X4Y151_SLICE_X4Y151_A2 = CLBLM_R_X3Y145_SLICE_X2Y145_CQ;
  assign CLBLL_L_X4Y151_SLICE_X4Y151_A3 = CLBLL_L_X4Y151_SLICE_X4Y151_AQ;
  assign CLBLL_L_X4Y151_SLICE_X4Y151_A4 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLL_L_X4Y151_SLICE_X4Y151_A5 = CLBLL_L_X4Y143_SLICE_X5Y143_CO5;
  assign CLBLL_L_X4Y151_SLICE_X4Y151_A6 = CLBLL_L_X4Y150_SLICE_X4Y150_A5Q;
  assign CLBLM_R_X11Y148_SLICE_X15Y148_D1 = CLBLM_R_X11Y147_SLICE_X15Y147_CO6;
  assign CLBLL_L_X4Y151_SLICE_X4Y151_AX = CLBLM_R_X3Y151_SLICE_X3Y151_DO6;
  assign CLBLM_R_X5Y152_SLICE_X7Y152_D1 = CLBLM_R_X3Y146_SLICE_X3Y146_AQ;
  assign CLBLL_L_X4Y151_SLICE_X4Y151_B1 = CLBLM_R_X3Y151_SLICE_X3Y151_A5Q;
  assign CLBLL_L_X4Y151_SLICE_X4Y151_B2 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLL_L_X4Y151_SLICE_X4Y151_B3 = CLBLM_L_X10Y153_SLICE_X13Y153_A5Q;
  assign CLBLL_L_X4Y151_SLICE_X4Y151_B4 = 1'b1;
  assign CLBLL_L_X4Y151_SLICE_X4Y151_B5 = RIOB33_X105Y107_IOB_X1Y107_I;
  assign CLBLL_L_X4Y151_SLICE_X4Y151_B6 = 1'b1;
  assign CLBLM_R_X5Y152_SLICE_X7Y152_D2 = CLBLM_R_X5Y151_SLICE_X7Y151_CO6;
  assign CLBLM_R_X11Y148_SLICE_X15Y148_D4 = CLBLM_R_X11Y150_SLICE_X15Y150_CO6;
  assign CLBLM_R_X5Y152_SLICE_X7Y152_D3 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLL_L_X4Y151_SLICE_X4Y151_C1 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLL_L_X4Y151_SLICE_X4Y151_C2 = CLBLL_L_X4Y143_SLICE_X4Y143_AQ;
  assign CLBLL_L_X4Y151_SLICE_X4Y151_C3 = CLBLM_R_X3Y147_SLICE_X3Y147_CQ;
  assign CLBLL_L_X4Y151_SLICE_X4Y151_C4 = CLBLM_L_X10Y150_SLICE_X12Y150_AQ;
  assign CLBLL_L_X4Y151_SLICE_X4Y151_C5 = CLBLM_R_X5Y152_SLICE_X7Y152_DQ;
  assign CLBLL_L_X4Y151_SLICE_X4Y151_C6 = 1'b1;
  assign CLBLM_R_X7Y150_SLICE_X8Y150_C4 = CLBLM_L_X10Y146_SLICE_X13Y146_DO6;
  assign CLBLM_R_X11Y148_SLICE_X14Y148_A1 = CLBLM_R_X7Y147_SLICE_X8Y147_DO6;
  assign CLBLM_L_X10Y152_SLICE_X12Y152_C6 = 1'b1;
  assign CLBLL_L_X4Y151_SLICE_X4Y151_CLK = CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O;
  assign CLBLM_R_X7Y150_SLICE_X8Y150_C5 = CLBLM_R_X7Y150_SLICE_X8Y150_DO6;
  assign CLBLM_R_X11Y148_SLICE_X14Y148_A5 = CLBLM_L_X12Y147_SLICE_X16Y147_DO6;
  assign CLBLM_R_X11Y148_SLICE_X14Y148_A6 = CLBLM_R_X7Y149_SLICE_X8Y149_CO6;
  assign CLBLL_L_X4Y151_SLICE_X4Y151_D1 = CLBLL_L_X4Y142_SLICE_X4Y142_AQ;
  assign CLBLL_L_X4Y151_SLICE_X4Y151_D2 = CLBLM_L_X12Y151_SLICE_X16Y151_AQ;
  assign CLBLL_L_X4Y151_SLICE_X4Y151_D3 = CLBLM_R_X3Y143_SLICE_X3Y143_BQ;
  assign CLBLL_L_X4Y151_SLICE_X4Y151_D4 = CLBLL_L_X4Y152_SLICE_X4Y152_AQ;
  assign CLBLL_L_X4Y151_SLICE_X4Y151_D5 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLL_L_X4Y151_SLICE_X4Y151_D6 = CLBLM_R_X7Y153_SLICE_X8Y153_CQ;
  assign CLBLM_R_X7Y150_SLICE_X8Y150_C6 = CLBLM_L_X10Y150_SLICE_X12Y150_BO6;
  assign CLBLM_R_X11Y148_SLICE_X14Y148_B5 = CLBLM_L_X12Y146_SLICE_X16Y146_DO6;
  assign CLBLM_R_X11Y148_SLICE_X14Y148_C1 = CLBLM_R_X13Y146_SLICE_X18Y146_BO6;
  assign CLBLM_R_X11Y148_SLICE_X14Y148_C2 = CLBLM_L_X12Y145_SLICE_X16Y145_BO6;
  assign CLBLM_R_X11Y148_SLICE_X14Y148_C3 = CLBLM_R_X3Y145_SLICE_X2Y145_AQ;
  assign CLBLM_R_X11Y148_SLICE_X14Y148_C4 = CLBLM_L_X12Y147_SLICE_X17Y147_BO6;
  assign CLBLM_R_X11Y148_SLICE_X14Y148_C5 = CLBLM_L_X10Y147_SLICE_X12Y147_DO6;
  assign CLBLM_R_X11Y148_SLICE_X14Y148_C6 = CLBLM_R_X11Y144_SLICE_X14Y144_DO6;
  assign CLBLM_R_X11Y148_SLICE_X14Y148_D1 = CLBLM_L_X12Y148_SLICE_X16Y148_BO6;
  assign CLBLM_R_X11Y148_SLICE_X14Y148_D2 = CLBLM_R_X13Y146_SLICE_X18Y146_BO6;
  assign CLBLM_R_X11Y148_SLICE_X14Y148_D3 = CLBLM_L_X10Y151_SLICE_X12Y151_AQ;
  assign CLBLM_R_X11Y148_SLICE_X14Y148_D4 = CLBLM_L_X12Y145_SLICE_X16Y145_BO6;
  assign CLBLM_R_X11Y148_SLICE_X14Y148_D5 = CLBLM_L_X8Y148_SLICE_X10Y148_CO6;
  assign CLBLM_R_X11Y148_SLICE_X14Y148_D6 = CLBLM_R_X11Y144_SLICE_X14Y144_DO6;
  assign CLBLL_L_X4Y151_SLICE_X5Y151_A1 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLL_L_X4Y151_SLICE_X5Y151_A2 = CLBLL_L_X4Y151_SLICE_X5Y151_DQ;
  assign CLBLL_L_X4Y151_SLICE_X5Y151_A3 = CLBLL_L_X4Y151_SLICE_X5Y151_AQ;
  assign CLBLL_L_X4Y151_SLICE_X5Y151_A4 = CLBLM_R_X7Y150_SLICE_X8Y150_AQ;
  assign CLBLL_L_X4Y151_SLICE_X5Y151_A5 = CLBLM_R_X7Y152_SLICE_X8Y152_D5Q;
  assign CLBLL_L_X4Y151_SLICE_X5Y151_A6 = CLBLM_R_X7Y142_SLICE_X8Y142_C5Q;
  assign CLBLL_L_X4Y151_SLICE_X5Y151_B1 = CLBLL_L_X4Y145_SLICE_X5Y145_AQ;
  assign CLBLL_L_X4Y151_SLICE_X5Y151_B2 = CLBLL_L_X4Y145_SLICE_X5Y145_BQ;
  assign CLBLL_L_X4Y151_SLICE_X5Y151_B3 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLL_L_X4Y151_SLICE_X5Y151_B4 = CLBLL_L_X4Y146_SLICE_X4Y146_CQ;
  assign CLBLL_L_X4Y151_SLICE_X5Y151_B5 = CLBLM_L_X10Y153_SLICE_X13Y153_A5Q;
  assign CLBLL_L_X4Y151_SLICE_X5Y151_B6 = 1'b1;
  assign CLBLL_L_X4Y151_SLICE_X5Y151_C1 = CLBLL_L_X4Y151_SLICE_X4Y151_AQ;
  assign CLBLL_L_X4Y151_SLICE_X5Y151_C2 = CLBLL_L_X4Y151_SLICE_X5Y151_CQ;
  assign CLBLL_L_X4Y151_SLICE_X5Y151_C3 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLL_L_X4Y151_SLICE_X5Y151_C4 = CLBLM_R_X3Y145_SLICE_X2Y145_CQ;
  assign CLBLL_L_X4Y151_SLICE_X5Y151_C5 = CLBLL_L_X4Y151_SLICE_X5Y151_B5Q;
  assign CLBLL_L_X4Y151_SLICE_X5Y151_C6 = CLBLL_L_X4Y143_SLICE_X5Y143_CO5;
  assign CLBLL_L_X4Y151_SLICE_X5Y151_CLK = CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O;
  assign CLBLM_R_X3Y143_SLICE_X2Y143_A4 = CLBLM_L_X10Y144_SLICE_X12Y144_AO6;
  assign CLBLL_L_X4Y151_SLICE_X5Y151_D1 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLL_L_X4Y151_SLICE_X5Y151_D2 = CLBLM_R_X5Y144_SLICE_X7Y144_CQ;
  assign CLBLL_L_X4Y151_SLICE_X5Y151_D3 = CLBLL_L_X4Y151_SLICE_X5Y151_DQ;
  assign CLBLL_L_X4Y151_SLICE_X5Y151_D4 = CLBLM_R_X3Y151_SLICE_X3Y151_BQ;
  assign CLBLL_L_X4Y151_SLICE_X5Y151_D5 = CLBLM_R_X3Y149_SLICE_X2Y149_C5Q;
  assign CLBLL_L_X4Y151_SLICE_X5Y151_D6 = 1'b1;
  assign CLBLM_R_X7Y150_SLICE_X8Y150_D5 = CLBLM_R_X7Y144_SLICE_X8Y144_D5Q;
  assign CLBLM_R_X3Y143_SLICE_X2Y143_A5 = CLBLM_R_X3Y143_SLICE_X2Y143_CO5;
  assign CLBLM_L_X10Y155_SLICE_X13Y155_A1 = CLBLM_R_X5Y147_SLICE_X6Y147_AQ;
  assign CLBLM_L_X10Y155_SLICE_X13Y155_A2 = CLBLM_R_X7Y146_SLICE_X8Y146_A5Q;
  assign CLBLM_L_X10Y155_SLICE_X13Y155_A3 = CLBLM_R_X11Y153_SLICE_X15Y153_DO6;
  assign CLBLM_L_X10Y155_SLICE_X13Y155_A4 = CLBLM_L_X10Y153_SLICE_X13Y153_BQ;
  assign CLBLM_L_X10Y155_SLICE_X13Y155_A5 = CLBLM_L_X10Y155_SLICE_X12Y155_AQ;
  assign CLBLM_L_X10Y155_SLICE_X13Y155_A6 = 1'b1;
  assign CLBLM_L_X10Y155_SLICE_X13Y155_B1 = CLBLM_L_X10Y154_SLICE_X12Y154_A5Q;
  assign CLBLM_L_X10Y155_SLICE_X13Y155_B2 = CLBLM_L_X10Y153_SLICE_X13Y153_BQ;
  assign CLBLM_L_X10Y155_SLICE_X13Y155_B3 = CLBLM_R_X11Y153_SLICE_X15Y153_DO6;
  assign CLBLM_L_X10Y155_SLICE_X13Y155_B4 = CLBLM_L_X10Y155_SLICE_X12Y155_BO5;
  assign CLBLM_L_X10Y155_SLICE_X13Y155_B5 = CLBLM_L_X10Y155_SLICE_X12Y155_AQ;
  assign CLBLM_L_X10Y155_SLICE_X13Y155_B6 = CLBLM_L_X10Y155_SLICE_X13Y155_AO5;
  assign CLBLM_R_X3Y143_SLICE_X2Y143_A6 = 1'b1;
  assign CLBLM_R_X5Y152_SLICE_X6Y152_B5 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X5Y152_SLICE_X6Y152_B6 = 1'b1;
  assign CLBLM_L_X8Y145_SLICE_X11Y145_A1 = CLBLM_R_X7Y145_SLICE_X8Y145_D5Q;
  assign CLBLM_L_X8Y145_SLICE_X11Y145_A2 = CLBLM_R_X7Y152_SLICE_X8Y152_D5Q;
  assign CLBLM_L_X8Y145_SLICE_X11Y145_A3 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_L_X10Y155_SLICE_X13Y155_C4 = CLBLM_L_X10Y153_SLICE_X13Y153_BQ;
  assign CLBLM_L_X10Y155_SLICE_X13Y155_C5 = CLBLM_R_X11Y153_SLICE_X15Y153_DO6;
  assign CLBLM_L_X10Y155_SLICE_X13Y155_C6 = CLBLM_R_X7Y146_SLICE_X8Y146_A5Q;
  assign CLBLM_L_X8Y145_SLICE_X11Y145_A4 = CLBLM_L_X8Y145_SLICE_X11Y145_AQ;
  assign CLBLM_L_X8Y145_SLICE_X11Y145_A5 = CLBLM_R_X7Y142_SLICE_X8Y142_C5Q;
  assign CLBLM_L_X8Y145_SLICE_X11Y145_A6 = CLBLM_L_X8Y145_SLICE_X10Y145_AQ;
  assign CLBLM_L_X10Y155_SLICE_X13Y155_C1 = CLBLM_L_X10Y155_SLICE_X12Y155_AQ;
  assign CLBLM_L_X10Y155_SLICE_X13Y155_C2 = CLBLM_L_X10Y153_SLICE_X13Y153_CQ;
  assign CLBLM_L_X8Y145_SLICE_X11Y145_B1 = CLBLM_L_X10Y144_SLICE_X13Y144_CQ;
  assign CLBLM_L_X8Y145_SLICE_X11Y145_B2 = CLBLM_L_X8Y145_SLICE_X11Y145_BQ;
  assign CLBLM_L_X8Y145_SLICE_X11Y145_B3 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_L_X8Y145_SLICE_X11Y145_B4 = CLBLL_L_X4Y146_SLICE_X5Y146_BQ;
  assign CLBLM_L_X8Y145_SLICE_X11Y145_B5 = CLBLM_L_X8Y147_SLICE_X10Y147_C5Q;
  assign CLBLM_L_X8Y145_SLICE_X11Y145_B6 = CLBLM_R_X3Y145_SLICE_X3Y145_DQ;
  assign CLBLM_L_X10Y155_SLICE_X13Y155_D5 = 1'b1;
  assign CLBLM_L_X10Y155_SLICE_X13Y155_D6 = 1'b1;
  assign CLBLM_L_X10Y155_SLICE_X13Y155_D1 = 1'b1;
  assign CLBLM_L_X10Y155_SLICE_X13Y155_D2 = 1'b1;
  assign CLBLM_L_X8Y145_SLICE_X11Y145_C1 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_L_X8Y145_SLICE_X11Y145_C2 = CLBLM_L_X10Y149_SLICE_X13Y149_AQ;
  assign CLBLM_L_X8Y145_SLICE_X11Y145_C3 = CLBLM_L_X8Y144_SLICE_X11Y144_DQ;
  assign CLBLM_L_X8Y145_SLICE_X11Y145_C4 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_L_X8Y145_SLICE_X11Y145_C5 = CLBLM_L_X8Y153_SLICE_X10Y153_D5Q;
  assign CLBLM_L_X8Y145_SLICE_X11Y145_C6 = 1'b1;
  assign CLBLM_L_X8Y145_SLICE_X11Y145_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X10Y155_SLICE_X12Y155_A1 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_L_X10Y155_SLICE_X12Y155_A2 = CLBLM_L_X10Y155_SLICE_X12Y155_BO5;
  assign CLBLM_L_X10Y155_SLICE_X12Y155_A3 = CLBLM_L_X10Y155_SLICE_X12Y155_AQ;
  assign CLBLM_L_X10Y155_SLICE_X12Y155_A4 = CLBLM_L_X10Y155_SLICE_X12Y155_BO6;
  assign CLBLM_L_X10Y155_SLICE_X12Y155_A5 = CLBLM_L_X10Y155_SLICE_X13Y155_AO6;
  assign CLBLM_L_X8Y145_SLICE_X11Y145_D1 = CLBLM_L_X10Y144_SLICE_X12Y144_CO6;
  assign CLBLM_L_X8Y145_SLICE_X11Y145_D2 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_L_X8Y145_SLICE_X11Y145_D3 = CLBLM_L_X8Y145_SLICE_X11Y145_DQ;
  assign CLBLM_L_X8Y145_SLICE_X11Y145_D4 = 1'b1;
  assign CLBLM_L_X8Y145_SLICE_X11Y145_D5 = CLBLM_R_X7Y152_SLICE_X9Y152_DO6;
  assign CLBLM_L_X10Y155_SLICE_X12Y155_B5 = CLBLM_R_X7Y146_SLICE_X8Y146_A5Q;
  assign CLBLM_L_X10Y155_SLICE_X12Y155_B6 = 1'b1;
  assign CLBLM_L_X8Y145_SLICE_X11Y145_D6 = CLBLM_L_X8Y145_SLICE_X11Y145_AQ;
  assign CLBLM_L_X10Y155_SLICE_X12Y155_B1 = CLBLM_R_X5Y147_SLICE_X6Y147_AQ;
  assign CLBLM_L_X10Y155_SLICE_X12Y155_B2 = CLBLM_L_X10Y153_SLICE_X13Y153_BQ;
  assign CLBLM_L_X10Y155_SLICE_X12Y155_C1 = 1'b1;
  assign CLBLM_L_X10Y155_SLICE_X12Y155_C2 = 1'b1;
  assign CLBLM_L_X10Y155_SLICE_X12Y155_C3 = 1'b1;
  assign CLBLM_L_X10Y155_SLICE_X12Y155_C4 = 1'b1;
  assign CLBLM_L_X10Y155_SLICE_X12Y155_C5 = 1'b1;
  assign CLBLM_L_X8Y145_SLICE_X10Y145_A1 = CLBLM_L_X10Y143_SLICE_X12Y143_BQ;
  assign CLBLM_L_X8Y145_SLICE_X10Y145_A2 = CLBLM_L_X8Y144_SLICE_X11Y144_B5Q;
endmodule
